magic
tech sky130A
magscale 1 2
timestamp 1694038050
<< pwell >>
rect -347 -448 347 448
<< mvnmos >>
rect -129 -200 -29 200
rect 29 -200 129 200
<< mvndiff >>
rect -187 187 -129 200
rect -187 153 -175 187
rect -141 153 -129 187
rect -187 119 -129 153
rect -187 85 -175 119
rect -141 85 -129 119
rect -187 51 -129 85
rect -187 17 -175 51
rect -141 17 -129 51
rect -187 -17 -129 17
rect -187 -51 -175 -17
rect -141 -51 -129 -17
rect -187 -85 -129 -51
rect -187 -119 -175 -85
rect -141 -119 -129 -85
rect -187 -153 -129 -119
rect -187 -187 -175 -153
rect -141 -187 -129 -153
rect -187 -200 -129 -187
rect -29 187 29 200
rect -29 153 -17 187
rect 17 153 29 187
rect -29 119 29 153
rect -29 85 -17 119
rect 17 85 29 119
rect -29 51 29 85
rect -29 17 -17 51
rect 17 17 29 51
rect -29 -17 29 17
rect -29 -51 -17 -17
rect 17 -51 29 -17
rect -29 -85 29 -51
rect -29 -119 -17 -85
rect 17 -119 29 -85
rect -29 -153 29 -119
rect -29 -187 -17 -153
rect 17 -187 29 -153
rect -29 -200 29 -187
rect 129 187 187 200
rect 129 153 141 187
rect 175 153 187 187
rect 129 119 187 153
rect 129 85 141 119
rect 175 85 187 119
rect 129 51 187 85
rect 129 17 141 51
rect 175 17 187 51
rect 129 -17 187 17
rect 129 -51 141 -17
rect 175 -51 187 -17
rect 129 -85 187 -51
rect 129 -119 141 -85
rect 175 -119 187 -85
rect 129 -153 187 -119
rect 129 -187 141 -153
rect 175 -187 187 -153
rect 129 -200 187 -187
<< mvndiffc >>
rect -175 153 -141 187
rect -175 85 -141 119
rect -175 17 -141 51
rect -175 -51 -141 -17
rect -175 -119 -141 -85
rect -175 -187 -141 -153
rect -17 153 17 187
rect -17 85 17 119
rect -17 17 17 51
rect -17 -51 17 -17
rect -17 -119 17 -85
rect -17 -187 17 -153
rect 141 153 175 187
rect 141 85 175 119
rect 141 17 175 51
rect 141 -51 175 -17
rect 141 -119 175 -85
rect 141 -187 175 -153
<< mvpsubdiff >>
rect -321 410 321 422
rect -321 376 -187 410
rect -153 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 153 410
rect 187 376 321 410
rect -321 364 321 376
rect -321 -364 -263 364
rect 263 -364 321 364
rect -321 -376 321 -364
rect -321 -410 -187 -376
rect -153 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 153 -376
rect 187 -410 321 -376
rect -321 -422 321 -410
<< mvpsubdiffcont >>
rect -187 376 -153 410
rect -119 376 -85 410
rect -51 376 -17 410
rect 17 376 51 410
rect 85 376 119 410
rect 153 376 187 410
rect -187 -410 -153 -376
rect -119 -410 -85 -376
rect -51 -410 -17 -376
rect 17 -410 51 -376
rect 85 -410 119 -376
rect 153 -410 187 -376
<< poly >>
rect -129 272 -29 288
rect -129 238 -96 272
rect -62 238 -29 272
rect -129 200 -29 238
rect 29 272 129 288
rect 29 238 62 272
rect 96 238 129 272
rect 29 200 129 238
rect -129 -238 -29 -200
rect -129 -272 -96 -238
rect -62 -272 -29 -238
rect -129 -288 -29 -272
rect 29 -238 129 -200
rect 29 -272 62 -238
rect 96 -272 129 -238
rect 29 -288 129 -272
<< polycont >>
rect -96 238 -62 272
rect 62 238 96 272
rect -96 -272 -62 -238
rect 62 -272 96 -238
<< locali >>
rect -309 376 -187 410
rect -153 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 153 410
rect 187 376 309 410
rect -309 -376 -275 376
rect -129 238 -96 272
rect -62 238 -29 272
rect 29 238 62 272
rect 96 238 129 272
rect -175 187 -141 204
rect -175 119 -141 127
rect -175 51 -141 55
rect -175 -55 -141 -51
rect -175 -127 -141 -119
rect -175 -204 -141 -187
rect -17 187 17 204
rect -17 119 17 127
rect -17 51 17 55
rect -17 -55 17 -51
rect -17 -127 17 -119
rect -17 -204 17 -187
rect 141 187 175 204
rect 141 119 175 127
rect 141 51 175 55
rect 141 -55 175 -51
rect 141 -127 175 -119
rect 141 -204 175 -187
rect -129 -272 -96 -238
rect -62 -272 -29 -238
rect 29 -272 62 -238
rect 96 -272 129 -238
rect 275 -376 309 376
rect -309 -410 -187 -376
rect -153 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 153 -376
rect 187 -410 309 -376
<< viali >>
rect -96 238 -62 272
rect 62 238 96 272
rect -175 153 -141 161
rect -175 127 -141 153
rect -175 85 -141 89
rect -175 55 -141 85
rect -175 -17 -141 17
rect -175 -85 -141 -55
rect -175 -89 -141 -85
rect -175 -153 -141 -127
rect -175 -161 -141 -153
rect -17 153 17 161
rect -17 127 17 153
rect -17 85 17 89
rect -17 55 17 85
rect -17 -17 17 17
rect -17 -85 17 -55
rect -17 -89 17 -85
rect -17 -153 17 -127
rect -17 -161 17 -153
rect 141 153 175 161
rect 141 127 175 153
rect 141 85 175 89
rect 141 55 175 85
rect 141 -17 175 17
rect 141 -85 175 -55
rect 141 -89 175 -85
rect 141 -153 175 -127
rect 141 -161 175 -153
rect -96 -272 -62 -238
rect 62 -272 96 -238
<< metal1 >>
rect -125 272 -33 278
rect -125 238 -96 272
rect -62 238 -33 272
rect -125 232 -33 238
rect 33 272 125 278
rect 33 238 62 272
rect 96 238 125 272
rect 33 232 125 238
rect -181 161 -135 200
rect -181 127 -175 161
rect -141 127 -135 161
rect -181 89 -135 127
rect -181 55 -175 89
rect -141 55 -135 89
rect -181 17 -135 55
rect -181 -17 -175 17
rect -141 -17 -135 17
rect -181 -55 -135 -17
rect -181 -89 -175 -55
rect -141 -89 -135 -55
rect -181 -127 -135 -89
rect -181 -161 -175 -127
rect -141 -161 -135 -127
rect -181 -200 -135 -161
rect -23 161 23 200
rect -23 127 -17 161
rect 17 127 23 161
rect -23 89 23 127
rect -23 55 -17 89
rect 17 55 23 89
rect -23 17 23 55
rect -23 -17 -17 17
rect 17 -17 23 17
rect -23 -55 23 -17
rect -23 -89 -17 -55
rect 17 -89 23 -55
rect -23 -127 23 -89
rect -23 -161 -17 -127
rect 17 -161 23 -127
rect -23 -200 23 -161
rect 135 161 181 200
rect 135 127 141 161
rect 175 127 181 161
rect 135 89 181 127
rect 135 55 141 89
rect 175 55 181 89
rect 135 17 181 55
rect 135 -17 141 17
rect 175 -17 181 17
rect 135 -55 181 -17
rect 135 -89 141 -55
rect 175 -89 181 -55
rect 135 -127 181 -89
rect 135 -161 141 -127
rect 175 -161 181 -127
rect 135 -200 181 -161
rect -125 -238 -33 -232
rect -125 -272 -96 -238
rect -62 -272 -33 -238
rect -125 -278 -33 -272
rect 33 -238 125 -232
rect 33 -272 62 -238
rect 96 -272 125 -238
rect 33 -278 125 -272
<< properties >>
string FIXED_BBOX -292 -393 292 393
<< end >>
