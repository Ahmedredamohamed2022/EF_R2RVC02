* NGSPICE file created from EF_R2RVC02.ext - technology: sky130A

.subckt EF_R2RVC02 VSS VO SELB A2 B2 B1 SELA DVSS A1 DVDD VDD
X0 a_1821_8526.t3 comparator_top_0.comparator_bias_0.VBN.t4 comparator_top_0.comparator_bias_0.VBN.t5 VDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=15
X1 VSS.t52 VSS.t51 VSS.t52 VSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X2 VSS.t50 VSS.t48 VSS.t49 VSS.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X3 a_2551_4880.t1 a_2151_4783.t8 VDD.t138 VDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 comparator_top_0.comparator_0.VOUT a_8881_1782.t2 VDD.t143 VDD.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=2
X5 a_570_n5724# a_470_n5812# DVSS.t117 DVSS.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X6 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 B1.t7 DVSS.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X7 DVSS.t74 a_570_n5724# a_1777_n6060# DVSS.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X8 VDD.t44 a_1821_8526.t6 a_2221_8623.t3 VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X9 a_2093_3714.t7 comparator_top_0.comparator_bias_0.VBP.t4 VDD.t124 VDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X10 VDD.t122 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 VDD.t121 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
D0 DVSS.t12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X11 a_6351_6657# a_10811_7187# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X12 VSS.t3 a_2151_594.t8 a_2551_620.t1 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X13 a_5299_3714.t7 comparator_top_0.VINP a_2093_3714.t3 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X14 DVSS.t187 a_3916_n5703# a_5123_n6039# DVSS.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X15 VSS.t60 comparator_top_0.comparator_bias_0.VBN.t9 a_2093_1782.t7 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X16 a_10542_n5707# a_10442_n5795# DVSS.t144 DVSS.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X17 a_2093_3714.t5 VDD.t101 VDD.t103 VDD.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X18 DVSS.t9 a_10965_3602# a_10975_4108# DVSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X19 a_7889_n6842# a_7464_n6798# DVSS.t185 DVSS.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X20 VDD.t100 VDD.t99 VDD.t100 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X21 DVSS.t175 a_10975_4108# VO.t1 DVSS.t174 sky130_fd_pr__nfet_01v8 ad=0.196 pd=2.01 as=0.196 ps=2.01 w=0.74 l=0.15
X22 DVSS.t84 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 DVSS.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X23 VDD.t9 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 VDD.t15 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X25 EF_AMUX21m_1.array_1ls_1tgm_0.l0 SELA.t0 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X26 DVSS.t183 a_7464_n6798# a_7889_n6842# DVSS.t182 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X27 DVDD.t21 EF_AMUX21m_2.array_1ls_1tgm_0.l0 a_10442_n5795# DVDD.t20 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X28 a_7464_n6798# a_7096_n5816# DVDD.t11 DVDD.t10 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_5123_n6039# DVSS.t62 DVSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X30 a_4184_n6773# a_3816_n5791# DVDD.t25 DVDD.t24 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X31 VSS.t47 VSS.t45 comparator_top_0.comparator_bias_0.VBN.t6 VSS.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X32 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 comparator_top_0.VINM DVSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=0.5
X33 a_2093_3714.t2 comparator_top_0.VINP a_5299_3714.t6 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X34 VSS.t1 a_5299_620.t8 a_8881_1782.t0 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
D1 DVSS.t47 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X35 DVSS.t14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 DVSS.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X36 a_4609_n6817# a_4184_n6773# DVSS.t72 DVSS.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X37 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_1777_n6060# VDD.t156 VDD.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X38 A1.t7 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 comparator_top_0.VINP VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X39 a_838_n6794# a_470_n5812# DVDD.t13 DVDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X40 DVSS.t60 comparator_top_0.comparator_0.VOUT a_11031_3400# DVSS.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X41 VSS.t44 VSS.t43 VSS.t44 VSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X42 VDD.t73 a_11235_n6821# a_10542_n5707# VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X43 VDD.t98 VDD.t96 VDD.t98 VDD.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X44 a_2151_594.t7 comparator_top_0.VINM a_2093_3714.t11 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
D2 DVSS.t81 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X45 comparator_top_0.comparator_bias_0.VBN.t0 a_2221_8623.t6 a_1821_8526.t0 VDD.t33 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X46 a_7464_n6798# a_7096_n5816# DVSS.t104 DVSS.t103 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVSS.t24 DVSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_11749_n6043# VDD.t116 VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X49 VDD.t109 a_570_n5724# a_1777_n6060# VDD.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X50 a_5299_1782.t7 a_5299_1782.t6 VDD.t11 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X51 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 A1.t6 VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X52 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 comparator_top_0.VINP VDD.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.32 ps=20.6 w=1 l=0.5
X53 a_7889_n6842# a_7464_n6798# DVSS.t181 DVSS.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X54 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD.t64 VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X55 comparator_top_0.comparator_0.VOUT a_8881_1782.t3 VSS.t67 VSS.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X56 EF_AMUX21m_1.array_1ls_1tgm_0.l0 SELA.t1 DVSS.t76 DVSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X57 DVSS.t46 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 DVSS.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X58 DVDD.t23 a_11271_4224# a_10975_4108# DVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.297 ps=2.77 w=1.12 l=0.15
X59 a_11271_4224# a_11031_3400# DVSS.t92 DVSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X60 B1.t5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 B1.t4 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X61 VDD.t30 a_10542_n5707# a_11749_n6043# VDD.t29 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X62 VDD.t139 a_2151_4783.t9 a_2551_4880.t0 VDD.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X63 a_2093_1782.t6 comparator_top_0.comparator_bias_0.VBN.t10 VSS.t59 VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X64 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 B2.t3 VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X65 a_838_n6794# a_470_n5812# DVSS.t115 DVSS.t114 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X66 a_2093_3714.t10 comparator_top_0.VINM a_2151_594.t6 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X67 a_11271_4224# a_10975_4108# DVDD.t28 DVDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.157 ps=1.4 w=1.12 l=0.15
X68 EF_AMUX21m_2.array_1ls_1tgm_0.l0 SELB.t0 DVDD.t9 DVDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X69 VDD.t159 a_3916_n5703# a_5123_n6039# VDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X70 a_3916_n5703# a_3816_n5791# DVSS.t173 DVSS.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X71 a_5299_1782.t3 comparator_top_0.VINP a_2093_1782.t0 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X72 VSS.t13 a_5299_3714.t8 a_5299_620.t2 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X73 DVSS.t171 a_3816_n5791# a_3916_n5703# DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X74 VDD.t95 VDD.t93 VDD.t94 VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X75 VDD.t105 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 VDD.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X76 VDD.t46 a_5299_1782.t4 a_5299_1782.t5 VDD.t45 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X77 comparator_top_0.comparator_bias_0.VBN.t3 comparator_top_0.comparator_bias_0.VBN.t2 VSS.t58 VSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X78 DVSS.t7 a_10965_3602# a_10975_4108# DVSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X79 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_5123_n6039# VDD.t75 VDD.t74 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X80 DVSS.t132 a_7196_n5728# a_8403_n6064# DVSS.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X81 a_2093_1782.t5 VSS.t41 VSS.t42 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X82 a_570_n5724# a_470_n5812# DVSS.t113 DVSS.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X83 a_10810_n6777# a_10442_n5795# DVSS.t142 DVSS.t141 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X84 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVSS.t55 DVSS.t54 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X85 a_6349_9307# a_10809_9307# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X86 A2.t5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 comparator_top_0.VINP VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X87 a_2151_4783.t3 a_2151_4783.t2 VDD.t3 VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X88 DVDD.t19 SELB.t1 EF_AMUX21m_2.array_1ls_1tgm_0.l0 DVDD.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X89 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD.t26 VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X90 a_6351_7717# a_10811_7187# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X91 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 VDD.t36 VDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X92 DVSS.t41 a_10810_n6777# a_11235_n6821# DVSS.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X93 DVSS.t179 a_7464_n6798# a_7889_n6842# DVSS.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X94 a_1821_8526.t1 a_2221_8623.t7 comparator_top_0.comparator_bias_0.VBN.t1 VDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X95 a_7889_n6842# a_7464_n6798# DVSS.t177 DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X96 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_8403_n6064# DVSS.t20 DVSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X97 B2.t5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 B2.t4 VDD.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X98 a_2093_1782.t3 comparator_top_0.VINP a_5299_1782.t2 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X99 DVSS.t189 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 DVSS.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X100 EF_AMUX21m_2.array_1ls_1tgm_0.l0 SELB.t2 DVSS.t149 DVSS.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X101 VSS.t40 VSS.t38 VSS.t40 VSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X102 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 B2.t7 DVSS.t44 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X103 DVDD.t27 a_10975_4108# VO.t0 DVDD.t26 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.4 as=0.297 ps=2.77 w=1.12 l=0.15
X104 a_2151_4783.t7 comparator_top_0.VINM a_2093_1782.t11 VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X105 A2.t7 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 A2.t6 DVSS.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X106 VDD.t111 a_2551_620.t4 a_2551_620.t5 VDD.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X107 DVSS.t91 a_11031_3400# a_10965_3602# DVSS.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X108 VSS.t64 a_5299_3714.t2 a_5299_3714.t3 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X109 a_2151_594.t5 comparator_top_0.VINM a_2093_3714.t9 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X110 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 VDD.t123 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X111 a_1263_n6838# a_838_n6794# DVSS.t161 DVSS.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X112 VDD.t92 VDD.t89 VDD.t91 VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X113 DVSS.t89 a_11031_3400# a_11271_4224# DVSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X114 a_570_n5724# a_470_n5812# DVSS.t111 DVSS.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X115 DVSS.t31 SELB.t3 EF_AMUX21m_2.array_1ls_1tgm_0.l0 DVSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X116 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD.t56 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X117 VDD.t66 a_1263_n6838# a_570_n5724# VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X118 VSS.t37 VSS.t35 VSS.t37 VSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X119 DVSS.t80 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 DVSS.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X120 VDD.t42 a_1821_8526.t7 a_2221_8623.t2 VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X121 a_6351_6657# a_1821_8526.t2 DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X122 a_11235_n6821# a_10810_n6777# DVSS.t39 DVSS.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X123 a_6349_9307# a_10811_8247# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X124 VDD.t88 VDD.t87 VDD.t88 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X125 a_2093_1782.t10 comparator_top_0.VINM a_2151_4783.t6 VSS.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X126 comparator_top_0.comparator_bias_0.VBP.t3 comparator_top_0.comparator_bias_0.VBP.t2 VDD.t113 VDD.t112 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=2
X127 VDD.t150 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 VDD.t149 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X128 a_10810_n6777# a_10442_n5795# DVDD.t17 DVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X129 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 VDD.t7 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X130 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 comparator_top_0.VINM DVSS.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X131 a_7196_n5728# a_7096_n5816# DVSS.t102 DVSS.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X132 VSS.t34 VSS.t31 VSS.t33 VSS.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
D3 DVSS.t17 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X133 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 comparator_top_0.VINM VDD.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.32 ps=20.6 w=1 l=0.5
X134 DVSS.t169 a_3816_n5791# a_3916_n5703# DVSS.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X135 A2.t1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 comparator_top_0.VINP DVSS.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X136 DVSS.t100 a_7096_n5816# a_7196_n5728# DVSS.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X137 comparator_top_0.comparator_bias_0.VBN.t7 a_2221_8623.t8 a_1821_8526.t4 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X138 VDD.t120 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 VDD.t119 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X139 DVSS.t159 a_838_n6794# a_1263_n6838# DVSS.t158 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X140 a_1263_n6838# a_838_n6794# DVSS.t157 DVSS.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X141 DVSS.t109 a_470_n5812# a_570_n5724# DVSS.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X142 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVSS.t51 DVSS.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X143 VSS.t56 comparator_top_0.comparator_bias_0.VBN.t11 a_2221_8623.t5 VSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X144 VDD.t52 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 VDD.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X145 DVSS.t37 a_10810_n6777# a_11235_n6821# DVSS.t36 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X146 a_2551_620.t3 a_2551_620.t2 VDD.t132 VDD.t129 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X147 a_2093_3714.t1 comparator_top_0.VINP a_5299_3714.t5 VDD.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X148 a_4609_n6817# a_4184_n6773# DVSS.t70 DVSS.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X149 DVDD.t5 SELA.t2 a_470_n5812# DVDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X150 a_11235_n6821# a_10810_n6777# DVSS.t35 DVSS.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X151 VSS.t68 a_2551_4880.t6 a_5299_620.t6 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X152 a_5299_620.t1 a_5299_3714.t9 VSS.t7 VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X153 VDD.t20 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 VDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X154 A1.t5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 A1.t4 DVSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X155 DVSS.t16 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 DVSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X156 A1.t3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 comparator_top_0.VINP DVSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X157 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 VDD.t50 VDD.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X158 VDD.t13 a_5299_1782.t8 a_5299_620.t0 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X159 B1.t0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 comparator_top_0.VINM VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X160 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 comparator_top_0.VINM VDD.t47 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X161 DVSS.t120 EF_AMUX21m_1.array_1ls_1tgm_0.l0 a_3816_n5791# DVSS.t119 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X162 DVSS.t98 a_7096_n5816# a_7196_n5728# DVSS.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X163 B1.t3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 B1.t2 DVSS.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X164 a_3916_n5703# a_3816_n5791# DVSS.t167 DVSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X165 a_2221_8623.t1 a_1821_8526.t8 VDD.t40 VDD.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X166 VDD.t86 VDD.t84 a_2093_3714.t4 VDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X167 a_2151_4783.t5 comparator_top_0.VINM a_2093_1782.t9 VSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X168 a_7196_n5728# a_7096_n5816# DVSS.t96 DVSS.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X169 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 A1.t2 DVSS.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X170 DVSS.t128 SELA.t3 a_470_n5812# DVSS.t127 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X171 VDD.t107 a_570_n5724# a_1263_n6838# VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X172 a_5299_620.t5 a_2551_4880.t7 VSS.t69 VSS.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X173 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 comparator_top_0.VINP VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X174 A1.t1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 A1.t0 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X175 a_1263_n6838# a_838_n6794# DVSS.t155 DVSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X176 DVSS.t107 a_470_n5812# a_570_n5724# DVSS.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X177 a_2093_3714.t8 comparator_top_0.VINM a_2151_594.t4 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X178 VDD.t54 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 VDD.t53 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X179 VDD.t28 a_10542_n5707# a_11235_n6821# VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X180 VSS.t30 VSS.t29 VSS.t30 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X181 a_11271_4224# a_11031_3400# DVSS.t88 DVSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X182 a_11235_n6821# a_10810_n6777# DVSS.t33 DVSS.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X183 DVSS.t68 a_4184_n6773# a_4609_n6817# DVSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X184 a_2151_594.t3 a_2151_594.t2 VSS.t11 VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X185 VSS.t65 a_2551_4880.t4 a_2551_4880.t5 VSS.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X186 a_10975_4108# a_10965_3602# DVSS.t5 DVSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X187 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 A2.t4 VDD.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X188 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_11749_n6043# DVSS.t78 DVSS.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X189 a_2221_8623.t4 VSS.t26 VSS.t28 VSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X190 VDD.t114 a_2551_620.t6 a_5299_620.t4 VDD.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X191 VDD.t58 a_7889_n6842# a_7196_n5728# VDD.t57 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X192 a_5299_3714.t4 comparator_top_0.VINP a_2093_3714.t0 VDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X193 B1.t6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 comparator_top_0.VINM DVSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X194 comparator_top_0.comparator_bias_0.VBP.t0 VSS.t23 VSS.t25 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X195 a_5299_3714.t1 a_5299_3714.t0 VSS.t63 VSS.t17 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X196 a_10542_n5707# a_10442_n5795# DVSS.t140 DVSS.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X197 DVSS.t26 a_10542_n5707# a_11749_n6043# DVSS.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X198 DVDD.t3 SELA.t4 EF_AMUX21m_1.array_1ls_1tgm_0.l0 DVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X199 DVDD.t1 SELB.t4 a_7096_n5816# DVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X200 a_1821_8526.t5 a_2221_8623.t9 comparator_top_0.comparator_bias_0.VBN.t8 VDD.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X201 a_10965_3602# a_11031_3400# VDD.t128 VDD.t127 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X202 a_11031_3400# comparator_top_0.comparator_0.VOUT VDD.t71 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X203 a_2093_1782.t2 comparator_top_0.VINP a_5299_1782.t1 VSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X204 a_2551_4880.t3 a_2551_4880.t2 VSS.t70 VSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X205 DVSS.t11 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 DVSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X206 DVSS.t49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 DVSS.t48 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X207 DVDD.t15 EF_AMUX21m_1.array_1ls_1tgm_0.l0 a_3816_n5791# DVDD.t14 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X208 a_5299_620.t7 a_5299_1782.t9 VDD.t144 VDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X209 VDD.t83 VDD.t82 VDD.t83 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X210 VDD.t147 a_7196_n5728# a_8403_n6064# VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X211 a_4609_n6817# a_4184_n6773# DVSS.t66 DVSS.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X212 DVSS.t64 a_4184_n6773# a_4609_n6817# DVSS.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X213 DVSS.t126 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 DVSS.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X214 VDD.t49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X215 VDD.t1 a_2151_4783.t0 a_2151_4783.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X216 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVSS.t124 DVSS.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X217 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_8403_n6064# VDD.t22 VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X218 a_2551_620.t0 a_2151_594.t9 VSS.t5 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X219 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 comparator_top_0.VINP DVSS.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=0.5
X220 DVSS.t22 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 DVSS.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X221 VSS.t22 VSS.t21 a_2093_1782.t4 VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X222 a_3916_n5703# a_3816_n5791# DVSS.t165 DVSS.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X223 DVSS.t43 SELB.t5 a_7096_n5816# DVSS.t42 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X224 VDD.t137 a_10809_9307# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X225 VDD.t126 comparator_top_0.comparator_bias_0.VBP.t5 a_2093_3714.t6 VDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X226 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 VDD.t32 VDD.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X227 B2.t2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 comparator_top_0.VINM VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X228 VDD.t62 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X229 a_7196_n5728# a_7096_n5816# DVSS.t94 DVSS.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X230 DVSS.t2 SELA.t5 EF_AMUX21m_1.array_1ls_1tgm_0.l0 DVSS.t1 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X231 DVSS.t86 a_11031_3400# a_11271_4224# DVSS.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X232 VSS.t9 a_2151_594.t0 a_2151_594.t1 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X233 a_5299_620.t3 a_2551_620.t7 VDD.t115 VDD.t59 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X234 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 B1.t1 VDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X235 a_2093_1782.t8 comparator_top_0.VINM a_2151_4783.t4 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X236 DVSS.t29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 DVSS.t28 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X237 DVSS.t153 a_838_n6794# a_1263_n6838# DVSS.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X238 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 comparator_top_0.VINP DVSS.t82 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X239 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 A2.t0 DVSS.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X240 VDD.t158 a_3916_n5703# a_4609_n6817# VDD.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X241 DVSS.t4 a_10965_3602# a_10975_4108# DVSS.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X242 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 VDD.t118 VDD.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X243 VSS.t20 VSS.t18 VSS.t20 VSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X244 a_6351_7717# a_10811_8247# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X245 VDD.t131 a_5299_620.t9 a_8881_1782.t1 VDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=2
X246 VDD.t81 VDD.t79 VDD.t81 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X247 VDD.t153 a_4609_n6817# a_3916_n5703# VDD.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X248 VDD.t136 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 VDD.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X249 a_2221_8623.t0 a_1821_8526.t9 VDD.t38 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X250 VDD.t78 VDD.t76 VDD.t78 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X251 a_5299_1782.t0 comparator_top_0.VINP a_2093_1782.t1 VSS.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X252 A2.t3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 A2.t2 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X253 DVSS.t138 a_10442_n5795# a_10542_n5707# DVSS.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X254 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD.t134 VDD.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X255 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 VDD.t18 VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X256 DVSS.t146 EF_AMUX21m_2.array_1ls_1tgm_0.l0 a_10442_n5795# DVSS.t145 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X257 DVSS.t53 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 DVSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X258 a_4184_n6773# a_3816_n5791# DVSS.t163 DVSS.t162 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X259 a_10542_n5707# a_10442_n5795# DVSS.t136 DVSS.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X260 VSS.t54 comparator_top_0.comparator_bias_0.VBN.t12 comparator_top_0.comparator_bias_0.VBP.t1 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X261 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_1777_n6060# DVSS.t151 DVSS.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X262 VDD.t24 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 VDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X263 VDD.t146 a_7196_n5728# a_7889_n6842# VDD.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X264 B2.t6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 comparator_top_0.VINM DVSS.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X265 B2.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 B2.t0 DVSS.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X266 DVSS.t134 a_10442_n5795# a_10542_n5707# DVSS.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
R0 comparator_top_0.comparator_bias_0.VBN.n263 comparator_top_0.comparator_bias_0.VBN.t2 60.2505
R1 comparator_top_0.comparator_bias_0.VBN.n284 comparator_top_0.comparator_bias_0.VBN.t11 60.2505
R2 comparator_top_0.comparator_bias_0.VBN.n304 comparator_top_0.comparator_bias_0.VBN.t12 60.2505
R3 comparator_top_0.comparator_bias_0.VBN.n306 comparator_top_0.comparator_bias_0.VBN.t10 60.2505
R4 comparator_top_0.comparator_bias_0.VBN.n318 comparator_top_0.comparator_bias_0.VBN.t9 60.2505
R5 comparator_top_0.comparator_bias_0.VBN.n97 comparator_top_0.comparator_bias_0.VBN.n95 41.8847
R6 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.t5 35.1154
R7 comparator_top_0.comparator_bias_0.VBN.n105 comparator_top_0.comparator_bias_0.VBN.n102 26.3366
R8 comparator_top_0.comparator_bias_0.VBN.n52 comparator_top_0.comparator_bias_0.VBN.n51 26.3366
R9 comparator_top_0.comparator_bias_0.VBN.n38 comparator_top_0.comparator_bias_0.VBN.n35 26.3366
R10 comparator_top_0.comparator_bias_0.VBN.n97 comparator_top_0.comparator_bias_0.VBN.n96 15.9528
R11 comparator_top_0.comparator_bias_0.VBN.n44 comparator_top_0.comparator_bias_0.VBN.n42 12.8005
R12 comparator_top_0.comparator_bias_0.VBN.n44 comparator_top_0.comparator_bias_0.VBN.n43 12.8005
R13 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n267 9.3005
R14 comparator_top_0.comparator_bias_0.VBN.n273 comparator_top_0.comparator_bias_0.VBN.n272 9.3005
R15 comparator_top_0.comparator_bias_0.VBN.n282 comparator_top_0.comparator_bias_0.VBN.n281 9.3005
R16 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n276 9.3005
R17 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n287 9.3005
R18 comparator_top_0.comparator_bias_0.VBN.n302 comparator_top_0.comparator_bias_0.VBN.n301 9.3005
R19 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n296 9.3005
R20 comparator_top_0.comparator_bias_0.VBN.n293 comparator_top_0.comparator_bias_0.VBN.n292 9.3005
R21 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.n23 9.3005
R22 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.n31 9.3005
R23 comparator_top_0.comparator_bias_0.VBN.n11 comparator_top_0.comparator_bias_0.VBN.n40 9.3005
R24 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n46 9.3005
R25 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n55 9.3005
R26 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n63 9.3005
R27 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n71 9.3005
R28 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n79 9.3005
R29 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n87 9.3005
R30 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n86 9.3005
R31 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n85 9.3005
R32 comparator_top_0.comparator_bias_0.VBN.n85 comparator_top_0.comparator_bias_0.VBN.n84 9.3005
R33 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n78 9.3005
R34 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n77 9.3005
R35 comparator_top_0.comparator_bias_0.VBN.n77 comparator_top_0.comparator_bias_0.VBN.n76 9.3005
R36 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n70 9.3005
R37 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n69 9.3005
R38 comparator_top_0.comparator_bias_0.VBN.n69 comparator_top_0.comparator_bias_0.VBN.n68 9.3005
R39 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n62 9.3005
R40 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n61 9.3005
R41 comparator_top_0.comparator_bias_0.VBN.n61 comparator_top_0.comparator_bias_0.VBN.n60 9.3005
R42 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n54 9.3005
R43 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n53 9.3005
R44 comparator_top_0.comparator_bias_0.VBN.n53 comparator_top_0.comparator_bias_0.VBN.n52 9.3005
R45 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n45 9.3005
R46 comparator_top_0.comparator_bias_0.VBN.n11 comparator_top_0.comparator_bias_0.VBN.n41 9.3005
R47 comparator_top_0.comparator_bias_0.VBN.n11 comparator_top_0.comparator_bias_0.VBN.n39 9.3005
R48 comparator_top_0.comparator_bias_0.VBN.n39 comparator_top_0.comparator_bias_0.VBN.n38 9.3005
R49 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.n32 9.3005
R50 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.n30 9.3005
R51 comparator_top_0.comparator_bias_0.VBN.n30 comparator_top_0.comparator_bias_0.VBN.n29 9.3005
R52 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.n24 9.3005
R53 comparator_top_0.comparator_bias_0.VBN.n14 comparator_top_0.comparator_bias_0.VBN.n22 9.3005
R54 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n155 9.3005
R55 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n147 9.3005
R56 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n139 9.3005
R57 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n131 9.3005
R58 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n123 9.3005
R59 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n115 9.3005
R60 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n107 9.3005
R61 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n98 9.3005
R62 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n106 9.3005
R63 comparator_top_0.comparator_bias_0.VBN.n106 comparator_top_0.comparator_bias_0.VBN.n105 9.3005
R64 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n99 9.3005
R65 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n108 9.3005
R66 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n114 9.3005
R67 comparator_top_0.comparator_bias_0.VBN.n114 comparator_top_0.comparator_bias_0.VBN.n113 9.3005
R68 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n122 9.3005
R69 comparator_top_0.comparator_bias_0.VBN.n122 comparator_top_0.comparator_bias_0.VBN.n121 9.3005
R70 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n116 9.3005
R71 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n124 9.3005
R72 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n130 9.3005
R73 comparator_top_0.comparator_bias_0.VBN.n130 comparator_top_0.comparator_bias_0.VBN.n129 9.3005
R74 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n138 9.3005
R75 comparator_top_0.comparator_bias_0.VBN.n138 comparator_top_0.comparator_bias_0.VBN.n137 9.3005
R76 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n132 9.3005
R77 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n140 9.3005
R78 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n146 9.3005
R79 comparator_top_0.comparator_bias_0.VBN.n146 comparator_top_0.comparator_bias_0.VBN.n145 9.3005
R80 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n154 9.3005
R81 comparator_top_0.comparator_bias_0.VBN.n154 comparator_top_0.comparator_bias_0.VBN.n153 9.3005
R82 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n148 9.3005
R83 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n156 9.3005
R84 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n162 9.3005
R85 comparator_top_0.comparator_bias_0.VBN.n162 comparator_top_0.comparator_bias_0.VBN.n161 9.3005
R86 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n170 9.3005
R87 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n171 9.3005
R88 comparator_top_0.comparator_bias_0.VBN.n177 comparator_top_0.comparator_bias_0.VBN.n176 9.3005
R89 comparator_top_0.comparator_bias_0.VBN.n92 comparator_top_0.comparator_bias_0.VBN.n91 9.3005
R90 comparator_top_0.comparator_bias_0.VBN.n167 comparator_top_0.comparator_bias_0.VBN.n166 9.3005
R91 comparator_top_0.comparator_bias_0.VBN.n20 comparator_top_0.comparator_bias_0.VBN.n315 9.3005
R92 comparator_top_0.comparator_bias_0.VBN.n20 comparator_top_0.comparator_bias_0.VBN.n313 9.3005
R93 comparator_top_0.comparator_bias_0.VBN.n313 comparator_top_0.comparator_bias_0.VBN.n312 9.3005
R94 comparator_top_0.comparator_bias_0.VBN.n20 comparator_top_0.comparator_bias_0.VBN.n314 9.3005
R95 comparator_top_0.comparator_bias_0.VBN.n17 comparator_top_0.comparator_bias_0.VBN.n327 9.3005
R96 comparator_top_0.comparator_bias_0.VBN.n17 comparator_top_0.comparator_bias_0.VBN.n326 9.3005
R97 comparator_top_0.comparator_bias_0.VBN.n17 comparator_top_0.comparator_bias_0.VBN.n325 9.3005
R98 comparator_top_0.comparator_bias_0.VBN.n325 comparator_top_0.comparator_bias_0.VBN.n324 9.3005
R99 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n246 9.3005
R100 comparator_top_0.comparator_bias_0.VBN.n252 comparator_top_0.comparator_bias_0.VBN.n251 9.3005
R101 comparator_top_0.comparator_bias_0.VBN.n261 comparator_top_0.comparator_bias_0.VBN.n260 9.3005
R102 comparator_top_0.comparator_bias_0.VBN.n18 comparator_top_0.comparator_bias_0.VBN.n255 9.3005
R103 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n242 9.3005
R104 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n241 9.3005
R105 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n243 9.3005
R106 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n197 9.3005
R107 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n192 9.3005
R108 comparator_top_0.comparator_bias_0.VBN.n285 comparator_top_0.comparator_bias_0.VBN.n284 8.76429
R109 comparator_top_0.comparator_bias_0.VBN.n305 comparator_top_0.comparator_bias_0.VBN.n304 8.76429
R110 comparator_top_0.comparator_bias_0.VBN.n264 comparator_top_0.comparator_bias_0.VBN.n263 8.76429
R111 comparator_top_0.comparator_bias_0.VBN.n271 comparator_top_0.comparator_bias_0.VBN.n270 8.21641
R112 comparator_top_0.comparator_bias_0.VBN.n280 comparator_top_0.comparator_bias_0.VBN.n279 8.21641
R113 comparator_top_0.comparator_bias_0.VBN.n291 comparator_top_0.comparator_bias_0.VBN.n290 8.21641
R114 comparator_top_0.comparator_bias_0.VBN.n300 comparator_top_0.comparator_bias_0.VBN.n299 8.21641
R115 comparator_top_0.comparator_bias_0.VBN.n311 comparator_top_0.comparator_bias_0.VBN.n310 8.21641
R116 comparator_top_0.comparator_bias_0.VBN.n323 comparator_top_0.comparator_bias_0.VBN.n322 8.21641
R117 comparator_top_0.comparator_bias_0.VBN.n250 comparator_top_0.comparator_bias_0.VBN.n249 8.21641
R118 comparator_top_0.comparator_bias_0.VBN.n259 comparator_top_0.comparator_bias_0.VBN.n258 8.21641
R119 comparator_top_0.comparator_bias_0.VBN.n160 comparator_top_0.comparator_bias_0.VBN.n159 7.95102
R120 comparator_top_0.comparator_bias_0.VBN.n165 comparator_top_0.comparator_bias_0.VBN.n164 7.95102
R121 comparator_top_0.comparator_bias_0.VBN.n105 comparator_top_0.comparator_bias_0.VBN.n104 7.45411
R122 comparator_top_0.comparator_bias_0.VBN.n52 comparator_top_0.comparator_bias_0.VBN.n50 7.45411
R123 comparator_top_0.comparator_bias_0.VBN.n38 comparator_top_0.comparator_bias_0.VBN.n37 7.45411
R124 comparator_top_0.comparator_bias_0.VBN.n152 comparator_top_0.comparator_bias_0.VBN.n151 6.9572
R125 comparator_top_0.comparator_bias_0.VBN.n175 comparator_top_0.comparator_bias_0.VBN.n174 6.9572
R126 comparator_top_0.comparator_bias_0.VBN.n319 comparator_top_0.comparator_bias_0.VBN.n318 6.92242
R127 comparator_top_0.comparator_bias_0.VBN.n307 comparator_top_0.comparator_bias_0.VBN.n306 6.92012
R128 comparator_top_0.comparator_bias_0.VBN.n113 comparator_top_0.comparator_bias_0.VBN.n112 6.46029
R129 comparator_top_0.comparator_bias_0.VBN.n60 comparator_top_0.comparator_bias_0.VBN.n59 6.46029
R130 comparator_top_0.comparator_bias_0.VBN.n29 comparator_top_0.comparator_bias_0.VBN.n28 6.46029
R131 comparator_top_0.comparator_bias_0.VBN.n158 comparator_top_0.comparator_bias_0.VBN.n157 6.02403
R132 comparator_top_0.comparator_bias_0.VBN.n144 comparator_top_0.comparator_bias_0.VBN.n143 5.96339
R133 comparator_top_0.comparator_bias_0.VBN.n90 comparator_top_0.comparator_bias_0.VBN.n89 5.96339
R134 comparator_top_0.comparator_bias_0.VBN.n269 comparator_top_0.comparator_bias_0.VBN.n268 5.64756
R135 comparator_top_0.comparator_bias_0.VBN.n278 comparator_top_0.comparator_bias_0.VBN.n277 5.64756
R136 comparator_top_0.comparator_bias_0.VBN.n289 comparator_top_0.comparator_bias_0.VBN.n288 5.64756
R137 comparator_top_0.comparator_bias_0.VBN.n298 comparator_top_0.comparator_bias_0.VBN.n297 5.64756
R138 comparator_top_0.comparator_bias_0.VBN.n106 comparator_top_0.comparator_bias_0.VBN.n101 5.64756
R139 comparator_top_0.comparator_bias_0.VBN.n53 comparator_top_0.comparator_bias_0.VBN.n48 5.64756
R140 comparator_top_0.comparator_bias_0.VBN.n39 comparator_top_0.comparator_bias_0.VBN.n34 5.64756
R141 comparator_top_0.comparator_bias_0.VBN.n309 comparator_top_0.comparator_bias_0.VBN.n308 5.64756
R142 comparator_top_0.comparator_bias_0.VBN.n321 comparator_top_0.comparator_bias_0.VBN.n320 5.64756
R143 comparator_top_0.comparator_bias_0.VBN.n248 comparator_top_0.comparator_bias_0.VBN.n247 5.64756
R144 comparator_top_0.comparator_bias_0.VBN.n257 comparator_top_0.comparator_bias_0.VBN.n256 5.64756
R145 comparator_top_0.comparator_bias_0.VBN.n210 comparator_top_0.comparator_bias_0.VBN.t1 5.5395
R146 comparator_top_0.comparator_bias_0.VBN.n210 comparator_top_0.comparator_bias_0.VBN.t7 5.5395
R147 comparator_top_0.comparator_bias_0.VBN.n227 comparator_top_0.comparator_bias_0.VBN.t8 5.5395
R148 comparator_top_0.comparator_bias_0.VBN.n227 comparator_top_0.comparator_bias_0.VBN.t0 5.5395
R149 comparator_top_0.comparator_bias_0.VBN.n121 comparator_top_0.comparator_bias_0.VBN.n120 5.46648
R150 comparator_top_0.comparator_bias_0.VBN.n68 comparator_top_0.comparator_bias_0.VBN.n67 5.46648
R151 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n244 5.28563
R152 comparator_top_0.comparator_bias_0.VBN.n150 comparator_top_0.comparator_bias_0.VBN.n149 5.27109
R153 comparator_top_0.comparator_bias_0.VBN.n136 comparator_top_0.comparator_bias_0.VBN.n135 4.96957
R154 comparator_top_0.comparator_bias_0.VBN.n83 comparator_top_0.comparator_bias_0.VBN.n82 4.96957
R155 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n266 4.911
R156 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n286 4.911
R157 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n275 4.91005
R158 comparator_top_0.comparator_bias_0.VBN.n18 comparator_top_0.comparator_bias_0.VBN.n254 4.91005
R159 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n295 4.90905
R160 comparator_top_0.comparator_bias_0.VBN.n114 comparator_top_0.comparator_bias_0.VBN.n110 4.89462
R161 comparator_top_0.comparator_bias_0.VBN.n61 comparator_top_0.comparator_bias_0.VBN.n57 4.89462
R162 comparator_top_0.comparator_bias_0.VBN.n30 comparator_top_0.comparator_bias_0.VBN.n26 4.89462
R163 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n245 4.76425
R164 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n44 4.6505
R165 comparator_top_0.comparator_bias_0.VBN.n142 comparator_top_0.comparator_bias_0.VBN.n141 4.51815
R166 comparator_top_0.comparator_bias_0.VBN.n169 comparator_top_0.comparator_bias_0.VBN.n163 4.51815
R167 comparator_top_0.comparator_bias_0.VBN.n195 comparator_top_0.comparator_bias_0.VBN.n194 4.51815
R168 comparator_top_0.comparator_bias_0.VBN.n206 comparator_top_0.comparator_bias_0.VBN.n205 4.51815
R169 comparator_top_0.comparator_bias_0.VBN.n236 comparator_top_0.comparator_bias_0.VBN.n235 4.51815
R170 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n94 4.5005
R171 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n182 4.5005
R172 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n179 4.5005
R173 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n169 4.5005
R174 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n274 4.5005
R175 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n283 4.5005
R176 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n303 4.5005
R177 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n294 4.5005
R178 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n253 4.5005
R179 comparator_top_0.comparator_bias_0.VBN.n18 comparator_top_0.comparator_bias_0.VBN.n262 4.5005
R180 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n195 4.5005
R181 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n190 4.5005
R182 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n185 4.5005
R183 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n239 4.5005
R184 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n200 4.5005
R185 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n216 4.5005
R186 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n204 4.5005
R187 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n213 4.5005
R188 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n209 4.5005
R189 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n226 4.5005
R190 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n231 4.5005
R191 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n234 4.5005
R192 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n220 4.5005
R193 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n224 4.5005
R194 comparator_top_0.comparator_bias_0.VBN.n129 comparator_top_0.comparator_bias_0.VBN.n128 4.47267
R195 comparator_top_0.comparator_bias_0.VBN.n76 comparator_top_0.comparator_bias_0.VBN.n75 4.47267
R196 comparator_top_0.comparator_bias_0.VBN.n21 comparator_top_0.comparator_bias_0.VBN.n7 4.44875
R197 comparator_top_0.comparator_bias_0.VBN.n7 comparator_top_0.comparator_bias_0.VBN.n316 7.3305
R198 comparator_top_0.comparator_bias_0.VBN.n17 comparator_top_0.comparator_bias_0.VBN.n329 4.24504
R199 comparator_top_0.comparator_bias_0.VBN.n122 comparator_top_0.comparator_bias_0.VBN.n118 4.14168
R200 comparator_top_0.comparator_bias_0.VBN.n69 comparator_top_0.comparator_bias_0.VBN.n65 4.14168
R201 comparator_top_0.comparator_bias_0.VBN.n128 comparator_top_0.comparator_bias_0.VBN.n127 3.97576
R202 comparator_top_0.comparator_bias_0.VBN.n75 comparator_top_0.comparator_bias_0.VBN.n74 3.97576
R203 comparator_top_0.comparator_bias_0.VBN.n134 comparator_top_0.comparator_bias_0.VBN.n133 3.76521
R204 comparator_top_0.comparator_bias_0.VBN.n179 comparator_top_0.comparator_bias_0.VBN.n173 3.76521
R205 comparator_top_0.comparator_bias_0.VBN.n182 comparator_top_0.comparator_bias_0.VBN.n180 3.76521
R206 comparator_top_0.comparator_bias_0.VBN.n81 comparator_top_0.comparator_bias_0.VBN.n80 3.76521
R207 comparator_top_0.comparator_bias_0.VBN.n239 comparator_top_0.comparator_bias_0.VBN.n238 3.76521
R208 comparator_top_0.comparator_bias_0.VBN.n137 comparator_top_0.comparator_bias_0.VBN.n136 3.47885
R209 comparator_top_0.comparator_bias_0.VBN.n84 comparator_top_0.comparator_bias_0.VBN.n83 3.47885
R210 comparator_top_0.comparator_bias_0.VBN.n20 comparator_top_0.comparator_bias_0.VBN.n307 3.47756
R211 comparator_top_0.comparator_bias_0.VBN.n17 comparator_top_0.comparator_bias_0.VBN.n319 3.4767
R212 comparator_top_0.comparator_bias_0.VBN.n130 comparator_top_0.comparator_bias_0.VBN.n126 3.38874
R213 comparator_top_0.comparator_bias_0.VBN.n77 comparator_top_0.comparator_bias_0.VBN.n73 3.38874
R214 comparator_top_0.comparator_bias_0.VBN.n186 comparator_top_0.comparator_bias_0.VBN.t6 3.3065
R215 comparator_top_0.comparator_bias_0.VBN.n186 comparator_top_0.comparator_bias_0.VBN.t3 3.3065
R216 comparator_top_0.comparator_bias_0.VBN.n190 comparator_top_0.comparator_bias_0.VBN.n188 3.74814
R217 comparator_top_0.comparator_bias_0.VBN.n15 comparator_top_0.comparator_bias_0.VBN.n187 3.15814
R218 comparator_top_0.comparator_bias_0.VBN.n3 comparator_top_0.comparator_bias_0.VBN.n285 3.03311
R219 comparator_top_0.comparator_bias_0.VBN.n2 comparator_top_0.comparator_bias_0.VBN.n305 3.03311
R220 comparator_top_0.comparator_bias_0.VBN.n18 comparator_top_0.comparator_bias_0.VBN.n264 3.03311
R221 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n206 3.03311
R222 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n236 3.03311
R223 comparator_top_0.comparator_bias_0.VBN.n126 comparator_top_0.comparator_bias_0.VBN.n125 3.01226
R224 comparator_top_0.comparator_bias_0.VBN.n94 comparator_top_0.comparator_bias_0.VBN.n88 3.01226
R225 comparator_top_0.comparator_bias_0.VBN.n73 comparator_top_0.comparator_bias_0.VBN.n72 3.01226
R226 comparator_top_0.comparator_bias_0.VBN.n190 comparator_top_0.comparator_bias_0.VBN.n189 3.01226
R227 comparator_top_0.comparator_bias_0.VBN.n120 comparator_top_0.comparator_bias_0.VBN.n119 2.98194
R228 comparator_top_0.comparator_bias_0.VBN.n67 comparator_top_0.comparator_bias_0.VBN.n66 2.98194
R229 comparator_top_0.comparator_bias_0.VBN.n138 comparator_top_0.comparator_bias_0.VBN.n134 2.63579
R230 comparator_top_0.comparator_bias_0.VBN.n85 comparator_top_0.comparator_bias_0.VBN.n81 2.63579
R231 comparator_top_0.comparator_bias_0.VBN.n239 comparator_top_0.comparator_bias_0.VBN.n237 2.63579
R232 comparator_top_0.comparator_bias_0.VBN.n204 comparator_top_0.comparator_bias_0.VBN.n202 2.63579
R233 comparator_top_0.comparator_bias_0.VBN.n224 comparator_top_0.comparator_bias_0.VBN.n222 2.63579
R234 comparator_top_0.comparator_bias_0.VBN.n192 comparator_top_0.comparator_bias_0.VBN.n191 2.61733
R235 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n198 2.60826
R236 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n218 2.60817
R237 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n183 2.53421
R238 comparator_top_0.comparator_bias_0.VBN.n145 comparator_top_0.comparator_bias_0.VBN.n144 2.48504
R239 comparator_top_0.comparator_bias_0.VBN.n91 comparator_top_0.comparator_bias_0.VBN.n90 2.48504
R240 comparator_top_0.comparator_bias_0.VBN.n7 comparator_top_0.comparator_bias_0.VBN.n17 2.42663
R241 comparator_top_0.comparator_bias_0.VBN.n7 comparator_top_0.comparator_bias_0.VBN.n20 2.39724
R242 comparator_top_0.comparator_bias_0.VBN.n118 comparator_top_0.comparator_bias_0.VBN.n117 2.25932
R243 comparator_top_0.comparator_bias_0.VBN.n65 comparator_top_0.comparator_bias_0.VBN.n64 2.25932
R244 comparator_top_0.comparator_bias_0.VBN.n216 comparator_top_0.comparator_bias_0.VBN.n214 2.25932
R245 comparator_top_0.comparator_bias_0.VBN.n208 comparator_top_0.comparator_bias_0.VBN.n207 2.25932
R246 comparator_top_0.comparator_bias_0.VBN.n234 comparator_top_0.comparator_bias_0.VBN.n232 2.25932
R247 comparator_top_0.comparator_bias_0.VBN.n230 comparator_top_0.comparator_bias_0.VBN.n229 2.25932
R248 comparator_top_0.comparator_bias_0.VBN.n216 comparator_top_0.comparator_bias_0.VBN.n215 2.25379
R249 comparator_top_0.comparator_bias_0.VBN.n234 comparator_top_0.comparator_bias_0.VBN.n233 2.25379
R250 comparator_top_0.comparator_bias_0.VBN.n7 comparator_top_0.comparator_bias_0.VBN.n317 2.2505
R251 comparator_top_0.comparator_bias_0.VBN.n197 comparator_top_0.comparator_bias_0.VBN.n196 2.24766
R252 comparator_top_0.comparator_bias_0.VBN.n265 comparator_top_0.comparator_bias_0.VBN.n18 2.073
R253 comparator_top_0.comparator_bias_0.VBN comparator_top_0.comparator_bias_0.VBN.n19 2.06925
R254 comparator_top_0.comparator_bias_0.VBN.n112 comparator_top_0.comparator_bias_0.VBN.n111 1.98813
R255 comparator_top_0.comparator_bias_0.VBN.n59 comparator_top_0.comparator_bias_0.VBN.n58 1.98813
R256 comparator_top_0.comparator_bias_0.VBN.n28 comparator_top_0.comparator_bias_0.VBN.n27 1.98813
R257 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n172 1.94045
R258 comparator_top_0.comparator_bias_0.VBN.n146 comparator_top_0.comparator_bias_0.VBN.n142 1.88285
R259 comparator_top_0.comparator_bias_0.VBN.n93 comparator_top_0.comparator_bias_0.VBN.n92 1.88285
R260 comparator_top_0.comparator_bias_0.VBN.n195 comparator_top_0.comparator_bias_0.VBN.n193 1.88285
R261 comparator_top_0.comparator_bias_0.VBN.n204 comparator_top_0.comparator_bias_0.VBN.n203 1.87949
R262 comparator_top_0.comparator_bias_0.VBN.n224 comparator_top_0.comparator_bias_0.VBN.n223 1.87949
R263 comparator_top_0.comparator_bias_0.VBN.n265 comparator_top_0.comparator_bias_0.VBN.n3 1.85011
R264 comparator_top_0.comparator_bias_0.VBN.n217 comparator_top_0.comparator_bias_0.VBN.n1 1.73899
R265 comparator_top_0.comparator_bias_0.VBN.n21 comparator_top_0.comparator_bias_0.VBN.n172 1.70776
R266 comparator_top_0.comparator_bias_0.VBN.n19 comparator_top_0.comparator_bias_0.VBN.n2 1.70567
R267 comparator_top_0.comparator_bias_0.VBN.n15 comparator_top_0.comparator_bias_0.VBN.n186 1.61779
R268 comparator_top_0.comparator_bias_0.VBN.n95 comparator_top_0.comparator_bias_0.VBN.t4 1.60717
R269 comparator_top_0.comparator_bias_0.VBN.n7 comparator_top_0.comparator_bias_0.VBN 1.60425
R270 comparator_top_0.comparator_bias_0.VBN.n110 comparator_top_0.comparator_bias_0.VBN.n109 1.50638
R271 comparator_top_0.comparator_bias_0.VBN.n169 comparator_top_0.comparator_bias_0.VBN.n168 1.50638
R272 comparator_top_0.comparator_bias_0.VBN.n179 comparator_top_0.comparator_bias_0.VBN.n178 1.50638
R273 comparator_top_0.comparator_bias_0.VBN.n94 comparator_top_0.comparator_bias_0.VBN.n93 1.50638
R274 comparator_top_0.comparator_bias_0.VBN.n57 comparator_top_0.comparator_bias_0.VBN.n56 1.50638
R275 comparator_top_0.comparator_bias_0.VBN.n26 comparator_top_0.comparator_bias_0.VBN.n25 1.50638
R276 comparator_top_0.comparator_bias_0.VBN.n213 comparator_top_0.comparator_bias_0.VBN.n212 1.50638
R277 comparator_top_0.comparator_bias_0.VBN.n226 comparator_top_0.comparator_bias_0.VBN.n225 1.50638
R278 comparator_top_0.comparator_bias_0.VBN.n228 comparator_top_0.comparator_bias_0.VBN.n227 1.50151
R279 comparator_top_0.comparator_bias_0.VBN.n211 comparator_top_0.comparator_bias_0.VBN.n210 1.50148
R280 comparator_top_0.comparator_bias_0.VBN.n153 comparator_top_0.comparator_bias_0.VBN.n152 1.49122
R281 comparator_top_0.comparator_bias_0.VBN.n176 comparator_top_0.comparator_bias_0.VBN.n175 1.49122
R282 comparator_top_0.comparator_bias_0.VBN.n19 comparator_top_0.comparator_bias_0.VBN.n265 1.26925
R283 comparator_top_0.comparator_bias_0.VBN.n217 comparator_top_0.comparator_bias_0.VBN.n0 1.1968
R284 comparator_top_0.comparator_bias_0.VBN.n19 comparator_top_0.comparator_bias_0.VBN.n21 1.1545
R285 comparator_top_0.comparator_bias_0.VBN.n154 comparator_top_0.comparator_bias_0.VBN.n150 1.12991
R286 comparator_top_0.comparator_bias_0.VBN.n178 comparator_top_0.comparator_bias_0.VBN.n177 1.12991
R287 comparator_top_0.comparator_bias_0.VBN.n185 comparator_top_0.comparator_bias_0.VBN.n184 1.12991
R288 comparator_top_0.comparator_bias_0.VBN.n272 comparator_top_0.comparator_bias_0.VBN.n271 1.09595
R289 comparator_top_0.comparator_bias_0.VBN.n281 comparator_top_0.comparator_bias_0.VBN.n280 1.09595
R290 comparator_top_0.comparator_bias_0.VBN.n292 comparator_top_0.comparator_bias_0.VBN.n291 1.09595
R291 comparator_top_0.comparator_bias_0.VBN.n301 comparator_top_0.comparator_bias_0.VBN.n300 1.09595
R292 comparator_top_0.comparator_bias_0.VBN.n312 comparator_top_0.comparator_bias_0.VBN.n311 1.09595
R293 comparator_top_0.comparator_bias_0.VBN.n324 comparator_top_0.comparator_bias_0.VBN.n323 1.09595
R294 comparator_top_0.comparator_bias_0.VBN.n251 comparator_top_0.comparator_bias_0.VBN.n250 1.09595
R295 comparator_top_0.comparator_bias_0.VBN.n260 comparator_top_0.comparator_bias_0.VBN.n259 1.09595
R296 comparator_top_0.comparator_bias_0.VBN.n13 comparator_top_0.comparator_bias_0.VBN.n97 1.03132
R297 comparator_top_0.comparator_bias_0.VBN.n104 comparator_top_0.comparator_bias_0.VBN.n103 0.994314
R298 comparator_top_0.comparator_bias_0.VBN.n50 comparator_top_0.comparator_bias_0.VBN.n49 0.994314
R299 comparator_top_0.comparator_bias_0.VBN.n37 comparator_top_0.comparator_bias_0.VBN.n36 0.994314
R300 comparator_top_0.comparator_bias_0.VBN.n183 comparator_top_0.comparator_bias_0.VBN.n217 0.890264
R301 comparator_top_0.comparator_bias_0.VBN.n0 comparator_top_0.comparator_bias_0.VBN.n228 0.833627
R302 comparator_top_0.comparator_bias_0.VBN.n1 comparator_top_0.comparator_bias_0.VBN.n211 0.833623
R303 comparator_top_0.comparator_bias_0.VBN.n6 comparator_top_0.comparator_bias_0.VBN.n16 0.766876
R304 comparator_top_0.comparator_bias_0.VBN.n274 comparator_top_0.comparator_bias_0.VBN.n273 0.753441
R305 comparator_top_0.comparator_bias_0.VBN.n273 comparator_top_0.comparator_bias_0.VBN.n269 0.753441
R306 comparator_top_0.comparator_bias_0.VBN.n282 comparator_top_0.comparator_bias_0.VBN.n278 0.753441
R307 comparator_top_0.comparator_bias_0.VBN.n283 comparator_top_0.comparator_bias_0.VBN.n282 0.753441
R308 comparator_top_0.comparator_bias_0.VBN.n294 comparator_top_0.comparator_bias_0.VBN.n293 0.753441
R309 comparator_top_0.comparator_bias_0.VBN.n293 comparator_top_0.comparator_bias_0.VBN.n289 0.753441
R310 comparator_top_0.comparator_bias_0.VBN.n302 comparator_top_0.comparator_bias_0.VBN.n298 0.753441
R311 comparator_top_0.comparator_bias_0.VBN.n303 comparator_top_0.comparator_bias_0.VBN.n302 0.753441
R312 comparator_top_0.comparator_bias_0.VBN.n101 comparator_top_0.comparator_bias_0.VBN.n100 0.753441
R313 comparator_top_0.comparator_bias_0.VBN.n48 comparator_top_0.comparator_bias_0.VBN.n47 0.753441
R314 comparator_top_0.comparator_bias_0.VBN.n34 comparator_top_0.comparator_bias_0.VBN.n33 0.753441
R315 comparator_top_0.comparator_bias_0.VBN.n313 comparator_top_0.comparator_bias_0.VBN.n309 0.753441
R316 comparator_top_0.comparator_bias_0.VBN.n325 comparator_top_0.comparator_bias_0.VBN.n321 0.753441
R317 comparator_top_0.comparator_bias_0.VBN.n253 comparator_top_0.comparator_bias_0.VBN.n252 0.753441
R318 comparator_top_0.comparator_bias_0.VBN.n252 comparator_top_0.comparator_bias_0.VBN.n248 0.753441
R319 comparator_top_0.comparator_bias_0.VBN.n261 comparator_top_0.comparator_bias_0.VBN.n257 0.753441
R320 comparator_top_0.comparator_bias_0.VBN.n262 comparator_top_0.comparator_bias_0.VBN.n261 0.753441
R321 comparator_top_0.comparator_bias_0.VBN.n200 comparator_top_0.comparator_bias_0.VBN.n199 0.753441
R322 comparator_top_0.comparator_bias_0.VBN.n209 comparator_top_0.comparator_bias_0.VBN.n208 0.753441
R323 comparator_top_0.comparator_bias_0.VBN.n220 comparator_top_0.comparator_bias_0.VBN.n219 0.753441
R324 comparator_top_0.comparator_bias_0.VBN.n231 comparator_top_0.comparator_bias_0.VBN.n230 0.753441
R325 comparator_top_0.comparator_bias_0.VBN.n329 comparator_top_0.comparator_bias_0.VBN.n328 0.738413
R326 comparator_top_0.comparator_bias_0.VBN.n5 comparator_top_0.comparator_bias_0.VBN.n4 0.700653
R327 comparator_top_0.comparator_bias_0.VBN.n4 comparator_top_0.comparator_bias_0.VBN.n10 0.571152
R328 comparator_top_0.comparator_bias_0.VBN.n18 comparator_top_0.comparator_bias_0.VBN.n6 0.498175
R329 comparator_top_0.comparator_bias_0.VBN.n161 comparator_top_0.comparator_bias_0.VBN.n160 0.497407
R330 comparator_top_0.comparator_bias_0.VBN.n166 comparator_top_0.comparator_bias_0.VBN.n165 0.497407
R331 comparator_top_0.comparator_bias_0.VBN.n16 comparator_top_0.comparator_bias_0.VBN.n15 0.48986
R332 comparator_top_0.comparator_bias_0.VBN.n241 comparator_top_0.comparator_bias_0.VBN.n240 0.461175
R333 comparator_top_0.comparator_bias_0.VBN.n12 comparator_top_0.comparator_bias_0.VBN.n11 0.42713
R334 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n5 0.387304
R335 comparator_top_0.comparator_bias_0.VBN.n11 comparator_top_0.comparator_bias_0.VBN.n14 0.380935
R336 comparator_top_0.comparator_bias_0.VBN.n9 comparator_top_0.comparator_bias_0.VBN.n8 0.380935
R337 comparator_top_0.comparator_bias_0.VBN.n10 comparator_top_0.comparator_bias_0.VBN.n13 0.380935
R338 comparator_top_0.comparator_bias_0.VBN.n8 comparator_top_0.comparator_bias_0.VBN.n12 0.380935
R339 comparator_top_0.comparator_bias_0.VBN.n162 comparator_top_0.comparator_bias_0.VBN.n158 0.376971
R340 comparator_top_0.comparator_bias_0.VBN.n168 comparator_top_0.comparator_bias_0.VBN.n167 0.376971
R341 comparator_top_0.comparator_bias_0.VBN.n182 comparator_top_0.comparator_bias_0.VBN.n181 0.376971
R342 comparator_top_0.comparator_bias_0.VBN.n202 comparator_top_0.comparator_bias_0.VBN.n201 0.376971
R343 comparator_top_0.comparator_bias_0.VBN.n222 comparator_top_0.comparator_bias_0.VBN.n221 0.376971
R344 a_1821_8526.t0 a_1821_8526.n12 121.124
R345 a_1821_8526.n171 a_1821_8526.t1 116.841
R346 a_1821_8526.n109 a_1821_8526.t6 60.2505
R347 a_1821_8526.n88 a_1821_8526.t9 60.2505
R348 a_1821_8526.n68 a_1821_8526.t7 60.2505
R349 a_1821_8526.n48 a_1821_8526.t8 60.2505
R350 a_1821_8526.n175 a_1821_8526.n174 52.6902
R351 a_1821_8526.n183 a_1821_8526.n182 46.104
R352 a_1821_8526.n199 a_1821_8526.n198 46.104
R353 a_1821_8526.n144 a_1821_8526.n143 39.5177
R354 a_1821_8526.n40 a_1821_8526.n39 39.5177
R355 a_1821_8526.n151 a_1821_8526.n150 32.9315
R356 a_1821_8526.n30 a_1821_8526.n29 32.9315
R357 a_1821_8526.n162 a_1821_8526.n161 29.6384
R358 a_1821_8526.n23 a_1821_8526.n22 29.6384
R359 a_1821_8526.n140 a_1821_8526.t3 27.6955
R360 a_1821_8526.n161 a_1821_8526.n160 26.3453
R361 a_1821_8526.n22 a_1821_8526.n21 26.3453
R362 a_1821_8526.n152 a_1821_8526.n151 23.0522
R363 a_1821_8526.n31 a_1821_8526.n30 23.0522
R364 a_1821_8526.n145 a_1821_8526.n144 16.466
R365 a_1821_8526.n41 a_1821_8526.n40 16.466
R366 a_1821_8526.n138 a_1821_8526.n137 13.177
R367 a_1821_8526.n184 a_1821_8526.n183 9.87981
R368 a_1821_8526.n200 a_1821_8526.n199 9.87981
R369 a_1821_8526.n10 a_1821_8526.n134 9.31646
R370 a_1821_8526.n3 a_1821_8526.n130 9.3005
R371 a_1821_8526.n3 a_1821_8526.n132 9.3005
R372 a_1821_8526.n11 a_1821_8526.n178 9.3005
R373 a_1821_8526.n1 a_1821_8526.n186 9.3005
R374 a_1821_8526.n11 a_1821_8526.n177 9.3005
R375 a_1821_8526.n177 a_1821_8526.n176 9.3005
R376 a_1821_8526.n11 a_1821_8526.n179 9.3005
R377 a_1821_8526.n1 a_1821_8526.n185 9.3005
R378 a_1821_8526.n185 a_1821_8526.n184 9.3005
R379 a_1821_8526.n1 a_1821_8526.n163 9.3005
R380 a_1821_8526.n163 a_1821_8526.n162 9.3005
R381 a_1821_8526.n1 a_1821_8526.n166 9.3005
R382 a_1821_8526.n153 a_1821_8526.n152 9.3005
R383 a_1821_8526.n146 a_1821_8526.n145 9.3005
R384 a_1821_8526.n10 a_1821_8526.n141 9.3005
R385 a_1821_8526.n9 a_1821_8526.n56 9.3005
R386 a_1821_8526.n9 a_1821_8526.n57 9.3005
R387 a_1821_8526.n9 a_1821_8526.n55 9.3005
R388 a_1821_8526.n55 a_1821_8526.n54 9.3005
R389 a_1821_8526.n7 a_1821_8526.n61 9.3005
R390 a_1821_8526.n8 a_1821_8526.n76 9.3005
R391 a_1821_8526.n8 a_1821_8526.n77 9.3005
R392 a_1821_8526.n8 a_1821_8526.n75 9.3005
R393 a_1821_8526.n75 a_1821_8526.n74 9.3005
R394 a_1821_8526.n7 a_1821_8526.n67 9.3005
R395 a_1821_8526.n67 a_1821_8526.n66 9.3005
R396 a_1821_8526.n7 a_1821_8526.n60 9.3005
R397 a_1821_8526.n5 a_1821_8526.n81 9.3005
R398 a_1821_8526.n6 a_1821_8526.n96 9.3005
R399 a_1821_8526.n6 a_1821_8526.n97 9.3005
R400 a_1821_8526.n6 a_1821_8526.n95 9.3005
R401 a_1821_8526.n95 a_1821_8526.n94 9.3005
R402 a_1821_8526.n5 a_1821_8526.n87 9.3005
R403 a_1821_8526.n87 a_1821_8526.n86 9.3005
R404 a_1821_8526.n5 a_1821_8526.n80 9.3005
R405 a_1821_8526.n4 a_1821_8526.n101 9.3005
R406 a_1821_8526.n13 a_1821_8526.n108 9.3005
R407 a_1821_8526.n13 a_1821_8526.n110 9.3005
R408 a_1821_8526.n4 a_1821_8526.n107 9.3005
R409 a_1821_8526.n107 a_1821_8526.n106 9.3005
R410 a_1821_8526.n4 a_1821_8526.n100 9.3005
R411 a_1821_8526.n117 a_1821_8526.n116 9.3005
R412 a_1821_8526.n12 a_1821_8526.n195 9.3005
R413 a_1821_8526.n12 a_1821_8526.n202 9.3005
R414 a_1821_8526.n2 a_1821_8526.n27 9.3005
R415 a_1821_8526.n12 a_1821_8526.n201 9.3005
R416 a_1821_8526.n201 a_1821_8526.n200 9.3005
R417 a_1821_8526.n42 a_1821_8526.n41 9.3005
R418 a_1821_8526.n2 a_1821_8526.n24 9.3005
R419 a_1821_8526.n24 a_1821_8526.n23 9.3005
R420 a_1821_8526.n32 a_1821_8526.n31 9.3005
R421 a_1821_8526.n141 a_1821_8526.n140 9.0206
R422 a_1821_8526.n69 a_1821_8526.n68 8.76429
R423 a_1821_8526.n89 a_1821_8526.n88 8.76429
R424 a_1821_8526.n110 a_1821_8526.n109 8.76429
R425 a_1821_8526.n14 a_1821_8526.t2 7.50197
R426 a_1821_8526.n115 a_1821_8526.n114 7.45411
R427 a_1821_8526.n105 a_1821_8526.n104 7.45411
R428 a_1821_8526.n93 a_1821_8526.n92 7.45411
R429 a_1821_8526.n85 a_1821_8526.n84 7.45411
R430 a_1821_8526.n73 a_1821_8526.n72 7.45411
R431 a_1821_8526.n65 a_1821_8526.n64 7.45411
R432 a_1821_8526.n53 a_1821_8526.n52 7.45411
R433 a_1821_8526.n49 a_1821_8526.n48 6.80105
R434 a_1821_8526.n173 a_1821_8526.n172 6.02403
R435 a_1821_8526.n103 a_1821_8526.n102 5.64756
R436 a_1821_8526.n91 a_1821_8526.n90 5.64756
R437 a_1821_8526.n83 a_1821_8526.n82 5.64756
R438 a_1821_8526.n71 a_1821_8526.n70 5.64756
R439 a_1821_8526.n63 a_1821_8526.n62 5.64756
R440 a_1821_8526.n51 a_1821_8526.n50 5.64756
R441 a_1821_8526.n192 a_1821_8526.t4 5.5395
R442 a_1821_8526.n192 a_1821_8526.t5 5.5395
R443 a_1821_8526.n181 a_1821_8526.n180 5.27109
R444 a_1821_8526.n197 a_1821_8526.n196 5.27109
R445 a_1821_8526.n2 a_1821_8526.n18 5.266
R446 a_1821_8526.n1 a_1821_8526.n159 5.266
R447 a_1821_8526.n4 a_1821_8526.n99 4.73575
R448 a_1821_8526.n6 a_1821_8526.n98 4.73575
R449 a_1821_8526.n5 a_1821_8526.n79 4.73575
R450 a_1821_8526.n8 a_1821_8526.n78 4.73575
R451 a_1821_8526.n7 a_1821_8526.n59 4.73575
R452 a_1821_8526.n9 a_1821_8526.n58 4.73575
R453 a_1821_8526.n7 a_1821_8526.n69 4.6505
R454 a_1821_8526.n5 a_1821_8526.n89 4.6505
R455 a_1821_8526.n15 a_1821_8526.n47 6.76219
R456 a_1821_8526.n191 a_1821_8526.n190 4.51815
R457 a_1821_8526.n170 a_1821_8526.n169 4.51815
R458 a_1821_8526.n37 a_1821_8526.n36 4.51815
R459 a_1821_8526.n3 a_1821_8526.n128 4.5005
R460 a_1821_8526.n1 a_1821_8526.n158 4.5005
R461 a_1821_8526.n1 a_1821_8526.n188 4.5005
R462 a_1821_8526.n10 a_1821_8526.n136 4.5005
R463 a_1821_8526.n10 a_1821_8526.n139 4.5005
R464 a_1821_8526.n13 a_1821_8526.n111 4.5005
R465 a_1821_8526.n112 a_1821_8526.n118 4.5005
R466 a_1821_8526.n3 a_1821_8526.n126 4.5005
R467 a_1821_8526.n3 a_1821_8526.n124 4.5005
R468 a_1821_8526.n1 a_1821_8526.n168 4.5005
R469 a_1821_8526.n1 a_1821_8526.n156 4.5005
R470 a_1821_8526.n1 a_1821_8526.n148 4.5005
R471 a_1821_8526.n2 a_1821_8526.n17 4.5005
R472 a_1821_8526.n2 a_1821_8526.n35 4.5005
R473 a_1821_8526.n2 a_1821_8526.n44 4.5005
R474 a_1821_8526.n12 a_1821_8526.n194 4.5005
R475 a_1821_8526.n2 a_1821_8526.n20 4.5005
R476 a_1821_8526.n11 a_1821_8526.n171 4.23684
R477 a_1821_8526.n148 a_1821_8526.n142 4.14168
R478 a_1821_8526.n118 a_1821_8526.n117 4.14168
R479 a_1821_8526.n44 a_1821_8526.n38 4.14168
R480 a_1821_8526.n47 a_1821_8526.n45 3.76521
R481 a_1821_8526.n9 a_1821_8526.n49 3.42768
R482 a_1821_8526.n124 a_1821_8526.n120 3.38874
R483 a_1821_8526.n156 a_1821_8526.n149 3.38874
R484 a_1821_8526.n35 a_1821_8526.n28 3.38874
R485 a_1821_8526.n132 a_1821_8526.n131 3.38537
R486 a_1821_8526.n176 a_1821_8526.n175 3.2936
R487 a_1821_8526.n0 a_1821_8526.n191 3.03311
R488 a_1821_8526.n1 a_1821_8526.n170 3.03311
R489 a_1821_8526.n2 a_1821_8526.n37 3.03311
R490 a_1821_8526.n165 a_1821_8526.n164 3.01226
R491 a_1821_8526.n26 a_1821_8526.n25 3.01226
R492 a_1821_8526.n3 a_1821_8526.n129 2.57905
R493 a_1821_8526.n123 a_1821_8526.n122 2.25932
R494 a_1821_8526.n155 a_1821_8526.n154 2.25932
R495 a_1821_8526.n118 a_1821_8526.n113 2.25932
R496 a_1821_8526.n34 a_1821_8526.n33 2.25932
R497 a_1821_8526.n15 a_1821_8526.n13 2.25727
R498 a_1821_8526.n15 a_1821_8526.n112 2.29192
R499 a_1821_8526.n189 a_1821_8526.n133 1.90999
R500 a_1821_8526.n147 a_1821_8526.n146 1.88285
R501 a_1821_8526.n166 a_1821_8526.n165 1.88285
R502 a_1821_8526.n47 a_1821_8526.n46 1.88285
R503 a_1821_8526.n43 a_1821_8526.n42 1.88285
R504 a_1821_8526.n27 a_1821_8526.n26 1.88285
R505 a_1821_8526.n0 a_1821_8526.n192 1.72048
R506 a_1821_8526.n133 a_1821_8526.n10 1.67144
R507 a_1821_8526.n128 a_1821_8526.n127 1.50638
R508 a_1821_8526.n158 a_1821_8526.n157 1.50638
R509 a_1821_8526.n20 a_1821_8526.n19 1.50638
R510 a_1821_8526.n14 a_1821_8526.n3 1.28885
R511 a_1821_8526.n14 a_1821_8526.n0 1.22346
R512 a_1821_8526.n185 a_1821_8526.n181 1.12991
R513 a_1821_8526.n201 a_1821_8526.n197 1.12991
R514 a_1821_8526.n189 a_1821_8526.n1 1.07918
R515 a_1821_8526.n116 a_1821_8526.n115 0.994314
R516 a_1821_8526.n106 a_1821_8526.n105 0.994314
R517 a_1821_8526.n94 a_1821_8526.n93 0.994314
R518 a_1821_8526.n86 a_1821_8526.n85 0.994314
R519 a_1821_8526.n74 a_1821_8526.n73 0.994314
R520 a_1821_8526.n66 a_1821_8526.n65 0.994314
R521 a_1821_8526.n54 a_1821_8526.n53 0.994314
R522 a_1821_8526.n126 a_1821_8526.n125 0.753441
R523 a_1821_8526.n188 a_1821_8526.n187 0.753441
R524 a_1821_8526.n168 a_1821_8526.n167 0.753441
R525 a_1821_8526.n107 a_1821_8526.n103 0.753441
R526 a_1821_8526.n95 a_1821_8526.n91 0.753441
R527 a_1821_8526.n87 a_1821_8526.n83 0.753441
R528 a_1821_8526.n75 a_1821_8526.n71 0.753441
R529 a_1821_8526.n67 a_1821_8526.n63 0.753441
R530 a_1821_8526.n55 a_1821_8526.n51 0.753441
R531 a_1821_8526.n194 a_1821_8526.n193 0.753441
R532 a_1821_8526.n17 a_1821_8526.n16 0.753441
R533 a_1821_8526.n12 a_1821_8526.n119 0.737441
R534 a_1821_8526.n119 a_1821_8526.n14 0.718062
R535 a_1821_8526.n1 a_1821_8526.n11 0.676808
R536 a_1821_8526.n7 a_1821_8526.n9 0.6634
R537 a_1821_8526.n5 a_1821_8526.n8 0.6634
R538 a_1821_8526.n4 a_1821_8526.n6 0.6634
R539 a_1821_8526.n12 a_1821_8526.n2 0.631263
R540 a_1821_8526.n8 a_1821_8526.n7 0.585981
R541 a_1821_8526.n6 a_1821_8526.n5 0.585981
R542 a_1821_8526.n14 a_1821_8526.n189 0.511626
R543 a_1821_8526.n13 a_1821_8526.n4 0.447235
R544 a_1821_8526.n119 a_1821_8526.n15 0.389962
R545 a_1821_8526.n124 a_1821_8526.n123 0.376971
R546 a_1821_8526.n122 a_1821_8526.n121 0.376971
R547 a_1821_8526.n177 a_1821_8526.n173 0.376971
R548 a_1821_8526.n148 a_1821_8526.n147 0.376971
R549 a_1821_8526.n156 a_1821_8526.n155 0.376971
R550 a_1821_8526.n154 a_1821_8526.n153 0.376971
R551 a_1821_8526.n136 a_1821_8526.n135 0.376971
R552 a_1821_8526.n139 a_1821_8526.n138 0.376971
R553 a_1821_8526.n44 a_1821_8526.n43 0.376971
R554 a_1821_8526.n35 a_1821_8526.n34 0.376971
R555 a_1821_8526.n33 a_1821_8526.n32 0.376971
R556 VDD.n3426 VDD.t70 840.188
R557 VDD.n3426 VDD.t127 840.188
R558 VDD.n3423 VDD.t71 403.574
R559 VDD.n3422 VDD.t128 403.574
R560 VDD.n1922 VDD.n1805 373.449
R561 VDD.n1828 VDD.n1802 373.449
R562 VDD.n2375 VDD.n2374 373.449
R563 VDD.n2391 VDD.n2217 373.449
R564 VDD.n1068 VDD.n951 373.449
R565 VDD.n974 VDD.n948 373.449
R566 VDD.n1521 VDD.n1520 373.449
R567 VDD.n1537 VDD.n1363 373.449
R568 VDD.n213 VDD.n96 373.449
R569 VDD.n119 VDD.n93 373.449
R570 VDD.n666 VDD.n665 373.449
R571 VDD.n682 VDD.n508 373.449
R572 VDD.n5235 VDD.n5234 357.288
R573 VDD.n3810 VDD.n3809 357.288
R574 VDD.n2304 VDD.n2233 351.829
R575 VDD.n2325 VDD.n2324 351.829
R576 VDD.n1935 VDD.n1824 351.829
R577 VDD.n1937 VDD.n1821 351.829
R578 VDD.n1450 VDD.n1379 351.829
R579 VDD.n1471 VDD.n1470 351.829
R580 VDD.n1081 VDD.n970 351.829
R581 VDD.n1083 VDD.n967 351.829
R582 VDD.n595 VDD.n524 351.829
R583 VDD.n616 VDD.n615 351.829
R584 VDD.n226 VDD.n115 351.829
R585 VDD.n228 VDD.n112 351.829
R586 VDD.n55 VDD.n37 321.882
R587 VDD.n41 VDD.n36 321.882
R588 VDD.n18 VDD.n10 321.882
R589 VDD.n31 VDD.n10 321.882
R590 VDD.n31 VDD.n8 321.882
R591 VDD.n60 VDD.n8 321.882
R592 VDD.n906 VDD.n899 321.882
R593 VDD.n898 VDD.n860 321.882
R594 VDD.n878 VDD.n869 321.882
R595 VDD.n881 VDD.n869 321.882
R596 VDD.n881 VDD.n862 321.882
R597 VDD.n894 VDD.n862 321.882
R598 VDD.n1764 VDD.n1746 321.882
R599 VDD.n1750 VDD.n1745 321.882
R600 VDD.n1727 VDD.n1719 321.882
R601 VDD.n1740 VDD.n1719 321.882
R602 VDD.n1740 VDD.n1717 321.882
R603 VDD.n1769 VDD.n1717 321.882
R604 VDD.n59 VDD.n58 266.731
R605 VDD.n896 VDD.n895 266.731
R606 VDD.n1768 VDD.n1767 266.731
R607 VDD.n915 VDD.t58 240.534
R608 VDD.n2624 VDD.t66 240.534
R609 VDD.n2270 VDD.n2246 239.793
R610 VDD.n2270 VDD.n2269 239.793
R611 VDD.n2260 VDD.n2243 239.793
R612 VDD.n2265 VDD.n2260 239.793
R613 VDD.n2353 VDD.n2251 239.793
R614 VDD.n2546 VDD.n1797 239.793
R615 VDD.n2351 VDD.n2284 239.793
R616 VDD.n2548 VDD.n1793 239.793
R617 VDD.n1416 VDD.n1392 239.793
R618 VDD.n1416 VDD.n1415 239.793
R619 VDD.n1406 VDD.n1389 239.793
R620 VDD.n1411 VDD.n1406 239.793
R621 VDD.n1499 VDD.n1397 239.793
R622 VDD.n1692 VDD.n943 239.793
R623 VDD.n1497 VDD.n1430 239.793
R624 VDD.n1694 VDD.n939 239.793
R625 VDD.n561 VDD.n537 239.793
R626 VDD.n561 VDD.n560 239.793
R627 VDD.n551 VDD.n534 239.793
R628 VDD.n556 VDD.n551 239.793
R629 VDD.n644 VDD.n542 239.793
R630 VDD.n837 VDD.n88 239.793
R631 VDD.n642 VDD.n575 239.793
R632 VDD.n839 VDD.n84 239.793
R633 VDD.n48 VDD.t73 239.697
R634 VDD.n1757 VDD.t153 239.697
R635 VDD.n2251 VDD.n2250 218.173
R636 VDD.n1827 VDD.n1797 218.173
R637 VDD.n2330 VDD.n2284 218.173
R638 VDD.n1927 VDD.n1793 218.173
R639 VDD.n1397 VDD.n1396 218.173
R640 VDD.n973 VDD.n943 218.173
R641 VDD.n1476 VDD.n1430 218.173
R642 VDD.n1073 VDD.n939 218.173
R643 VDD.n542 VDD.n541 218.173
R644 VDD.n118 VDD.n88 218.173
R645 VDD.n621 VDD.n575 218.173
R646 VDD.n218 VDD.n84 218.173
R647 VDD.n57 VDD.t72 217.947
R648 VDD.n908 VDD.t57 217.947
R649 VDD.n1766 VDD.t152 217.947
R650 VDD.n2617 VDD.t65 217.947
R651 VDD.n2106 VDD.n2076 205.079
R652 VDD.n2106 VDD.n2105 205.079
R653 VDD.n2105 VDD.n2104 205.079
R654 VDD.n2104 VDD.n2077 205.079
R655 VDD.n2098 VDD.n2077 205.079
R656 VDD.n2098 VDD.n2097 205.079
R657 VDD.n2097 VDD.n2096 205.079
R658 VDD.n2096 VDD.n2081 205.079
R659 VDD.n2090 VDD.n2081 205.079
R660 VDD.n2090 VDD.n2089 205.079
R661 VDD.n2089 VDD.n2088 205.079
R662 VDD.n2088 VDD.n1813 205.079
R663 VDD.n2531 VDD.n1813 205.079
R664 VDD.n2185 VDD.n2034 205.079
R665 VDD.n2191 VDD.n2034 205.079
R666 VDD.n2192 VDD.n2191 205.079
R667 VDD.n2193 VDD.n2192 205.079
R668 VDD.n2193 VDD.n2030 205.079
R669 VDD.n2199 VDD.n2030 205.079
R670 VDD.n2200 VDD.n2199 205.079
R671 VDD.n2201 VDD.n2200 205.079
R672 VDD.n2201 VDD.n2026 205.079
R673 VDD.n2207 VDD.n2026 205.079
R674 VDD.n2208 VDD.n2207 205.079
R675 VDD.n2210 VDD.n2208 205.079
R676 VDD.n2210 VDD.n2209 205.079
R677 VDD.n2529 VDD.n1815 205.079
R678 VDD.n2523 VDD.n1815 205.079
R679 VDD.n2523 VDD.n2522 205.079
R680 VDD.n2522 VDD.n2521 205.079
R681 VDD.n2521 VDD.n1943 205.079
R682 VDD.n2515 VDD.n1943 205.079
R683 VDD.n2515 VDD.n2514 205.079
R684 VDD.n2514 VDD.n2513 205.079
R685 VDD.n2513 VDD.n1947 205.079
R686 VDD.n2507 VDD.n1947 205.079
R687 VDD.n2507 VDD.n2506 205.079
R688 VDD.n2506 VDD.n2505 205.079
R689 VDD.n2505 VDD.n1951 205.079
R690 VDD.n2407 VDD.n2000 205.079
R691 VDD.n2408 VDD.n2407 205.079
R692 VDD.n2409 VDD.n2408 205.079
R693 VDD.n2409 VDD.n1996 205.079
R694 VDD.n2415 VDD.n1996 205.079
R695 VDD.n2416 VDD.n2415 205.079
R696 VDD.n2417 VDD.n2416 205.079
R697 VDD.n2417 VDD.n1992 205.079
R698 VDD.n2423 VDD.n1992 205.079
R699 VDD.n2424 VDD.n2423 205.079
R700 VDD.n2425 VDD.n2424 205.079
R701 VDD.n2425 VDD.n1987 205.079
R702 VDD.n2432 VDD.n1987 205.079
R703 VDD.n1252 VDD.n1222 205.079
R704 VDD.n1252 VDD.n1251 205.079
R705 VDD.n1251 VDD.n1250 205.079
R706 VDD.n1250 VDD.n1223 205.079
R707 VDD.n1244 VDD.n1223 205.079
R708 VDD.n1244 VDD.n1243 205.079
R709 VDD.n1243 VDD.n1242 205.079
R710 VDD.n1242 VDD.n1227 205.079
R711 VDD.n1236 VDD.n1227 205.079
R712 VDD.n1236 VDD.n1235 205.079
R713 VDD.n1235 VDD.n1234 205.079
R714 VDD.n1234 VDD.n959 205.079
R715 VDD.n1677 VDD.n959 205.079
R716 VDD.n1331 VDD.n1180 205.079
R717 VDD.n1337 VDD.n1180 205.079
R718 VDD.n1338 VDD.n1337 205.079
R719 VDD.n1339 VDD.n1338 205.079
R720 VDD.n1339 VDD.n1176 205.079
R721 VDD.n1345 VDD.n1176 205.079
R722 VDD.n1346 VDD.n1345 205.079
R723 VDD.n1347 VDD.n1346 205.079
R724 VDD.n1347 VDD.n1172 205.079
R725 VDD.n1353 VDD.n1172 205.079
R726 VDD.n1354 VDD.n1353 205.079
R727 VDD.n1356 VDD.n1354 205.079
R728 VDD.n1356 VDD.n1355 205.079
R729 VDD.n1675 VDD.n961 205.079
R730 VDD.n1669 VDD.n961 205.079
R731 VDD.n1669 VDD.n1668 205.079
R732 VDD.n1668 VDD.n1667 205.079
R733 VDD.n1667 VDD.n1089 205.079
R734 VDD.n1661 VDD.n1089 205.079
R735 VDD.n1661 VDD.n1660 205.079
R736 VDD.n1660 VDD.n1659 205.079
R737 VDD.n1659 VDD.n1093 205.079
R738 VDD.n1653 VDD.n1093 205.079
R739 VDD.n1653 VDD.n1652 205.079
R740 VDD.n1652 VDD.n1651 205.079
R741 VDD.n1651 VDD.n1097 205.079
R742 VDD.n1553 VDD.n1146 205.079
R743 VDD.n1554 VDD.n1553 205.079
R744 VDD.n1555 VDD.n1554 205.079
R745 VDD.n1555 VDD.n1142 205.079
R746 VDD.n1561 VDD.n1142 205.079
R747 VDD.n1562 VDD.n1561 205.079
R748 VDD.n1563 VDD.n1562 205.079
R749 VDD.n1563 VDD.n1138 205.079
R750 VDD.n1569 VDD.n1138 205.079
R751 VDD.n1570 VDD.n1569 205.079
R752 VDD.n1571 VDD.n1570 205.079
R753 VDD.n1571 VDD.n1133 205.079
R754 VDD.n1578 VDD.n1133 205.079
R755 VDD.n397 VDD.n367 205.079
R756 VDD.n397 VDD.n396 205.079
R757 VDD.n396 VDD.n395 205.079
R758 VDD.n395 VDD.n368 205.079
R759 VDD.n389 VDD.n368 205.079
R760 VDD.n389 VDD.n388 205.079
R761 VDD.n388 VDD.n387 205.079
R762 VDD.n387 VDD.n372 205.079
R763 VDD.n381 VDD.n372 205.079
R764 VDD.n381 VDD.n380 205.079
R765 VDD.n380 VDD.n379 205.079
R766 VDD.n379 VDD.n104 205.079
R767 VDD.n822 VDD.n104 205.079
R768 VDD.n476 VDD.n325 205.079
R769 VDD.n482 VDD.n325 205.079
R770 VDD.n483 VDD.n482 205.079
R771 VDD.n484 VDD.n483 205.079
R772 VDD.n484 VDD.n321 205.079
R773 VDD.n490 VDD.n321 205.079
R774 VDD.n491 VDD.n490 205.079
R775 VDD.n492 VDD.n491 205.079
R776 VDD.n492 VDD.n317 205.079
R777 VDD.n498 VDD.n317 205.079
R778 VDD.n499 VDD.n498 205.079
R779 VDD.n501 VDD.n499 205.079
R780 VDD.n501 VDD.n500 205.079
R781 VDD.n820 VDD.n106 205.079
R782 VDD.n814 VDD.n106 205.079
R783 VDD.n814 VDD.n813 205.079
R784 VDD.n813 VDD.n812 205.079
R785 VDD.n812 VDD.n234 205.079
R786 VDD.n806 VDD.n234 205.079
R787 VDD.n806 VDD.n805 205.079
R788 VDD.n805 VDD.n804 205.079
R789 VDD.n804 VDD.n238 205.079
R790 VDD.n798 VDD.n238 205.079
R791 VDD.n798 VDD.n797 205.079
R792 VDD.n797 VDD.n796 205.079
R793 VDD.n796 VDD.n242 205.079
R794 VDD.n698 VDD.n291 205.079
R795 VDD.n699 VDD.n698 205.079
R796 VDD.n700 VDD.n699 205.079
R797 VDD.n700 VDD.n287 205.079
R798 VDD.n706 VDD.n287 205.079
R799 VDD.n707 VDD.n706 205.079
R800 VDD.n708 VDD.n707 205.079
R801 VDD.n708 VDD.n283 205.079
R802 VDD.n714 VDD.n283 205.079
R803 VDD.n715 VDD.n714 205.079
R804 VDD.n716 VDD.n715 205.079
R805 VDD.n716 VDD.n278 205.079
R806 VDD.n723 VDD.n278 205.079
R807 VDD.n2440 VDD.n1982 203.786
R808 VDD.n2441 VDD.n2440 203.786
R809 VDD.n2442 VDD.n2441 203.786
R810 VDD.n2442 VDD.n1978 203.786
R811 VDD.n2448 VDD.n1978 203.786
R812 VDD.n2449 VDD.n2448 203.786
R813 VDD.n2450 VDD.n2449 203.786
R814 VDD.n2450 VDD.n1974 203.786
R815 VDD.n2456 VDD.n1974 203.786
R816 VDD.n2457 VDD.n2456 203.786
R817 VDD.n2458 VDD.n2457 203.786
R818 VDD.n2458 VDD.n1970 203.786
R819 VDD.n2464 VDD.n1970 203.786
R820 VDD.n2465 VDD.n2464 203.786
R821 VDD.n2466 VDD.n2465 203.786
R822 VDD.n2466 VDD.n1966 203.786
R823 VDD.n2472 VDD.n1966 203.786
R824 VDD.n2473 VDD.n2472 203.786
R825 VDD.n2474 VDD.n2473 203.786
R826 VDD.n2474 VDD.n1962 203.786
R827 VDD.n2480 VDD.n1962 203.786
R828 VDD.n2481 VDD.n2480 203.786
R829 VDD.n2482 VDD.n2481 203.786
R830 VDD.n2482 VDD.n1958 203.786
R831 VDD.n2488 VDD.n1958 203.786
R832 VDD.n2489 VDD.n2488 203.786
R833 VDD.n2492 VDD.n2489 203.786
R834 VDD.n2492 VDD.n2491 203.786
R835 VDD.n1586 VDD.n1128 203.786
R836 VDD.n1587 VDD.n1586 203.786
R837 VDD.n1588 VDD.n1587 203.786
R838 VDD.n1588 VDD.n1124 203.786
R839 VDD.n1594 VDD.n1124 203.786
R840 VDD.n1595 VDD.n1594 203.786
R841 VDD.n1596 VDD.n1595 203.786
R842 VDD.n1596 VDD.n1120 203.786
R843 VDD.n1602 VDD.n1120 203.786
R844 VDD.n1603 VDD.n1602 203.786
R845 VDD.n1604 VDD.n1603 203.786
R846 VDD.n1604 VDD.n1116 203.786
R847 VDD.n1610 VDD.n1116 203.786
R848 VDD.n1611 VDD.n1610 203.786
R849 VDD.n1612 VDD.n1611 203.786
R850 VDD.n1612 VDD.n1112 203.786
R851 VDD.n1618 VDD.n1112 203.786
R852 VDD.n1619 VDD.n1618 203.786
R853 VDD.n1620 VDD.n1619 203.786
R854 VDD.n1620 VDD.n1108 203.786
R855 VDD.n1626 VDD.n1108 203.786
R856 VDD.n1627 VDD.n1626 203.786
R857 VDD.n1628 VDD.n1627 203.786
R858 VDD.n1628 VDD.n1104 203.786
R859 VDD.n1634 VDD.n1104 203.786
R860 VDD.n1635 VDD.n1634 203.786
R861 VDD.n1638 VDD.n1635 203.786
R862 VDD.n1638 VDD.n1637 203.786
R863 VDD.n731 VDD.n273 203.786
R864 VDD.n732 VDD.n731 203.786
R865 VDD.n733 VDD.n732 203.786
R866 VDD.n733 VDD.n269 203.786
R867 VDD.n739 VDD.n269 203.786
R868 VDD.n740 VDD.n739 203.786
R869 VDD.n741 VDD.n740 203.786
R870 VDD.n741 VDD.n265 203.786
R871 VDD.n747 VDD.n265 203.786
R872 VDD.n748 VDD.n747 203.786
R873 VDD.n749 VDD.n748 203.786
R874 VDD.n749 VDD.n261 203.786
R875 VDD.n755 VDD.n261 203.786
R876 VDD.n756 VDD.n755 203.786
R877 VDD.n757 VDD.n756 203.786
R878 VDD.n757 VDD.n257 203.786
R879 VDD.n763 VDD.n257 203.786
R880 VDD.n764 VDD.n763 203.786
R881 VDD.n765 VDD.n764 203.786
R882 VDD.n765 VDD.n253 203.786
R883 VDD.n771 VDD.n253 203.786
R884 VDD.n772 VDD.n771 203.786
R885 VDD.n773 VDD.n772 203.786
R886 VDD.n773 VDD.n249 203.786
R887 VDD.n779 VDD.n249 203.786
R888 VDD.n780 VDD.n779 203.786
R889 VDD.n783 VDD.n780 203.786
R890 VDD.n783 VDD.n782 203.786
R891 VDD.n32 VDD.n9 175.386
R892 VDD.n59 VDD.n33 175.386
R893 VDD.n880 VDD.n879 175.386
R894 VDD.n895 VDD.n861 175.386
R895 VDD.n1741 VDD.n1718 175.386
R896 VDD.n1768 VDD.n1742 175.386
R897 VDD.n18 VDD.t53 171.452
R898 VDD.t23 VDD.n878 171.452
R899 VDD.n1727 VDD.t61 171.452
R900 VDD.n2530 VDD.n2529 168.889
R901 VDD.n2004 VDD.n2000 168.889
R902 VDD.n1676 VDD.n1675 168.889
R903 VDD.n1150 VDD.n1146 168.889
R904 VDD.n821 VDD.n820 168.889
R905 VDD.n295 VDD.n291 168.889
R906 VDD.n2434 VDD.n2433 164.827
R907 VDD.n1580 VDD.n1579 164.827
R908 VDD.n725 VDD.n724 164.827
R909 VDD.n2490 VDD.n1951 162.857
R910 VDD.n2433 VDD.n2432 162.857
R911 VDD.n1636 VDD.n1097 162.857
R912 VDD.n1579 VDD.n1578 162.857
R913 VDD.n781 VDD.n242 162.857
R914 VDD.n724 VDD.n723 162.857
R915 VDD.n2490 VDD.n1954 161.831
R916 VDD.n1636 VDD.n1100 161.831
R917 VDD.n781 VDD.n245 161.831
R918 VDD.n21 VDD.t54 160.743
R919 VDD.n870 VDD.t24 160.743
R920 VDD.n1730 VDD.t62 160.743
R921 VDD.n2573 VDD.t136 160.743
R922 VDD.n2389 VDD.n2004 160.256
R923 VDD.n1535 VDD.n1150 160.256
R924 VDD.n680 VDD.n295 160.256
R925 VDD.n2183 VDD.n2039 159.113
R926 VDD.n2169 VDD.n2039 159.113
R927 VDD.n2169 VDD.n2168 159.113
R928 VDD.n2168 VDD.n2167 159.113
R929 VDD.n2167 VDD.n2044 159.113
R930 VDD.n2161 VDD.n2044 159.113
R931 VDD.n2161 VDD.n2160 159.113
R932 VDD.n2160 VDD.n2159 159.113
R933 VDD.n2159 VDD.n2048 159.113
R934 VDD.n2153 VDD.n2048 159.113
R935 VDD.n2153 VDD.n2152 159.113
R936 VDD.n2152 VDD.n2151 159.113
R937 VDD.n2151 VDD.n2052 159.113
R938 VDD.n2145 VDD.n2052 159.113
R939 VDD.n2145 VDD.n2144 159.113
R940 VDD.n2144 VDD.n2143 159.113
R941 VDD.n2143 VDD.n2056 159.113
R942 VDD.n2137 VDD.n2056 159.113
R943 VDD.n2137 VDD.n2136 159.113
R944 VDD.n2136 VDD.n2135 159.113
R945 VDD.n2135 VDD.n2060 159.113
R946 VDD.n2129 VDD.n2060 159.113
R947 VDD.n2129 VDD.n2128 159.113
R948 VDD.n2128 VDD.n2127 159.113
R949 VDD.n2127 VDD.n2064 159.113
R950 VDD.n2121 VDD.n2064 159.113
R951 VDD.n2121 VDD.n2120 159.113
R952 VDD.n2120 VDD.n2119 159.113
R953 VDD.n1329 VDD.n1185 159.113
R954 VDD.n1315 VDD.n1185 159.113
R955 VDD.n1315 VDD.n1314 159.113
R956 VDD.n1314 VDD.n1313 159.113
R957 VDD.n1313 VDD.n1190 159.113
R958 VDD.n1307 VDD.n1190 159.113
R959 VDD.n1307 VDD.n1306 159.113
R960 VDD.n1306 VDD.n1305 159.113
R961 VDD.n1305 VDD.n1194 159.113
R962 VDD.n1299 VDD.n1194 159.113
R963 VDD.n1299 VDD.n1298 159.113
R964 VDD.n1298 VDD.n1297 159.113
R965 VDD.n1297 VDD.n1198 159.113
R966 VDD.n1291 VDD.n1198 159.113
R967 VDD.n1291 VDD.n1290 159.113
R968 VDD.n1290 VDD.n1289 159.113
R969 VDD.n1289 VDD.n1202 159.113
R970 VDD.n1283 VDD.n1202 159.113
R971 VDD.n1283 VDD.n1282 159.113
R972 VDD.n1282 VDD.n1281 159.113
R973 VDD.n1281 VDD.n1206 159.113
R974 VDD.n1275 VDD.n1206 159.113
R975 VDD.n1275 VDD.n1274 159.113
R976 VDD.n1274 VDD.n1273 159.113
R977 VDD.n1273 VDD.n1210 159.113
R978 VDD.n1267 VDD.n1210 159.113
R979 VDD.n1267 VDD.n1266 159.113
R980 VDD.n1266 VDD.n1265 159.113
R981 VDD.n474 VDD.n330 159.113
R982 VDD.n460 VDD.n330 159.113
R983 VDD.n460 VDD.n459 159.113
R984 VDD.n459 VDD.n458 159.113
R985 VDD.n458 VDD.n335 159.113
R986 VDD.n452 VDD.n335 159.113
R987 VDD.n452 VDD.n451 159.113
R988 VDD.n451 VDD.n450 159.113
R989 VDD.n450 VDD.n339 159.113
R990 VDD.n444 VDD.n339 159.113
R991 VDD.n444 VDD.n443 159.113
R992 VDD.n443 VDD.n442 159.113
R993 VDD.n442 VDD.n343 159.113
R994 VDD.n436 VDD.n343 159.113
R995 VDD.n436 VDD.n435 159.113
R996 VDD.n435 VDD.n434 159.113
R997 VDD.n434 VDD.n347 159.113
R998 VDD.n428 VDD.n347 159.113
R999 VDD.n428 VDD.n427 159.113
R1000 VDD.n427 VDD.n426 159.113
R1001 VDD.n426 VDD.n351 159.113
R1002 VDD.n420 VDD.n351 159.113
R1003 VDD.n420 VDD.n419 159.113
R1004 VDD.n419 VDD.n418 159.113
R1005 VDD.n418 VDD.n355 159.113
R1006 VDD.n412 VDD.n355 159.113
R1007 VDD.n412 VDD.n411 159.113
R1008 VDD.n411 VDD.n410 159.113
R1009 VDD.n13 VDD.t56 158.225
R1010 VDD.n891 VDD.t26 158.225
R1011 VDD.n1722 VDD.t64 158.225
R1012 VDD.n2571 VDD.t134 158.225
R1013 VDD.n2530 VDD.n1814 154.488
R1014 VDD.n1676 VDD.n960 154.488
R1015 VDD.n821 VDD.n105 154.488
R1016 VDD.t10 VDD.t60 151.181
R1017 VDD.t110 VDD.t129 151.181
R1018 VDD.t129 VDD.t0 151.181
R1019 VDD.t102 VDD.t2 151.181
R1020 VDD.t125 VDD.t102 151.181
R1021 VDD.t97 VDD.t125 151.181
R1022 VDD.t90 VDD.t97 151.181
R1023 VDD.n2182 VDD.n2040 141.731
R1024 VDD.n2118 VDD.n2069 141.731
R1025 VDD.n1328 VDD.n1186 141.731
R1026 VDD.n1264 VDD.n1215 141.731
R1027 VDD.n473 VDD.n331 141.731
R1028 VDD.n409 VDD.n360 141.731
R1029 VDD.n2435 VDD.n1983 140.19
R1030 VDD.n2497 VDD.n1955 140.19
R1031 VDD.n1581 VDD.n1129 140.19
R1032 VDD.n1643 VDD.n1101 140.19
R1033 VDD.n726 VDD.n274 140.19
R1034 VDD.n788 VDD.n246 140.19
R1035 VDD.n2662 VDD.n2658 133.655
R1036 VDD.n2917 VDD.n2916 133.655
R1037 VDD.n3045 VDD.n3044 133.655
R1038 VDD.n2645 VDD.n2644 133.655
R1039 VDD.n3398 VDD.n3395 133.655
R1040 VDD.n3314 VDD.n3313 133.655
R1041 VDD.n2335 VDD.n2251 133.655
R1042 VDD.n2346 VDD.n2284 133.655
R1043 VDD.n2281 VDD.n2260 133.655
R1044 VDD.n2277 VDD.n2259 133.655
R1045 VDD.n2275 VDD.n2274 133.655
R1046 VDD.n2271 VDD.n2270 133.655
R1047 VDD.n1836 VDD.n1828 133.655
R1048 VDD.n2374 VDD.n2229 133.655
R1049 VDD.n2366 VDD.n2229 133.655
R1050 VDD.n2366 VDD.n2236 133.655
R1051 VDD.n2358 VDD.n2236 133.655
R1052 VDD.n2358 VDD.n2246 133.655
R1053 VDD.n2269 VDD.n2268 133.655
R1054 VDD.n2268 VDD.n1801 133.655
R1055 VDD.n2543 VDD.n1801 133.655
R1056 VDD.n2543 VDD.n2542 133.655
R1057 VDD.n2542 VDD.n1802 133.655
R1058 VDD.n2387 VDD.n2218 133.655
R1059 VDD.n2379 VDD.n2224 133.655
R1060 VDD.n2239 VDD.n2217 133.655
R1061 VDD.n2364 VDD.n2239 133.655
R1062 VDD.n2364 VDD.n2240 133.655
R1063 VDD.n2360 VDD.n2240 133.655
R1064 VDD.n2360 VDD.n2243 133.655
R1065 VDD.n2265 VDD.n2264 133.655
R1066 VDD.n2264 VDD.n2263 133.655
R1067 VDD.n2263 VDD.n1804 133.655
R1068 VDD.n2540 VDD.n1804 133.655
R1069 VDD.n2540 VDD.n1805 133.655
R1070 VDD.n2310 VDD.n2309 133.655
R1071 VDD.n2316 VDD.n2315 133.655
R1072 VDD.n2371 VDD.n2233 133.655
R1073 VDD.n2371 VDD.n2234 133.655
R1074 VDD.n2250 VDD.n2234 133.655
R1075 VDD.n2353 VDD.n2255 133.655
R1076 VDD.n2255 VDD.n1785 133.655
R1077 VDD.n2554 VDD.n1785 133.655
R1078 VDD.n2554 VDD.n1786 133.655
R1079 VDD.n2546 VDD.n1786 133.655
R1080 VDD.n1932 VDD.n1827 133.655
R1081 VDD.n1935 VDD.n1823 133.655
R1082 VDD.n1867 VDD.n1866 133.655
R1083 VDD.n1858 VDD.n1856 133.655
R1084 VDD.n2325 VDD.n2232 133.655
R1085 VDD.n2329 VDD.n2232 133.655
R1086 VDD.n2330 VDD.n2329 133.655
R1087 VDD.n2351 VDD.n2287 133.655
R1088 VDD.n2287 VDD.n1789 133.655
R1089 VDD.n2552 VDD.n1789 133.655
R1090 VDD.n2552 VDD.n1790 133.655
R1091 VDD.n2548 VDD.n1790 133.655
R1092 VDD.n1930 VDD.n1927 133.655
R1093 VDD.n1930 VDD.n1820 133.655
R1094 VDD.n1937 VDD.n1820 133.655
R1095 VDD.n1893 VDD.n1797 133.655
R1096 VDD.n1882 VDD.n1793 133.655
R1097 VDD.n1481 VDD.n1397 133.655
R1098 VDD.n1492 VDD.n1430 133.655
R1099 VDD.n1427 VDD.n1406 133.655
R1100 VDD.n1423 VDD.n1405 133.655
R1101 VDD.n1421 VDD.n1420 133.655
R1102 VDD.n1417 VDD.n1416 133.655
R1103 VDD.n982 VDD.n974 133.655
R1104 VDD.n1520 VDD.n1375 133.655
R1105 VDD.n1512 VDD.n1375 133.655
R1106 VDD.n1512 VDD.n1382 133.655
R1107 VDD.n1504 VDD.n1382 133.655
R1108 VDD.n1504 VDD.n1392 133.655
R1109 VDD.n1415 VDD.n1414 133.655
R1110 VDD.n1414 VDD.n947 133.655
R1111 VDD.n1689 VDD.n947 133.655
R1112 VDD.n1689 VDD.n1688 133.655
R1113 VDD.n1688 VDD.n948 133.655
R1114 VDD.n1533 VDD.n1364 133.655
R1115 VDD.n1525 VDD.n1370 133.655
R1116 VDD.n1385 VDD.n1363 133.655
R1117 VDD.n1510 VDD.n1385 133.655
R1118 VDD.n1510 VDD.n1386 133.655
R1119 VDD.n1506 VDD.n1386 133.655
R1120 VDD.n1506 VDD.n1389 133.655
R1121 VDD.n1411 VDD.n1410 133.655
R1122 VDD.n1410 VDD.n1409 133.655
R1123 VDD.n1409 VDD.n950 133.655
R1124 VDD.n1686 VDD.n950 133.655
R1125 VDD.n1686 VDD.n951 133.655
R1126 VDD.n1456 VDD.n1455 133.655
R1127 VDD.n1462 VDD.n1461 133.655
R1128 VDD.n1517 VDD.n1379 133.655
R1129 VDD.n1517 VDD.n1380 133.655
R1130 VDD.n1396 VDD.n1380 133.655
R1131 VDD.n1499 VDD.n1401 133.655
R1132 VDD.n1401 VDD.n931 133.655
R1133 VDD.n1700 VDD.n931 133.655
R1134 VDD.n1700 VDD.n932 133.655
R1135 VDD.n1692 VDD.n932 133.655
R1136 VDD.n1078 VDD.n973 133.655
R1137 VDD.n1081 VDD.n969 133.655
R1138 VDD.n1013 VDD.n1012 133.655
R1139 VDD.n1004 VDD.n1002 133.655
R1140 VDD.n1471 VDD.n1378 133.655
R1141 VDD.n1475 VDD.n1378 133.655
R1142 VDD.n1476 VDD.n1475 133.655
R1143 VDD.n1497 VDD.n1433 133.655
R1144 VDD.n1433 VDD.n935 133.655
R1145 VDD.n1698 VDD.n935 133.655
R1146 VDD.n1698 VDD.n936 133.655
R1147 VDD.n1694 VDD.n936 133.655
R1148 VDD.n1076 VDD.n1073 133.655
R1149 VDD.n1076 VDD.n966 133.655
R1150 VDD.n1083 VDD.n966 133.655
R1151 VDD.n1039 VDD.n943 133.655
R1152 VDD.n1028 VDD.n939 133.655
R1153 VDD.n626 VDD.n542 133.655
R1154 VDD.n637 VDD.n575 133.655
R1155 VDD.n572 VDD.n551 133.655
R1156 VDD.n568 VDD.n550 133.655
R1157 VDD.n566 VDD.n565 133.655
R1158 VDD.n562 VDD.n561 133.655
R1159 VDD.n127 VDD.n119 133.655
R1160 VDD.n665 VDD.n520 133.655
R1161 VDD.n657 VDD.n520 133.655
R1162 VDD.n657 VDD.n527 133.655
R1163 VDD.n649 VDD.n527 133.655
R1164 VDD.n649 VDD.n537 133.655
R1165 VDD.n560 VDD.n559 133.655
R1166 VDD.n559 VDD.n92 133.655
R1167 VDD.n834 VDD.n92 133.655
R1168 VDD.n834 VDD.n833 133.655
R1169 VDD.n833 VDD.n93 133.655
R1170 VDD.n678 VDD.n509 133.655
R1171 VDD.n670 VDD.n515 133.655
R1172 VDD.n530 VDD.n508 133.655
R1173 VDD.n655 VDD.n530 133.655
R1174 VDD.n655 VDD.n531 133.655
R1175 VDD.n651 VDD.n531 133.655
R1176 VDD.n651 VDD.n534 133.655
R1177 VDD.n556 VDD.n555 133.655
R1178 VDD.n555 VDD.n554 133.655
R1179 VDD.n554 VDD.n95 133.655
R1180 VDD.n831 VDD.n95 133.655
R1181 VDD.n831 VDD.n96 133.655
R1182 VDD.n601 VDD.n600 133.655
R1183 VDD.n607 VDD.n606 133.655
R1184 VDD.n662 VDD.n524 133.655
R1185 VDD.n662 VDD.n525 133.655
R1186 VDD.n541 VDD.n525 133.655
R1187 VDD.n644 VDD.n546 133.655
R1188 VDD.n546 VDD.n76 133.655
R1189 VDD.n845 VDD.n76 133.655
R1190 VDD.n845 VDD.n77 133.655
R1191 VDD.n837 VDD.n77 133.655
R1192 VDD.n223 VDD.n118 133.655
R1193 VDD.n226 VDD.n114 133.655
R1194 VDD.n158 VDD.n157 133.655
R1195 VDD.n149 VDD.n147 133.655
R1196 VDD.n616 VDD.n523 133.655
R1197 VDD.n620 VDD.n523 133.655
R1198 VDD.n621 VDD.n620 133.655
R1199 VDD.n642 VDD.n578 133.655
R1200 VDD.n578 VDD.n80 133.655
R1201 VDD.n843 VDD.n80 133.655
R1202 VDD.n843 VDD.n81 133.655
R1203 VDD.n839 VDD.n81 133.655
R1204 VDD.n221 VDD.n218 133.655
R1205 VDD.n221 VDD.n111 133.655
R1206 VDD.n228 VDD.n111 133.655
R1207 VDD.n184 VDD.n88 133.655
R1208 VDD.n173 VDD.n84 133.655
R1209 VDD.n2184 VDD.n2038 128.696
R1210 VDD.n1330 VDD.n1184 128.696
R1211 VDD.n475 VDD.n329 128.696
R1212 VDD.n3761 VDD.t90 126.425
R1213 VDD.n2072 VDD.n2068 126.356
R1214 VDD.n1218 VDD.n1214 126.356
R1215 VDD.n363 VDD.n359 126.356
R1216 VDD.t27 VDD.n57 117.838
R1217 VDD.n908 VDD.t145 117.838
R1218 VDD.t157 VDD.n1766 117.838
R1219 VDD.n2617 VDD.t106 117.838
R1220 VDD.n7114 VDD.n7113 117.62
R1221 VDD.n5307 VDD.t95 116.841
R1222 VDD.n8611 VDD.t44 116.841
R1223 VDD.n8973 VDD.t40 116.841
R1224 VDD.n5157 VDD.t92 116.841
R1225 VDD.n8883 VDD.t113 116.841
R1226 VDD.n2170 VDD.n2041 104.757
R1227 VDD.n2170 VDD.n2043 104.757
R1228 VDD.n2166 VDD.n2043 104.757
R1229 VDD.n2166 VDD.n2045 104.757
R1230 VDD.n2162 VDD.n2045 104.757
R1231 VDD.n2162 VDD.n2047 104.757
R1232 VDD.n2158 VDD.n2047 104.757
R1233 VDD.n2158 VDD.n2049 104.757
R1234 VDD.n2154 VDD.n2049 104.757
R1235 VDD.n2154 VDD.n2051 104.757
R1236 VDD.n2150 VDD.n2051 104.757
R1237 VDD.n2150 VDD.n2053 104.757
R1238 VDD.n2146 VDD.n2053 104.757
R1239 VDD.n2146 VDD.n2055 104.757
R1240 VDD.n2142 VDD.n2055 104.757
R1241 VDD.n2142 VDD.n2057 104.757
R1242 VDD.n2138 VDD.n2057 104.757
R1243 VDD.n2138 VDD.n2059 104.757
R1244 VDD.n2134 VDD.n2059 104.757
R1245 VDD.n2134 VDD.n2061 104.757
R1246 VDD.n2130 VDD.n2061 104.757
R1247 VDD.n2130 VDD.n2063 104.757
R1248 VDD.n2126 VDD.n2063 104.757
R1249 VDD.n2126 VDD.n2065 104.757
R1250 VDD.n2122 VDD.n2065 104.757
R1251 VDD.n2122 VDD.n2067 104.757
R1252 VDD.n2118 VDD.n2067 104.757
R1253 VDD.n2186 VDD.n2037 104.757
R1254 VDD.n2186 VDD.n2035 104.757
R1255 VDD.n2190 VDD.n2035 104.757
R1256 VDD.n2190 VDD.n2033 104.757
R1257 VDD.n2194 VDD.n2033 104.757
R1258 VDD.n2194 VDD.n2031 104.757
R1259 VDD.n2198 VDD.n2031 104.757
R1260 VDD.n2198 VDD.n2029 104.757
R1261 VDD.n2202 VDD.n2029 104.757
R1262 VDD.n2202 VDD.n2027 104.757
R1263 VDD.n2206 VDD.n2027 104.757
R1264 VDD.n2206 VDD.n2025 104.757
R1265 VDD.n2211 VDD.n2025 104.757
R1266 VDD.n2211 VDD.n2023 104.757
R1267 VDD.n2398 VDD.n2023 104.757
R1268 VDD.n2377 VDD.n2015 104.757
R1269 VDD.n2294 VDD.n2015 104.757
R1270 VDD.n2298 VDD.n2297 104.757
R1271 VDD.n2402 VDD.n2001 104.757
R1272 VDD.n2406 VDD.n2001 104.757
R1273 VDD.n2406 VDD.n1999 104.757
R1274 VDD.n2410 VDD.n1999 104.757
R1275 VDD.n2410 VDD.n1997 104.757
R1276 VDD.n2414 VDD.n1997 104.757
R1277 VDD.n2414 VDD.n1995 104.757
R1278 VDD.n2418 VDD.n1995 104.757
R1279 VDD.n2418 VDD.n1993 104.757
R1280 VDD.n2422 VDD.n1993 104.757
R1281 VDD.n2422 VDD.n1991 104.757
R1282 VDD.n2426 VDD.n1991 104.757
R1283 VDD.n2426 VDD.n1988 104.757
R1284 VDD.n2431 VDD.n1988 104.757
R1285 VDD.n2431 VDD.n1989 104.757
R1286 VDD.n2435 VDD.n1985 104.757
R1287 VDD.n2439 VDD.n1983 104.757
R1288 VDD.n2439 VDD.n1981 104.757
R1289 VDD.n2443 VDD.n1981 104.757
R1290 VDD.n2443 VDD.n1979 104.757
R1291 VDD.n2447 VDD.n1979 104.757
R1292 VDD.n2447 VDD.n1977 104.757
R1293 VDD.n2451 VDD.n1977 104.757
R1294 VDD.n2451 VDD.n1975 104.757
R1295 VDD.n2455 VDD.n1975 104.757
R1296 VDD.n2455 VDD.n1973 104.757
R1297 VDD.n2459 VDD.n1973 104.757
R1298 VDD.n2459 VDD.n1971 104.757
R1299 VDD.n2463 VDD.n1971 104.757
R1300 VDD.n2463 VDD.n1969 104.757
R1301 VDD.n2467 VDD.n1969 104.757
R1302 VDD.n2467 VDD.n1967 104.757
R1303 VDD.n2471 VDD.n1967 104.757
R1304 VDD.n2471 VDD.n1965 104.757
R1305 VDD.n2475 VDD.n1965 104.757
R1306 VDD.n2475 VDD.n1963 104.757
R1307 VDD.n2479 VDD.n1963 104.757
R1308 VDD.n2479 VDD.n1961 104.757
R1309 VDD.n2483 VDD.n1961 104.757
R1310 VDD.n2483 VDD.n1959 104.757
R1311 VDD.n2487 VDD.n1959 104.757
R1312 VDD.n2487 VDD.n1957 104.757
R1313 VDD.n2493 VDD.n1957 104.757
R1314 VDD.n2493 VDD.n1955 104.757
R1315 VDD.n2114 VDD.n2113 104.757
R1316 VDD.n2111 VDD.n2073 104.757
R1317 VDD.n2107 VDD.n2073 104.757
R1318 VDD.n2107 VDD.n2075 104.757
R1319 VDD.n2103 VDD.n2075 104.757
R1320 VDD.n2103 VDD.n2078 104.757
R1321 VDD.n2099 VDD.n2078 104.757
R1322 VDD.n2099 VDD.n2080 104.757
R1323 VDD.n2095 VDD.n2080 104.757
R1324 VDD.n2095 VDD.n2082 104.757
R1325 VDD.n2091 VDD.n2082 104.757
R1326 VDD.n2091 VDD.n2084 104.757
R1327 VDD.n2087 VDD.n2084 104.757
R1328 VDD.n2087 VDD.n1811 104.757
R1329 VDD.n2532 VDD.n1811 104.757
R1330 VDD.n2533 VDD.n2532 104.757
R1331 VDD.n1919 VDD.n1834 104.757
R1332 VDD.n1917 VDD.n1835 104.757
R1333 VDD.n1909 VDD.n1908 104.757
R1334 VDD.n1904 VDD.n1903 104.757
R1335 VDD.n1872 VDD.n1841 104.757
R1336 VDD.n1863 VDD.n1847 104.757
R1337 VDD.n1861 VDD.n1848 104.757
R1338 VDD.n1852 VDD.n1851 104.757
R1339 VDD.n2528 VDD.n1816 104.757
R1340 VDD.n2528 VDD.n1817 104.757
R1341 VDD.n2524 VDD.n1817 104.757
R1342 VDD.n2524 VDD.n1942 104.757
R1343 VDD.n2520 VDD.n1942 104.757
R1344 VDD.n2520 VDD.n1944 104.757
R1345 VDD.n2516 VDD.n1944 104.757
R1346 VDD.n2516 VDD.n1946 104.757
R1347 VDD.n2512 VDD.n1946 104.757
R1348 VDD.n2512 VDD.n1948 104.757
R1349 VDD.n2508 VDD.n1948 104.757
R1350 VDD.n2508 VDD.n1950 104.757
R1351 VDD.n2504 VDD.n1950 104.757
R1352 VDD.n2504 VDD.n1952 104.757
R1353 VDD.n2500 VDD.n1952 104.757
R1354 VDD.n2498 VDD.n2497 104.757
R1355 VDD.n1316 VDD.n1187 104.757
R1356 VDD.n1316 VDD.n1189 104.757
R1357 VDD.n1312 VDD.n1189 104.757
R1358 VDD.n1312 VDD.n1191 104.757
R1359 VDD.n1308 VDD.n1191 104.757
R1360 VDD.n1308 VDD.n1193 104.757
R1361 VDD.n1304 VDD.n1193 104.757
R1362 VDD.n1304 VDD.n1195 104.757
R1363 VDD.n1300 VDD.n1195 104.757
R1364 VDD.n1300 VDD.n1197 104.757
R1365 VDD.n1296 VDD.n1197 104.757
R1366 VDD.n1296 VDD.n1199 104.757
R1367 VDD.n1292 VDD.n1199 104.757
R1368 VDD.n1292 VDD.n1201 104.757
R1369 VDD.n1288 VDD.n1201 104.757
R1370 VDD.n1288 VDD.n1203 104.757
R1371 VDD.n1284 VDD.n1203 104.757
R1372 VDD.n1284 VDD.n1205 104.757
R1373 VDD.n1280 VDD.n1205 104.757
R1374 VDD.n1280 VDD.n1207 104.757
R1375 VDD.n1276 VDD.n1207 104.757
R1376 VDD.n1276 VDD.n1209 104.757
R1377 VDD.n1272 VDD.n1209 104.757
R1378 VDD.n1272 VDD.n1211 104.757
R1379 VDD.n1268 VDD.n1211 104.757
R1380 VDD.n1268 VDD.n1213 104.757
R1381 VDD.n1264 VDD.n1213 104.757
R1382 VDD.n1332 VDD.n1183 104.757
R1383 VDD.n1332 VDD.n1181 104.757
R1384 VDD.n1336 VDD.n1181 104.757
R1385 VDD.n1336 VDD.n1179 104.757
R1386 VDD.n1340 VDD.n1179 104.757
R1387 VDD.n1340 VDD.n1177 104.757
R1388 VDD.n1344 VDD.n1177 104.757
R1389 VDD.n1344 VDD.n1175 104.757
R1390 VDD.n1348 VDD.n1175 104.757
R1391 VDD.n1348 VDD.n1173 104.757
R1392 VDD.n1352 VDD.n1173 104.757
R1393 VDD.n1352 VDD.n1171 104.757
R1394 VDD.n1357 VDD.n1171 104.757
R1395 VDD.n1357 VDD.n1169 104.757
R1396 VDD.n1544 VDD.n1169 104.757
R1397 VDD.n1523 VDD.n1161 104.757
R1398 VDD.n1440 VDD.n1161 104.757
R1399 VDD.n1444 VDD.n1443 104.757
R1400 VDD.n1548 VDD.n1147 104.757
R1401 VDD.n1552 VDD.n1147 104.757
R1402 VDD.n1552 VDD.n1145 104.757
R1403 VDD.n1556 VDD.n1145 104.757
R1404 VDD.n1556 VDD.n1143 104.757
R1405 VDD.n1560 VDD.n1143 104.757
R1406 VDD.n1560 VDD.n1141 104.757
R1407 VDD.n1564 VDD.n1141 104.757
R1408 VDD.n1564 VDD.n1139 104.757
R1409 VDD.n1568 VDD.n1139 104.757
R1410 VDD.n1568 VDD.n1137 104.757
R1411 VDD.n1572 VDD.n1137 104.757
R1412 VDD.n1572 VDD.n1134 104.757
R1413 VDD.n1577 VDD.n1134 104.757
R1414 VDD.n1577 VDD.n1135 104.757
R1415 VDD.n1581 VDD.n1131 104.757
R1416 VDD.n1585 VDD.n1129 104.757
R1417 VDD.n1585 VDD.n1127 104.757
R1418 VDD.n1589 VDD.n1127 104.757
R1419 VDD.n1589 VDD.n1125 104.757
R1420 VDD.n1593 VDD.n1125 104.757
R1421 VDD.n1593 VDD.n1123 104.757
R1422 VDD.n1597 VDD.n1123 104.757
R1423 VDD.n1597 VDD.n1121 104.757
R1424 VDD.n1601 VDD.n1121 104.757
R1425 VDD.n1601 VDD.n1119 104.757
R1426 VDD.n1605 VDD.n1119 104.757
R1427 VDD.n1605 VDD.n1117 104.757
R1428 VDD.n1609 VDD.n1117 104.757
R1429 VDD.n1609 VDD.n1115 104.757
R1430 VDD.n1613 VDD.n1115 104.757
R1431 VDD.n1613 VDD.n1113 104.757
R1432 VDD.n1617 VDD.n1113 104.757
R1433 VDD.n1617 VDD.n1111 104.757
R1434 VDD.n1621 VDD.n1111 104.757
R1435 VDD.n1621 VDD.n1109 104.757
R1436 VDD.n1625 VDD.n1109 104.757
R1437 VDD.n1625 VDD.n1107 104.757
R1438 VDD.n1629 VDD.n1107 104.757
R1439 VDD.n1629 VDD.n1105 104.757
R1440 VDD.n1633 VDD.n1105 104.757
R1441 VDD.n1633 VDD.n1103 104.757
R1442 VDD.n1639 VDD.n1103 104.757
R1443 VDD.n1639 VDD.n1101 104.757
R1444 VDD.n1260 VDD.n1259 104.757
R1445 VDD.n1257 VDD.n1219 104.757
R1446 VDD.n1253 VDD.n1219 104.757
R1447 VDD.n1253 VDD.n1221 104.757
R1448 VDD.n1249 VDD.n1221 104.757
R1449 VDD.n1249 VDD.n1224 104.757
R1450 VDD.n1245 VDD.n1224 104.757
R1451 VDD.n1245 VDD.n1226 104.757
R1452 VDD.n1241 VDD.n1226 104.757
R1453 VDD.n1241 VDD.n1228 104.757
R1454 VDD.n1237 VDD.n1228 104.757
R1455 VDD.n1237 VDD.n1230 104.757
R1456 VDD.n1233 VDD.n1230 104.757
R1457 VDD.n1233 VDD.n957 104.757
R1458 VDD.n1678 VDD.n957 104.757
R1459 VDD.n1679 VDD.n1678 104.757
R1460 VDD.n1065 VDD.n980 104.757
R1461 VDD.n1063 VDD.n981 104.757
R1462 VDD.n1055 VDD.n1054 104.757
R1463 VDD.n1050 VDD.n1049 104.757
R1464 VDD.n1018 VDD.n987 104.757
R1465 VDD.n1009 VDD.n993 104.757
R1466 VDD.n1007 VDD.n994 104.757
R1467 VDD.n998 VDD.n997 104.757
R1468 VDD.n1674 VDD.n962 104.757
R1469 VDD.n1674 VDD.n963 104.757
R1470 VDD.n1670 VDD.n963 104.757
R1471 VDD.n1670 VDD.n1088 104.757
R1472 VDD.n1666 VDD.n1088 104.757
R1473 VDD.n1666 VDD.n1090 104.757
R1474 VDD.n1662 VDD.n1090 104.757
R1475 VDD.n1662 VDD.n1092 104.757
R1476 VDD.n1658 VDD.n1092 104.757
R1477 VDD.n1658 VDD.n1094 104.757
R1478 VDD.n1654 VDD.n1094 104.757
R1479 VDD.n1654 VDD.n1096 104.757
R1480 VDD.n1650 VDD.n1096 104.757
R1481 VDD.n1650 VDD.n1098 104.757
R1482 VDD.n1646 VDD.n1098 104.757
R1483 VDD.n1644 VDD.n1643 104.757
R1484 VDD.n461 VDD.n332 104.757
R1485 VDD.n461 VDD.n334 104.757
R1486 VDD.n457 VDD.n334 104.757
R1487 VDD.n457 VDD.n336 104.757
R1488 VDD.n453 VDD.n336 104.757
R1489 VDD.n453 VDD.n338 104.757
R1490 VDD.n449 VDD.n338 104.757
R1491 VDD.n449 VDD.n340 104.757
R1492 VDD.n445 VDD.n340 104.757
R1493 VDD.n445 VDD.n342 104.757
R1494 VDD.n441 VDD.n342 104.757
R1495 VDD.n441 VDD.n344 104.757
R1496 VDD.n437 VDD.n344 104.757
R1497 VDD.n437 VDD.n346 104.757
R1498 VDD.n433 VDD.n346 104.757
R1499 VDD.n433 VDD.n348 104.757
R1500 VDD.n429 VDD.n348 104.757
R1501 VDD.n429 VDD.n350 104.757
R1502 VDD.n425 VDD.n350 104.757
R1503 VDD.n425 VDD.n352 104.757
R1504 VDD.n421 VDD.n352 104.757
R1505 VDD.n421 VDD.n354 104.757
R1506 VDD.n417 VDD.n354 104.757
R1507 VDD.n417 VDD.n356 104.757
R1508 VDD.n413 VDD.n356 104.757
R1509 VDD.n413 VDD.n358 104.757
R1510 VDD.n409 VDD.n358 104.757
R1511 VDD.n477 VDD.n328 104.757
R1512 VDD.n477 VDD.n326 104.757
R1513 VDD.n481 VDD.n326 104.757
R1514 VDD.n481 VDD.n324 104.757
R1515 VDD.n485 VDD.n324 104.757
R1516 VDD.n485 VDD.n322 104.757
R1517 VDD.n489 VDD.n322 104.757
R1518 VDD.n489 VDD.n320 104.757
R1519 VDD.n493 VDD.n320 104.757
R1520 VDD.n493 VDD.n318 104.757
R1521 VDD.n497 VDD.n318 104.757
R1522 VDD.n497 VDD.n316 104.757
R1523 VDD.n502 VDD.n316 104.757
R1524 VDD.n502 VDD.n314 104.757
R1525 VDD.n689 VDD.n314 104.757
R1526 VDD.n668 VDD.n306 104.757
R1527 VDD.n585 VDD.n306 104.757
R1528 VDD.n589 VDD.n588 104.757
R1529 VDD.n693 VDD.n292 104.757
R1530 VDD.n697 VDD.n292 104.757
R1531 VDD.n697 VDD.n290 104.757
R1532 VDD.n701 VDD.n290 104.757
R1533 VDD.n701 VDD.n288 104.757
R1534 VDD.n705 VDD.n288 104.757
R1535 VDD.n705 VDD.n286 104.757
R1536 VDD.n709 VDD.n286 104.757
R1537 VDD.n709 VDD.n284 104.757
R1538 VDD.n713 VDD.n284 104.757
R1539 VDD.n713 VDD.n282 104.757
R1540 VDD.n717 VDD.n282 104.757
R1541 VDD.n717 VDD.n279 104.757
R1542 VDD.n722 VDD.n279 104.757
R1543 VDD.n722 VDD.n280 104.757
R1544 VDD.n726 VDD.n276 104.757
R1545 VDD.n730 VDD.n274 104.757
R1546 VDD.n730 VDD.n272 104.757
R1547 VDD.n734 VDD.n272 104.757
R1548 VDD.n734 VDD.n270 104.757
R1549 VDD.n738 VDD.n270 104.757
R1550 VDD.n738 VDD.n268 104.757
R1551 VDD.n742 VDD.n268 104.757
R1552 VDD.n742 VDD.n266 104.757
R1553 VDD.n746 VDD.n266 104.757
R1554 VDD.n746 VDD.n264 104.757
R1555 VDD.n750 VDD.n264 104.757
R1556 VDD.n750 VDD.n262 104.757
R1557 VDD.n754 VDD.n262 104.757
R1558 VDD.n754 VDD.n260 104.757
R1559 VDD.n758 VDD.n260 104.757
R1560 VDD.n758 VDD.n258 104.757
R1561 VDD.n762 VDD.n258 104.757
R1562 VDD.n762 VDD.n256 104.757
R1563 VDD.n766 VDD.n256 104.757
R1564 VDD.n766 VDD.n254 104.757
R1565 VDD.n770 VDD.n254 104.757
R1566 VDD.n770 VDD.n252 104.757
R1567 VDD.n774 VDD.n252 104.757
R1568 VDD.n774 VDD.n250 104.757
R1569 VDD.n778 VDD.n250 104.757
R1570 VDD.n778 VDD.n248 104.757
R1571 VDD.n784 VDD.n248 104.757
R1572 VDD.n784 VDD.n246 104.757
R1573 VDD.n405 VDD.n404 104.757
R1574 VDD.n402 VDD.n364 104.757
R1575 VDD.n398 VDD.n364 104.757
R1576 VDD.n398 VDD.n366 104.757
R1577 VDD.n394 VDD.n366 104.757
R1578 VDD.n394 VDD.n369 104.757
R1579 VDD.n390 VDD.n369 104.757
R1580 VDD.n390 VDD.n371 104.757
R1581 VDD.n386 VDD.n371 104.757
R1582 VDD.n386 VDD.n373 104.757
R1583 VDD.n382 VDD.n373 104.757
R1584 VDD.n382 VDD.n375 104.757
R1585 VDD.n378 VDD.n375 104.757
R1586 VDD.n378 VDD.n102 104.757
R1587 VDD.n823 VDD.n102 104.757
R1588 VDD.n824 VDD.n823 104.757
R1589 VDD.n210 VDD.n125 104.757
R1590 VDD.n208 VDD.n126 104.757
R1591 VDD.n200 VDD.n199 104.757
R1592 VDD.n195 VDD.n194 104.757
R1593 VDD.n163 VDD.n132 104.757
R1594 VDD.n154 VDD.n138 104.757
R1595 VDD.n152 VDD.n139 104.757
R1596 VDD.n143 VDD.n142 104.757
R1597 VDD.n819 VDD.n107 104.757
R1598 VDD.n819 VDD.n108 104.757
R1599 VDD.n815 VDD.n108 104.757
R1600 VDD.n815 VDD.n233 104.757
R1601 VDD.n811 VDD.n233 104.757
R1602 VDD.n811 VDD.n235 104.757
R1603 VDD.n807 VDD.n235 104.757
R1604 VDD.n807 VDD.n237 104.757
R1605 VDD.n803 VDD.n237 104.757
R1606 VDD.n803 VDD.n239 104.757
R1607 VDD.n799 VDD.n239 104.757
R1608 VDD.n799 VDD.n241 104.757
R1609 VDD.n795 VDD.n241 104.757
R1610 VDD.n795 VDD.n243 104.757
R1611 VDD.n791 VDD.n243 104.757
R1612 VDD.n789 VDD.n788 104.757
R1613 VDD.n3109 VDD.n3066 96.8641
R1614 VDD.n2118 VDD.n2117 96.8641
R1615 VDD.n1264 VDD.n1263 96.8641
R1616 VDD.n409 VDD.n408 96.8641
R1617 VDD.t55 VDD.n32 96.8274
R1618 VDD.n880 VDD.t25 96.8274
R1619 VDD.t63 VDD.n1741 96.8274
R1620 VDD.n2076 VDD.n2068 96.5084
R1621 VDD.n2185 VDD.n2184 96.5084
R1622 VDD.n1222 VDD.n1214 96.5084
R1623 VDD.n1331 VDD.n1330 96.5084
R1624 VDD.n367 VDD.n359 96.5084
R1625 VDD.n476 VDD.n475 96.5084
R1626 VDD.n8854 VDD.n8853 92.5005
R1627 VDD.n8852 VDD.n8851 92.5005
R1628 VDD.n6495 VDD.n6494 92.5005
R1629 VDD.n3599 VDD.n3598 92.5005
R1630 VDD.n6822 VDD.n6821 92.5005
R1631 VDD.n6818 VDD.n6817 92.5005
R1632 VDD.n6814 VDD.n6813 92.5005
R1633 VDD.n6810 VDD.n6809 92.5005
R1634 VDD.n6806 VDD.n6805 92.5005
R1635 VDD.n6802 VDD.n6801 92.5005
R1636 VDD.n6801 VDD.n6800 92.5005
R1637 VDD.n6797 VDD.n6796 92.5005
R1638 VDD.n6796 VDD.n6795 92.5005
R1639 VDD.n6789 VDD.n6788 92.5005
R1640 VDD.n6788 VDD.n6787 92.5005
R1641 VDD.n6792 VDD.n6791 92.5005
R1642 VDD.n6791 VDD.n6790 92.5005
R1643 VDD.n6784 VDD.n6783 92.5005
R1644 VDD.n6783 VDD.n6782 92.5005
R1645 VDD.n6779 VDD.n6778 92.5005
R1646 VDD.n6778 VDD.n6777 92.5005
R1647 VDD.n6774 VDD.n6773 92.5005
R1648 VDD.n6773 VDD.n6772 92.5005
R1649 VDD.n6769 VDD.n6768 92.5005
R1650 VDD.n6768 VDD.n6767 92.5005
R1651 VDD.n6764 VDD.n6763 92.5005
R1652 VDD.n6763 VDD.n6762 92.5005
R1653 VDD.n6759 VDD.n6758 92.5005
R1654 VDD.n6758 VDD.n6757 92.5005
R1655 VDD.n6754 VDD.n6753 92.5005
R1656 VDD.n6753 VDD.n6752 92.5005
R1657 VDD.n6749 VDD.n6748 92.5005
R1658 VDD.n6748 VDD.n6747 92.5005
R1659 VDD.n6744 VDD.n6743 92.5005
R1660 VDD.n6743 VDD.n6742 92.5005
R1661 VDD.n6739 VDD.n6738 92.5005
R1662 VDD.n6738 VDD.n6737 92.5005
R1663 VDD.n6734 VDD.n6733 92.5005
R1664 VDD.n6733 VDD.n6732 92.5005
R1665 VDD.n6729 VDD.n6728 92.5005
R1666 VDD.n6728 VDD.n6727 92.5005
R1667 VDD.n6724 VDD.n6723 92.5005
R1668 VDD.n6723 VDD.n6722 92.5005
R1669 VDD.n6719 VDD.n6718 92.5005
R1670 VDD.n6718 VDD.n6717 92.5005
R1671 VDD.n6714 VDD.n6713 92.5005
R1672 VDD.n6713 VDD.n6712 92.5005
R1673 VDD.n6709 VDD.n6708 92.5005
R1674 VDD.n6708 VDD.n6707 92.5005
R1675 VDD.n6701 VDD.n6700 92.5005
R1676 VDD.n6700 VDD.n6699 92.5005
R1677 VDD.n6704 VDD.n6703 92.5005
R1678 VDD.n6703 VDD.n6702 92.5005
R1679 VDD.n6696 VDD.n6695 92.5005
R1680 VDD.n6692 VDD.n6691 92.5005
R1681 VDD.n6688 VDD.n6687 92.5005
R1682 VDD.n6684 VDD.n6683 92.5005
R1683 VDD.n6680 VDD.n6679 92.5005
R1684 VDD.n6676 VDD.n6675 92.5005
R1685 VDD.n6672 VDD.n6671 92.5005
R1686 VDD.n6651 VDD.n6650 92.5005
R1687 VDD.n6647 VDD.n6646 92.5005
R1688 VDD.n6643 VDD.n6642 92.5005
R1689 VDD.n6639 VDD.n6638 92.5005
R1690 VDD.n6635 VDD.n6634 92.5005
R1691 VDD.n6631 VDD.n6630 92.5005
R1692 VDD.n6627 VDD.n6626 92.5005
R1693 VDD.n6626 VDD.n6625 92.5005
R1694 VDD.n6622 VDD.n6621 92.5005
R1695 VDD.n6621 VDD.n6620 92.5005
R1696 VDD.n6617 VDD.n6616 92.5005
R1697 VDD.n6616 VDD.n6615 92.5005
R1698 VDD.n6609 VDD.n6608 92.5005
R1699 VDD.n6608 VDD.n6607 92.5005
R1700 VDD.n6612 VDD.n6611 92.5005
R1701 VDD.n6611 VDD.n6610 92.5005
R1702 VDD.n6604 VDD.n6603 92.5005
R1703 VDD.n6603 VDD.n6602 92.5005
R1704 VDD.n6599 VDD.n6598 92.5005
R1705 VDD.n6598 VDD.n6597 92.5005
R1706 VDD.n6594 VDD.n6593 92.5005
R1707 VDD.n6593 VDD.n6592 92.5005
R1708 VDD.n6589 VDD.n6588 92.5005
R1709 VDD.n6588 VDD.n6587 92.5005
R1710 VDD.n6584 VDD.n6583 92.5005
R1711 VDD.n6583 VDD.n6582 92.5005
R1712 VDD.n6579 VDD.n6578 92.5005
R1713 VDD.n6578 VDD.n6577 92.5005
R1714 VDD.n6574 VDD.n6573 92.5005
R1715 VDD.n6573 VDD.n6572 92.5005
R1716 VDD.n6569 VDD.n6568 92.5005
R1717 VDD.n6568 VDD.n6567 92.5005
R1718 VDD.n6564 VDD.n6563 92.5005
R1719 VDD.n6563 VDD.n6562 92.5005
R1720 VDD.n6559 VDD.n6558 92.5005
R1721 VDD.n6558 VDD.n6557 92.5005
R1722 VDD.n6554 VDD.n6553 92.5005
R1723 VDD.n6553 VDD.n6552 92.5005
R1724 VDD.n6549 VDD.n6548 92.5005
R1725 VDD.n6548 VDD.n6547 92.5005
R1726 VDD.n6544 VDD.n6543 92.5005
R1727 VDD.n6543 VDD.n6542 92.5005
R1728 VDD.n6539 VDD.n6538 92.5005
R1729 VDD.n6538 VDD.n6537 92.5005
R1730 VDD.n6534 VDD.n6533 92.5005
R1731 VDD.n6533 VDD.n6532 92.5005
R1732 VDD.n6529 VDD.n6528 92.5005
R1733 VDD.n6528 VDD.n6527 92.5005
R1734 VDD.n6522 VDD.n6521 92.5005
R1735 VDD.n6524 VDD.n6523 92.5005
R1736 VDD.n6518 VDD.n6517 92.5005
R1737 VDD.n6514 VDD.n6513 92.5005
R1738 VDD.n6510 VDD.n6509 92.5005
R1739 VDD.n8847 VDD.n8846 92.5005
R1740 VDD.n8850 VDD.n8849 92.5005
R1741 VDD.n8857 VDD.n8856 92.5005
R1742 VDD.n7607 VDD.n7606 92.5005
R1743 VDD.n7609 VDD.n7608 92.5005
R1744 VDD.n7611 VDD.n7610 92.5005
R1745 VDD.n7613 VDD.n7612 92.5005
R1746 VDD.n7615 VDD.n7614 92.5005
R1747 VDD.n7618 VDD.n7617 92.5005
R1748 VDD.n8568 VDD.n8556 92.5005
R1749 VDD.n8064 VDD.n8063 92.5005
R1750 VDD.n8070 VDD.n8069 92.5005
R1751 VDD.n8077 VDD.n8076 92.5005
R1752 VDD.n8084 VDD.n8083 92.5005
R1753 VDD.n8086 VDD.n8085 92.5005
R1754 VDD.n8093 VDD.n8092 92.5005
R1755 VDD.n8100 VDD.n8099 92.5005
R1756 VDD.n8107 VDD.n8106 92.5005
R1757 VDD.n8114 VDD.n8113 92.5005
R1758 VDD.n8121 VDD.n8120 92.5005
R1759 VDD.n8128 VDD.n8127 92.5005
R1760 VDD.n8140 VDD.n8139 92.5005
R1761 VDD.n8056 VDD.n8055 92.5005
R1762 VDD.n8061 VDD.n8060 92.5005
R1763 VDD.n8068 VDD.n8067 92.5005
R1764 VDD.n8072 VDD.n8071 92.5005
R1765 VDD.n8080 VDD.n8079 92.5005
R1766 VDD.n8088 VDD.n8087 92.5005
R1767 VDD.n8096 VDD.n8095 92.5005
R1768 VDD.n8102 VDD.n8101 92.5005
R1769 VDD.n8110 VDD.n8109 92.5005
R1770 VDD.n8116 VDD.n8115 92.5005
R1771 VDD.n8124 VDD.n8123 92.5005
R1772 VDD.n8131 VDD.n8130 92.5005
R1773 VDD.n8135 VDD.n8134 92.5005
R1774 VDD.n8144 VDD.n8143 92.5005
R1775 VDD.n8053 VDD.n8052 92.5005
R1776 VDD.n8036 VDD.n8035 92.5005
R1777 VDD.n8035 VDD.n8034 92.5005
R1778 VDD.n8028 VDD.n8027 92.5005
R1779 VDD.n8027 VDD.n8026 92.5005
R1780 VDD.n8020 VDD.n8019 92.5005
R1781 VDD.n8019 VDD.n8018 92.5005
R1782 VDD.n8012 VDD.n8011 92.5005
R1783 VDD.n8011 VDD.n8010 92.5005
R1784 VDD.n8004 VDD.n8003 92.5005
R1785 VDD.n8003 VDD.n8002 92.5005
R1786 VDD.n7996 VDD.n7995 92.5005
R1787 VDD.n7995 VDD.n7994 92.5005
R1788 VDD.n7988 VDD.n7987 92.5005
R1789 VDD.n7987 VDD.n7986 92.5005
R1790 VDD.n7980 VDD.n7979 92.5005
R1791 VDD.n7979 VDD.n7978 92.5005
R1792 VDD.n7969 VDD.n7968 92.5005
R1793 VDD.n7968 VDD.n7967 92.5005
R1794 VDD.n7975 VDD.n7974 92.5005
R1795 VDD.n7974 VDD.n7973 92.5005
R1796 VDD.n7964 VDD.n7963 92.5005
R1797 VDD.n7963 VDD.n7962 92.5005
R1798 VDD.n7956 VDD.n7955 92.5005
R1799 VDD.n7955 VDD.n7954 92.5005
R1800 VDD.n7945 VDD.n7944 92.5005
R1801 VDD.n7944 VDD.n7943 92.5005
R1802 VDD.n7937 VDD.n7936 92.5005
R1803 VDD.n7936 VDD.n7935 92.5005
R1804 VDD.n7929 VDD.n7928 92.5005
R1805 VDD.n7928 VDD.n7927 92.5005
R1806 VDD.n7921 VDD.n7920 92.5005
R1807 VDD.n7920 VDD.n7919 92.5005
R1808 VDD.n7913 VDD.n7912 92.5005
R1809 VDD.n7912 VDD.n7911 92.5005
R1810 VDD.n7905 VDD.n7904 92.5005
R1811 VDD.n7904 VDD.n7903 92.5005
R1812 VDD.n7894 VDD.n7893 92.5005
R1813 VDD.n7893 VDD.n7892 92.5005
R1814 VDD.n7886 VDD.n7885 92.5005
R1815 VDD.n7885 VDD.n7884 92.5005
R1816 VDD.n7878 VDD.n7877 92.5005
R1817 VDD.n7877 VDD.n7876 92.5005
R1818 VDD.n7870 VDD.n7869 92.5005
R1819 VDD.n7869 VDD.n7868 92.5005
R1820 VDD.n7862 VDD.n7861 92.5005
R1821 VDD.n7861 VDD.n7860 92.5005
R1822 VDD.n7854 VDD.n7853 92.5005
R1823 VDD.n7853 VDD.n7852 92.5005
R1824 VDD.n7846 VDD.n7845 92.5005
R1825 VDD.n7845 VDD.n7844 92.5005
R1826 VDD.n7838 VDD.n7837 92.5005
R1827 VDD.n7837 VDD.n7836 92.5005
R1828 VDD.n7828 VDD.n7827 92.5005
R1829 VDD.n7827 VDD.n7826 92.5005
R1830 VDD.n7833 VDD.n7832 92.5005
R1831 VDD.n7823 VDD.n7822 92.5005
R1832 VDD.n7817 VDD.n7816 92.5005
R1833 VDD.n7809 VDD.n7808 92.5005
R1834 VDD.n7803 VDD.n7802 92.5005
R1835 VDD.n7797 VDD.n7796 92.5005
R1836 VDD.n7796 VDD.n7795 92.5005
R1837 VDD.n7789 VDD.n7788 92.5005
R1838 VDD.n7788 VDD.n7787 92.5005
R1839 VDD.n7781 VDD.n7780 92.5005
R1840 VDD.n7780 VDD.n7779 92.5005
R1841 VDD.n7773 VDD.n7772 92.5005
R1842 VDD.n7772 VDD.n7771 92.5005
R1843 VDD.n7762 VDD.n7761 92.5005
R1844 VDD.n7761 VDD.n7760 92.5005
R1845 VDD.n7754 VDD.n7753 92.5005
R1846 VDD.n7753 VDD.n7752 92.5005
R1847 VDD.n7746 VDD.n7745 92.5005
R1848 VDD.n7745 VDD.n7744 92.5005
R1849 VDD.n7738 VDD.n7737 92.5005
R1850 VDD.n7737 VDD.n7736 92.5005
R1851 VDD.n7730 VDD.n7729 92.5005
R1852 VDD.n7729 VDD.n7728 92.5005
R1853 VDD.n7722 VDD.n7721 92.5005
R1854 VDD.n7721 VDD.n7720 92.5005
R1855 VDD.n7714 VDD.n7713 92.5005
R1856 VDD.n7713 VDD.n7712 92.5005
R1857 VDD.n7706 VDD.n7705 92.5005
R1858 VDD.n7705 VDD.n7704 92.5005
R1859 VDD.n7695 VDD.n7694 92.5005
R1860 VDD.n7694 VDD.n7693 92.5005
R1861 VDD.n7701 VDD.n7700 92.5005
R1862 VDD.n7700 VDD.n7699 92.5005
R1863 VDD.n7690 VDD.n7689 92.5005
R1864 VDD.n7689 VDD.n7688 92.5005
R1865 VDD.n7682 VDD.n7681 92.5005
R1866 VDD.n7681 VDD.n7680 92.5005
R1867 VDD.n7671 VDD.n7670 92.5005
R1868 VDD.n7670 VDD.n7669 92.5005
R1869 VDD.n7663 VDD.n7662 92.5005
R1870 VDD.n7662 VDD.n7661 92.5005
R1871 VDD.n7655 VDD.n7654 92.5005
R1872 VDD.n7654 VDD.n7653 92.5005
R1873 VDD.n7647 VDD.n7646 92.5005
R1874 VDD.n7646 VDD.n7645 92.5005
R1875 VDD.n7634 VDD.n7633 92.5005
R1876 VDD.n7633 VDD.n7632 92.5005
R1877 VDD.n7639 VDD.n7638 92.5005
R1878 VDD.n7638 VDD.n7637 92.5005
R1879 VDD.n7644 VDD.n7643 92.5005
R1880 VDD.n7643 VDD.n7642 92.5005
R1881 VDD.n7652 VDD.n7651 92.5005
R1882 VDD.n7651 VDD.n7650 92.5005
R1883 VDD.n7660 VDD.n7659 92.5005
R1884 VDD.n7659 VDD.n7658 92.5005
R1885 VDD.n7668 VDD.n7667 92.5005
R1886 VDD.n7667 VDD.n7666 92.5005
R1887 VDD.n7679 VDD.n7678 92.5005
R1888 VDD.n7678 VDD.n7677 92.5005
R1889 VDD.n7676 VDD.n7675 92.5005
R1890 VDD.n7675 VDD.n7674 92.5005
R1891 VDD.n7687 VDD.n7686 92.5005
R1892 VDD.n7686 VDD.n7685 92.5005
R1893 VDD.n7698 VDD.n7697 92.5005
R1894 VDD.n7697 VDD.n7696 92.5005
R1895 VDD.n7709 VDD.n7708 92.5005
R1896 VDD.n7708 VDD.n7707 92.5005
R1897 VDD.n7717 VDD.n7716 92.5005
R1898 VDD.n7716 VDD.n7715 92.5005
R1899 VDD.n7725 VDD.n7724 92.5005
R1900 VDD.n7724 VDD.n7723 92.5005
R1901 VDD.n7733 VDD.n7732 92.5005
R1902 VDD.n7732 VDD.n7731 92.5005
R1903 VDD.n7741 VDD.n7740 92.5005
R1904 VDD.n7740 VDD.n7739 92.5005
R1905 VDD.n7749 VDD.n7748 92.5005
R1906 VDD.n7748 VDD.n7747 92.5005
R1907 VDD.n7757 VDD.n7756 92.5005
R1908 VDD.n7756 VDD.n7755 92.5005
R1909 VDD.n7765 VDD.n7764 92.5005
R1910 VDD.n7764 VDD.n7763 92.5005
R1911 VDD.n7770 VDD.n7769 92.5005
R1912 VDD.n7769 VDD.n7768 92.5005
R1913 VDD.n7778 VDD.n7777 92.5005
R1914 VDD.n7777 VDD.n7776 92.5005
R1915 VDD.n7786 VDD.n7785 92.5005
R1916 VDD.n7785 VDD.n7784 92.5005
R1917 VDD.n7794 VDD.n7793 92.5005
R1918 VDD.n7793 VDD.n7792 92.5005
R1919 VDD.n7801 VDD.n7800 92.5005
R1920 VDD.n7807 VDD.n7806 92.5005
R1921 VDD.n7815 VDD.n7814 92.5005
R1922 VDD.n7813 VDD.n7812 92.5005
R1923 VDD.n7821 VDD.n7820 92.5005
R1924 VDD.n7831 VDD.n7830 92.5005
R1925 VDD.n7830 VDD.n7829 92.5005
R1926 VDD.n7841 VDD.n7840 92.5005
R1927 VDD.n7840 VDD.n7839 92.5005
R1928 VDD.n7849 VDD.n7848 92.5005
R1929 VDD.n7848 VDD.n7847 92.5005
R1930 VDD.n7857 VDD.n7856 92.5005
R1931 VDD.n7856 VDD.n7855 92.5005
R1932 VDD.n7865 VDD.n7864 92.5005
R1933 VDD.n7864 VDD.n7863 92.5005
R1934 VDD.n7873 VDD.n7872 92.5005
R1935 VDD.n7872 VDD.n7871 92.5005
R1936 VDD.n7881 VDD.n7880 92.5005
R1937 VDD.n7880 VDD.n7879 92.5005
R1938 VDD.n7889 VDD.n7888 92.5005
R1939 VDD.n7888 VDD.n7887 92.5005
R1940 VDD.n7897 VDD.n7896 92.5005
R1941 VDD.n7896 VDD.n7895 92.5005
R1942 VDD.n7902 VDD.n7901 92.5005
R1943 VDD.n7901 VDD.n7900 92.5005
R1944 VDD.n7910 VDD.n7909 92.5005
R1945 VDD.n7909 VDD.n7908 92.5005
R1946 VDD.n7918 VDD.n7917 92.5005
R1947 VDD.n7917 VDD.n7916 92.5005
R1948 VDD.n7926 VDD.n7925 92.5005
R1949 VDD.n7925 VDD.n7924 92.5005
R1950 VDD.n7934 VDD.n7933 92.5005
R1951 VDD.n7933 VDD.n7932 92.5005
R1952 VDD.n7942 VDD.n7941 92.5005
R1953 VDD.n7941 VDD.n7940 92.5005
R1954 VDD.n7953 VDD.n7952 92.5005
R1955 VDD.n7952 VDD.n7951 92.5005
R1956 VDD.n7950 VDD.n7949 92.5005
R1957 VDD.n7949 VDD.n7948 92.5005
R1958 VDD.n7961 VDD.n7960 92.5005
R1959 VDD.n7960 VDD.n7959 92.5005
R1960 VDD.n7972 VDD.n7971 92.5005
R1961 VDD.n7971 VDD.n7970 92.5005
R1962 VDD.n7983 VDD.n7982 92.5005
R1963 VDD.n7982 VDD.n7981 92.5005
R1964 VDD.n7991 VDD.n7990 92.5005
R1965 VDD.n7990 VDD.n7989 92.5005
R1966 VDD.n7999 VDD.n7998 92.5005
R1967 VDD.n7998 VDD.n7997 92.5005
R1968 VDD.n8007 VDD.n8006 92.5005
R1969 VDD.n8006 VDD.n8005 92.5005
R1970 VDD.n8015 VDD.n8014 92.5005
R1971 VDD.n8014 VDD.n8013 92.5005
R1972 VDD.n8023 VDD.n8022 92.5005
R1973 VDD.n8022 VDD.n8021 92.5005
R1974 VDD.n8031 VDD.n8030 92.5005
R1975 VDD.n8030 VDD.n8029 92.5005
R1976 VDD.n8042 VDD.n8041 92.5005
R1977 VDD.n8041 VDD.n8040 92.5005
R1978 VDD.n8039 VDD.n8038 92.5005
R1979 VDD.n8038 VDD.n8037 92.5005
R1980 VDD.n8051 VDD.n8050 92.5005
R1981 VDD.n7579 VDD.n7578 92.5005
R1982 VDD.n7578 VDD.n7577 92.5005
R1983 VDD.n7567 VDD.n7566 92.5005
R1984 VDD.n7566 VDD.n7565 92.5005
R1985 VDD.n7584 VDD.n7583 92.5005
R1986 VDD.n7583 VDD.n7582 92.5005
R1987 VDD.n7589 VDD.n7588 92.5005
R1988 VDD.n7588 VDD.n7587 92.5005
R1989 VDD.n7594 VDD.n7593 92.5005
R1990 VDD.n7593 VDD.n7592 92.5005
R1991 VDD.n7599 VDD.n7598 92.5005
R1992 VDD.n7598 VDD.n7597 92.5005
R1993 VDD.n7500 VDD.n7499 92.5005
R1994 VDD.n7504 VDD.n7503 92.5005
R1995 VDD.n7509 VDD.n7508 92.5005
R1996 VDD.n7514 VDD.n7513 92.5005
R1997 VDD.n7519 VDD.n7518 92.5005
R1998 VDD.n7524 VDD.n7523 92.5005
R1999 VDD.n7529 VDD.n7528 92.5005
R2000 VDD.n7535 VDD.n7534 92.5005
R2001 VDD.n7540 VDD.n7539 92.5005
R2002 VDD.n7545 VDD.n7544 92.5005
R2003 VDD.n7550 VDD.n7549 92.5005
R2004 VDD.n7555 VDD.n7554 92.5005
R2005 VDD.n7562 VDD.n7561 92.5005
R2006 VDD.n7559 VDD.n7558 92.5005
R2007 VDD.n7575 VDD.n7574 92.5005
R2008 VDD.n7569 VDD.n7568 92.5005
R2009 VDD.n7571 VDD.n7570 92.5005
R2010 VDD.n6501 VDD.n6500 92.5005
R2011 VDD.n6491 VDD.n6490 92.5005
R2012 VDD.n6486 VDD.n6485 92.5005
R2013 VDD.n6482 VDD.n6481 92.5005
R2014 VDD.n6477 VDD.n6476 92.5005
R2015 VDD.n6473 VDD.n6472 92.5005
R2016 VDD.n6468 VDD.n6467 92.5005
R2017 VDD.n6461 VDD.n6460 92.5005
R2018 VDD.n6464 VDD.n6463 92.5005
R2019 VDD.n6457 VDD.n6456 92.5005
R2020 VDD.n6453 VDD.n6452 92.5005
R2021 VDD.n6448 VDD.n6447 92.5005
R2022 VDD.n6444 VDD.n6443 92.5005
R2023 VDD.n6439 VDD.n6438 92.5005
R2024 VDD.n6435 VDD.n6434 92.5005
R2025 VDD.n6430 VDD.n6429 92.5005
R2026 VDD.n6426 VDD.n6425 92.5005
R2027 VDD.n6421 VDD.n6420 92.5005
R2028 VDD.n6416 VDD.n6415 92.5005
R2029 VDD.n6412 VDD.n6411 92.5005
R2030 VDD.n6407 VDD.n6406 92.5005
R2031 VDD.n6403 VDD.n6402 92.5005
R2032 VDD.n6398 VDD.n6397 92.5005
R2033 VDD.n6394 VDD.n6393 92.5005
R2034 VDD.n6389 VDD.n6388 92.5005
R2035 VDD.n6382 VDD.n6381 92.5005
R2036 VDD.n6385 VDD.n6384 92.5005
R2037 VDD.n6378 VDD.n6377 92.5005
R2038 VDD.n6374 VDD.n6373 92.5005
R2039 VDD.n6369 VDD.n6368 92.5005
R2040 VDD.n6368 VDD.n6367 92.5005
R2041 VDD.n6364 VDD.n6363 92.5005
R2042 VDD.n6363 VDD.n6362 92.5005
R2043 VDD.n6359 VDD.n6358 92.5005
R2044 VDD.n6358 VDD.n6357 92.5005
R2045 VDD.n6354 VDD.n6353 92.5005
R2046 VDD.n6353 VDD.n6352 92.5005
R2047 VDD.n6349 VDD.n6348 92.5005
R2048 VDD.n6348 VDD.n6347 92.5005
R2049 VDD.n6344 VDD.n6343 92.5005
R2050 VDD.n6343 VDD.n6342 92.5005
R2051 VDD.n6339 VDD.n6338 92.5005
R2052 VDD.n6338 VDD.n6337 92.5005
R2053 VDD.n6334 VDD.n6333 92.5005
R2054 VDD.n6333 VDD.n6332 92.5005
R2055 VDD.n6329 VDD.n6328 92.5005
R2056 VDD.n6328 VDD.n6327 92.5005
R2057 VDD.n6324 VDD.n6323 92.5005
R2058 VDD.n6323 VDD.n6322 92.5005
R2059 VDD.n6319 VDD.n6318 92.5005
R2060 VDD.n6318 VDD.n6317 92.5005
R2061 VDD.n6314 VDD.n6313 92.5005
R2062 VDD.n6313 VDD.n6312 92.5005
R2063 VDD.n6309 VDD.n6308 92.5005
R2064 VDD.n6308 VDD.n6307 92.5005
R2065 VDD.n6304 VDD.n6303 92.5005
R2066 VDD.n6303 VDD.n6302 92.5005
R2067 VDD.n6296 VDD.n6295 92.5005
R2068 VDD.n6295 VDD.n6294 92.5005
R2069 VDD.n6299 VDD.n6298 92.5005
R2070 VDD.n6298 VDD.n6297 92.5005
R2071 VDD.n6291 VDD.n6290 92.5005
R2072 VDD.n6290 VDD.n6289 92.5005
R2073 VDD.n6286 VDD.n6285 92.5005
R2074 VDD.n6285 VDD.n6284 92.5005
R2075 VDD.n6281 VDD.n6280 92.5005
R2076 VDD.n6280 VDD.n6279 92.5005
R2077 VDD.n6276 VDD.n6275 92.5005
R2078 VDD.n6275 VDD.n6274 92.5005
R2079 VDD.n6271 VDD.n6270 92.5005
R2080 VDD.n6270 VDD.n6269 92.5005
R2081 VDD.n6266 VDD.n6265 92.5005
R2082 VDD.n6265 VDD.n6264 92.5005
R2083 VDD.n6261 VDD.n6260 92.5005
R2084 VDD.n6260 VDD.n6259 92.5005
R2085 VDD.n6256 VDD.n6255 92.5005
R2086 VDD.n6255 VDD.n6254 92.5005
R2087 VDD.n6251 VDD.n6250 92.5005
R2088 VDD.n6250 VDD.n6249 92.5005
R2089 VDD.n6246 VDD.n6245 92.5005
R2090 VDD.n6245 VDD.n6244 92.5005
R2091 VDD.n6241 VDD.n6240 92.5005
R2092 VDD.n6240 VDD.n6239 92.5005
R2093 VDD.n6236 VDD.n6235 92.5005
R2094 VDD.n6235 VDD.n6234 92.5005
R2095 VDD.n6231 VDD.n6230 92.5005
R2096 VDD.n6230 VDD.n6229 92.5005
R2097 VDD.n6226 VDD.n6225 92.5005
R2098 VDD.n6225 VDD.n6224 92.5005
R2099 VDD.n6063 VDD.n6062 92.5005
R2100 VDD.n6221 VDD.n6220 92.5005
R2101 VDD.n6217 VDD.n6216 92.5005
R2102 VDD.n6211 VDD.n6210 92.5005
R2103 VDD.n6213 VDD.n6212 92.5005
R2104 VDD.n6207 VDD.n6206 92.5005
R2105 VDD.n6203 VDD.n6202 92.5005
R2106 VDD.n6199 VDD.n6198 92.5005
R2107 VDD.n6195 VDD.n6194 92.5005
R2108 VDD.n6191 VDD.n6190 92.5005
R2109 VDD.n6187 VDD.n6186 92.5005
R2110 VDD.n6183 VDD.n6182 92.5005
R2111 VDD.n6179 VDD.n6178 92.5005
R2112 VDD.n6175 VDD.n6174 92.5005
R2113 VDD.n6171 VDD.n6170 92.5005
R2114 VDD.n6167 VDD.n6166 92.5005
R2115 VDD.n6163 VDD.n6162 92.5005
R2116 VDD.n6159 VDD.n6158 92.5005
R2117 VDD.n6155 VDD.n6154 92.5005
R2118 VDD.n6151 VDD.n6150 92.5005
R2119 VDD.n6147 VDD.n6146 92.5005
R2120 VDD.n6141 VDD.n6140 92.5005
R2121 VDD.n6143 VDD.n6142 92.5005
R2122 VDD.n6137 VDD.n6136 92.5005
R2123 VDD.n6133 VDD.n6132 92.5005
R2124 VDD.n6129 VDD.n6128 92.5005
R2125 VDD.n6125 VDD.n6124 92.5005
R2126 VDD.n6121 VDD.n6120 92.5005
R2127 VDD.n6117 VDD.n6116 92.5005
R2128 VDD.n6113 VDD.n6112 92.5005
R2129 VDD.n6109 VDD.n6108 92.5005
R2130 VDD.n6105 VDD.n6104 92.5005
R2131 VDD.n6101 VDD.n6100 92.5005
R2132 VDD.n6097 VDD.n6096 92.5005
R2133 VDD.n6093 VDD.n6092 92.5005
R2134 VDD.n6089 VDD.n6088 92.5005
R2135 VDD.n6085 VDD.n6084 92.5005
R2136 VDD.n6081 VDD.n6080 92.5005
R2137 VDD.n6077 VDD.n6076 92.5005
R2138 VDD.n6071 VDD.n6070 92.5005
R2139 VDD.n6073 VDD.n6072 92.5005
R2140 VDD.n6067 VDD.n6066 92.5005
R2141 VDD.n6059 VDD.n6058 92.5005
R2142 VDD.n6055 VDD.n6054 92.5005
R2143 VDD.n6054 VDD.n6053 92.5005
R2144 VDD.n6050 VDD.n6049 92.5005
R2145 VDD.n6049 VDD.n6048 92.5005
R2146 VDD.n6045 VDD.n6044 92.5005
R2147 VDD.n6044 VDD.n6043 92.5005
R2148 VDD.n6040 VDD.n6039 92.5005
R2149 VDD.n6039 VDD.n6038 92.5005
R2150 VDD.n6035 VDD.n6034 92.5005
R2151 VDD.n6034 VDD.n6033 92.5005
R2152 VDD.n6030 VDD.n6029 92.5005
R2153 VDD.n6029 VDD.n6028 92.5005
R2154 VDD.n6025 VDD.n6024 92.5005
R2155 VDD.n6024 VDD.n6023 92.5005
R2156 VDD.n6020 VDD.n6019 92.5005
R2157 VDD.n6019 VDD.n6018 92.5005
R2158 VDD.n6015 VDD.n6014 92.5005
R2159 VDD.n6014 VDD.n6013 92.5005
R2160 VDD.n6010 VDD.n6009 92.5005
R2161 VDD.n6009 VDD.n6008 92.5005
R2162 VDD.n6005 VDD.n6004 92.5005
R2163 VDD.n6004 VDD.n6003 92.5005
R2164 VDD.n6000 VDD.n5999 92.5005
R2165 VDD.n5999 VDD.n5998 92.5005
R2166 VDD.n5995 VDD.n5994 92.5005
R2167 VDD.n5994 VDD.n5993 92.5005
R2168 VDD.n5987 VDD.n5986 92.5005
R2169 VDD.n5986 VDD.n5985 92.5005
R2170 VDD.n5990 VDD.n5989 92.5005
R2171 VDD.n5989 VDD.n5988 92.5005
R2172 VDD.n5982 VDD.n5981 92.5005
R2173 VDD.n5981 VDD.n5980 92.5005
R2174 VDD.n5977 VDD.n5976 92.5005
R2175 VDD.n5976 VDD.n5975 92.5005
R2176 VDD.n5972 VDD.n5971 92.5005
R2177 VDD.n5971 VDD.n5970 92.5005
R2178 VDD.n5967 VDD.n5966 92.5005
R2179 VDD.n5966 VDD.n5965 92.5005
R2180 VDD.n5962 VDD.n5961 92.5005
R2181 VDD.n5961 VDD.n5960 92.5005
R2182 VDD.n5957 VDD.n5956 92.5005
R2183 VDD.n5956 VDD.n5955 92.5005
R2184 VDD.n5952 VDD.n5951 92.5005
R2185 VDD.n5951 VDD.n5950 92.5005
R2186 VDD.n5947 VDD.n5946 92.5005
R2187 VDD.n5946 VDD.n5945 92.5005
R2188 VDD.n5942 VDD.n5941 92.5005
R2189 VDD.n5941 VDD.n5940 92.5005
R2190 VDD.n5937 VDD.n5936 92.5005
R2191 VDD.n5936 VDD.n5935 92.5005
R2192 VDD.n5932 VDD.n5931 92.5005
R2193 VDD.n5931 VDD.n5930 92.5005
R2194 VDD.n5927 VDD.n5926 92.5005
R2195 VDD.n5926 VDD.n5925 92.5005
R2196 VDD.n5922 VDD.n5921 92.5005
R2197 VDD.n5921 VDD.n5920 92.5005
R2198 VDD.n5917 VDD.n5916 92.5005
R2199 VDD.n5916 VDD.n5915 92.5005
R2200 VDD.n5912 VDD.n5911 92.5005
R2201 VDD.n5911 VDD.n5910 92.5005
R2202 VDD.n5907 VDD.n5906 92.5005
R2203 VDD.n5906 VDD.n5905 92.5005
R2204 VDD.n5899 VDD.n5898 92.5005
R2205 VDD.n5898 VDD.n5897 92.5005
R2206 VDD.n5902 VDD.n5901 92.5005
R2207 VDD.n5901 VDD.n5900 92.5005
R2208 VDD.n5894 VDD.n5893 92.5005
R2209 VDD.n5893 VDD.n5892 92.5005
R2210 VDD.n5889 VDD.n5888 92.5005
R2211 VDD.n5888 VDD.n5887 92.5005
R2212 VDD.n5884 VDD.n5883 92.5005
R2213 VDD.n5883 VDD.n5882 92.5005
R2214 VDD.n5879 VDD.n5878 92.5005
R2215 VDD.n5878 VDD.n5877 92.5005
R2216 VDD.n5874 VDD.n5873 92.5005
R2217 VDD.n5873 VDD.n5872 92.5005
R2218 VDD.n5869 VDD.n5868 92.5005
R2219 VDD.n5868 VDD.n5867 92.5005
R2220 VDD.n5864 VDD.n5863 92.5005
R2221 VDD.n5863 VDD.n5862 92.5005
R2222 VDD.n5859 VDD.n5858 92.5005
R2223 VDD.n5858 VDD.n5857 92.5005
R2224 VDD.n5854 VDD.n5853 92.5005
R2225 VDD.n5853 VDD.n5852 92.5005
R2226 VDD.n5849 VDD.n5848 92.5005
R2227 VDD.n5848 VDD.n5847 92.5005
R2228 VDD.n5836 VDD.n5835 92.5005
R2229 VDD.n5835 VDD.n5834 92.5005
R2230 VDD.n7119 VDD.n7118 92.5005
R2231 VDD.n7127 VDD.n7126 92.5005
R2232 VDD.n7131 VDD.n7130 92.5005
R2233 VDD.n5842 VDD.n5841 92.5005
R2234 VDD.n5839 VDD.n5838 92.5005
R2235 VDD.n5838 VDD.n5837 92.5005
R2236 VDD.n5830 VDD.n5829 92.5005
R2237 VDD.n5829 VDD.n5828 92.5005
R2238 VDD.n5825 VDD.n5824 92.5005
R2239 VDD.n5824 VDD.n5823 92.5005
R2240 VDD.n5820 VDD.n5819 92.5005
R2241 VDD.n5819 VDD.n5818 92.5005
R2242 VDD.n5815 VDD.n5814 92.5005
R2243 VDD.n5814 VDD.n5813 92.5005
R2244 VDD.n5810 VDD.n5809 92.5005
R2245 VDD.n5809 VDD.n5808 92.5005
R2246 VDD.n5805 VDD.n5804 92.5005
R2247 VDD.n5804 VDD.n5803 92.5005
R2248 VDD.n5800 VDD.n5799 92.5005
R2249 VDD.n5799 VDD.n5798 92.5005
R2250 VDD.n5795 VDD.n5794 92.5005
R2251 VDD.n5794 VDD.n5793 92.5005
R2252 VDD.n5790 VDD.n5789 92.5005
R2253 VDD.n5789 VDD.n5788 92.5005
R2254 VDD.n5785 VDD.n5784 92.5005
R2255 VDD.n5784 VDD.n5783 92.5005
R2256 VDD.n5780 VDD.n5779 92.5005
R2257 VDD.n5779 VDD.n5778 92.5005
R2258 VDD.n5777 VDD.n5776 92.5005
R2259 VDD.n5776 VDD.n5775 92.5005
R2260 VDD.n5772 VDD.n5771 92.5005
R2261 VDD.n5771 VDD.n5770 92.5005
R2262 VDD.n5767 VDD.n5766 92.5005
R2263 VDD.n5766 VDD.n5765 92.5005
R2264 VDD.n5762 VDD.n5761 92.5005
R2265 VDD.n5761 VDD.n5760 92.5005
R2266 VDD.n5757 VDD.n5756 92.5005
R2267 VDD.n5756 VDD.n5755 92.5005
R2268 VDD.n5752 VDD.n5751 92.5005
R2269 VDD.n5751 VDD.n5750 92.5005
R2270 VDD.n5747 VDD.n5746 92.5005
R2271 VDD.n5746 VDD.n5745 92.5005
R2272 VDD.n5742 VDD.n5741 92.5005
R2273 VDD.n5741 VDD.n5740 92.5005
R2274 VDD.n5737 VDD.n5736 92.5005
R2275 VDD.n5736 VDD.n5735 92.5005
R2276 VDD.n5732 VDD.n5731 92.5005
R2277 VDD.n5731 VDD.n5730 92.5005
R2278 VDD.n5727 VDD.n5726 92.5005
R2279 VDD.n5726 VDD.n5725 92.5005
R2280 VDD.n5722 VDD.n5721 92.5005
R2281 VDD.n5721 VDD.n5720 92.5005
R2282 VDD.n5717 VDD.n5716 92.5005
R2283 VDD.n5716 VDD.n5715 92.5005
R2284 VDD.n5712 VDD.n5711 92.5005
R2285 VDD.n5711 VDD.n5710 92.5005
R2286 VDD.n5707 VDD.n5706 92.5005
R2287 VDD.n5706 VDD.n5705 92.5005
R2288 VDD.n5702 VDD.n5701 92.5005
R2289 VDD.n5701 VDD.n5700 92.5005
R2290 VDD.n5697 VDD.n5696 92.5005
R2291 VDD.n5696 VDD.n5695 92.5005
R2292 VDD.n5692 VDD.n5691 92.5005
R2293 VDD.n5691 VDD.n5690 92.5005
R2294 VDD.n5689 VDD.n5688 92.5005
R2295 VDD.n5688 VDD.n5687 92.5005
R2296 VDD.n5684 VDD.n5683 92.5005
R2297 VDD.n5683 VDD.n5682 92.5005
R2298 VDD.n5679 VDD.n5678 92.5005
R2299 VDD.n5678 VDD.n5677 92.5005
R2300 VDD.n5674 VDD.n5673 92.5005
R2301 VDD.n5673 VDD.n5672 92.5005
R2302 VDD.n5669 VDD.n5668 92.5005
R2303 VDD.n5668 VDD.n5667 92.5005
R2304 VDD.n5664 VDD.n5663 92.5005
R2305 VDD.n5663 VDD.n5662 92.5005
R2306 VDD.n5659 VDD.n5658 92.5005
R2307 VDD.n5658 VDD.n5657 92.5005
R2308 VDD.n5654 VDD.n5653 92.5005
R2309 VDD.n5653 VDD.n5652 92.5005
R2310 VDD.n5649 VDD.n5648 92.5005
R2311 VDD.n5648 VDD.n5647 92.5005
R2312 VDD.n5644 VDD.n5643 92.5005
R2313 VDD.n5643 VDD.n5642 92.5005
R2314 VDD.n5639 VDD.n5638 92.5005
R2315 VDD.n5638 VDD.n5637 92.5005
R2316 VDD.n5634 VDD.n5633 92.5005
R2317 VDD.n5633 VDD.n5632 92.5005
R2318 VDD.n5629 VDD.n5628 92.5005
R2319 VDD.n5628 VDD.n5627 92.5005
R2320 VDD.n5624 VDD.n5623 92.5005
R2321 VDD.n5623 VDD.n5622 92.5005
R2322 VDD.n5619 VDD.n5618 92.5005
R2323 VDD.n5618 VDD.n5617 92.5005
R2324 VDD.n5614 VDD.n5613 92.5005
R2325 VDD.n5613 VDD.n5612 92.5005
R2326 VDD.n5609 VDD.n5608 92.5005
R2327 VDD.n5608 VDD.n5607 92.5005
R2328 VDD.n5604 VDD.n5603 92.5005
R2329 VDD.n5603 VDD.n5602 92.5005
R2330 VDD.n5601 VDD.n5600 92.5005
R2331 VDD.n5600 VDD.n5599 92.5005
R2332 VDD.n5596 VDD.n5595 92.5005
R2333 VDD.n5595 VDD.n5594 92.5005
R2334 VDD.n5591 VDD.n5590 92.5005
R2335 VDD.n5590 VDD.n5589 92.5005
R2336 VDD.n5586 VDD.n5585 92.5005
R2337 VDD.n5585 VDD.n5584 92.5005
R2338 VDD.n5581 VDD.n5580 92.5005
R2339 VDD.n5580 VDD.n5579 92.5005
R2340 VDD.n5576 VDD.n5575 92.5005
R2341 VDD.n5575 VDD.n5574 92.5005
R2342 VDD.n5571 VDD.n5570 92.5005
R2343 VDD.n5570 VDD.n5569 92.5005
R2344 VDD.n5566 VDD.n5565 92.5005
R2345 VDD.n5565 VDD.n5564 92.5005
R2346 VDD.n5561 VDD.n5560 92.5005
R2347 VDD.n5560 VDD.n5559 92.5005
R2348 VDD.n5556 VDD.n5555 92.5005
R2349 VDD.n5555 VDD.n5554 92.5005
R2350 VDD.n5551 VDD.n5550 92.5005
R2351 VDD.n5550 VDD.n5549 92.5005
R2352 VDD.n5546 VDD.n5545 92.5005
R2353 VDD.n5545 VDD.n5544 92.5005
R2354 VDD.n5541 VDD.n5540 92.5005
R2355 VDD.n5540 VDD.n5539 92.5005
R2356 VDD.n5536 VDD.n5535 92.5005
R2357 VDD.n5535 VDD.n5534 92.5005
R2358 VDD.n5531 VDD.n5530 92.5005
R2359 VDD.n5530 VDD.n5529 92.5005
R2360 VDD.n5526 VDD.n5525 92.5005
R2361 VDD.n5525 VDD.n5524 92.5005
R2362 VDD.n5521 VDD.n5520 92.5005
R2363 VDD.n5520 VDD.n5519 92.5005
R2364 VDD.n5516 VDD.n5515 92.5005
R2365 VDD.n5515 VDD.n5514 92.5005
R2366 VDD.n5513 VDD.n5512 92.5005
R2367 VDD.n5512 VDD.n5511 92.5005
R2368 VDD.n5508 VDD.n5507 92.5005
R2369 VDD.n5507 VDD.n5506 92.5005
R2370 VDD.n5503 VDD.n5502 92.5005
R2371 VDD.n5502 VDD.n5501 92.5005
R2372 VDD.n5498 VDD.n5497 92.5005
R2373 VDD.n5497 VDD.n5496 92.5005
R2374 VDD.n5493 VDD.n5492 92.5005
R2375 VDD.n5492 VDD.n5491 92.5005
R2376 VDD.n5488 VDD.n5487 92.5005
R2377 VDD.n5487 VDD.n5486 92.5005
R2378 VDD.n5483 VDD.n5482 92.5005
R2379 VDD.n5482 VDD.n5481 92.5005
R2380 VDD.n5478 VDD.n5477 92.5005
R2381 VDD.n5477 VDD.n5476 92.5005
R2382 VDD.n5473 VDD.n5472 92.5005
R2383 VDD.n5472 VDD.n5471 92.5005
R2384 VDD.n5468 VDD.n5467 92.5005
R2385 VDD.n5467 VDD.n5466 92.5005
R2386 VDD.n5463 VDD.n5462 92.5005
R2387 VDD.n5462 VDD.n5461 92.5005
R2388 VDD.n5458 VDD.n5457 92.5005
R2389 VDD.n5457 VDD.n5456 92.5005
R2390 VDD.n5453 VDD.n5452 92.5005
R2391 VDD.n5452 VDD.n5451 92.5005
R2392 VDD.n6829 VDD.n6828 92.5005
R2393 VDD.n6828 VDD.n6827 92.5005
R2394 VDD.n6834 VDD.n6833 92.5005
R2395 VDD.n6833 VDD.n6832 92.5005
R2396 VDD.n6839 VDD.n6838 92.5005
R2397 VDD.n6838 VDD.n6837 92.5005
R2398 VDD.n6844 VDD.n6843 92.5005
R2399 VDD.n6843 VDD.n6842 92.5005
R2400 VDD.n6852 VDD.n6851 92.5005
R2401 VDD.n6851 VDD.n6850 92.5005
R2402 VDD.n6849 VDD.n6848 92.5005
R2403 VDD.n6848 VDD.n6847 92.5005
R2404 VDD.n6857 VDD.n6856 92.5005
R2405 VDD.n6856 VDD.n6855 92.5005
R2406 VDD.n6862 VDD.n6861 92.5005
R2407 VDD.n6861 VDD.n6860 92.5005
R2408 VDD.n6867 VDD.n6866 92.5005
R2409 VDD.n6866 VDD.n6865 92.5005
R2410 VDD.n6872 VDD.n6871 92.5005
R2411 VDD.n6871 VDD.n6870 92.5005
R2412 VDD.n6877 VDD.n6876 92.5005
R2413 VDD.n6876 VDD.n6875 92.5005
R2414 VDD.n6882 VDD.n6881 92.5005
R2415 VDD.n6881 VDD.n6880 92.5005
R2416 VDD.n6887 VDD.n6886 92.5005
R2417 VDD.n6886 VDD.n6885 92.5005
R2418 VDD.n6892 VDD.n6891 92.5005
R2419 VDD.n6891 VDD.n6890 92.5005
R2420 VDD.n6897 VDD.n6896 92.5005
R2421 VDD.n6896 VDD.n6895 92.5005
R2422 VDD.n6902 VDD.n6901 92.5005
R2423 VDD.n6901 VDD.n6900 92.5005
R2424 VDD.n6907 VDD.n6906 92.5005
R2425 VDD.n6906 VDD.n6905 92.5005
R2426 VDD.n6912 VDD.n6911 92.5005
R2427 VDD.n6911 VDD.n6910 92.5005
R2428 VDD.n6917 VDD.n6916 92.5005
R2429 VDD.n6916 VDD.n6915 92.5005
R2430 VDD.n6922 VDD.n6921 92.5005
R2431 VDD.n6921 VDD.n6920 92.5005
R2432 VDD.n6927 VDD.n6926 92.5005
R2433 VDD.n6926 VDD.n6925 92.5005
R2434 VDD.n6932 VDD.n6931 92.5005
R2435 VDD.n6931 VDD.n6930 92.5005
R2436 VDD.n6940 VDD.n6939 92.5005
R2437 VDD.n6939 VDD.n6938 92.5005
R2438 VDD.n6937 VDD.n6936 92.5005
R2439 VDD.n6936 VDD.n6935 92.5005
R2440 VDD.n6945 VDD.n6944 92.5005
R2441 VDD.n6944 VDD.n6943 92.5005
R2442 VDD.n6950 VDD.n6949 92.5005
R2443 VDD.n6949 VDD.n6948 92.5005
R2444 VDD.n6955 VDD.n6954 92.5005
R2445 VDD.n6954 VDD.n6953 92.5005
R2446 VDD.n6960 VDD.n6959 92.5005
R2447 VDD.n6959 VDD.n6958 92.5005
R2448 VDD.n6965 VDD.n6964 92.5005
R2449 VDD.n6964 VDD.n6963 92.5005
R2450 VDD.n6970 VDD.n6969 92.5005
R2451 VDD.n6969 VDD.n6968 92.5005
R2452 VDD.n6975 VDD.n6974 92.5005
R2453 VDD.n6974 VDD.n6973 92.5005
R2454 VDD.n6980 VDD.n6979 92.5005
R2455 VDD.n6979 VDD.n6978 92.5005
R2456 VDD.n6985 VDD.n6984 92.5005
R2457 VDD.n6984 VDD.n6983 92.5005
R2458 VDD.n6990 VDD.n6989 92.5005
R2459 VDD.n6989 VDD.n6988 92.5005
R2460 VDD.n6995 VDD.n6994 92.5005
R2461 VDD.n6994 VDD.n6993 92.5005
R2462 VDD.n7000 VDD.n6999 92.5005
R2463 VDD.n6999 VDD.n6998 92.5005
R2464 VDD.n7005 VDD.n7004 92.5005
R2465 VDD.n7004 VDD.n7003 92.5005
R2466 VDD.n7010 VDD.n7009 92.5005
R2467 VDD.n7009 VDD.n7008 92.5005
R2468 VDD.n7015 VDD.n7014 92.5005
R2469 VDD.n7014 VDD.n7013 92.5005
R2470 VDD.n7020 VDD.n7019 92.5005
R2471 VDD.n7019 VDD.n7018 92.5005
R2472 VDD.n7028 VDD.n7027 92.5005
R2473 VDD.n7027 VDD.n7026 92.5005
R2474 VDD.n7025 VDD.n7024 92.5005
R2475 VDD.n7024 VDD.n7023 92.5005
R2476 VDD.n7033 VDD.n7032 92.5005
R2477 VDD.n7032 VDD.n7031 92.5005
R2478 VDD.n7038 VDD.n7037 92.5005
R2479 VDD.n7037 VDD.n7036 92.5005
R2480 VDD.n7043 VDD.n7042 92.5005
R2481 VDD.n7042 VDD.n7041 92.5005
R2482 VDD.n7048 VDD.n7047 92.5005
R2483 VDD.n7047 VDD.n7046 92.5005
R2484 VDD.n7053 VDD.n7052 92.5005
R2485 VDD.n7052 VDD.n7051 92.5005
R2486 VDD.n7058 VDD.n7057 92.5005
R2487 VDD.n7057 VDD.n7056 92.5005
R2488 VDD.n7063 VDD.n7062 92.5005
R2489 VDD.n7062 VDD.n7061 92.5005
R2490 VDD.n7068 VDD.n7067 92.5005
R2491 VDD.n7067 VDD.n7066 92.5005
R2492 VDD.n7073 VDD.n7072 92.5005
R2493 VDD.n7072 VDD.n7071 92.5005
R2494 VDD.n7078 VDD.n7077 92.5005
R2495 VDD.n7077 VDD.n7076 92.5005
R2496 VDD.n7083 VDD.n7082 92.5005
R2497 VDD.n7082 VDD.n7081 92.5005
R2498 VDD.n7088 VDD.n7087 92.5005
R2499 VDD.n7087 VDD.n7086 92.5005
R2500 VDD.n7093 VDD.n7092 92.5005
R2501 VDD.n7092 VDD.n7091 92.5005
R2502 VDD.n7098 VDD.n7097 92.5005
R2503 VDD.n7097 VDD.n7096 92.5005
R2504 VDD.n7103 VDD.n7102 92.5005
R2505 VDD.n7102 VDD.n7101 92.5005
R2506 VDD.n7108 VDD.n7107 92.5005
R2507 VDD.n7107 VDD.n7106 92.5005
R2508 VDD.n7123 VDD.n7122 92.5005
R2509 VDD.n7122 VDD.n7121 92.5005
R2510 VDD.n7112 VDD.n7111 92.5005
R2511 VDD.n7115 VDD.n7114 92.5005
R2512 VDD.n7136 VDD.n7135 92.5005
R2513 VDD.n7135 VDD.n7134 92.5005
R2514 VDD.n7141 VDD.n7140 92.5005
R2515 VDD.n7140 VDD.n7139 92.5005
R2516 VDD.n7146 VDD.n7145 92.5005
R2517 VDD.n7145 VDD.n7144 92.5005
R2518 VDD.n7151 VDD.n7150 92.5005
R2519 VDD.n7150 VDD.n7149 92.5005
R2520 VDD.n7156 VDD.n7155 92.5005
R2521 VDD.n7155 VDD.n7154 92.5005
R2522 VDD.n7161 VDD.n7160 92.5005
R2523 VDD.n7160 VDD.n7159 92.5005
R2524 VDD.n7166 VDD.n7165 92.5005
R2525 VDD.n7165 VDD.n7164 92.5005
R2526 VDD.n7174 VDD.n7173 92.5005
R2527 VDD.n7173 VDD.n7172 92.5005
R2528 VDD.n7171 VDD.n7170 92.5005
R2529 VDD.n7170 VDD.n7169 92.5005
R2530 VDD.n7179 VDD.n7178 92.5005
R2531 VDD.n7178 VDD.n7177 92.5005
R2532 VDD.n7184 VDD.n7183 92.5005
R2533 VDD.n7183 VDD.n7182 92.5005
R2534 VDD.n7189 VDD.n7188 92.5005
R2535 VDD.n7188 VDD.n7187 92.5005
R2536 VDD.n7194 VDD.n7193 92.5005
R2537 VDD.n7193 VDD.n7192 92.5005
R2538 VDD.n7199 VDD.n7198 92.5005
R2539 VDD.n7198 VDD.n7197 92.5005
R2540 VDD.n7204 VDD.n7203 92.5005
R2541 VDD.n7203 VDD.n7202 92.5005
R2542 VDD.n7209 VDD.n7208 92.5005
R2543 VDD.n7208 VDD.n7207 92.5005
R2544 VDD.n7214 VDD.n7213 92.5005
R2545 VDD.n7213 VDD.n7212 92.5005
R2546 VDD.n7218 VDD.n7217 92.5005
R2547 VDD.n7217 VDD.n7216 92.5005
R2548 VDD.n7223 VDD.n7222 92.5005
R2549 VDD.n7222 VDD.n7221 92.5005
R2550 VDD.n7228 VDD.n7227 92.5005
R2551 VDD.n7227 VDD.n7226 92.5005
R2552 VDD.n7233 VDD.n7232 92.5005
R2553 VDD.n7232 VDD.n7231 92.5005
R2554 VDD.n7238 VDD.n7237 92.5005
R2555 VDD.n7237 VDD.n7236 92.5005
R2556 VDD.n7243 VDD.n7242 92.5005
R2557 VDD.n7242 VDD.n7241 92.5005
R2558 VDD.n7248 VDD.n7247 92.5005
R2559 VDD.n7247 VDD.n7246 92.5005
R2560 VDD.n7253 VDD.n7252 92.5005
R2561 VDD.n7252 VDD.n7251 92.5005
R2562 VDD.n7261 VDD.n7260 92.5005
R2563 VDD.n7260 VDD.n7259 92.5005
R2564 VDD.n7258 VDD.n7257 92.5005
R2565 VDD.n7257 VDD.n7256 92.5005
R2566 VDD.n7266 VDD.n7265 92.5005
R2567 VDD.n7265 VDD.n7264 92.5005
R2568 VDD.n7271 VDD.n7270 92.5005
R2569 VDD.n7270 VDD.n7269 92.5005
R2570 VDD.n7276 VDD.n7275 92.5005
R2571 VDD.n7275 VDD.n7274 92.5005
R2572 VDD.n7281 VDD.n7280 92.5005
R2573 VDD.n7280 VDD.n7279 92.5005
R2574 VDD.n7286 VDD.n7285 92.5005
R2575 VDD.n7285 VDD.n7284 92.5005
R2576 VDD.n7291 VDD.n7290 92.5005
R2577 VDD.n7290 VDD.n7289 92.5005
R2578 VDD.n7296 VDD.n7295 92.5005
R2579 VDD.n7295 VDD.n7294 92.5005
R2580 VDD.n7301 VDD.n7300 92.5005
R2581 VDD.n7300 VDD.n7299 92.5005
R2582 VDD.n7305 VDD.n7304 92.5005
R2583 VDD.n7304 VDD.n7303 92.5005
R2584 VDD.n7310 VDD.n7309 92.5005
R2585 VDD.n7309 VDD.n7308 92.5005
R2586 VDD.n7315 VDD.n7314 92.5005
R2587 VDD.n7314 VDD.n7313 92.5005
R2588 VDD.n7320 VDD.n7319 92.5005
R2589 VDD.n7319 VDD.n7318 92.5005
R2590 VDD.n7325 VDD.n7324 92.5005
R2591 VDD.n7324 VDD.n7323 92.5005
R2592 VDD.n7330 VDD.n7329 92.5005
R2593 VDD.n7329 VDD.n7328 92.5005
R2594 VDD.n7335 VDD.n7334 92.5005
R2595 VDD.n7334 VDD.n7333 92.5005
R2596 VDD.n7340 VDD.n7339 92.5005
R2597 VDD.n7339 VDD.n7338 92.5005
R2598 VDD.n7346 VDD.n7345 92.5005
R2599 VDD.n3471 VDD.n3470 92.5005
R2600 VDD.n3473 VDD.n3472 92.5005
R2601 VDD.n3475 VDD.n3474 92.5005
R2602 VDD.n3477 VDD.n3476 92.5005
R2603 VDD.n3479 VDD.n3478 92.5005
R2604 VDD.n3482 VDD.n3481 92.5005
R2605 VDD.n3485 VDD.n3484 92.5005
R2606 VDD.n3488 VDD.n3487 92.5005
R2607 VDD.n3491 VDD.n3490 92.5005
R2608 VDD.n3494 VDD.n3493 92.5005
R2609 VDD.n3497 VDD.n3496 92.5005
R2610 VDD.n3500 VDD.n3499 92.5005
R2611 VDD.n3503 VDD.n3502 92.5005
R2612 VDD.n3506 VDD.n3505 92.5005
R2613 VDD.n3509 VDD.n3508 92.5005
R2614 VDD.n3512 VDD.n3511 92.5005
R2615 VDD.n3515 VDD.n3514 92.5005
R2616 VDD.n3518 VDD.n3517 92.5005
R2617 VDD.n3521 VDD.n3520 92.5005
R2618 VDD.n3524 VDD.n3523 92.5005
R2619 VDD.n3527 VDD.n3526 92.5005
R2620 VDD.n3530 VDD.n3529 92.5005
R2621 VDD.n3533 VDD.n3532 92.5005
R2622 VDD.n3536 VDD.n3535 92.5005
R2623 VDD.n3540 VDD.n3539 92.5005
R2624 VDD.n3454 VDD.n3453 92.5005
R2625 VDD.n3451 VDD.n3450 92.5005
R2626 VDD.n3448 VDD.n3447 92.5005
R2627 VDD.n3445 VDD.n3444 92.5005
R2628 VDD.n3442 VDD.n3441 92.5005
R2629 VDD.n3439 VDD.n3438 92.5005
R2630 VDD.n3577 VDD.n3576 92.5005
R2631 VDD.n3580 VDD.n3579 92.5005
R2632 VDD.n3583 VDD.n3582 92.5005
R2633 VDD.n3586 VDD.n3585 92.5005
R2634 VDD.n3589 VDD.n3588 92.5005
R2635 VDD.n3592 VDD.n3591 92.5005
R2636 VDD.n3595 VDD.n3594 92.5005
R2637 VDD.n3575 VDD.n3574 92.5005
R2638 VDD.n3571 VDD.n3570 92.5005
R2639 VDD.n3568 VDD.n3567 92.5005
R2640 VDD.n3565 VDD.n3564 92.5005
R2641 VDD.n3562 VDD.n3561 92.5005
R2642 VDD.n3559 VDD.n3558 92.5005
R2643 VDD.n3556 VDD.n3555 92.5005
R2644 VDD.n3604 VDD.n3603 92.5005
R2645 VDD.n3607 VDD.n3606 92.5005
R2646 VDD.n3610 VDD.n3609 92.5005
R2647 VDD.n3613 VDD.n3612 92.5005
R2648 VDD.n3616 VDD.n3615 92.5005
R2649 VDD.n3619 VDD.n3618 92.5005
R2650 VDD.n3469 VDD.n3468 92.5005
R2651 VDD.n3467 VDD.n3466 92.5005
R2652 VDD.n3465 VDD.n3464 92.5005
R2653 VDD.n3463 VDD.n3462 92.5005
R2654 VDD.n8517 VDD.n8516 92.5005
R2655 VDD.n8508 VDD.n8507 92.5005
R2656 VDD.n8499 VDD.n8498 92.5005
R2657 VDD.n8491 VDD.n8490 92.5005
R2658 VDD.n8482 VDD.n8481 92.5005
R2659 VDD.n8470 VDD.n8469 92.5005
R2660 VDD.n8461 VDD.n8460 92.5005
R2661 VDD.n8451 VDD.n8450 92.5005
R2662 VDD.n8452 VDD.n8451 92.5005
R2663 VDD.n8441 VDD.n8440 92.5005
R2664 VDD.n8442 VDD.n8441 92.5005
R2665 VDD.n8431 VDD.n8430 92.5005
R2666 VDD.n8432 VDD.n8431 92.5005
R2667 VDD.n8421 VDD.n8420 92.5005
R2668 VDD.n8422 VDD.n8421 92.5005
R2669 VDD.n8411 VDD.n8410 92.5005
R2670 VDD.n8412 VDD.n8411 92.5005
R2671 VDD.n4119 VDD.n4118 92.5005
R2672 VDD.n4120 VDD.n4119 92.5005
R2673 VDD.n4123 VDD.n4122 92.5005
R2674 VDD.n4124 VDD.n4123 92.5005
R2675 VDD.n4127 VDD.n4126 92.5005
R2676 VDD.n4128 VDD.n4127 92.5005
R2677 VDD.n4131 VDD.n4130 92.5005
R2678 VDD.n4132 VDD.n4131 92.5005
R2679 VDD.n4135 VDD.n4134 92.5005
R2680 VDD.n4136 VDD.n4135 92.5005
R2681 VDD.n4139 VDD.n4138 92.5005
R2682 VDD.n4140 VDD.n4139 92.5005
R2683 VDD.n4143 VDD.n4142 92.5005
R2684 VDD.n4144 VDD.n4143 92.5005
R2685 VDD.n4147 VDD.n4146 92.5005
R2686 VDD.n4148 VDD.n4147 92.5005
R2687 VDD.n4151 VDD.n4150 92.5005
R2688 VDD.n4152 VDD.n4151 92.5005
R2689 VDD.n4155 VDD.n4154 92.5005
R2690 VDD.n4156 VDD.n4155 92.5005
R2691 VDD.n4159 VDD.n4158 92.5005
R2692 VDD.n4160 VDD.n4159 92.5005
R2693 VDD.n4163 VDD.n4162 92.5005
R2694 VDD.n4164 VDD.n4163 92.5005
R2695 VDD.n4167 VDD.n4166 92.5005
R2696 VDD.n4168 VDD.n4167 92.5005
R2697 VDD.n4171 VDD.n4170 92.5005
R2698 VDD.n4172 VDD.n4171 92.5005
R2699 VDD.n4175 VDD.n4174 92.5005
R2700 VDD.n4176 VDD.n4175 92.5005
R2701 VDD.n4179 VDD.n4178 92.5005
R2702 VDD.n4180 VDD.n4179 92.5005
R2703 VDD.n4183 VDD.n4182 92.5005
R2704 VDD.n4184 VDD.n4183 92.5005
R2705 VDD.n4187 VDD.n4186 92.5005
R2706 VDD.n4188 VDD.n4187 92.5005
R2707 VDD.n4191 VDD.n4190 92.5005
R2708 VDD.n4192 VDD.n4191 92.5005
R2709 VDD.n4195 VDD.n4194 92.5005
R2710 VDD.n4196 VDD.n4195 92.5005
R2711 VDD.n4107 VDD.n4106 92.5005
R2712 VDD.n4108 VDD.n4107 92.5005
R2713 VDD.n4102 VDD.n4101 92.5005
R2714 VDD.n4103 VDD.n4102 92.5005
R2715 VDD.n4098 VDD.n4097 92.5005
R2716 VDD.n4099 VDD.n4098 92.5005
R2717 VDD.n4094 VDD.n4093 92.5005
R2718 VDD.n4095 VDD.n4094 92.5005
R2719 VDD.n4090 VDD.n4089 92.5005
R2720 VDD.n4091 VDD.n4090 92.5005
R2721 VDD.n4086 VDD.n4085 92.5005
R2722 VDD.n4087 VDD.n4086 92.5005
R2723 VDD.n4082 VDD.n4081 92.5005
R2724 VDD.n4083 VDD.n4082 92.5005
R2725 VDD.n4224 VDD.n4223 92.5005
R2726 VDD.n4225 VDD.n4224 92.5005
R2727 VDD.n4228 VDD.n4227 92.5005
R2728 VDD.n4229 VDD.n4228 92.5005
R2729 VDD.n4232 VDD.n4231 92.5005
R2730 VDD.n4233 VDD.n4232 92.5005
R2731 VDD.n4221 VDD.n4220 92.5005
R2732 VDD.n4222 VDD.n4221 92.5005
R2733 VDD.n4217 VDD.n4216 92.5005
R2734 VDD.n4218 VDD.n4217 92.5005
R2735 VDD.n4213 VDD.n4212 92.5005
R2736 VDD.n4214 VDD.n4213 92.5005
R2737 VDD.n4035 VDD.n4034 92.5005
R2738 VDD.n4036 VDD.n4035 92.5005
R2739 VDD.n4039 VDD.n4038 92.5005
R2740 VDD.n4040 VDD.n4039 92.5005
R2741 VDD.n4043 VDD.n4042 92.5005
R2742 VDD.n4044 VDD.n4043 92.5005
R2743 VDD.n4047 VDD.n4046 92.5005
R2744 VDD.n4048 VDD.n4047 92.5005
R2745 VDD.n4051 VDD.n4050 92.5005
R2746 VDD.n4052 VDD.n4051 92.5005
R2747 VDD.n4055 VDD.n4054 92.5005
R2748 VDD.n4056 VDD.n4055 92.5005
R2749 VDD.n4032 VDD.n4031 92.5005
R2750 VDD.n4033 VDD.n4032 92.5005
R2751 VDD.n4027 VDD.n4026 92.5005
R2752 VDD.n4028 VDD.n4027 92.5005
R2753 VDD.n4023 VDD.n4022 92.5005
R2754 VDD.n4024 VDD.n4023 92.5005
R2755 VDD.n4019 VDD.n4018 92.5005
R2756 VDD.n4020 VDD.n4019 92.5005
R2757 VDD.n4014 VDD.n4013 92.5005
R2758 VDD.n4015 VDD.n4014 92.5005
R2759 VDD.n3973 VDD.n3972 92.5005
R2760 VDD.n3974 VDD.n3973 92.5005
R2761 VDD.n3969 VDD.n3968 92.5005
R2762 VDD.n3970 VDD.n3969 92.5005
R2763 VDD.n7344 VDD.n7343 92.5005
R2764 VDD.n7350 VDD.n7349 92.5005
R2765 VDD.n7354 VDD.n7353 92.5005
R2766 VDD.n7358 VDD.n7357 92.5005
R2767 VDD.n7362 VDD.n7361 92.5005
R2768 VDD.n7366 VDD.n7365 92.5005
R2769 VDD.n7370 VDD.n7369 92.5005
R2770 VDD.n7374 VDD.n7373 92.5005
R2771 VDD.n7378 VDD.n7377 92.5005
R2772 VDD.n7381 VDD.n7380 92.5005
R2773 VDD.n7385 VDD.n7384 92.5005
R2774 VDD.n7389 VDD.n7388 92.5005
R2775 VDD.n7393 VDD.n7392 92.5005
R2776 VDD.n7397 VDD.n7396 92.5005
R2777 VDD.n7401 VDD.n7400 92.5005
R2778 VDD.n7405 VDD.n7404 92.5005
R2779 VDD.n7409 VDD.n7408 92.5005
R2780 VDD.n7415 VDD.n7414 92.5005
R2781 VDD.n7413 VDD.n7412 92.5005
R2782 VDD.n7419 VDD.n7418 92.5005
R2783 VDD.n7423 VDD.n7422 92.5005
R2784 VDD.n7427 VDD.n7426 92.5005
R2785 VDD.n7431 VDD.n7430 92.5005
R2786 VDD.n7435 VDD.n7434 92.5005
R2787 VDD.n7439 VDD.n7438 92.5005
R2788 VDD.n7443 VDD.n7442 92.5005
R2789 VDD.n7447 VDD.n7446 92.5005
R2790 VDD.n7450 VDD.n7449 92.5005
R2791 VDD.n7454 VDD.n7453 92.5005
R2792 VDD.n7458 VDD.n7457 92.5005
R2793 VDD.n7462 VDD.n7461 92.5005
R2794 VDD.n7466 VDD.n7465 92.5005
R2795 VDD.n7470 VDD.n7469 92.5005
R2796 VDD.n7474 VDD.n7473 92.5005
R2797 VDD.n7478 VDD.n7477 92.5005
R2798 VDD.n7484 VDD.n7483 92.5005
R2799 VDD.n7482 VDD.n7481 92.5005
R2800 VDD.n7494 VDD.n7493 92.5005
R2801 VDD.n8146 VDD.n8145 92.5005
R2802 VDD.n8151 VDD.n8150 92.5005
R2803 VDD.n8157 VDD.n8156 92.5005
R2804 VDD.n8163 VDD.n8162 92.5005
R2805 VDD.n8169 VDD.n8168 92.5005
R2806 VDD.n8175 VDD.n8174 92.5005
R2807 VDD.n8181 VDD.n8180 92.5005
R2808 VDD.n8187 VDD.n8186 92.5005
R2809 VDD.n8193 VDD.n8192 92.5005
R2810 VDD.n8199 VDD.n8198 92.5005
R2811 VDD.n8201 VDD.n8200 92.5005
R2812 VDD.n8207 VDD.n8206 92.5005
R2813 VDD.n8213 VDD.n8212 92.5005
R2814 VDD.n8219 VDD.n8218 92.5005
R2815 VDD.n8225 VDD.n8224 92.5005
R2816 VDD.n8231 VDD.n8230 92.5005
R2817 VDD.n8237 VDD.n8236 92.5005
R2818 VDD.n8245 VDD.n8244 92.5005
R2819 VDD.n8251 VDD.n8250 92.5005
R2820 VDD.n8256 VDD.n8255 92.5005
R2821 VDD.n8262 VDD.n8261 92.5005
R2822 VDD.n8268 VDD.n8267 92.5005
R2823 VDD.n8274 VDD.n8273 92.5005
R2824 VDD.n8280 VDD.n8279 92.5005
R2825 VDD.n8286 VDD.n8285 92.5005
R2826 VDD.n8292 VDD.n8291 92.5005
R2827 VDD.n8298 VDD.n8297 92.5005
R2828 VDD.n8304 VDD.n8303 92.5005
R2829 VDD.n8306 VDD.n8305 92.5005
R2830 VDD.n8312 VDD.n8311 92.5005
R2831 VDD.n8318 VDD.n8317 92.5005
R2832 VDD.n8324 VDD.n8323 92.5005
R2833 VDD.n8330 VDD.n8329 92.5005
R2834 VDD.n8336 VDD.n8335 92.5005
R2835 VDD.n8342 VDD.n8341 92.5005
R2836 VDD.n8350 VDD.n8349 92.5005
R2837 VDD.n8356 VDD.n8355 92.5005
R2838 VDD.n8361 VDD.n8360 92.5005
R2839 VDD.n8367 VDD.n8366 92.5005
R2840 VDD.n8373 VDD.n8372 92.5005
R2841 VDD.n8379 VDD.n8378 92.5005
R2842 VDD.n8385 VDD.n8384 92.5005
R2843 VDD.n8391 VDD.n8390 92.5005
R2844 VDD.n8397 VDD.n8396 92.5005
R2845 VDD.n8403 VDD.n8402 92.5005
R2846 VDD.n8409 VDD.n8408 92.5005
R2847 VDD.n8414 VDD.n8413 92.5005
R2848 VDD.n8413 VDD.n8412 92.5005
R2849 VDD.n8424 VDD.n8423 92.5005
R2850 VDD.n8423 VDD.n8422 92.5005
R2851 VDD.n8434 VDD.n8433 92.5005
R2852 VDD.n8433 VDD.n8432 92.5005
R2853 VDD.n8444 VDD.n8443 92.5005
R2854 VDD.n8443 VDD.n8442 92.5005
R2855 VDD.n8454 VDD.n8453 92.5005
R2856 VDD.n8453 VDD.n8452 92.5005
R2857 VDD.n8463 VDD.n8462 92.5005
R2858 VDD.n8462 VDD.n8461 92.5005
R2859 VDD.n8472 VDD.n8471 92.5005
R2860 VDD.n8471 VDD.n8470 92.5005
R2861 VDD.n8484 VDD.n8483 92.5005
R2862 VDD.n8483 VDD.n8482 92.5005
R2863 VDD.n8493 VDD.n8492 92.5005
R2864 VDD.n8492 VDD.n8491 92.5005
R2865 VDD.n8501 VDD.n8500 92.5005
R2866 VDD.n8500 VDD.n8499 92.5005
R2867 VDD.n8510 VDD.n8509 92.5005
R2868 VDD.n8509 VDD.n8508 92.5005
R2869 VDD.n8519 VDD.n8518 92.5005
R2870 VDD.n8518 VDD.n8517 92.5005
R2871 VDD.n8527 VDD.n8526 92.5005
R2872 VDD.n8526 VDD.n8525 92.5005
R2873 VDD.n8535 VDD.n8534 92.5005
R2874 VDD.n8534 VDD.n8533 92.5005
R2875 VDD.n8541 VDD.n8540 92.5005
R2876 VDD.n8149 VDD.n8148 92.5005
R2877 VDD.n8155 VDD.n8154 92.5005
R2878 VDD.n8161 VDD.n8160 92.5005
R2879 VDD.n8167 VDD.n8166 92.5005
R2880 VDD.n8173 VDD.n8172 92.5005
R2881 VDD.n8179 VDD.n8178 92.5005
R2882 VDD.n8185 VDD.n8184 92.5005
R2883 VDD.n8189 VDD.n8188 92.5005
R2884 VDD.n8195 VDD.n8194 92.5005
R2885 VDD.n8203 VDD.n8202 92.5005
R2886 VDD.n8209 VDD.n8208 92.5005
R2887 VDD.n8215 VDD.n8214 92.5005
R2888 VDD.n8221 VDD.n8220 92.5005
R2889 VDD.n8227 VDD.n8226 92.5005
R2890 VDD.n8233 VDD.n8232 92.5005
R2891 VDD.n8239 VDD.n8238 92.5005
R2892 VDD.n8243 VDD.n8242 92.5005
R2893 VDD.n8249 VDD.n8248 92.5005
R2894 VDD.n8254 VDD.n8253 92.5005
R2895 VDD.n8260 VDD.n8259 92.5005
R2896 VDD.n8266 VDD.n8265 92.5005
R2897 VDD.n8272 VDD.n8271 92.5005
R2898 VDD.n8278 VDD.n8277 92.5005
R2899 VDD.n8284 VDD.n8283 92.5005
R2900 VDD.n8290 VDD.n8289 92.5005
R2901 VDD.n8294 VDD.n8293 92.5005
R2902 VDD.n8300 VDD.n8299 92.5005
R2903 VDD.n8308 VDD.n8307 92.5005
R2904 VDD.n8314 VDD.n8313 92.5005
R2905 VDD.n8320 VDD.n8319 92.5005
R2906 VDD.n8326 VDD.n8325 92.5005
R2907 VDD.n8332 VDD.n8331 92.5005
R2908 VDD.n8338 VDD.n8337 92.5005
R2909 VDD.n8344 VDD.n8343 92.5005
R2910 VDD.n8348 VDD.n8347 92.5005
R2911 VDD.n8354 VDD.n8353 92.5005
R2912 VDD.n8359 VDD.n8358 92.5005
R2913 VDD.n8365 VDD.n8364 92.5005
R2914 VDD.n8371 VDD.n8370 92.5005
R2915 VDD.n8377 VDD.n8376 92.5005
R2916 VDD.n8383 VDD.n8382 92.5005
R2917 VDD.n8389 VDD.n8388 92.5005
R2918 VDD.n8395 VDD.n8394 92.5005
R2919 VDD.n8399 VDD.n8398 92.5005
R2920 VDD.n8405 VDD.n8404 92.5005
R2921 VDD.n8417 VDD.n8416 92.5005
R2922 VDD.n8416 VDD.n8415 92.5005
R2923 VDD.n8427 VDD.n8426 92.5005
R2924 VDD.n8426 VDD.n8425 92.5005
R2925 VDD.n8437 VDD.n8436 92.5005
R2926 VDD.n8436 VDD.n8435 92.5005
R2927 VDD.n8447 VDD.n8446 92.5005
R2928 VDD.n8446 VDD.n8445 92.5005
R2929 VDD.n8457 VDD.n8456 92.5005
R2930 VDD.n8456 VDD.n8455 92.5005
R2931 VDD.n8466 VDD.n8465 92.5005
R2932 VDD.n8465 VDD.n8464 92.5005
R2933 VDD.n8475 VDD.n8474 92.5005
R2934 VDD.n8474 VDD.n8473 92.5005
R2935 VDD.n8480 VDD.n8479 92.5005
R2936 VDD.n8479 VDD.n8478 92.5005
R2937 VDD.n8489 VDD.n8488 92.5005
R2938 VDD.n8488 VDD.n8487 92.5005
R2939 VDD.n8497 VDD.n8496 92.5005
R2940 VDD.n8496 VDD.n8495 92.5005
R2941 VDD.n8506 VDD.n8505 92.5005
R2942 VDD.n8505 VDD.n8504 92.5005
R2943 VDD.n8515 VDD.n8514 92.5005
R2944 VDD.n8514 VDD.n8513 92.5005
R2945 VDD.n8524 VDD.n8523 92.5005
R2946 VDD.n8523 VDD.n8522 92.5005
R2947 VDD.n8532 VDD.n8531 92.5005
R2948 VDD.n8531 VDD.n8530 92.5005
R2949 VDD.n8539 VDD.n8538 92.5005
R2950 VDD.n8570 VDD.n8569 92.5005
R2951 VDD.n8566 VDD.n8565 92.5005
R2952 VDD.n2671 VDD.n2670 92.5005
R2953 VDD.n3063 VDD.n3062 92.5005
R2954 VDD.n3061 VDD.n3060 92.5005
R2955 VDD.n3059 VDD.n3058 92.5005
R2956 VDD.n3057 VDD.n3056 92.5005
R2957 VDD.n3055 VDD.n3054 92.5005
R2958 VDD.n3053 VDD.n3052 92.5005
R2959 VDD.n3043 VDD.n3042 92.5005
R2960 VDD.n2635 VDD.n2634 92.5005
R2961 VDD.n2638 VDD.n2637 92.5005
R2962 VDD.n2640 VDD.n2639 92.5005
R2963 VDD.n2646 VDD.n2645 92.5005
R2964 VDD.n3046 VDD.n3045 92.5005
R2965 VDD.n3050 VDD.n3049 92.5005
R2966 VDD.n3048 VDD.n3047 92.5005
R2967 VDD.n2665 VDD.n2664 92.5005
R2968 VDD.n2667 VDD.n2666 92.5005
R2969 VDD.n2669 VDD.n2668 92.5005
R2970 VDD.n2910 VDD.n2909 92.5005
R2971 VDD.n2909 VDD.n2908 92.5005
R2972 VDD.n2877 VDD.n2876 92.5005
R2973 VDD.n2876 VDD.n2875 92.5005
R2974 VDD.n2880 VDD.n2879 92.5005
R2975 VDD.n2879 VDD.n2878 92.5005
R2976 VDD.n2883 VDD.n2882 92.5005
R2977 VDD.n2882 VDD.n2881 92.5005
R2978 VDD.n2886 VDD.n2885 92.5005
R2979 VDD.n2885 VDD.n2884 92.5005
R2980 VDD.n2889 VDD.n2888 92.5005
R2981 VDD.n2888 VDD.n2887 92.5005
R2982 VDD.n2892 VDD.n2891 92.5005
R2983 VDD.n2891 VDD.n2890 92.5005
R2984 VDD.n2895 VDD.n2894 92.5005
R2985 VDD.n2894 VDD.n2893 92.5005
R2986 VDD.n2898 VDD.n2897 92.5005
R2987 VDD.n2897 VDD.n2896 92.5005
R2988 VDD.n2901 VDD.n2900 92.5005
R2989 VDD.n2900 VDD.n2899 92.5005
R2990 VDD.n2904 VDD.n2903 92.5005
R2991 VDD.n2903 VDD.n2902 92.5005
R2992 VDD.n2907 VDD.n2906 92.5005
R2993 VDD.n2906 VDD.n2905 92.5005
R2994 VDD.n2874 VDD.n2873 92.5005
R2995 VDD.n2873 VDD.n2872 92.5005
R2996 VDD.n2871 VDD.n2870 92.5005
R2997 VDD.n2870 VDD.n2869 92.5005
R2998 VDD.n2868 VDD.n2867 92.5005
R2999 VDD.n2864 VDD.n2863 92.5005
R3000 VDD.n2862 VDD.n2861 92.5005
R3001 VDD.n2856 VDD.n2855 92.5005
R3002 VDD.n2855 VDD.n2854 92.5005
R3003 VDD.n2853 VDD.n2852 92.5005
R3004 VDD.n2852 VDD.n2851 92.5005
R3005 VDD.n2850 VDD.n2849 92.5005
R3006 VDD.n2849 VDD.n2848 92.5005
R3007 VDD.n2847 VDD.n2846 92.5005
R3008 VDD.n2846 VDD.n2845 92.5005
R3009 VDD.n2844 VDD.n2843 92.5005
R3010 VDD.n2843 VDD.n2842 92.5005
R3011 VDD.n2841 VDD.n2840 92.5005
R3012 VDD.n2840 VDD.n2839 92.5005
R3013 VDD.n2838 VDD.n2837 92.5005
R3014 VDD.n2837 VDD.n2836 92.5005
R3015 VDD.n2835 VDD.n2834 92.5005
R3016 VDD.n2834 VDD.n2833 92.5005
R3017 VDD.n2832 VDD.n2831 92.5005
R3018 VDD.n2831 VDD.n2830 92.5005
R3019 VDD.n2829 VDD.n2828 92.5005
R3020 VDD.n2828 VDD.n2827 92.5005
R3021 VDD.n2826 VDD.n2825 92.5005
R3022 VDD.n2825 VDD.n2824 92.5005
R3023 VDD.n2823 VDD.n2822 92.5005
R3024 VDD.n2822 VDD.n2821 92.5005
R3025 VDD.n2820 VDD.n2819 92.5005
R3026 VDD.n2819 VDD.n2818 92.5005
R3027 VDD.n3214 VDD.n3213 92.5005
R3028 VDD.n3213 VDD.n3212 92.5005
R3029 VDD.n3217 VDD.n3216 92.5005
R3030 VDD.n3216 VDD.n3215 92.5005
R3031 VDD.n3220 VDD.n3219 92.5005
R3032 VDD.n3219 VDD.n3218 92.5005
R3033 VDD.n3223 VDD.n3222 92.5005
R3034 VDD.n3222 VDD.n3221 92.5005
R3035 VDD.n3226 VDD.n3225 92.5005
R3036 VDD.n3225 VDD.n3224 92.5005
R3037 VDD.n3229 VDD.n3228 92.5005
R3038 VDD.n3228 VDD.n3227 92.5005
R3039 VDD.n3232 VDD.n3231 92.5005
R3040 VDD.n3231 VDD.n3230 92.5005
R3041 VDD.n3235 VDD.n3234 92.5005
R3042 VDD.n3234 VDD.n3233 92.5005
R3043 VDD.n3238 VDD.n3237 92.5005
R3044 VDD.n3237 VDD.n3236 92.5005
R3045 VDD.n3241 VDD.n3240 92.5005
R3046 VDD.n3240 VDD.n3239 92.5005
R3047 VDD.n3244 VDD.n3243 92.5005
R3048 VDD.n3243 VDD.n3242 92.5005
R3049 VDD.n3247 VDD.n3246 92.5005
R3050 VDD.n3246 VDD.n3245 92.5005
R3051 VDD.n3250 VDD.n3249 92.5005
R3052 VDD.n3249 VDD.n3248 92.5005
R3053 VDD.n3253 VDD.n3252 92.5005
R3054 VDD.n3252 VDD.n3251 92.5005
R3055 VDD.n3257 VDD.n3256 92.5005
R3056 VDD.n3256 VDD.n3255 92.5005
R3057 VDD.n2860 VDD.n2859 92.5005
R3058 VDD.n2859 VDD.n2858 92.5005
R3059 VDD.n3277 VDD.n3276 92.5005
R3060 VDD.n3276 VDD.n3275 92.5005
R3061 VDD.n3280 VDD.n3279 92.5005
R3062 VDD.n3279 VDD.n3278 92.5005
R3063 VDD.n3283 VDD.n3282 92.5005
R3064 VDD.n3282 VDD.n3281 92.5005
R3065 VDD.n3286 VDD.n3285 92.5005
R3066 VDD.n3285 VDD.n3284 92.5005
R3067 VDD.n3289 VDD.n3288 92.5005
R3068 VDD.n3288 VDD.n3287 92.5005
R3069 VDD.n3292 VDD.n3291 92.5005
R3070 VDD.n3291 VDD.n3290 92.5005
R3071 VDD.n3295 VDD.n3294 92.5005
R3072 VDD.n3294 VDD.n3293 92.5005
R3073 VDD.n3298 VDD.n3297 92.5005
R3074 VDD.n3297 VDD.n3296 92.5005
R3075 VDD.n3301 VDD.n3300 92.5005
R3076 VDD.n3300 VDD.n3299 92.5005
R3077 VDD.n3304 VDD.n3303 92.5005
R3078 VDD.n3303 VDD.n3302 92.5005
R3079 VDD.n3307 VDD.n3306 92.5005
R3080 VDD.n3306 VDD.n3305 92.5005
R3081 VDD.n3271 VDD.n3270 92.5005
R3082 VDD.n3270 VDD.n3269 92.5005
R3083 VDD.n3268 VDD.n3267 92.5005
R3084 VDD.n3267 VDD.n3266 92.5005
R3085 VDD.n3265 VDD.n3264 92.5005
R3086 VDD.n3261 VDD.n3260 92.5005
R3087 VDD.n3259 VDD.n3258 92.5005
R3088 VDD.n3274 VDD.n3273 92.5005
R3089 VDD.n3273 VDD.n3272 92.5005
R3090 VDD.n3309 VDD.n3308 92.5005
R3091 VDD.n3372 VDD.n3371 92.5005
R3092 VDD.n3365 VDD.n3364 92.5005
R3093 VDD.n3360 VDD.n3359 92.5005
R3094 VDD.n3355 VDD.n3354 92.5005
R3095 VDD.n3350 VDD.n3349 92.5005
R3096 VDD.n3345 VDD.n3344 92.5005
R3097 VDD.n3340 VDD.n3339 92.5005
R3098 VDD.n3338 VDD.n3337 92.5005
R3099 VDD.n3374 VDD.n3373 92.5005
R3100 VDD.n3385 VDD.n3384 92.5005
R3101 VDD.n3211 VDD.n3210 92.5005
R3102 VDD.n3171 VDD.n3170 92.5005
R3103 VDD.n3176 VDD.n3175 92.5005
R3104 VDD.n3181 VDD.n3180 92.5005
R3105 VDD.n3186 VDD.n3185 92.5005
R3106 VDD.n3192 VDD.n3191 92.5005
R3107 VDD.n3198 VDD.n3197 92.5005
R3108 VDD.n3196 VDD.n3195 92.5005
R3109 VDD.n3189 VDD.n3188 92.5005
R3110 VDD.n3184 VDD.n3183 92.5005
R3111 VDD.n3178 VDD.n3177 92.5005
R3112 VDD.n3174 VDD.n3173 92.5005
R3113 VDD.n3165 VDD.n3164 92.5005
R3114 VDD.n3168 VDD.n3167 92.5005
R3115 VDD.n3200 VDD.n3199 92.5005
R3116 VDD.n3205 VDD.n3204 92.5005
R3117 VDD.n3208 VDD.n3207 92.5005
R3118 VDD.n3066 VDD.n3065 92.5005
R3119 VDD.n3111 VDD.n3110 92.5005
R3120 VDD.n3114 VDD.n3113 92.5005
R3121 VDD.n3116 VDD.n3115 92.5005
R3122 VDD.n3120 VDD.n3119 92.5005
R3123 VDD.n3123 VDD.n3122 92.5005
R3124 VDD.n3122 VDD.n3121 92.5005
R3125 VDD.n3126 VDD.n3125 92.5005
R3126 VDD.n3125 VDD.n3124 92.5005
R3127 VDD.n3129 VDD.n3128 92.5005
R3128 VDD.n3128 VDD.n3127 92.5005
R3129 VDD.n3132 VDD.n3131 92.5005
R3130 VDD.n3131 VDD.n3130 92.5005
R3131 VDD.n3135 VDD.n3134 92.5005
R3132 VDD.n3134 VDD.n3133 92.5005
R3133 VDD.n3138 VDD.n3137 92.5005
R3134 VDD.n3137 VDD.n3136 92.5005
R3135 VDD.n3141 VDD.n3140 92.5005
R3136 VDD.n3140 VDD.n3139 92.5005
R3137 VDD.n3144 VDD.n3143 92.5005
R3138 VDD.n3143 VDD.n3142 92.5005
R3139 VDD.n3147 VDD.n3146 92.5005
R3140 VDD.n3146 VDD.n3145 92.5005
R3141 VDD.n3150 VDD.n3149 92.5005
R3142 VDD.n3149 VDD.n3148 92.5005
R3143 VDD.n3153 VDD.n3152 92.5005
R3144 VDD.n3152 VDD.n3151 92.5005
R3145 VDD.n3156 VDD.n3155 92.5005
R3146 VDD.n3155 VDD.n3154 92.5005
R3147 VDD.n3159 VDD.n3158 92.5005
R3148 VDD.n3158 VDD.n3157 92.5005
R3149 VDD.n3162 VDD.n3161 92.5005
R3150 VDD.n3161 VDD.n3160 92.5005
R3151 VDD.n2707 VDD.n2706 92.5005
R3152 VDD.n2706 VDD.n2705 92.5005
R3153 VDD.n2704 VDD.n2703 92.5005
R3154 VDD.n2703 VDD.n2702 92.5005
R3155 VDD.n2701 VDD.n2700 92.5005
R3156 VDD.n2700 VDD.n2699 92.5005
R3157 VDD.n2698 VDD.n2697 92.5005
R3158 VDD.n2697 VDD.n2696 92.5005
R3159 VDD.n2695 VDD.n2694 92.5005
R3160 VDD.n2694 VDD.n2693 92.5005
R3161 VDD.n2692 VDD.n2691 92.5005
R3162 VDD.n2691 VDD.n2690 92.5005
R3163 VDD.n2689 VDD.n2688 92.5005
R3164 VDD.n2688 VDD.n2687 92.5005
R3165 VDD.n2686 VDD.n2685 92.5005
R3166 VDD.n2685 VDD.n2684 92.5005
R3167 VDD.n2683 VDD.n2682 92.5005
R3168 VDD.n2682 VDD.n2681 92.5005
R3169 VDD.n2680 VDD.n2679 92.5005
R3170 VDD.n2679 VDD.n2678 92.5005
R3171 VDD.n2677 VDD.n2676 92.5005
R3172 VDD.n2676 VDD.n2675 92.5005
R3173 VDD.n2674 VDD.n2673 92.5005
R3174 VDD.n2673 VDD.n2672 92.5005
R3175 VDD.n3069 VDD.n3068 92.5005
R3176 VDD.n3068 VDD.n3067 92.5005
R3177 VDD.n3072 VDD.n3071 92.5005
R3178 VDD.n3071 VDD.n3070 92.5005
R3179 VDD.n3075 VDD.n3074 92.5005
R3180 VDD.n3074 VDD.n3073 92.5005
R3181 VDD.n3078 VDD.n3077 92.5005
R3182 VDD.n3077 VDD.n3076 92.5005
R3183 VDD.n3081 VDD.n3080 92.5005
R3184 VDD.n3080 VDD.n3079 92.5005
R3185 VDD.n3084 VDD.n3083 92.5005
R3186 VDD.n3083 VDD.n3082 92.5005
R3187 VDD.n3087 VDD.n3086 92.5005
R3188 VDD.n3086 VDD.n3085 92.5005
R3189 VDD.n3090 VDD.n3089 92.5005
R3190 VDD.n3089 VDD.n3088 92.5005
R3191 VDD.n3093 VDD.n3092 92.5005
R3192 VDD.n3092 VDD.n3091 92.5005
R3193 VDD.n3096 VDD.n3095 92.5005
R3194 VDD.n3095 VDD.n3094 92.5005
R3195 VDD.n3099 VDD.n3098 92.5005
R3196 VDD.n3098 VDD.n3097 92.5005
R3197 VDD.n3102 VDD.n3101 92.5005
R3198 VDD.n3101 VDD.n3100 92.5005
R3199 VDD.n3105 VDD.n3104 92.5005
R3200 VDD.n3104 VDD.n3103 92.5005
R3201 VDD.n3108 VDD.n3107 92.5005
R3202 VDD.n3107 VDD.n3106 92.5005
R3203 VDD.n2717 VDD.n2716 92.5005
R3204 VDD.n2710 VDD.n2709 92.5005
R3205 VDD.n2712 VDD.n2711 92.5005
R3206 VDD.n2768 VDD.n2767 92.5005
R3207 VDD.n2767 VDD.n2766 92.5005
R3208 VDD.n2765 VDD.n2764 92.5005
R3209 VDD.n2764 VDD.n2763 92.5005
R3210 VDD.n2762 VDD.n2761 92.5005
R3211 VDD.n2761 VDD.n2760 92.5005
R3212 VDD.n2759 VDD.n2758 92.5005
R3213 VDD.n2758 VDD.n2757 92.5005
R3214 VDD.n2756 VDD.n2755 92.5005
R3215 VDD.n2755 VDD.n2754 92.5005
R3216 VDD.n2753 VDD.n2752 92.5005
R3217 VDD.n2752 VDD.n2751 92.5005
R3218 VDD.n2750 VDD.n2749 92.5005
R3219 VDD.n2749 VDD.n2748 92.5005
R3220 VDD.n2747 VDD.n2746 92.5005
R3221 VDD.n2746 VDD.n2745 92.5005
R3222 VDD.n2744 VDD.n2743 92.5005
R3223 VDD.n2743 VDD.n2742 92.5005
R3224 VDD.n2741 VDD.n2740 92.5005
R3225 VDD.n2740 VDD.n2739 92.5005
R3226 VDD.n2738 VDD.n2737 92.5005
R3227 VDD.n2737 VDD.n2736 92.5005
R3228 VDD.n2735 VDD.n2734 92.5005
R3229 VDD.n2734 VDD.n2733 92.5005
R3230 VDD.n2732 VDD.n2731 92.5005
R3231 VDD.n2731 VDD.n2730 92.5005
R3232 VDD.n2729 VDD.n2728 92.5005
R3233 VDD.n2728 VDD.n2727 92.5005
R3234 VDD.n2726 VDD.n2725 92.5005
R3235 VDD.n2722 VDD.n2721 92.5005
R3236 VDD.n2719 VDD.n2718 92.5005
R3237 VDD.n2913 VDD.n2912 92.5005
R3238 VDD.n2930 VDD.n2929 92.5005
R3239 VDD.n2933 VDD.n2932 92.5005
R3240 VDD.n2938 VDD.n2937 92.5005
R3241 VDD.n2944 VDD.n2943 92.5005
R3242 VDD.n2949 VDD.n2948 92.5005
R3243 VDD.n2955 VDD.n2954 92.5005
R3244 VDD.n2960 VDD.n2959 92.5005
R3245 VDD.n2966 VDD.n2965 92.5005
R3246 VDD.n2969 VDD.n2968 92.5005
R3247 VDD.n2804 VDD.n2803 92.5005
R3248 VDD.n2799 VDD.n2798 92.5005
R3249 VDD.n2793 VDD.n2792 92.5005
R3250 VDD.n2788 VDD.n2787 92.5005
R3251 VDD.n2782 VDD.n2781 92.5005
R3252 VDD.n2777 VDD.n2776 92.5005
R3253 VDD.n2774 VDD.n2773 92.5005
R3254 VDD.n2771 VDD.n2770 92.5005
R3255 VDD.n2779 VDD.n2778 92.5005
R3256 VDD.n2785 VDD.n2784 92.5005
R3257 VDD.n2790 VDD.n2789 92.5005
R3258 VDD.n2796 VDD.n2795 92.5005
R3259 VDD.n2801 VDD.n2800 92.5005
R3260 VDD.n2810 VDD.n2809 92.5005
R3261 VDD.n2808 VDD.n2807 92.5005
R3262 VDD.n2812 VDD.n2811 92.5005
R3263 VDD.n2817 VDD.n2816 92.5005
R3264 VDD.n2972 VDD.n2971 92.5005
R3265 VDD.n2963 VDD.n2962 92.5005
R3266 VDD.n2935 VDD.n2934 92.5005
R3267 VDD.n2941 VDD.n2940 92.5005
R3268 VDD.n2946 VDD.n2945 92.5005
R3269 VDD.n2952 VDD.n2951 92.5005
R3270 VDD.n2957 VDD.n2956 92.5005
R3271 VDD.n3376 VDD.n3375 92.5005
R3272 VDD.n3378 VDD.n3377 92.5005
R3273 VDD.n3382 VDD.n3381 92.5005
R3274 VDD.n3381 VDD.n3380 92.5005
R3275 VDD.n3362 VDD.n3361 92.5005
R3276 VDD.n3358 VDD.n3357 92.5005
R3277 VDD.n3352 VDD.n3351 92.5005
R3278 VDD.n3348 VDD.n3347 92.5005
R3279 VDD.n3342 VDD.n3341 92.5005
R3280 VDD.n3369 VDD.n3368 92.5005
R3281 VDD.n3315 VDD.n3314 92.5005
R3282 VDD.n3311 VDD.n3310 92.5005
R3283 VDD.n3388 VDD.n3387 92.5005
R3284 VDD.n3391 VDD.n3390 92.5005
R3285 VDD.n3394 VDD.n3393 92.5005
R3286 VDD.n3399 VDD.n3398 92.5005
R3287 VDD.n3334 VDD.n3333 92.5005
R3288 VDD.n3332 VDD.n3331 92.5005
R3289 VDD.n3330 VDD.n3329 92.5005
R3290 VDD.n3328 VDD.n3327 92.5005
R3291 VDD.n3325 VDD.n3324 92.5005
R3292 VDD.n3323 VDD.n3322 92.5005
R3293 VDD.n3321 VDD.n3320 92.5005
R3294 VDD.n3319 VDD.n3318 92.5005
R3295 VDD.n3317 VDD.n3316 92.5005
R3296 VDD.n2915 VDD.n2914 92.5005
R3297 VDD.n2921 VDD.n2920 92.5005
R3298 VDD.n2923 VDD.n2922 92.5005
R3299 VDD.n2925 VDD.n2924 92.5005
R3300 VDD.n2927 VDD.n2926 92.5005
R3301 VDD.n2918 VDD.n2917 92.5005
R3302 VDD.n2648 VDD.n2647 92.5005
R3303 VDD.n2651 VDD.n2650 92.5005
R3304 VDD.n2654 VDD.n2653 92.5005
R3305 VDD.n2657 VDD.n2656 92.5005
R3306 VDD.n2663 VDD.n2662 92.5005
R3307 VDD.n2976 VDD.n2975 92.5005
R3308 VDD.n2975 VDD.n2974 92.5005
R3309 VDD.n2982 VDD.n2981 92.5005
R3310 VDD.n2981 VDD.n2980 92.5005
R3311 VDD.n2988 VDD.n2987 92.5005
R3312 VDD.n2987 VDD.n2986 92.5005
R3313 VDD.n2994 VDD.n2993 92.5005
R3314 VDD.n2993 VDD.n2992 92.5005
R3315 VDD.n3007 VDD.n3006 92.5005
R3316 VDD.n3006 VDD.n3005 92.5005
R3317 VDD.n3011 VDD.n3010 92.5005
R3318 VDD.n3010 VDD.n3009 92.5005
R3319 VDD.n3016 VDD.n3015 92.5005
R3320 VDD.n3015 VDD.n3014 92.5005
R3321 VDD.n3037 VDD.n3036 92.5005
R3322 VDD.n3036 VDD.n3035 92.5005
R3323 VDD.n3031 VDD.n3030 92.5005
R3324 VDD.n3030 VDD.n3029 92.5005
R3325 VDD.n3025 VDD.n3024 92.5005
R3326 VDD.n3024 VDD.n3023 92.5005
R3327 VDD.n3409 VDD.n3408 92.5005
R3328 VDD.n3408 VDD.n3407 92.5005
R3329 VDD.n2985 VDD.n2984 92.5005
R3330 VDD.n2984 VDD.n2983 92.5005
R3331 VDD.n2991 VDD.n2990 92.5005
R3332 VDD.n2990 VDD.n2989 92.5005
R3333 VDD.n2997 VDD.n2996 92.5005
R3334 VDD.n2996 VDD.n2995 92.5005
R3335 VDD.n3000 VDD.n2999 92.5005
R3336 VDD.n2999 VDD.n2998 92.5005
R3337 VDD.n3004 VDD.n3003 92.5005
R3338 VDD.n3003 VDD.n3002 92.5005
R3339 VDD.n3019 VDD.n3018 92.5005
R3340 VDD.n3018 VDD.n3017 92.5005
R3341 VDD.n3034 VDD.n3033 92.5005
R3342 VDD.n3033 VDD.n3032 92.5005
R3343 VDD.n3028 VDD.n3027 92.5005
R3344 VDD.n3027 VDD.n3026 92.5005
R3345 VDD.n3022 VDD.n3021 92.5005
R3346 VDD.n3021 VDD.n3020 92.5005
R3347 VDD.n3402 VDD.n3401 92.5005
R3348 VDD.n3401 VDD.n3400 92.5005
R3349 VDD.n3406 VDD.n3405 92.5005
R3350 VDD.n3405 VDD.n3404 92.5005
R3351 VDD.n2979 VDD.n2978 92.5005
R3352 VDD.n2978 VDD.n2977 92.5005
R3353 VDD.n2217 VDD.n2214 92.5005
R3354 VDD.n2373 VDD.n2217 92.5005
R3355 VDD.n2538 VDD.n1805 92.5005
R3356 VDD.n1925 VDD.n1805 92.5005
R3357 VDD.n2540 VDD.n2539 92.5005
R3358 VDD.n2541 VDD.n2540 92.5005
R3359 VDD.n1806 VDD.n1804 92.5005
R3360 VDD.n1804 VDD.n1796 92.5005
R3361 VDD.n2263 VDD.n2262 92.5005
R3362 VDD.n2263 VDD.n1795 92.5005
R3363 VDD.n2264 VDD.n2261 92.5005
R3364 VDD.n2264 VDD.n1788 92.5005
R3365 VDD.n2266 VDD.n2265 92.5005
R3366 VDD.n2265 VDD.n1787 92.5005
R3367 VDD.n2279 VDD.n2259 92.5005
R3368 VDD.n2278 VDD.n2277 92.5005
R3369 VDD.n2276 VDD.n2275 92.5005
R3370 VDD.n2274 VDD.n2273 92.5005
R3371 VDD.n2272 VDD.n2271 92.5005
R3372 VDD.n2281 VDD.n2280 92.5005
R3373 VDD.n2243 VDD.n2242 92.5005
R3374 VDD.n2256 VDD.n2243 92.5005
R3375 VDD.n2361 VDD.n2360 92.5005
R3376 VDD.n2360 VDD.n2359 92.5005
R3377 VDD.n2362 VDD.n2240 92.5005
R3378 VDD.n2244 VDD.n2240 92.5005
R3379 VDD.n2364 VDD.n2363 92.5005
R3380 VDD.n2365 VDD.n2364 92.5005
R3381 VDD.n2241 VDD.n2239 92.5005
R3382 VDD.n2239 VDD.n2231 92.5005
R3383 VDD.n2404 VDD.n2001 92.5005
R3384 VDD.n2001 VDD.n2000 92.5005
R3385 VDD.n2427 VDD.n2426 92.5005
R3386 VDD.n2426 VDD.n2425 92.5005
R3387 VDD.n1991 VDD.n1990 92.5005
R3388 VDD.n2424 VDD.n1991 92.5005
R3389 VDD.n2422 VDD.n2421 92.5005
R3390 VDD.n2423 VDD.n2422 92.5005
R3391 VDD.n2420 VDD.n1993 92.5005
R3392 VDD.n1993 VDD.n1992 92.5005
R3393 VDD.n2419 VDD.n2418 92.5005
R3394 VDD.n2418 VDD.n2417 92.5005
R3395 VDD.n1995 VDD.n1994 92.5005
R3396 VDD.n2416 VDD.n1995 92.5005
R3397 VDD.n2414 VDD.n2413 92.5005
R3398 VDD.n2415 VDD.n2414 92.5005
R3399 VDD.n2412 VDD.n1997 92.5005
R3400 VDD.n1997 VDD.n1996 92.5005
R3401 VDD.n2411 VDD.n2410 92.5005
R3402 VDD.n2410 VDD.n2409 92.5005
R3403 VDD.n1999 VDD.n1998 92.5005
R3404 VDD.n2408 VDD.n1999 92.5005
R3405 VDD.n2406 VDD.n2405 92.5005
R3406 VDD.n2407 VDD.n2406 92.5005
R3407 VDD.n2428 VDD.n1988 92.5005
R3408 VDD.n1988 VDD.n1987 92.5005
R3409 VDD.n2431 VDD.n2430 92.5005
R3410 VDD.n2432 VDD.n2431 92.5005
R3411 VDD.n2429 VDD.n1989 92.5005
R3412 VDD.n1985 VDD.n1984 92.5005
R3413 VDD.n2436 VDD.n2435 92.5005
R3414 VDD.n2435 VDD.n2434 92.5005
R3415 VDD.n2439 VDD.n2438 92.5005
R3416 VDD.n2440 VDD.n2439 92.5005
R3417 VDD.n1981 VDD.n1980 92.5005
R3418 VDD.n2441 VDD.n1981 92.5005
R3419 VDD.n2444 VDD.n2443 92.5005
R3420 VDD.n2443 VDD.n2442 92.5005
R3421 VDD.n2445 VDD.n1979 92.5005
R3422 VDD.n1979 VDD.n1978 92.5005
R3423 VDD.n2447 VDD.n2446 92.5005
R3424 VDD.n2448 VDD.n2447 92.5005
R3425 VDD.n1977 VDD.n1976 92.5005
R3426 VDD.n2449 VDD.n1977 92.5005
R3427 VDD.n2452 VDD.n2451 92.5005
R3428 VDD.n2451 VDD.n2450 92.5005
R3429 VDD.n2453 VDD.n1975 92.5005
R3430 VDD.n1975 VDD.n1974 92.5005
R3431 VDD.n2455 VDD.n2454 92.5005
R3432 VDD.n2456 VDD.n2455 92.5005
R3433 VDD.n1973 VDD.n1972 92.5005
R3434 VDD.n2457 VDD.n1973 92.5005
R3435 VDD.n2460 VDD.n2459 92.5005
R3436 VDD.n2459 VDD.n2458 92.5005
R3437 VDD.n2461 VDD.n1971 92.5005
R3438 VDD.n1971 VDD.n1970 92.5005
R3439 VDD.n2463 VDD.n2462 92.5005
R3440 VDD.n2464 VDD.n2463 92.5005
R3441 VDD.n1969 VDD.n1968 92.5005
R3442 VDD.n2465 VDD.n1969 92.5005
R3443 VDD.n2468 VDD.n2467 92.5005
R3444 VDD.n2467 VDD.n2466 92.5005
R3445 VDD.n2469 VDD.n1967 92.5005
R3446 VDD.n1967 VDD.n1966 92.5005
R3447 VDD.n2471 VDD.n2470 92.5005
R3448 VDD.n2472 VDD.n2471 92.5005
R3449 VDD.n1965 VDD.n1964 92.5005
R3450 VDD.n2473 VDD.n1965 92.5005
R3451 VDD.n2476 VDD.n2475 92.5005
R3452 VDD.n2475 VDD.n2474 92.5005
R3453 VDD.n2477 VDD.n1963 92.5005
R3454 VDD.n1963 VDD.n1962 92.5005
R3455 VDD.n2479 VDD.n2478 92.5005
R3456 VDD.n2480 VDD.n2479 92.5005
R3457 VDD.n1961 VDD.n1960 92.5005
R3458 VDD.n2481 VDD.n1961 92.5005
R3459 VDD.n2484 VDD.n2483 92.5005
R3460 VDD.n2483 VDD.n2482 92.5005
R3461 VDD.n2485 VDD.n1959 92.5005
R3462 VDD.n1959 VDD.n1958 92.5005
R3463 VDD.n2487 VDD.n2486 92.5005
R3464 VDD.n2488 VDD.n2487 92.5005
R3465 VDD.n1957 VDD.n1956 92.5005
R3466 VDD.n2489 VDD.n1957 92.5005
R3467 VDD.n2494 VDD.n2493 92.5005
R3468 VDD.n2493 VDD.n2492 92.5005
R3469 VDD.n2495 VDD.n1955 92.5005
R3470 VDD.n2491 VDD.n1955 92.5005
R3471 VDD.n2437 VDD.n1983 92.5005
R3472 VDD.n1983 VDD.n1982 92.5005
R3473 VDD.n2509 VDD.n2508 92.5005
R3474 VDD.n2508 VDD.n2507 92.5005
R3475 VDD.n2510 VDD.n1948 92.5005
R3476 VDD.n1948 VDD.n1947 92.5005
R3477 VDD.n2512 VDD.n2511 92.5005
R3478 VDD.n2513 VDD.n2512 92.5005
R3479 VDD.n1946 VDD.n1945 92.5005
R3480 VDD.n2514 VDD.n1946 92.5005
R3481 VDD.n2517 VDD.n2516 92.5005
R3482 VDD.n2516 VDD.n2515 92.5005
R3483 VDD.n2518 VDD.n1944 92.5005
R3484 VDD.n1944 VDD.n1943 92.5005
R3485 VDD.n2520 VDD.n2519 92.5005
R3486 VDD.n2521 VDD.n2520 92.5005
R3487 VDD.n1942 VDD.n1941 92.5005
R3488 VDD.n2522 VDD.n1942 92.5005
R3489 VDD.n2525 VDD.n2524 92.5005
R3490 VDD.n2524 VDD.n2523 92.5005
R3491 VDD.n2526 VDD.n1817 92.5005
R3492 VDD.n1817 VDD.n1815 92.5005
R3493 VDD.n2528 VDD.n2527 92.5005
R3494 VDD.n2529 VDD.n2528 92.5005
R3495 VDD.n2504 VDD.n2503 92.5005
R3496 VDD.n2505 VDD.n2504 92.5005
R3497 VDD.n2502 VDD.n1952 92.5005
R3498 VDD.n1952 VDD.n1951 92.5005
R3499 VDD.n2501 VDD.n2500 92.5005
R3500 VDD.n2498 VDD.n1953 92.5005
R3501 VDD.n2497 VDD.n2496 92.5005
R3502 VDD.n2497 VDD.n1954 92.5005
R3503 VDD.n1950 VDD.n1949 92.5005
R3504 VDD.n2506 VDD.n1950 92.5005
R3505 VDD.n1940 VDD.n1816 92.5005
R3506 VDD.n1872 VDD.n1871 92.5005
R3507 VDD.n1869 VDD.n1841 92.5005
R3508 VDD.n1847 VDD.n1842 92.5005
R3509 VDD.n1864 VDD.n1863 92.5005
R3510 VDD.n1861 VDD.n1860 92.5005
R3511 VDD.n1855 VDD.n1848 92.5005
R3512 VDD.n1853 VDD.n1852 92.5005
R3513 VDD.n1851 VDD.n1818 92.5005
R3514 VDD.n1874 VDD.n1826 92.5005
R3515 VDD.n1876 VDD.n1825 92.5005
R3516 VDD.n1901 VDD.n1900 92.5005
R3517 VDD.n1834 VDD.n1808 92.5005
R3518 VDD.n1920 VDD.n1919 92.5005
R3519 VDD.n1917 VDD.n1916 92.5005
R3520 VDD.n1913 VDD.n1835 92.5005
R3521 VDD.n1910 VDD.n1909 92.5005
R3522 VDD.n1908 VDD.n1907 92.5005
R3523 VDD.n1837 VDD.n1836 92.5005
R3524 VDD.n1912 VDD.n1911 92.5005
R3525 VDD.n1915 VDD.n1914 92.5005
R3526 VDD.n1833 VDD.n1832 92.5005
R3527 VDD.n1922 VDD.n1921 92.5005
R3528 VDD.n2533 VDD.n1807 92.5005
R3529 VDD.n2536 VDD.n2535 92.5005
R3530 VDD.n1906 VDD.n1828 92.5005
R3531 VDD.n1924 VDD.n1828 92.5005
R3532 VDD.n1905 VDD.n1904 92.5005
R3533 VDD.n1903 VDD.n1840 92.5005
R3534 VDD.n2119 VDD.n2118 92.5005
R3535 VDD.n2116 VDD.n2069 92.5005
R3536 VDD.n2115 VDD.n2114 92.5005
R3537 VDD.n2113 VDD.n2070 92.5005
R3538 VDD.n2111 VDD.n2110 92.5005
R3539 VDD.n2109 VDD.n2073 92.5005
R3540 VDD.n2076 VDD.n2073 92.5005
R3541 VDD.n2108 VDD.n2107 92.5005
R3542 VDD.n2107 VDD.n2106 92.5005
R3543 VDD.n2075 VDD.n2074 92.5005
R3544 VDD.n2105 VDD.n2075 92.5005
R3545 VDD.n2103 VDD.n2102 92.5005
R3546 VDD.n2104 VDD.n2103 92.5005
R3547 VDD.n2101 VDD.n2078 92.5005
R3548 VDD.n2078 VDD.n2077 92.5005
R3549 VDD.n2100 VDD.n2099 92.5005
R3550 VDD.n2099 VDD.n2098 92.5005
R3551 VDD.n2080 VDD.n2079 92.5005
R3552 VDD.n2097 VDD.n2080 92.5005
R3553 VDD.n2095 VDD.n2094 92.5005
R3554 VDD.n2096 VDD.n2095 92.5005
R3555 VDD.n2093 VDD.n2082 92.5005
R3556 VDD.n2082 VDD.n2081 92.5005
R3557 VDD.n2092 VDD.n2091 92.5005
R3558 VDD.n2091 VDD.n2090 92.5005
R3559 VDD.n2084 VDD.n2083 92.5005
R3560 VDD.n2089 VDD.n2084 92.5005
R3561 VDD.n2087 VDD.n2086 92.5005
R3562 VDD.n2088 VDD.n2087 92.5005
R3563 VDD.n2085 VDD.n1811 92.5005
R3564 VDD.n1813 VDD.n1811 92.5005
R3565 VDD.n2532 VDD.n1812 92.5005
R3566 VDD.n2532 VDD.n2531 92.5005
R3567 VDD.n2171 VDD.n2170 92.5005
R3568 VDD.n2170 VDD.n2169 92.5005
R3569 VDD.n2043 VDD.n2042 92.5005
R3570 VDD.n2168 VDD.n2043 92.5005
R3571 VDD.n2166 VDD.n2165 92.5005
R3572 VDD.n2167 VDD.n2166 92.5005
R3573 VDD.n2164 VDD.n2045 92.5005
R3574 VDD.n2045 VDD.n2044 92.5005
R3575 VDD.n2163 VDD.n2162 92.5005
R3576 VDD.n2162 VDD.n2161 92.5005
R3577 VDD.n2047 VDD.n2046 92.5005
R3578 VDD.n2160 VDD.n2047 92.5005
R3579 VDD.n2158 VDD.n2157 92.5005
R3580 VDD.n2159 VDD.n2158 92.5005
R3581 VDD.n2156 VDD.n2049 92.5005
R3582 VDD.n2049 VDD.n2048 92.5005
R3583 VDD.n2155 VDD.n2154 92.5005
R3584 VDD.n2154 VDD.n2153 92.5005
R3585 VDD.n2051 VDD.n2050 92.5005
R3586 VDD.n2152 VDD.n2051 92.5005
R3587 VDD.n2150 VDD.n2149 92.5005
R3588 VDD.n2151 VDD.n2150 92.5005
R3589 VDD.n2148 VDD.n2053 92.5005
R3590 VDD.n2053 VDD.n2052 92.5005
R3591 VDD.n2147 VDD.n2146 92.5005
R3592 VDD.n2146 VDD.n2145 92.5005
R3593 VDD.n2055 VDD.n2054 92.5005
R3594 VDD.n2144 VDD.n2055 92.5005
R3595 VDD.n2142 VDD.n2141 92.5005
R3596 VDD.n2143 VDD.n2142 92.5005
R3597 VDD.n2140 VDD.n2057 92.5005
R3598 VDD.n2057 VDD.n2056 92.5005
R3599 VDD.n2139 VDD.n2138 92.5005
R3600 VDD.n2138 VDD.n2137 92.5005
R3601 VDD.n2059 VDD.n2058 92.5005
R3602 VDD.n2136 VDD.n2059 92.5005
R3603 VDD.n2134 VDD.n2133 92.5005
R3604 VDD.n2135 VDD.n2134 92.5005
R3605 VDD.n2132 VDD.n2061 92.5005
R3606 VDD.n2061 VDD.n2060 92.5005
R3607 VDD.n2131 VDD.n2130 92.5005
R3608 VDD.n2130 VDD.n2129 92.5005
R3609 VDD.n2063 VDD.n2062 92.5005
R3610 VDD.n2128 VDD.n2063 92.5005
R3611 VDD.n2126 VDD.n2125 92.5005
R3612 VDD.n2127 VDD.n2126 92.5005
R3613 VDD.n2124 VDD.n2065 92.5005
R3614 VDD.n2065 VDD.n2064 92.5005
R3615 VDD.n2123 VDD.n2122 92.5005
R3616 VDD.n2122 VDD.n2121 92.5005
R3617 VDD.n2067 VDD.n2066 92.5005
R3618 VDD.n2120 VDD.n2067 92.5005
R3619 VDD.n2179 VDD.n2040 92.5005
R3620 VDD.n2183 VDD.n2182 92.5005
R3621 VDD.n2041 VDD.n2039 92.5005
R3622 VDD.n2213 VDD.n2023 92.5005
R3623 VDD.n2209 VDD.n2023 92.5005
R3624 VDD.n2212 VDD.n2211 92.5005
R3625 VDD.n2211 VDD.n2210 92.5005
R3626 VDD.n2025 VDD.n2024 92.5005
R3627 VDD.n2208 VDD.n2025 92.5005
R3628 VDD.n2206 VDD.n2205 92.5005
R3629 VDD.n2207 VDD.n2206 92.5005
R3630 VDD.n2204 VDD.n2027 92.5005
R3631 VDD.n2027 VDD.n2026 92.5005
R3632 VDD.n2203 VDD.n2202 92.5005
R3633 VDD.n2202 VDD.n2201 92.5005
R3634 VDD.n2029 VDD.n2028 92.5005
R3635 VDD.n2200 VDD.n2029 92.5005
R3636 VDD.n2198 VDD.n2197 92.5005
R3637 VDD.n2199 VDD.n2198 92.5005
R3638 VDD.n2196 VDD.n2031 92.5005
R3639 VDD.n2031 VDD.n2030 92.5005
R3640 VDD.n2195 VDD.n2194 92.5005
R3641 VDD.n2194 VDD.n2193 92.5005
R3642 VDD.n2033 VDD.n2032 92.5005
R3643 VDD.n2192 VDD.n2033 92.5005
R3644 VDD.n2190 VDD.n2189 92.5005
R3645 VDD.n2191 VDD.n2190 92.5005
R3646 VDD.n2188 VDD.n2035 92.5005
R3647 VDD.n2035 VDD.n2034 92.5005
R3648 VDD.n2187 VDD.n2186 92.5005
R3649 VDD.n2186 VDD.n2185 92.5005
R3650 VDD.n2037 VDD.n2036 92.5005
R3651 VDD.n2175 VDD.n2172 92.5005
R3652 VDD.n2178 VDD.n2177 92.5005
R3653 VDD.n2403 VDD.n2402 92.5005
R3654 VDD.n2320 VDD.n2003 92.5005
R3655 VDD.n2322 VDD.n2321 92.5005
R3656 VDD.n2319 VDD.n2318 92.5005
R3657 VDD.n2289 VDD.n2288 92.5005
R3658 VDD.n2313 VDD.n2312 92.5005
R3659 VDD.n2291 VDD.n2290 92.5005
R3660 VDD.n2307 VDD.n2306 92.5005
R3661 VDD.n2303 VDD.n2302 92.5005
R3662 VDD.n2301 VDD.n2300 92.5005
R3663 VDD.n2378 VDD.n2377 92.5005
R3664 VDD.n2382 VDD.n2381 92.5005
R3665 VDD.n2385 VDD.n2384 92.5005
R3666 VDD.n2227 VDD.n2226 92.5005
R3667 VDD.n2216 VDD.n2215 92.5005
R3668 VDD.n2394 VDD.n2393 92.5005
R3669 VDD.n2395 VDD.n2022 92.5005
R3670 VDD.n2398 VDD.n2397 92.5005
R3671 VDD.n2392 VDD.n2391 92.5005
R3672 VDD.n2225 VDD.n2218 92.5005
R3673 VDD.n2387 VDD.n2386 92.5005
R3674 VDD.n2383 VDD.n2224 92.5005
R3675 VDD.n2380 VDD.n2379 92.5005
R3676 VDD.n2228 VDD.n2015 92.5005
R3677 VDD.n2400 VDD.n2015 92.5005
R3678 VDD.n2376 VDD.n2375 92.5005
R3679 VDD.n2295 VDD.n2294 92.5005
R3680 VDD.n2297 VDD.n2296 92.5005
R3681 VDD.n2299 VDD.n2298 92.5005
R3682 VDD.n2305 VDD.n2304 92.5005
R3683 VDD.n2324 VDD.n2323 92.5005
R3684 VDD.n2317 VDD.n2316 92.5005
R3685 VDD.n2315 VDD.n2314 92.5005
R3686 VDD.n2311 VDD.n2310 92.5005
R3687 VDD.n2309 VDD.n2308 92.5005
R3688 VDD.n1932 VDD.n1931 92.5005
R3689 VDD.n1823 VDD.n1822 92.5005
R3690 VDD.n1935 VDD.n1934 92.5005
R3691 VDD.n1936 VDD.n1935 92.5005
R3692 VDD.n1868 VDD.n1867 92.5005
R3693 VDD.n1866 VDD.n1865 92.5005
R3694 VDD.n1856 VDD.n1845 92.5005
R3695 VDD.n1859 VDD.n1858 92.5005
R3696 VDD.n1854 VDD.n1821 92.5005
R3697 VDD.n1870 VDD.n1824 92.5005
R3698 VDD.n1882 VDD.n1881 92.5005
R3699 VDD.n1884 VDD.n1880 92.5005
R3700 VDD.n1887 VDD.n1886 92.5005
R3701 VDD.n1889 VDD.n1888 92.5005
R3702 VDD.n1891 VDD.n1878 92.5005
R3703 VDD.n1894 VDD.n1893 92.5005
R3704 VDD.n1938 VDD.n1937 92.5005
R3705 VDD.n1937 VDD.n1936 92.5005
R3706 VDD.n1820 VDD.n1819 92.5005
R3707 VDD.n1822 VDD.n1820 92.5005
R3708 VDD.n1930 VDD.n1929 92.5005
R3709 VDD.n1931 VDD.n1930 92.5005
R3710 VDD.n1928 VDD.n1927 92.5005
R3711 VDD.n1927 VDD.n1926 92.5005
R3712 VDD.n2549 VDD.n2548 92.5005
R3713 VDD.n2548 VDD.n2547 92.5005
R3714 VDD.n2550 VDD.n1790 92.5005
R3715 VDD.n1794 VDD.n1790 92.5005
R3716 VDD.n2552 VDD.n2551 92.5005
R3717 VDD.n2553 VDD.n2552 92.5005
R3718 VDD.n1791 VDD.n1789 92.5005
R3719 VDD.n2285 VDD.n1789 92.5005
R3720 VDD.n2349 VDD.n2287 92.5005
R3721 VDD.n2287 VDD.n2286 92.5005
R3722 VDD.n2351 VDD.n2350 92.5005
R3723 VDD.n2352 VDD.n2351 92.5005
R3724 VDD.n2331 VDD.n2330 92.5005
R3725 VDD.n2330 VDD.n2238 92.5005
R3726 VDD.n2329 VDD.n2328 92.5005
R3727 VDD.n2329 VDD.n2237 92.5005
R3728 VDD.n2327 VDD.n2232 92.5005
R3729 VDD.n2372 VDD.n2232 92.5005
R3730 VDD.n2326 VDD.n2325 92.5005
R3731 VDD.n2325 VDD.n2219 92.5005
R3732 VDD.n2347 VDD.n2346 92.5005
R3733 VDD.n2344 VDD.n2332 92.5005
R3734 VDD.n2342 VDD.n2341 92.5005
R3735 VDD.n2340 VDD.n2339 92.5005
R3736 VDD.n2337 VDD.n2334 92.5005
R3737 VDD.n2335 VDD.n2248 92.5005
R3738 VDD.n2292 VDD.n2233 92.5005
R3739 VDD.n2233 VDD.n2219 92.5005
R3740 VDD.n2371 VDD.n2370 92.5005
R3741 VDD.n2372 VDD.n2371 92.5005
R3742 VDD.n2368 VDD.n2234 92.5005
R3743 VDD.n2237 VDD.n2234 92.5005
R3744 VDD.n2250 VDD.n2235 92.5005
R3745 VDD.n2250 VDD.n2238 92.5005
R3746 VDD.n2354 VDD.n2353 92.5005
R3747 VDD.n2353 VDD.n2352 92.5005
R3748 VDD.n2255 VDD.n2254 92.5005
R3749 VDD.n2286 VDD.n2255 92.5005
R3750 VDD.n2253 VDD.n1785 92.5005
R3751 VDD.n2285 VDD.n1785 92.5005
R3752 VDD.n2555 VDD.n2554 92.5005
R3753 VDD.n2554 VDD.n2553 92.5005
R3754 VDD.n1798 VDD.n1786 92.5005
R3755 VDD.n1794 VDD.n1786 92.5005
R3756 VDD.n2546 VDD.n2545 92.5005
R3757 VDD.n2547 VDD.n2546 92.5005
R3758 VDD.n1897 VDD.n1827 92.5005
R3759 VDD.n1926 VDD.n1827 92.5005
R3760 VDD.n2369 VDD.n2229 92.5005
R3761 VDD.n2231 VDD.n2229 92.5005
R3762 VDD.n2367 VDD.n2366 92.5005
R3763 VDD.n2366 VDD.n2365 92.5005
R3764 VDD.n2247 VDD.n2236 92.5005
R3765 VDD.n2244 VDD.n2236 92.5005
R3766 VDD.n2358 VDD.n2357 92.5005
R3767 VDD.n2359 VDD.n2358 92.5005
R3768 VDD.n2355 VDD.n2246 92.5005
R3769 VDD.n2256 VDD.n2246 92.5005
R3770 VDD.n2269 VDD.n1783 92.5005
R3771 VDD.n2269 VDD.n1787 92.5005
R3772 VDD.n2268 VDD.n1784 92.5005
R3773 VDD.n2268 VDD.n1788 92.5005
R3774 VDD.n1801 VDD.n1799 92.5005
R3775 VDD.n1801 VDD.n1795 92.5005
R3776 VDD.n2544 VDD.n2543 92.5005
R3777 VDD.n2543 VDD.n1796 92.5005
R3778 VDD.n2542 VDD.n1800 92.5005
R3779 VDD.n2542 VDD.n2541 92.5005
R3780 VDD.n1896 VDD.n1802 92.5005
R3781 VDD.n1925 VDD.n1802 92.5005
R3782 VDD.n2374 VDD.n2230 92.5005
R3783 VDD.n2374 VDD.n2373 92.5005
R3784 VDD.n1363 VDD.n1360 92.5005
R3785 VDD.n1519 VDD.n1363 92.5005
R3786 VDD.n1684 VDD.n951 92.5005
R3787 VDD.n1071 VDD.n951 92.5005
R3788 VDD.n1686 VDD.n1685 92.5005
R3789 VDD.n1687 VDD.n1686 92.5005
R3790 VDD.n952 VDD.n950 92.5005
R3791 VDD.n950 VDD.n942 92.5005
R3792 VDD.n1409 VDD.n1408 92.5005
R3793 VDD.n1409 VDD.n941 92.5005
R3794 VDD.n1410 VDD.n1407 92.5005
R3795 VDD.n1410 VDD.n934 92.5005
R3796 VDD.n1412 VDD.n1411 92.5005
R3797 VDD.n1411 VDD.n933 92.5005
R3798 VDD.n1425 VDD.n1405 92.5005
R3799 VDD.n1424 VDD.n1423 92.5005
R3800 VDD.n1422 VDD.n1421 92.5005
R3801 VDD.n1420 VDD.n1419 92.5005
R3802 VDD.n1418 VDD.n1417 92.5005
R3803 VDD.n1427 VDD.n1426 92.5005
R3804 VDD.n1389 VDD.n1388 92.5005
R3805 VDD.n1402 VDD.n1389 92.5005
R3806 VDD.n1507 VDD.n1506 92.5005
R3807 VDD.n1506 VDD.n1505 92.5005
R3808 VDD.n1508 VDD.n1386 92.5005
R3809 VDD.n1390 VDD.n1386 92.5005
R3810 VDD.n1510 VDD.n1509 92.5005
R3811 VDD.n1511 VDD.n1510 92.5005
R3812 VDD.n1387 VDD.n1385 92.5005
R3813 VDD.n1385 VDD.n1377 92.5005
R3814 VDD.n1550 VDD.n1147 92.5005
R3815 VDD.n1147 VDD.n1146 92.5005
R3816 VDD.n1573 VDD.n1572 92.5005
R3817 VDD.n1572 VDD.n1571 92.5005
R3818 VDD.n1137 VDD.n1136 92.5005
R3819 VDD.n1570 VDD.n1137 92.5005
R3820 VDD.n1568 VDD.n1567 92.5005
R3821 VDD.n1569 VDD.n1568 92.5005
R3822 VDD.n1566 VDD.n1139 92.5005
R3823 VDD.n1139 VDD.n1138 92.5005
R3824 VDD.n1565 VDD.n1564 92.5005
R3825 VDD.n1564 VDD.n1563 92.5005
R3826 VDD.n1141 VDD.n1140 92.5005
R3827 VDD.n1562 VDD.n1141 92.5005
R3828 VDD.n1560 VDD.n1559 92.5005
R3829 VDD.n1561 VDD.n1560 92.5005
R3830 VDD.n1558 VDD.n1143 92.5005
R3831 VDD.n1143 VDD.n1142 92.5005
R3832 VDD.n1557 VDD.n1556 92.5005
R3833 VDD.n1556 VDD.n1555 92.5005
R3834 VDD.n1145 VDD.n1144 92.5005
R3835 VDD.n1554 VDD.n1145 92.5005
R3836 VDD.n1552 VDD.n1551 92.5005
R3837 VDD.n1553 VDD.n1552 92.5005
R3838 VDD.n1574 VDD.n1134 92.5005
R3839 VDD.n1134 VDD.n1133 92.5005
R3840 VDD.n1577 VDD.n1576 92.5005
R3841 VDD.n1578 VDD.n1577 92.5005
R3842 VDD.n1575 VDD.n1135 92.5005
R3843 VDD.n1131 VDD.n1130 92.5005
R3844 VDD.n1582 VDD.n1581 92.5005
R3845 VDD.n1581 VDD.n1580 92.5005
R3846 VDD.n1585 VDD.n1584 92.5005
R3847 VDD.n1586 VDD.n1585 92.5005
R3848 VDD.n1127 VDD.n1126 92.5005
R3849 VDD.n1587 VDD.n1127 92.5005
R3850 VDD.n1590 VDD.n1589 92.5005
R3851 VDD.n1589 VDD.n1588 92.5005
R3852 VDD.n1591 VDD.n1125 92.5005
R3853 VDD.n1125 VDD.n1124 92.5005
R3854 VDD.n1593 VDD.n1592 92.5005
R3855 VDD.n1594 VDD.n1593 92.5005
R3856 VDD.n1123 VDD.n1122 92.5005
R3857 VDD.n1595 VDD.n1123 92.5005
R3858 VDD.n1598 VDD.n1597 92.5005
R3859 VDD.n1597 VDD.n1596 92.5005
R3860 VDD.n1599 VDD.n1121 92.5005
R3861 VDD.n1121 VDD.n1120 92.5005
R3862 VDD.n1601 VDD.n1600 92.5005
R3863 VDD.n1602 VDD.n1601 92.5005
R3864 VDD.n1119 VDD.n1118 92.5005
R3865 VDD.n1603 VDD.n1119 92.5005
R3866 VDD.n1606 VDD.n1605 92.5005
R3867 VDD.n1605 VDD.n1604 92.5005
R3868 VDD.n1607 VDD.n1117 92.5005
R3869 VDD.n1117 VDD.n1116 92.5005
R3870 VDD.n1609 VDD.n1608 92.5005
R3871 VDD.n1610 VDD.n1609 92.5005
R3872 VDD.n1115 VDD.n1114 92.5005
R3873 VDD.n1611 VDD.n1115 92.5005
R3874 VDD.n1614 VDD.n1613 92.5005
R3875 VDD.n1613 VDD.n1612 92.5005
R3876 VDD.n1615 VDD.n1113 92.5005
R3877 VDD.n1113 VDD.n1112 92.5005
R3878 VDD.n1617 VDD.n1616 92.5005
R3879 VDD.n1618 VDD.n1617 92.5005
R3880 VDD.n1111 VDD.n1110 92.5005
R3881 VDD.n1619 VDD.n1111 92.5005
R3882 VDD.n1622 VDD.n1621 92.5005
R3883 VDD.n1621 VDD.n1620 92.5005
R3884 VDD.n1623 VDD.n1109 92.5005
R3885 VDD.n1109 VDD.n1108 92.5005
R3886 VDD.n1625 VDD.n1624 92.5005
R3887 VDD.n1626 VDD.n1625 92.5005
R3888 VDD.n1107 VDD.n1106 92.5005
R3889 VDD.n1627 VDD.n1107 92.5005
R3890 VDD.n1630 VDD.n1629 92.5005
R3891 VDD.n1629 VDD.n1628 92.5005
R3892 VDD.n1631 VDD.n1105 92.5005
R3893 VDD.n1105 VDD.n1104 92.5005
R3894 VDD.n1633 VDD.n1632 92.5005
R3895 VDD.n1634 VDD.n1633 92.5005
R3896 VDD.n1103 VDD.n1102 92.5005
R3897 VDD.n1635 VDD.n1103 92.5005
R3898 VDD.n1640 VDD.n1639 92.5005
R3899 VDD.n1639 VDD.n1638 92.5005
R3900 VDD.n1641 VDD.n1101 92.5005
R3901 VDD.n1637 VDD.n1101 92.5005
R3902 VDD.n1583 VDD.n1129 92.5005
R3903 VDD.n1129 VDD.n1128 92.5005
R3904 VDD.n1655 VDD.n1654 92.5005
R3905 VDD.n1654 VDD.n1653 92.5005
R3906 VDD.n1656 VDD.n1094 92.5005
R3907 VDD.n1094 VDD.n1093 92.5005
R3908 VDD.n1658 VDD.n1657 92.5005
R3909 VDD.n1659 VDD.n1658 92.5005
R3910 VDD.n1092 VDD.n1091 92.5005
R3911 VDD.n1660 VDD.n1092 92.5005
R3912 VDD.n1663 VDD.n1662 92.5005
R3913 VDD.n1662 VDD.n1661 92.5005
R3914 VDD.n1664 VDD.n1090 92.5005
R3915 VDD.n1090 VDD.n1089 92.5005
R3916 VDD.n1666 VDD.n1665 92.5005
R3917 VDD.n1667 VDD.n1666 92.5005
R3918 VDD.n1088 VDD.n1087 92.5005
R3919 VDD.n1668 VDD.n1088 92.5005
R3920 VDD.n1671 VDD.n1670 92.5005
R3921 VDD.n1670 VDD.n1669 92.5005
R3922 VDD.n1672 VDD.n963 92.5005
R3923 VDD.n963 VDD.n961 92.5005
R3924 VDD.n1674 VDD.n1673 92.5005
R3925 VDD.n1675 VDD.n1674 92.5005
R3926 VDD.n1650 VDD.n1649 92.5005
R3927 VDD.n1651 VDD.n1650 92.5005
R3928 VDD.n1648 VDD.n1098 92.5005
R3929 VDD.n1098 VDD.n1097 92.5005
R3930 VDD.n1647 VDD.n1646 92.5005
R3931 VDD.n1644 VDD.n1099 92.5005
R3932 VDD.n1643 VDD.n1642 92.5005
R3933 VDD.n1643 VDD.n1100 92.5005
R3934 VDD.n1096 VDD.n1095 92.5005
R3935 VDD.n1652 VDD.n1096 92.5005
R3936 VDD.n1086 VDD.n962 92.5005
R3937 VDD.n1018 VDD.n1017 92.5005
R3938 VDD.n1015 VDD.n987 92.5005
R3939 VDD.n993 VDD.n988 92.5005
R3940 VDD.n1010 VDD.n1009 92.5005
R3941 VDD.n1007 VDD.n1006 92.5005
R3942 VDD.n1001 VDD.n994 92.5005
R3943 VDD.n999 VDD.n998 92.5005
R3944 VDD.n997 VDD.n964 92.5005
R3945 VDD.n1020 VDD.n972 92.5005
R3946 VDD.n1022 VDD.n971 92.5005
R3947 VDD.n1047 VDD.n1046 92.5005
R3948 VDD.n980 VDD.n954 92.5005
R3949 VDD.n1066 VDD.n1065 92.5005
R3950 VDD.n1063 VDD.n1062 92.5005
R3951 VDD.n1059 VDD.n981 92.5005
R3952 VDD.n1056 VDD.n1055 92.5005
R3953 VDD.n1054 VDD.n1053 92.5005
R3954 VDD.n983 VDD.n982 92.5005
R3955 VDD.n1058 VDD.n1057 92.5005
R3956 VDD.n1061 VDD.n1060 92.5005
R3957 VDD.n979 VDD.n978 92.5005
R3958 VDD.n1068 VDD.n1067 92.5005
R3959 VDD.n1679 VDD.n953 92.5005
R3960 VDD.n1682 VDD.n1681 92.5005
R3961 VDD.n1052 VDD.n974 92.5005
R3962 VDD.n1070 VDD.n974 92.5005
R3963 VDD.n1051 VDD.n1050 92.5005
R3964 VDD.n1049 VDD.n986 92.5005
R3965 VDD.n1265 VDD.n1264 92.5005
R3966 VDD.n1262 VDD.n1215 92.5005
R3967 VDD.n1261 VDD.n1260 92.5005
R3968 VDD.n1259 VDD.n1216 92.5005
R3969 VDD.n1257 VDD.n1256 92.5005
R3970 VDD.n1255 VDD.n1219 92.5005
R3971 VDD.n1222 VDD.n1219 92.5005
R3972 VDD.n1254 VDD.n1253 92.5005
R3973 VDD.n1253 VDD.n1252 92.5005
R3974 VDD.n1221 VDD.n1220 92.5005
R3975 VDD.n1251 VDD.n1221 92.5005
R3976 VDD.n1249 VDD.n1248 92.5005
R3977 VDD.n1250 VDD.n1249 92.5005
R3978 VDD.n1247 VDD.n1224 92.5005
R3979 VDD.n1224 VDD.n1223 92.5005
R3980 VDD.n1246 VDD.n1245 92.5005
R3981 VDD.n1245 VDD.n1244 92.5005
R3982 VDD.n1226 VDD.n1225 92.5005
R3983 VDD.n1243 VDD.n1226 92.5005
R3984 VDD.n1241 VDD.n1240 92.5005
R3985 VDD.n1242 VDD.n1241 92.5005
R3986 VDD.n1239 VDD.n1228 92.5005
R3987 VDD.n1228 VDD.n1227 92.5005
R3988 VDD.n1238 VDD.n1237 92.5005
R3989 VDD.n1237 VDD.n1236 92.5005
R3990 VDD.n1230 VDD.n1229 92.5005
R3991 VDD.n1235 VDD.n1230 92.5005
R3992 VDD.n1233 VDD.n1232 92.5005
R3993 VDD.n1234 VDD.n1233 92.5005
R3994 VDD.n1231 VDD.n957 92.5005
R3995 VDD.n959 VDD.n957 92.5005
R3996 VDD.n1678 VDD.n958 92.5005
R3997 VDD.n1678 VDD.n1677 92.5005
R3998 VDD.n1317 VDD.n1316 92.5005
R3999 VDD.n1316 VDD.n1315 92.5005
R4000 VDD.n1189 VDD.n1188 92.5005
R4001 VDD.n1314 VDD.n1189 92.5005
R4002 VDD.n1312 VDD.n1311 92.5005
R4003 VDD.n1313 VDD.n1312 92.5005
R4004 VDD.n1310 VDD.n1191 92.5005
R4005 VDD.n1191 VDD.n1190 92.5005
R4006 VDD.n1309 VDD.n1308 92.5005
R4007 VDD.n1308 VDD.n1307 92.5005
R4008 VDD.n1193 VDD.n1192 92.5005
R4009 VDD.n1306 VDD.n1193 92.5005
R4010 VDD.n1304 VDD.n1303 92.5005
R4011 VDD.n1305 VDD.n1304 92.5005
R4012 VDD.n1302 VDD.n1195 92.5005
R4013 VDD.n1195 VDD.n1194 92.5005
R4014 VDD.n1301 VDD.n1300 92.5005
R4015 VDD.n1300 VDD.n1299 92.5005
R4016 VDD.n1197 VDD.n1196 92.5005
R4017 VDD.n1298 VDD.n1197 92.5005
R4018 VDD.n1296 VDD.n1295 92.5005
R4019 VDD.n1297 VDD.n1296 92.5005
R4020 VDD.n1294 VDD.n1199 92.5005
R4021 VDD.n1199 VDD.n1198 92.5005
R4022 VDD.n1293 VDD.n1292 92.5005
R4023 VDD.n1292 VDD.n1291 92.5005
R4024 VDD.n1201 VDD.n1200 92.5005
R4025 VDD.n1290 VDD.n1201 92.5005
R4026 VDD.n1288 VDD.n1287 92.5005
R4027 VDD.n1289 VDD.n1288 92.5005
R4028 VDD.n1286 VDD.n1203 92.5005
R4029 VDD.n1203 VDD.n1202 92.5005
R4030 VDD.n1285 VDD.n1284 92.5005
R4031 VDD.n1284 VDD.n1283 92.5005
R4032 VDD.n1205 VDD.n1204 92.5005
R4033 VDD.n1282 VDD.n1205 92.5005
R4034 VDD.n1280 VDD.n1279 92.5005
R4035 VDD.n1281 VDD.n1280 92.5005
R4036 VDD.n1278 VDD.n1207 92.5005
R4037 VDD.n1207 VDD.n1206 92.5005
R4038 VDD.n1277 VDD.n1276 92.5005
R4039 VDD.n1276 VDD.n1275 92.5005
R4040 VDD.n1209 VDD.n1208 92.5005
R4041 VDD.n1274 VDD.n1209 92.5005
R4042 VDD.n1272 VDD.n1271 92.5005
R4043 VDD.n1273 VDD.n1272 92.5005
R4044 VDD.n1270 VDD.n1211 92.5005
R4045 VDD.n1211 VDD.n1210 92.5005
R4046 VDD.n1269 VDD.n1268 92.5005
R4047 VDD.n1268 VDD.n1267 92.5005
R4048 VDD.n1213 VDD.n1212 92.5005
R4049 VDD.n1266 VDD.n1213 92.5005
R4050 VDD.n1325 VDD.n1186 92.5005
R4051 VDD.n1329 VDD.n1328 92.5005
R4052 VDD.n1187 VDD.n1185 92.5005
R4053 VDD.n1359 VDD.n1169 92.5005
R4054 VDD.n1355 VDD.n1169 92.5005
R4055 VDD.n1358 VDD.n1357 92.5005
R4056 VDD.n1357 VDD.n1356 92.5005
R4057 VDD.n1171 VDD.n1170 92.5005
R4058 VDD.n1354 VDD.n1171 92.5005
R4059 VDD.n1352 VDD.n1351 92.5005
R4060 VDD.n1353 VDD.n1352 92.5005
R4061 VDD.n1350 VDD.n1173 92.5005
R4062 VDD.n1173 VDD.n1172 92.5005
R4063 VDD.n1349 VDD.n1348 92.5005
R4064 VDD.n1348 VDD.n1347 92.5005
R4065 VDD.n1175 VDD.n1174 92.5005
R4066 VDD.n1346 VDD.n1175 92.5005
R4067 VDD.n1344 VDD.n1343 92.5005
R4068 VDD.n1345 VDD.n1344 92.5005
R4069 VDD.n1342 VDD.n1177 92.5005
R4070 VDD.n1177 VDD.n1176 92.5005
R4071 VDD.n1341 VDD.n1340 92.5005
R4072 VDD.n1340 VDD.n1339 92.5005
R4073 VDD.n1179 VDD.n1178 92.5005
R4074 VDD.n1338 VDD.n1179 92.5005
R4075 VDD.n1336 VDD.n1335 92.5005
R4076 VDD.n1337 VDD.n1336 92.5005
R4077 VDD.n1334 VDD.n1181 92.5005
R4078 VDD.n1181 VDD.n1180 92.5005
R4079 VDD.n1333 VDD.n1332 92.5005
R4080 VDD.n1332 VDD.n1331 92.5005
R4081 VDD.n1183 VDD.n1182 92.5005
R4082 VDD.n1321 VDD.n1318 92.5005
R4083 VDD.n1324 VDD.n1323 92.5005
R4084 VDD.n1549 VDD.n1548 92.5005
R4085 VDD.n1466 VDD.n1149 92.5005
R4086 VDD.n1468 VDD.n1467 92.5005
R4087 VDD.n1465 VDD.n1464 92.5005
R4088 VDD.n1435 VDD.n1434 92.5005
R4089 VDD.n1459 VDD.n1458 92.5005
R4090 VDD.n1437 VDD.n1436 92.5005
R4091 VDD.n1453 VDD.n1452 92.5005
R4092 VDD.n1449 VDD.n1448 92.5005
R4093 VDD.n1447 VDD.n1446 92.5005
R4094 VDD.n1524 VDD.n1523 92.5005
R4095 VDD.n1528 VDD.n1527 92.5005
R4096 VDD.n1531 VDD.n1530 92.5005
R4097 VDD.n1373 VDD.n1372 92.5005
R4098 VDD.n1362 VDD.n1361 92.5005
R4099 VDD.n1540 VDD.n1539 92.5005
R4100 VDD.n1541 VDD.n1168 92.5005
R4101 VDD.n1544 VDD.n1543 92.5005
R4102 VDD.n1538 VDD.n1537 92.5005
R4103 VDD.n1371 VDD.n1364 92.5005
R4104 VDD.n1533 VDD.n1532 92.5005
R4105 VDD.n1529 VDD.n1370 92.5005
R4106 VDD.n1526 VDD.n1525 92.5005
R4107 VDD.n1374 VDD.n1161 92.5005
R4108 VDD.n1546 VDD.n1161 92.5005
R4109 VDD.n1522 VDD.n1521 92.5005
R4110 VDD.n1441 VDD.n1440 92.5005
R4111 VDD.n1443 VDD.n1442 92.5005
R4112 VDD.n1445 VDD.n1444 92.5005
R4113 VDD.n1451 VDD.n1450 92.5005
R4114 VDD.n1470 VDD.n1469 92.5005
R4115 VDD.n1463 VDD.n1462 92.5005
R4116 VDD.n1461 VDD.n1460 92.5005
R4117 VDD.n1457 VDD.n1456 92.5005
R4118 VDD.n1455 VDD.n1454 92.5005
R4119 VDD.n1078 VDD.n1077 92.5005
R4120 VDD.n969 VDD.n968 92.5005
R4121 VDD.n1081 VDD.n1080 92.5005
R4122 VDD.n1082 VDD.n1081 92.5005
R4123 VDD.n1014 VDD.n1013 92.5005
R4124 VDD.n1012 VDD.n1011 92.5005
R4125 VDD.n1002 VDD.n991 92.5005
R4126 VDD.n1005 VDD.n1004 92.5005
R4127 VDD.n1000 VDD.n967 92.5005
R4128 VDD.n1016 VDD.n970 92.5005
R4129 VDD.n1028 VDD.n1027 92.5005
R4130 VDD.n1030 VDD.n1026 92.5005
R4131 VDD.n1033 VDD.n1032 92.5005
R4132 VDD.n1035 VDD.n1034 92.5005
R4133 VDD.n1037 VDD.n1024 92.5005
R4134 VDD.n1040 VDD.n1039 92.5005
R4135 VDD.n1084 VDD.n1083 92.5005
R4136 VDD.n1083 VDD.n1082 92.5005
R4137 VDD.n966 VDD.n965 92.5005
R4138 VDD.n968 VDD.n966 92.5005
R4139 VDD.n1076 VDD.n1075 92.5005
R4140 VDD.n1077 VDD.n1076 92.5005
R4141 VDD.n1074 VDD.n1073 92.5005
R4142 VDD.n1073 VDD.n1072 92.5005
R4143 VDD.n1695 VDD.n1694 92.5005
R4144 VDD.n1694 VDD.n1693 92.5005
R4145 VDD.n1696 VDD.n936 92.5005
R4146 VDD.n940 VDD.n936 92.5005
R4147 VDD.n1698 VDD.n1697 92.5005
R4148 VDD.n1699 VDD.n1698 92.5005
R4149 VDD.n937 VDD.n935 92.5005
R4150 VDD.n1431 VDD.n935 92.5005
R4151 VDD.n1495 VDD.n1433 92.5005
R4152 VDD.n1433 VDD.n1432 92.5005
R4153 VDD.n1497 VDD.n1496 92.5005
R4154 VDD.n1498 VDD.n1497 92.5005
R4155 VDD.n1477 VDD.n1476 92.5005
R4156 VDD.n1476 VDD.n1384 92.5005
R4157 VDD.n1475 VDD.n1474 92.5005
R4158 VDD.n1475 VDD.n1383 92.5005
R4159 VDD.n1473 VDD.n1378 92.5005
R4160 VDD.n1518 VDD.n1378 92.5005
R4161 VDD.n1472 VDD.n1471 92.5005
R4162 VDD.n1471 VDD.n1365 92.5005
R4163 VDD.n1493 VDD.n1492 92.5005
R4164 VDD.n1490 VDD.n1478 92.5005
R4165 VDD.n1488 VDD.n1487 92.5005
R4166 VDD.n1486 VDD.n1485 92.5005
R4167 VDD.n1483 VDD.n1480 92.5005
R4168 VDD.n1481 VDD.n1394 92.5005
R4169 VDD.n1438 VDD.n1379 92.5005
R4170 VDD.n1379 VDD.n1365 92.5005
R4171 VDD.n1517 VDD.n1516 92.5005
R4172 VDD.n1518 VDD.n1517 92.5005
R4173 VDD.n1514 VDD.n1380 92.5005
R4174 VDD.n1383 VDD.n1380 92.5005
R4175 VDD.n1396 VDD.n1381 92.5005
R4176 VDD.n1396 VDD.n1384 92.5005
R4177 VDD.n1500 VDD.n1499 92.5005
R4178 VDD.n1499 VDD.n1498 92.5005
R4179 VDD.n1401 VDD.n1400 92.5005
R4180 VDD.n1432 VDD.n1401 92.5005
R4181 VDD.n1399 VDD.n931 92.5005
R4182 VDD.n1431 VDD.n931 92.5005
R4183 VDD.n1701 VDD.n1700 92.5005
R4184 VDD.n1700 VDD.n1699 92.5005
R4185 VDD.n944 VDD.n932 92.5005
R4186 VDD.n940 VDD.n932 92.5005
R4187 VDD.n1692 VDD.n1691 92.5005
R4188 VDD.n1693 VDD.n1692 92.5005
R4189 VDD.n1043 VDD.n973 92.5005
R4190 VDD.n1072 VDD.n973 92.5005
R4191 VDD.n1515 VDD.n1375 92.5005
R4192 VDD.n1377 VDD.n1375 92.5005
R4193 VDD.n1513 VDD.n1512 92.5005
R4194 VDD.n1512 VDD.n1511 92.5005
R4195 VDD.n1393 VDD.n1382 92.5005
R4196 VDD.n1390 VDD.n1382 92.5005
R4197 VDD.n1504 VDD.n1503 92.5005
R4198 VDD.n1505 VDD.n1504 92.5005
R4199 VDD.n1501 VDD.n1392 92.5005
R4200 VDD.n1402 VDD.n1392 92.5005
R4201 VDD.n1415 VDD.n929 92.5005
R4202 VDD.n1415 VDD.n933 92.5005
R4203 VDD.n1414 VDD.n930 92.5005
R4204 VDD.n1414 VDD.n934 92.5005
R4205 VDD.n947 VDD.n945 92.5005
R4206 VDD.n947 VDD.n941 92.5005
R4207 VDD.n1690 VDD.n1689 92.5005
R4208 VDD.n1689 VDD.n942 92.5005
R4209 VDD.n1688 VDD.n946 92.5005
R4210 VDD.n1688 VDD.n1687 92.5005
R4211 VDD.n1042 VDD.n948 92.5005
R4212 VDD.n1071 VDD.n948 92.5005
R4213 VDD.n1520 VDD.n1376 92.5005
R4214 VDD.n1520 VDD.n1519 92.5005
R4215 VDD.n508 VDD.n505 92.5005
R4216 VDD.n664 VDD.n508 92.5005
R4217 VDD.n829 VDD.n96 92.5005
R4218 VDD.n216 VDD.n96 92.5005
R4219 VDD.n831 VDD.n830 92.5005
R4220 VDD.n832 VDD.n831 92.5005
R4221 VDD.n97 VDD.n95 92.5005
R4222 VDD.n95 VDD.n87 92.5005
R4223 VDD.n554 VDD.n553 92.5005
R4224 VDD.n554 VDD.n86 92.5005
R4225 VDD.n555 VDD.n552 92.5005
R4226 VDD.n555 VDD.n79 92.5005
R4227 VDD.n557 VDD.n556 92.5005
R4228 VDD.n556 VDD.n78 92.5005
R4229 VDD.n570 VDD.n550 92.5005
R4230 VDD.n569 VDD.n568 92.5005
R4231 VDD.n567 VDD.n566 92.5005
R4232 VDD.n565 VDD.n564 92.5005
R4233 VDD.n563 VDD.n562 92.5005
R4234 VDD.n572 VDD.n571 92.5005
R4235 VDD.n534 VDD.n533 92.5005
R4236 VDD.n547 VDD.n534 92.5005
R4237 VDD.n652 VDD.n651 92.5005
R4238 VDD.n651 VDD.n650 92.5005
R4239 VDD.n653 VDD.n531 92.5005
R4240 VDD.n535 VDD.n531 92.5005
R4241 VDD.n655 VDD.n654 92.5005
R4242 VDD.n656 VDD.n655 92.5005
R4243 VDD.n532 VDD.n530 92.5005
R4244 VDD.n530 VDD.n522 92.5005
R4245 VDD.n695 VDD.n292 92.5005
R4246 VDD.n292 VDD.n291 92.5005
R4247 VDD.n718 VDD.n717 92.5005
R4248 VDD.n717 VDD.n716 92.5005
R4249 VDD.n282 VDD.n281 92.5005
R4250 VDD.n715 VDD.n282 92.5005
R4251 VDD.n713 VDD.n712 92.5005
R4252 VDD.n714 VDD.n713 92.5005
R4253 VDD.n711 VDD.n284 92.5005
R4254 VDD.n284 VDD.n283 92.5005
R4255 VDD.n710 VDD.n709 92.5005
R4256 VDD.n709 VDD.n708 92.5005
R4257 VDD.n286 VDD.n285 92.5005
R4258 VDD.n707 VDD.n286 92.5005
R4259 VDD.n705 VDD.n704 92.5005
R4260 VDD.n706 VDD.n705 92.5005
R4261 VDD.n703 VDD.n288 92.5005
R4262 VDD.n288 VDD.n287 92.5005
R4263 VDD.n702 VDD.n701 92.5005
R4264 VDD.n701 VDD.n700 92.5005
R4265 VDD.n290 VDD.n289 92.5005
R4266 VDD.n699 VDD.n290 92.5005
R4267 VDD.n697 VDD.n696 92.5005
R4268 VDD.n698 VDD.n697 92.5005
R4269 VDD.n719 VDD.n279 92.5005
R4270 VDD.n279 VDD.n278 92.5005
R4271 VDD.n722 VDD.n721 92.5005
R4272 VDD.n723 VDD.n722 92.5005
R4273 VDD.n720 VDD.n280 92.5005
R4274 VDD.n276 VDD.n275 92.5005
R4275 VDD.n727 VDD.n726 92.5005
R4276 VDD.n726 VDD.n725 92.5005
R4277 VDD.n730 VDD.n729 92.5005
R4278 VDD.n731 VDD.n730 92.5005
R4279 VDD.n272 VDD.n271 92.5005
R4280 VDD.n732 VDD.n272 92.5005
R4281 VDD.n735 VDD.n734 92.5005
R4282 VDD.n734 VDD.n733 92.5005
R4283 VDD.n736 VDD.n270 92.5005
R4284 VDD.n270 VDD.n269 92.5005
R4285 VDD.n738 VDD.n737 92.5005
R4286 VDD.n739 VDD.n738 92.5005
R4287 VDD.n268 VDD.n267 92.5005
R4288 VDD.n740 VDD.n268 92.5005
R4289 VDD.n743 VDD.n742 92.5005
R4290 VDD.n742 VDD.n741 92.5005
R4291 VDD.n744 VDD.n266 92.5005
R4292 VDD.n266 VDD.n265 92.5005
R4293 VDD.n746 VDD.n745 92.5005
R4294 VDD.n747 VDD.n746 92.5005
R4295 VDD.n264 VDD.n263 92.5005
R4296 VDD.n748 VDD.n264 92.5005
R4297 VDD.n751 VDD.n750 92.5005
R4298 VDD.n750 VDD.n749 92.5005
R4299 VDD.n752 VDD.n262 92.5005
R4300 VDD.n262 VDD.n261 92.5005
R4301 VDD.n754 VDD.n753 92.5005
R4302 VDD.n755 VDD.n754 92.5005
R4303 VDD.n260 VDD.n259 92.5005
R4304 VDD.n756 VDD.n260 92.5005
R4305 VDD.n759 VDD.n758 92.5005
R4306 VDD.n758 VDD.n757 92.5005
R4307 VDD.n760 VDD.n258 92.5005
R4308 VDD.n258 VDD.n257 92.5005
R4309 VDD.n762 VDD.n761 92.5005
R4310 VDD.n763 VDD.n762 92.5005
R4311 VDD.n256 VDD.n255 92.5005
R4312 VDD.n764 VDD.n256 92.5005
R4313 VDD.n767 VDD.n766 92.5005
R4314 VDD.n766 VDD.n765 92.5005
R4315 VDD.n768 VDD.n254 92.5005
R4316 VDD.n254 VDD.n253 92.5005
R4317 VDD.n770 VDD.n769 92.5005
R4318 VDD.n771 VDD.n770 92.5005
R4319 VDD.n252 VDD.n251 92.5005
R4320 VDD.n772 VDD.n252 92.5005
R4321 VDD.n775 VDD.n774 92.5005
R4322 VDD.n774 VDD.n773 92.5005
R4323 VDD.n776 VDD.n250 92.5005
R4324 VDD.n250 VDD.n249 92.5005
R4325 VDD.n778 VDD.n777 92.5005
R4326 VDD.n779 VDD.n778 92.5005
R4327 VDD.n248 VDD.n247 92.5005
R4328 VDD.n780 VDD.n248 92.5005
R4329 VDD.n785 VDD.n784 92.5005
R4330 VDD.n784 VDD.n783 92.5005
R4331 VDD.n786 VDD.n246 92.5005
R4332 VDD.n782 VDD.n246 92.5005
R4333 VDD.n728 VDD.n274 92.5005
R4334 VDD.n274 VDD.n273 92.5005
R4335 VDD.n800 VDD.n799 92.5005
R4336 VDD.n799 VDD.n798 92.5005
R4337 VDD.n801 VDD.n239 92.5005
R4338 VDD.n239 VDD.n238 92.5005
R4339 VDD.n803 VDD.n802 92.5005
R4340 VDD.n804 VDD.n803 92.5005
R4341 VDD.n237 VDD.n236 92.5005
R4342 VDD.n805 VDD.n237 92.5005
R4343 VDD.n808 VDD.n807 92.5005
R4344 VDD.n807 VDD.n806 92.5005
R4345 VDD.n809 VDD.n235 92.5005
R4346 VDD.n235 VDD.n234 92.5005
R4347 VDD.n811 VDD.n810 92.5005
R4348 VDD.n812 VDD.n811 92.5005
R4349 VDD.n233 VDD.n232 92.5005
R4350 VDD.n813 VDD.n233 92.5005
R4351 VDD.n816 VDD.n815 92.5005
R4352 VDD.n815 VDD.n814 92.5005
R4353 VDD.n817 VDD.n108 92.5005
R4354 VDD.n108 VDD.n106 92.5005
R4355 VDD.n819 VDD.n818 92.5005
R4356 VDD.n820 VDD.n819 92.5005
R4357 VDD.n795 VDD.n794 92.5005
R4358 VDD.n796 VDD.n795 92.5005
R4359 VDD.n793 VDD.n243 92.5005
R4360 VDD.n243 VDD.n242 92.5005
R4361 VDD.n792 VDD.n791 92.5005
R4362 VDD.n789 VDD.n244 92.5005
R4363 VDD.n788 VDD.n787 92.5005
R4364 VDD.n788 VDD.n245 92.5005
R4365 VDD.n241 VDD.n240 92.5005
R4366 VDD.n797 VDD.n241 92.5005
R4367 VDD.n231 VDD.n107 92.5005
R4368 VDD.n163 VDD.n162 92.5005
R4369 VDD.n160 VDD.n132 92.5005
R4370 VDD.n138 VDD.n133 92.5005
R4371 VDD.n155 VDD.n154 92.5005
R4372 VDD.n152 VDD.n151 92.5005
R4373 VDD.n146 VDD.n139 92.5005
R4374 VDD.n144 VDD.n143 92.5005
R4375 VDD.n142 VDD.n109 92.5005
R4376 VDD.n165 VDD.n117 92.5005
R4377 VDD.n167 VDD.n116 92.5005
R4378 VDD.n192 VDD.n191 92.5005
R4379 VDD.n125 VDD.n99 92.5005
R4380 VDD.n211 VDD.n210 92.5005
R4381 VDD.n208 VDD.n207 92.5005
R4382 VDD.n204 VDD.n126 92.5005
R4383 VDD.n201 VDD.n200 92.5005
R4384 VDD.n199 VDD.n198 92.5005
R4385 VDD.n128 VDD.n127 92.5005
R4386 VDD.n203 VDD.n202 92.5005
R4387 VDD.n206 VDD.n205 92.5005
R4388 VDD.n124 VDD.n123 92.5005
R4389 VDD.n213 VDD.n212 92.5005
R4390 VDD.n824 VDD.n98 92.5005
R4391 VDD.n827 VDD.n826 92.5005
R4392 VDD.n197 VDD.n119 92.5005
R4393 VDD.n215 VDD.n119 92.5005
R4394 VDD.n196 VDD.n195 92.5005
R4395 VDD.n194 VDD.n131 92.5005
R4396 VDD.n410 VDD.n409 92.5005
R4397 VDD.n407 VDD.n360 92.5005
R4398 VDD.n406 VDD.n405 92.5005
R4399 VDD.n404 VDD.n361 92.5005
R4400 VDD.n402 VDD.n401 92.5005
R4401 VDD.n400 VDD.n364 92.5005
R4402 VDD.n367 VDD.n364 92.5005
R4403 VDD.n399 VDD.n398 92.5005
R4404 VDD.n398 VDD.n397 92.5005
R4405 VDD.n366 VDD.n365 92.5005
R4406 VDD.n396 VDD.n366 92.5005
R4407 VDD.n394 VDD.n393 92.5005
R4408 VDD.n395 VDD.n394 92.5005
R4409 VDD.n392 VDD.n369 92.5005
R4410 VDD.n369 VDD.n368 92.5005
R4411 VDD.n391 VDD.n390 92.5005
R4412 VDD.n390 VDD.n389 92.5005
R4413 VDD.n371 VDD.n370 92.5005
R4414 VDD.n388 VDD.n371 92.5005
R4415 VDD.n386 VDD.n385 92.5005
R4416 VDD.n387 VDD.n386 92.5005
R4417 VDD.n384 VDD.n373 92.5005
R4418 VDD.n373 VDD.n372 92.5005
R4419 VDD.n383 VDD.n382 92.5005
R4420 VDD.n382 VDD.n381 92.5005
R4421 VDD.n375 VDD.n374 92.5005
R4422 VDD.n380 VDD.n375 92.5005
R4423 VDD.n378 VDD.n377 92.5005
R4424 VDD.n379 VDD.n378 92.5005
R4425 VDD.n376 VDD.n102 92.5005
R4426 VDD.n104 VDD.n102 92.5005
R4427 VDD.n823 VDD.n103 92.5005
R4428 VDD.n823 VDD.n822 92.5005
R4429 VDD.n462 VDD.n461 92.5005
R4430 VDD.n461 VDD.n460 92.5005
R4431 VDD.n334 VDD.n333 92.5005
R4432 VDD.n459 VDD.n334 92.5005
R4433 VDD.n457 VDD.n456 92.5005
R4434 VDD.n458 VDD.n457 92.5005
R4435 VDD.n455 VDD.n336 92.5005
R4436 VDD.n336 VDD.n335 92.5005
R4437 VDD.n454 VDD.n453 92.5005
R4438 VDD.n453 VDD.n452 92.5005
R4439 VDD.n338 VDD.n337 92.5005
R4440 VDD.n451 VDD.n338 92.5005
R4441 VDD.n449 VDD.n448 92.5005
R4442 VDD.n450 VDD.n449 92.5005
R4443 VDD.n447 VDD.n340 92.5005
R4444 VDD.n340 VDD.n339 92.5005
R4445 VDD.n446 VDD.n445 92.5005
R4446 VDD.n445 VDD.n444 92.5005
R4447 VDD.n342 VDD.n341 92.5005
R4448 VDD.n443 VDD.n342 92.5005
R4449 VDD.n441 VDD.n440 92.5005
R4450 VDD.n442 VDD.n441 92.5005
R4451 VDD.n439 VDD.n344 92.5005
R4452 VDD.n344 VDD.n343 92.5005
R4453 VDD.n438 VDD.n437 92.5005
R4454 VDD.n437 VDD.n436 92.5005
R4455 VDD.n346 VDD.n345 92.5005
R4456 VDD.n435 VDD.n346 92.5005
R4457 VDD.n433 VDD.n432 92.5005
R4458 VDD.n434 VDD.n433 92.5005
R4459 VDD.n431 VDD.n348 92.5005
R4460 VDD.n348 VDD.n347 92.5005
R4461 VDD.n430 VDD.n429 92.5005
R4462 VDD.n429 VDD.n428 92.5005
R4463 VDD.n350 VDD.n349 92.5005
R4464 VDD.n427 VDD.n350 92.5005
R4465 VDD.n425 VDD.n424 92.5005
R4466 VDD.n426 VDD.n425 92.5005
R4467 VDD.n423 VDD.n352 92.5005
R4468 VDD.n352 VDD.n351 92.5005
R4469 VDD.n422 VDD.n421 92.5005
R4470 VDD.n421 VDD.n420 92.5005
R4471 VDD.n354 VDD.n353 92.5005
R4472 VDD.n419 VDD.n354 92.5005
R4473 VDD.n417 VDD.n416 92.5005
R4474 VDD.n418 VDD.n417 92.5005
R4475 VDD.n415 VDD.n356 92.5005
R4476 VDD.n356 VDD.n355 92.5005
R4477 VDD.n414 VDD.n413 92.5005
R4478 VDD.n413 VDD.n412 92.5005
R4479 VDD.n358 VDD.n357 92.5005
R4480 VDD.n411 VDD.n358 92.5005
R4481 VDD.n470 VDD.n331 92.5005
R4482 VDD.n474 VDD.n473 92.5005
R4483 VDD.n332 VDD.n330 92.5005
R4484 VDD.n504 VDD.n314 92.5005
R4485 VDD.n500 VDD.n314 92.5005
R4486 VDD.n503 VDD.n502 92.5005
R4487 VDD.n502 VDD.n501 92.5005
R4488 VDD.n316 VDD.n315 92.5005
R4489 VDD.n499 VDD.n316 92.5005
R4490 VDD.n497 VDD.n496 92.5005
R4491 VDD.n498 VDD.n497 92.5005
R4492 VDD.n495 VDD.n318 92.5005
R4493 VDD.n318 VDD.n317 92.5005
R4494 VDD.n494 VDD.n493 92.5005
R4495 VDD.n493 VDD.n492 92.5005
R4496 VDD.n320 VDD.n319 92.5005
R4497 VDD.n491 VDD.n320 92.5005
R4498 VDD.n489 VDD.n488 92.5005
R4499 VDD.n490 VDD.n489 92.5005
R4500 VDD.n487 VDD.n322 92.5005
R4501 VDD.n322 VDD.n321 92.5005
R4502 VDD.n486 VDD.n485 92.5005
R4503 VDD.n485 VDD.n484 92.5005
R4504 VDD.n324 VDD.n323 92.5005
R4505 VDD.n483 VDD.n324 92.5005
R4506 VDD.n481 VDD.n480 92.5005
R4507 VDD.n482 VDD.n481 92.5005
R4508 VDD.n479 VDD.n326 92.5005
R4509 VDD.n326 VDD.n325 92.5005
R4510 VDD.n478 VDD.n477 92.5005
R4511 VDD.n477 VDD.n476 92.5005
R4512 VDD.n328 VDD.n327 92.5005
R4513 VDD.n466 VDD.n463 92.5005
R4514 VDD.n469 VDD.n468 92.5005
R4515 VDD.n694 VDD.n693 92.5005
R4516 VDD.n611 VDD.n294 92.5005
R4517 VDD.n613 VDD.n612 92.5005
R4518 VDD.n610 VDD.n609 92.5005
R4519 VDD.n580 VDD.n579 92.5005
R4520 VDD.n604 VDD.n603 92.5005
R4521 VDD.n582 VDD.n581 92.5005
R4522 VDD.n598 VDD.n597 92.5005
R4523 VDD.n594 VDD.n593 92.5005
R4524 VDD.n592 VDD.n591 92.5005
R4525 VDD.n669 VDD.n668 92.5005
R4526 VDD.n673 VDD.n672 92.5005
R4527 VDD.n676 VDD.n675 92.5005
R4528 VDD.n518 VDD.n517 92.5005
R4529 VDD.n507 VDD.n506 92.5005
R4530 VDD.n685 VDD.n684 92.5005
R4531 VDD.n686 VDD.n313 92.5005
R4532 VDD.n689 VDD.n688 92.5005
R4533 VDD.n683 VDD.n682 92.5005
R4534 VDD.n516 VDD.n509 92.5005
R4535 VDD.n678 VDD.n677 92.5005
R4536 VDD.n674 VDD.n515 92.5005
R4537 VDD.n671 VDD.n670 92.5005
R4538 VDD.n519 VDD.n306 92.5005
R4539 VDD.n691 VDD.n306 92.5005
R4540 VDD.n667 VDD.n666 92.5005
R4541 VDD.n586 VDD.n585 92.5005
R4542 VDD.n588 VDD.n587 92.5005
R4543 VDD.n590 VDD.n589 92.5005
R4544 VDD.n596 VDD.n595 92.5005
R4545 VDD.n615 VDD.n614 92.5005
R4546 VDD.n608 VDD.n607 92.5005
R4547 VDD.n606 VDD.n605 92.5005
R4548 VDD.n602 VDD.n601 92.5005
R4549 VDD.n600 VDD.n599 92.5005
R4550 VDD.n223 VDD.n222 92.5005
R4551 VDD.n114 VDD.n113 92.5005
R4552 VDD.n226 VDD.n225 92.5005
R4553 VDD.n227 VDD.n226 92.5005
R4554 VDD.n159 VDD.n158 92.5005
R4555 VDD.n157 VDD.n156 92.5005
R4556 VDD.n147 VDD.n136 92.5005
R4557 VDD.n150 VDD.n149 92.5005
R4558 VDD.n145 VDD.n112 92.5005
R4559 VDD.n161 VDD.n115 92.5005
R4560 VDD.n173 VDD.n172 92.5005
R4561 VDD.n175 VDD.n171 92.5005
R4562 VDD.n178 VDD.n177 92.5005
R4563 VDD.n180 VDD.n179 92.5005
R4564 VDD.n182 VDD.n169 92.5005
R4565 VDD.n185 VDD.n184 92.5005
R4566 VDD.n229 VDD.n228 92.5005
R4567 VDD.n228 VDD.n227 92.5005
R4568 VDD.n111 VDD.n110 92.5005
R4569 VDD.n113 VDD.n111 92.5005
R4570 VDD.n221 VDD.n220 92.5005
R4571 VDD.n222 VDD.n221 92.5005
R4572 VDD.n219 VDD.n218 92.5005
R4573 VDD.n218 VDD.n217 92.5005
R4574 VDD.n840 VDD.n839 92.5005
R4575 VDD.n839 VDD.n838 92.5005
R4576 VDD.n841 VDD.n81 92.5005
R4577 VDD.n85 VDD.n81 92.5005
R4578 VDD.n843 VDD.n842 92.5005
R4579 VDD.n844 VDD.n843 92.5005
R4580 VDD.n82 VDD.n80 92.5005
R4581 VDD.n576 VDD.n80 92.5005
R4582 VDD.n640 VDD.n578 92.5005
R4583 VDD.n578 VDD.n577 92.5005
R4584 VDD.n642 VDD.n641 92.5005
R4585 VDD.n643 VDD.n642 92.5005
R4586 VDD.n622 VDD.n621 92.5005
R4587 VDD.n621 VDD.n529 92.5005
R4588 VDD.n620 VDD.n619 92.5005
R4589 VDD.n620 VDD.n528 92.5005
R4590 VDD.n618 VDD.n523 92.5005
R4591 VDD.n663 VDD.n523 92.5005
R4592 VDD.n617 VDD.n616 92.5005
R4593 VDD.n616 VDD.n510 92.5005
R4594 VDD.n638 VDD.n637 92.5005
R4595 VDD.n635 VDD.n623 92.5005
R4596 VDD.n633 VDD.n632 92.5005
R4597 VDD.n631 VDD.n630 92.5005
R4598 VDD.n628 VDD.n625 92.5005
R4599 VDD.n626 VDD.n539 92.5005
R4600 VDD.n583 VDD.n524 92.5005
R4601 VDD.n524 VDD.n510 92.5005
R4602 VDD.n662 VDD.n661 92.5005
R4603 VDD.n663 VDD.n662 92.5005
R4604 VDD.n659 VDD.n525 92.5005
R4605 VDD.n528 VDD.n525 92.5005
R4606 VDD.n541 VDD.n526 92.5005
R4607 VDD.n541 VDD.n529 92.5005
R4608 VDD.n645 VDD.n644 92.5005
R4609 VDD.n644 VDD.n643 92.5005
R4610 VDD.n546 VDD.n545 92.5005
R4611 VDD.n577 VDD.n546 92.5005
R4612 VDD.n544 VDD.n76 92.5005
R4613 VDD.n576 VDD.n76 92.5005
R4614 VDD.n846 VDD.n845 92.5005
R4615 VDD.n845 VDD.n844 92.5005
R4616 VDD.n89 VDD.n77 92.5005
R4617 VDD.n85 VDD.n77 92.5005
R4618 VDD.n837 VDD.n836 92.5005
R4619 VDD.n838 VDD.n837 92.5005
R4620 VDD.n188 VDD.n118 92.5005
R4621 VDD.n217 VDD.n118 92.5005
R4622 VDD.n660 VDD.n520 92.5005
R4623 VDD.n522 VDD.n520 92.5005
R4624 VDD.n658 VDD.n657 92.5005
R4625 VDD.n657 VDD.n656 92.5005
R4626 VDD.n538 VDD.n527 92.5005
R4627 VDD.n535 VDD.n527 92.5005
R4628 VDD.n649 VDD.n648 92.5005
R4629 VDD.n650 VDD.n649 92.5005
R4630 VDD.n646 VDD.n537 92.5005
R4631 VDD.n547 VDD.n537 92.5005
R4632 VDD.n560 VDD.n74 92.5005
R4633 VDD.n560 VDD.n78 92.5005
R4634 VDD.n559 VDD.n75 92.5005
R4635 VDD.n559 VDD.n79 92.5005
R4636 VDD.n92 VDD.n90 92.5005
R4637 VDD.n92 VDD.n86 92.5005
R4638 VDD.n835 VDD.n834 92.5005
R4639 VDD.n834 VDD.n87 92.5005
R4640 VDD.n833 VDD.n91 92.5005
R4641 VDD.n833 VDD.n832 92.5005
R4642 VDD.n187 VDD.n93 92.5005
R4643 VDD.n216 VDD.n93 92.5005
R4644 VDD.n665 VDD.n521 92.5005
R4645 VDD.n665 VDD.n664 92.5005
R4646 VDD.n44 VDD.t28 91.8719
R4647 VDD.n913 VDD.t146 91.8719
R4648 VDD.n1753 VDD.t158 91.8719
R4649 VDD.n2622 VDD.t107 91.8719
R4650 VDD.n58 VDD.t29 84.4681
R4651 VDD.n896 VDD.t21 84.4681
R4652 VDD.n1767 VDD.t74 84.4681
R4653 VDD.n2614 VDD.t108 84.4681
R4654 VDD.n44 VDD.n43 83.1021
R4655 VDD.n913 VDD.n912 83.1021
R4656 VDD.n1753 VDD.n1752 83.1021
R4657 VDD.n2622 VDD.n2621 83.1021
R4658 VDD.n33 VDD.t55 78.5582
R4659 VDD.t25 VDD.n861 78.5582
R4660 VDD.n1742 VDD.t63 78.5582
R4661 VDD.n2593 VDD.t133 78.5582
R4662 VDD.n2531 VDD.n2530 78.4132
R4663 VDD.n2209 VDD.n2004 78.4132
R4664 VDD.n1677 VDD.n1676 78.4132
R4665 VDD.n1355 VDD.n1150 78.4132
R4666 VDD.n822 VDD.n821 78.4132
R4667 VDD.n500 VDD.n295 78.4132
R4668 VDD.n3807 VDD.t59 75.5912
R4669 VDD.n3807 VDD.t110 75.5912
R4670 VDD.n3804 VDD.n3803 74.6009
R4671 VDD.n4011 VDD.n3976 72.0905
R4672 VDD.n4011 VDD.n3977 72.0905
R4673 VDD.n4011 VDD.n3978 72.0905
R4674 VDD.n4011 VDD.n3979 72.0905
R4675 VDD.n4011 VDD.n3980 72.0905
R4676 VDD.n4011 VDD.n3981 72.0905
R4677 VDD.n4011 VDD.n3982 72.0905
R4678 VDD.n4011 VDD.n3983 72.0905
R4679 VDD.n4011 VDD.n3984 72.0905
R4680 VDD.n4011 VDD.n3985 72.0905
R4681 VDD.n4011 VDD.n3986 72.0905
R4682 VDD.n4011 VDD.n3987 72.0905
R4683 VDD.n4011 VDD.n3988 72.0905
R4684 VDD.n4011 VDD.n3989 72.0905
R4685 VDD.n4011 VDD.n3990 72.0905
R4686 VDD.n4011 VDD.n3991 72.0905
R4687 VDD.n4011 VDD.n3992 72.0905
R4688 VDD.n4011 VDD.n3993 72.0905
R4689 VDD.n4011 VDD.n3994 72.0905
R4690 VDD.n4011 VDD.n3995 72.0905
R4691 VDD.n4011 VDD.n3996 72.0905
R4692 VDD.n4011 VDD.n3997 72.0905
R4693 VDD.n4011 VDD.n3998 72.0905
R4694 VDD.n4011 VDD.n3999 72.0905
R4695 VDD.n4011 VDD.n4000 72.0905
R4696 VDD.n4011 VDD.n4001 72.0905
R4697 VDD.n4011 VDD.n4002 72.0905
R4698 VDD.n4011 VDD.n4003 72.0905
R4699 VDD.n4011 VDD.n4004 72.0905
R4700 VDD.n4011 VDD.n4005 72.0905
R4701 VDD.n4011 VDD.n4006 72.0905
R4702 VDD.n4011 VDD.n4007 72.0905
R4703 VDD.n4011 VDD.n4008 72.0905
R4704 VDD.n4011 VDD.n4009 72.0905
R4705 VDD.n1875 VDD.n1810 72.0905
R4706 VDD.n1877 VDD.n1810 72.0905
R4707 VDD.n2176 VDD.n2038 72.0905
R4708 VDD.n2400 VDD.n2005 72.0905
R4709 VDD.n2400 VDD.n2006 72.0905
R4710 VDD.n2400 VDD.n2007 72.0905
R4711 VDD.n2400 VDD.n2008 72.0905
R4712 VDD.n2400 VDD.n2009 72.0905
R4713 VDD.n2400 VDD.n2010 72.0905
R4714 VDD.n2400 VDD.n2011 72.0905
R4715 VDD.n2400 VDD.n2012 72.0905
R4716 VDD.n2400 VDD.n2017 72.0905
R4717 VDD.n2400 VDD.n2018 72.0905
R4718 VDD.n2400 VDD.n2019 72.0905
R4719 VDD.n2400 VDD.n2020 72.0905
R4720 VDD.n2400 VDD.n2021 72.0905
R4721 VDD.n1021 VDD.n956 72.0905
R4722 VDD.n1023 VDD.n956 72.0905
R4723 VDD.n1322 VDD.n1184 72.0905
R4724 VDD.n1546 VDD.n1151 72.0905
R4725 VDD.n1546 VDD.n1152 72.0905
R4726 VDD.n1546 VDD.n1153 72.0905
R4727 VDD.n1546 VDD.n1154 72.0905
R4728 VDD.n1546 VDD.n1155 72.0905
R4729 VDD.n1546 VDD.n1156 72.0905
R4730 VDD.n1546 VDD.n1157 72.0905
R4731 VDD.n1546 VDD.n1158 72.0905
R4732 VDD.n1546 VDD.n1163 72.0905
R4733 VDD.n1546 VDD.n1164 72.0905
R4734 VDD.n1546 VDD.n1165 72.0905
R4735 VDD.n1546 VDD.n1166 72.0905
R4736 VDD.n1546 VDD.n1167 72.0905
R4737 VDD.n166 VDD.n101 72.0905
R4738 VDD.n168 VDD.n101 72.0905
R4739 VDD.n467 VDD.n329 72.0905
R4740 VDD.n691 VDD.n296 72.0905
R4741 VDD.n691 VDD.n297 72.0905
R4742 VDD.n691 VDD.n298 72.0905
R4743 VDD.n691 VDD.n299 72.0905
R4744 VDD.n691 VDD.n300 72.0905
R4745 VDD.n691 VDD.n301 72.0905
R4746 VDD.n691 VDD.n302 72.0905
R4747 VDD.n691 VDD.n303 72.0905
R4748 VDD.n691 VDD.n308 72.0905
R4749 VDD.n691 VDD.n309 72.0905
R4750 VDD.n691 VDD.n310 72.0905
R4751 VDD.n691 VDD.n311 72.0905
R4752 VDD.n691 VDD.n312 72.0905
R4753 VDD.n2389 VDD.n2219 71.1543
R4754 VDD.n1936 VDD.n1814 71.1543
R4755 VDD.n1535 VDD.n1365 71.1543
R4756 VDD.n1082 VDD.n960 71.1543
R4757 VDD.n680 VDD.n510 71.1543
R4758 VDD.n227 VDD.n105 71.1543
R4759 VDD.n3558 VDD.n3557 70.5361
R4760 VDD.n3561 VDD.n3560 70.5361
R4761 VDD.n3564 VDD.n3563 70.5361
R4762 VDD.n3567 VDD.n3566 70.5361
R4763 VDD.n3570 VDD.n3569 70.5361
R4764 VDD.n3574 VDD.n3572 70.5361
R4765 VDD.n3438 VDD.n3437 70.5361
R4766 VDD.n3441 VDD.n3440 70.5361
R4767 VDD.n3444 VDD.n3443 70.5361
R4768 VDD.n3447 VDD.n3446 70.5361
R4769 VDD.n3450 VDD.n3449 70.5361
R4770 VDD.n3453 VDD.n3452 70.5361
R4771 VDD.n3539 VDD.n3537 70.5361
R4772 VDD.n3481 VDD.n3480 70.5361
R4773 VDD.n3484 VDD.n3483 70.5361
R4774 VDD.n3487 VDD.n3486 70.5361
R4775 VDD.n3490 VDD.n3489 70.5361
R4776 VDD.n3493 VDD.n3492 70.5361
R4777 VDD.n3496 VDD.n3495 70.5361
R4778 VDD.n3499 VDD.n3498 70.5361
R4779 VDD.n3502 VDD.n3501 70.5361
R4780 VDD.n3505 VDD.n3504 70.5361
R4781 VDD.n3508 VDD.n3507 70.5361
R4782 VDD.n3511 VDD.n3510 70.5361
R4783 VDD.n3514 VDD.n3513 70.5361
R4784 VDD.n3517 VDD.n3516 70.5361
R4785 VDD.n3520 VDD.n3519 70.5361
R4786 VDD.n3523 VDD.n3522 70.5361
R4787 VDD.n3526 VDD.n3525 70.5361
R4788 VDD.n3529 VDD.n3528 70.5361
R4789 VDD.n3532 VDD.n3531 70.5361
R4790 VDD.n3535 VDD.n3534 70.5361
R4791 VDD.n3539 VDD.n3538 70.5361
R4792 VDD.n3579 VDD.n3578 70.5361
R4793 VDD.n3582 VDD.n3581 70.5361
R4794 VDD.n3585 VDD.n3584 70.5361
R4795 VDD.n3588 VDD.n3587 70.5361
R4796 VDD.n3591 VDD.n3590 70.5361
R4797 VDD.n3594 VDD.n3593 70.5361
R4798 VDD.n3574 VDD.n3573 70.5361
R4799 VDD.n3603 VDD.n3602 70.5361
R4800 VDD.n3606 VDD.n3605 70.5361
R4801 VDD.n3609 VDD.n3608 70.5361
R4802 VDD.n3612 VDD.n3611 70.5361
R4803 VDD.n3615 VDD.n3614 70.5361
R4804 VDD.n1924 VDD.n1830 67.9542
R4805 VDD.n1924 VDD.n1831 67.9542
R4806 VDD.n1885 VDD.n1803 67.9542
R4807 VDD.n1879 VDD.n1803 67.9542
R4808 VDD.n1890 VDD.n1803 67.9542
R4809 VDD.n2343 VDD.n2245 67.9542
R4810 VDD.n2333 VDD.n2245 67.9542
R4811 VDD.n2338 VDD.n2245 67.9542
R4812 VDD.n1070 VDD.n976 67.9542
R4813 VDD.n1070 VDD.n977 67.9542
R4814 VDD.n1031 VDD.n949 67.9542
R4815 VDD.n1025 VDD.n949 67.9542
R4816 VDD.n1036 VDD.n949 67.9542
R4817 VDD.n1489 VDD.n1391 67.9542
R4818 VDD.n1479 VDD.n1391 67.9542
R4819 VDD.n1484 VDD.n1391 67.9542
R4820 VDD.n215 VDD.n121 67.9542
R4821 VDD.n215 VDD.n122 67.9542
R4822 VDD.n176 VDD.n94 67.9542
R4823 VDD.n170 VDD.n94 67.9542
R4824 VDD.n181 VDD.n94 67.9542
R4825 VDD.n634 VDD.n536 67.9542
R4826 VDD.n624 VDD.n536 67.9542
R4827 VDD.n629 VDD.n536 67.9542
R4828 VDD.n6498 VDD.n6497 66.8858
R4829 VDD.n8049 VDD.n8048 66.8856
R4830 VDD.n4687 VDD.t79 60.2505
R4831 VDD.n4703 VDD.t99 60.2505
R4832 VDD.n5028 VDD.t96 60.2505
R4833 VDD.n5044 VDD.t89 60.2505
R4834 VDD.n4340 VDD.t76 60.2505
R4835 VDD.n4325 VDD.t82 60.2505
R4836 VDD.n4506 VDD.t84 60.2505
R4837 VDD.n4435 VDD.t87 60.2505
R4838 VDD.n3645 VDD.t101 60.2505
R4839 VDD.n5262 VDD.t93 60.2505
R4840 VDD.n1923 VDD.n1832 60.14
R4841 VDD.n1892 VDD.n1891 60.14
R4842 VDD.n2337 VDD.n2336 60.14
R4843 VDD.n1069 VDD.n978 60.14
R4844 VDD.n1038 VDD.n1037 60.14
R4845 VDD.n1483 VDD.n1482 60.14
R4846 VDD.n214 VDD.n123 60.14
R4847 VDD.n183 VDD.n182 60.14
R4848 VDD.n628 VDD.n627 60.14
R4849 VDD.n1911 VDD.n1829 60.1394
R4850 VDD.n1884 VDD.n1883 60.1394
R4851 VDD.n2345 VDD.n2344 60.1394
R4852 VDD.n1057 VDD.n975 60.1394
R4853 VDD.n1030 VDD.n1029 60.1394
R4854 VDD.n1491 VDD.n1490 60.1394
R4855 VDD.n202 VDD.n120 60.1394
R4856 VDD.n175 VDD.n174 60.1394
R4857 VDD.n636 VDD.n635 60.1394
R4858 VDD.t83 VDD.n4379 59.2764
R4859 VDD.n8564 VDD.n8561 57.2334
R4860 VDD.n8564 VDD.n8562 57.2334
R4861 VDD.n8564 VDD.n8563 57.2334
R4862 VDD.n2352 VDD.n2256 55.1287
R4863 VDD.n1498 VDD.n1402 55.1287
R4864 VDD.n643 VDD.n547 55.1287
R4865 VDD.n8047 VDD.n8046 54.6255
R4866 VDD.n4629 VDD.n4628 52.6902
R4867 VDD.n5161 VDD.n5160 52.6902
R4868 VDD.n5311 VDD.n5310 52.6902
R4869 VDD.n8615 VDD.n8614 52.6902
R4870 VDD.n8977 VDD.n8976 52.6902
R4871 VDD.n8887 VDD.n8886 52.6902
R4872 VDD.n8063 VDD.n8062 51.067
R4873 VDD.n8076 VDD.n8075 51.067
R4874 VDD.n8092 VDD.n8091 51.0665
R4875 VDD.n8106 VDD.n8105 51.0665
R4876 VDD.n8120 VDD.n8119 51.0665
R4877 VDD.n8139 VDD.n8138 51.0665
R4878 VDD.n7617 VDD.n7616 51.0664
R4879 VDD.n7624 VDD.n7622 51.0664
R4880 VDD.n7627 VDD.n7625 51.0664
R4881 VDD.n7630 VDD.n7628 51.0664
R4882 VDD.n7630 VDD.n7629 51.0664
R4883 VDD.n7627 VDD.n7626 51.0664
R4884 VDD.n7624 VDD.n7623 51.0664
R4885 VDD.n1902 VDD.n1901 50.7006
R4886 VDD.n2399 VDD.n2022 50.7006
R4887 VDD.n2300 VDD.n2013 50.7006
R4888 VDD.n1048 VDD.n1047 50.7006
R4889 VDD.n1545 VDD.n1168 50.7006
R4890 VDD.n1446 VDD.n1159 50.7006
R4891 VDD.n193 VDD.n192 50.7006
R4892 VDD.n690 VDD.n313 50.7006
R4893 VDD.n591 VDD.n304 50.7006
R4894 VDD.n8549 VDD.n8547 50.6999
R4895 VDD.n1874 VDD.n1873 50.6999
R4896 VDD.n2535 VDD.n1809 50.6999
R4897 VDD.n2535 VDD.n2534 50.6999
R4898 VDD.n2177 VDD.n2173 50.6999
R4899 VDD.n2175 VDD.n2174 50.6999
R4900 VDD.n2401 VDD.n2003 50.6999
R4901 VDD.n2381 VDD.n2016 50.6999
R4902 VDD.n1020 VDD.n1019 50.6999
R4903 VDD.n1681 VDD.n955 50.6999
R4904 VDD.n1681 VDD.n1680 50.6999
R4905 VDD.n1323 VDD.n1319 50.6999
R4906 VDD.n1321 VDD.n1320 50.6999
R4907 VDD.n1547 VDD.n1149 50.6999
R4908 VDD.n1527 VDD.n1162 50.6999
R4909 VDD.n165 VDD.n164 50.6999
R4910 VDD.n826 VDD.n100 50.6999
R4911 VDD.n826 VDD.n825 50.6999
R4912 VDD.n468 VDD.n464 50.6999
R4913 VDD.n466 VDD.n465 50.6999
R4914 VDD.n692 VDD.n294 50.6999
R4915 VDD.n672 VDD.n307 50.6999
R4916 VDD.n3183 VDD.n3182 49.0945
R4917 VDD.n3188 VDD.n3187 49.0945
R4918 VDD.n3387 VDD.n3386 49.0945
R4919 VDD.n3390 VDD.n3389 49.0945
R4920 VDD.n3393 VDD.n3392 49.0945
R4921 VDD.n2650 VDD.n2649 49.0945
R4922 VDD.n2653 VDD.n2652 49.0945
R4923 VDD.n2656 VDD.n2655 49.0945
R4924 VDD.n2339 VDD.n2338 49.0945
R4925 VDD.n2342 VDD.n2333 49.0945
R4926 VDD.n2344 VDD.n2343 49.0945
R4927 VDD.n1914 VDD.n1831 49.0945
R4928 VDD.n1911 VDD.n1830 49.0945
R4929 VDD.n1914 VDD.n1830 49.0945
R4930 VDD.n1832 VDD.n1831 49.0945
R4931 VDD.n1890 VDD.n1889 49.0945
R4932 VDD.n1886 VDD.n1879 49.0945
R4933 VDD.n1885 VDD.n1884 49.0945
R4934 VDD.n1886 VDD.n1885 49.0945
R4935 VDD.n1889 VDD.n1879 49.0945
R4936 VDD.n1891 VDD.n1890 49.0945
R4937 VDD.n2343 VDD.n2342 49.0945
R4938 VDD.n2339 VDD.n2333 49.0945
R4939 VDD.n2338 VDD.n2337 49.0945
R4940 VDD.n1485 VDD.n1484 49.0945
R4941 VDD.n1488 VDD.n1479 49.0945
R4942 VDD.n1490 VDD.n1489 49.0945
R4943 VDD.n1060 VDD.n977 49.0945
R4944 VDD.n1057 VDD.n976 49.0945
R4945 VDD.n1060 VDD.n976 49.0945
R4946 VDD.n978 VDD.n977 49.0945
R4947 VDD.n1036 VDD.n1035 49.0945
R4948 VDD.n1032 VDD.n1025 49.0945
R4949 VDD.n1031 VDD.n1030 49.0945
R4950 VDD.n1032 VDD.n1031 49.0945
R4951 VDD.n1035 VDD.n1025 49.0945
R4952 VDD.n1037 VDD.n1036 49.0945
R4953 VDD.n1489 VDD.n1488 49.0945
R4954 VDD.n1485 VDD.n1479 49.0945
R4955 VDD.n1484 VDD.n1483 49.0945
R4956 VDD.n630 VDD.n629 49.0945
R4957 VDD.n633 VDD.n624 49.0945
R4958 VDD.n635 VDD.n634 49.0945
R4959 VDD.n205 VDD.n122 49.0945
R4960 VDD.n202 VDD.n121 49.0945
R4961 VDD.n205 VDD.n121 49.0945
R4962 VDD.n123 VDD.n122 49.0945
R4963 VDD.n181 VDD.n180 49.0945
R4964 VDD.n177 VDD.n170 49.0945
R4965 VDD.n176 VDD.n175 49.0945
R4966 VDD.n177 VDD.n176 49.0945
R4967 VDD.n180 VDD.n170 49.0945
R4968 VDD.n182 VDD.n181 49.0945
R4969 VDD.n634 VDD.n633 49.0945
R4970 VDD.n630 VDD.n624 49.0945
R4971 VDD.n629 VDD.n628 49.0945
R4972 VDD.n3957 VDD.n3956 49.0838
R4973 VDD.n3959 VDD.n3958 49.0838
R4974 VDD.n3964 VDD.n3963 49.0838
R4975 VDD.n3962 VDD.n3961 49.0838
R4976 VDD.n3425 VDD.n3424 48.3613
R4977 VDD.n1926 VDD.n1925 48.0774
R4978 VDD.n1072 VDD.n1071 48.0774
R4979 VDD.n217 VDD.n216 48.0774
R4980 VDD.n3469 VDD.n3467 46.4193
R4981 VDD.n4640 VDD.n4639 46.104
R4982 VDD.n5172 VDD.n5171 46.104
R4983 VDD.n4293 VDD.n4292 46.104
R4984 VDD.n5322 VDD.n5321 46.104
R4985 VDD.n8626 VDD.n8625 46.104
R4986 VDD.n8988 VDD.n8987 46.104
R4987 VDD.n8898 VDD.n8897 46.104
R4988 VDD.n4674 VDD.n4673 44.9671
R4989 VDD.n5214 VDD.n5213 44.9671
R4990 VDD.n7129 VDD.n7128 44.7682
R4991 VDD.n4011 VDD.n4010 44.7682
R4992 VDD.n1902 VDD.n1810 44.7682
R4993 VDD.n2400 VDD.n2013 44.7682
R4994 VDD.n2400 VDD.n2399 44.7682
R4995 VDD.n1048 VDD.n956 44.7682
R4996 VDD.n1546 VDD.n1159 44.7682
R4997 VDD.n1546 VDD.n1545 44.7682
R4998 VDD.n193 VDD.n101 44.7682
R4999 VDD.n691 VDD.n304 44.7682
R5000 VDD.n691 VDD.n690 44.7682
R5001 VDD.n8568 VDD.n8549 44.768
R5002 VDD.n7498 VDD.n7497 44.768
R5003 VDD.n4011 VDD.n3975 44.768
R5004 VDD.n8568 VDD.n8567 44.768
R5005 VDD.n2724 VDD.n2723 44.768
R5006 VDD.n1873 VDD.n1810 44.768
R5007 VDD.n1810 VDD.n1809 44.768
R5008 VDD.n2534 VDD.n1810 44.768
R5009 VDD.n2173 VDD.n2038 44.768
R5010 VDD.n2174 VDD.n2038 44.768
R5011 VDD.n2401 VDD.n2400 44.768
R5012 VDD.n2400 VDD.n2016 44.768
R5013 VDD.n1019 VDD.n956 44.768
R5014 VDD.n956 VDD.n955 44.768
R5015 VDD.n1680 VDD.n956 44.768
R5016 VDD.n1319 VDD.n1184 44.768
R5017 VDD.n1320 VDD.n1184 44.768
R5018 VDD.n1547 VDD.n1546 44.768
R5019 VDD.n1546 VDD.n1162 44.768
R5020 VDD.n164 VDD.n101 44.768
R5021 VDD.n101 VDD.n100 44.768
R5022 VDD.n825 VDD.n101 44.768
R5023 VDD.n464 VDD.n329 44.768
R5024 VDD.n465 VDD.n329 44.768
R5025 VDD.n692 VDD.n691 44.768
R5026 VDD.n691 VDD.n307 44.768
R5027 VDD.n1936 VDD.n1822 43.5902
R5028 VDD.n1082 VDD.n968 43.5902
R5029 VDD.n227 VDD.n113 43.5902
R5030 VDD.n3259 VDD.n3257 41.7887
R5031 VDD.n2862 VDD.n2860 41.7887
R5032 VDD.n2496 VDD.n2495 41.7887
R5033 VDD.n2437 VDD.n2436 41.7887
R5034 VDD.n1642 VDD.n1641 41.7887
R5035 VDD.n1583 VDD.n1582 41.7887
R5036 VDD.n787 VDD.n786 41.7887
R5037 VDD.n728 VDD.n727 41.7887
R5038 VDD.n3618 VDD.n3617 41.7222
R5039 VDD.n3397 VDD.n3396 41.6217
R5040 VDD.n2661 VDD.n2660 41.6217
R5041 VDD.n1924 VDD.n1923 41.6217
R5042 VDD.n1892 VDD.n1803 41.6217
R5043 VDD.n2336 VDD.n2245 41.6217
R5044 VDD.n1070 VDD.n1069 41.6217
R5045 VDD.n1038 VDD.n949 41.6217
R5046 VDD.n1482 VDD.n1391 41.6217
R5047 VDD.n215 VDD.n214 41.6217
R5048 VDD.n183 VDD.n94 41.6217
R5049 VDD.n627 VDD.n536 41.6217
R5050 VDD.n3194 VDD.n3193 41.6215
R5051 VDD.n2660 VDD.n2659 41.6215
R5052 VDD.n1924 VDD.n1829 41.6215
R5053 VDD.n1883 VDD.n1803 41.6215
R5054 VDD.n2345 VDD.n2245 41.6215
R5055 VDD.n1070 VDD.n975 41.6215
R5056 VDD.n1029 VDD.n949 41.6215
R5057 VDD.n1491 VDD.n1391 41.6215
R5058 VDD.n215 VDD.n120 41.6215
R5059 VDD.n174 VDD.n94 41.6215
R5060 VDD.n636 VDD.n536 41.6215
R5061 VDD.n7561 VDD.n7560 40.8219
R5062 VDD.n7554 VDD.n7553 40.8219
R5063 VDD.n7549 VDD.n7548 40.8219
R5064 VDD.n7544 VDD.n7543 40.8219
R5065 VDD.n7539 VDD.n7538 40.8219
R5066 VDD.n7534 VDD.n7532 40.8219
R5067 VDD.n7508 VDD.n7507 40.8219
R5068 VDD.n7513 VDD.n7512 40.8219
R5069 VDD.n7518 VDD.n7517 40.8219
R5070 VDD.n7523 VDD.n7522 40.8219
R5071 VDD.n7528 VDD.n7527 40.8219
R5072 VDD.n7534 VDD.n7533 40.8219
R5073 VDD.n2721 VDD.n2720 40.8219
R5074 VDD.n2776 VDD.n2775 40.8219
R5075 VDD.n2781 VDD.n2780 40.8219
R5076 VDD.n2787 VDD.n2786 40.8219
R5077 VDD.n2792 VDD.n2791 40.8219
R5078 VDD.n2798 VDD.n2797 40.8219
R5079 VDD.n3384 VDD.n3383 40.8219
R5080 VDD.n3210 VDD.n3209 40.8219
R5081 VDD.n2968 VDD.n2967 40.8219
R5082 VDD.n2965 VDD.n2964 40.8219
R5083 VDD.n2959 VDD.n2958 40.8219
R5084 VDD.n2954 VDD.n2953 40.8219
R5085 VDD.n2948 VDD.n2947 40.8219
R5086 VDD.n2943 VDD.n2942 40.8219
R5087 VDD.n2937 VDD.n2936 40.8219
R5088 VDD.n2932 VDD.n2931 40.8219
R5089 VDD.n2176 VDD.n2175 40.8219
R5090 VDD.n2393 VDD.n2021 40.8219
R5091 VDD.n2215 VDD.n2020 40.8219
R5092 VDD.n2226 VDD.n2019 40.8219
R5093 VDD.n2384 VDD.n2018 40.8219
R5094 VDD.n2381 VDD.n2017 40.8219
R5095 VDD.n2302 VDD.n2012 40.8219
R5096 VDD.n2306 VDD.n2011 40.8219
R5097 VDD.n2290 VDD.n2010 40.8219
R5098 VDD.n2312 VDD.n2009 40.8219
R5099 VDD.n2288 VDD.n2008 40.8219
R5100 VDD.n2318 VDD.n2007 40.8219
R5101 VDD.n2321 VDD.n2006 40.8219
R5102 VDD.n2005 VDD.n2003 40.8219
R5103 VDD.n1877 VDD.n1876 40.8219
R5104 VDD.n1875 VDD.n1874 40.8219
R5105 VDD.n1876 VDD.n1875 40.8219
R5106 VDD.n1901 VDD.n1877 40.8219
R5107 VDD.n2177 VDD.n2176 40.8219
R5108 VDD.n2300 VDD.n2012 40.8219
R5109 VDD.n2302 VDD.n2011 40.8219
R5110 VDD.n2306 VDD.n2010 40.8219
R5111 VDD.n2290 VDD.n2009 40.8219
R5112 VDD.n2312 VDD.n2008 40.8219
R5113 VDD.n2288 VDD.n2007 40.8219
R5114 VDD.n2318 VDD.n2006 40.8219
R5115 VDD.n2321 VDD.n2005 40.8219
R5116 VDD.n2022 VDD.n2021 40.8219
R5117 VDD.n2393 VDD.n2020 40.8219
R5118 VDD.n2215 VDD.n2019 40.8219
R5119 VDD.n2226 VDD.n2018 40.8219
R5120 VDD.n2384 VDD.n2017 40.8219
R5121 VDD.n1322 VDD.n1321 40.8219
R5122 VDD.n1539 VDD.n1167 40.8219
R5123 VDD.n1361 VDD.n1166 40.8219
R5124 VDD.n1372 VDD.n1165 40.8219
R5125 VDD.n1530 VDD.n1164 40.8219
R5126 VDD.n1527 VDD.n1163 40.8219
R5127 VDD.n1448 VDD.n1158 40.8219
R5128 VDD.n1452 VDD.n1157 40.8219
R5129 VDD.n1436 VDD.n1156 40.8219
R5130 VDD.n1458 VDD.n1155 40.8219
R5131 VDD.n1434 VDD.n1154 40.8219
R5132 VDD.n1464 VDD.n1153 40.8219
R5133 VDD.n1467 VDD.n1152 40.8219
R5134 VDD.n1151 VDD.n1149 40.8219
R5135 VDD.n1023 VDD.n1022 40.8219
R5136 VDD.n1021 VDD.n1020 40.8219
R5137 VDD.n1022 VDD.n1021 40.8219
R5138 VDD.n1047 VDD.n1023 40.8219
R5139 VDD.n1323 VDD.n1322 40.8219
R5140 VDD.n1446 VDD.n1158 40.8219
R5141 VDD.n1448 VDD.n1157 40.8219
R5142 VDD.n1452 VDD.n1156 40.8219
R5143 VDD.n1436 VDD.n1155 40.8219
R5144 VDD.n1458 VDD.n1154 40.8219
R5145 VDD.n1434 VDD.n1153 40.8219
R5146 VDD.n1464 VDD.n1152 40.8219
R5147 VDD.n1467 VDD.n1151 40.8219
R5148 VDD.n1168 VDD.n1167 40.8219
R5149 VDD.n1539 VDD.n1166 40.8219
R5150 VDD.n1361 VDD.n1165 40.8219
R5151 VDD.n1372 VDD.n1164 40.8219
R5152 VDD.n1530 VDD.n1163 40.8219
R5153 VDD.n467 VDD.n466 40.8219
R5154 VDD.n684 VDD.n312 40.8219
R5155 VDD.n506 VDD.n311 40.8219
R5156 VDD.n517 VDD.n310 40.8219
R5157 VDD.n675 VDD.n309 40.8219
R5158 VDD.n672 VDD.n308 40.8219
R5159 VDD.n593 VDD.n303 40.8219
R5160 VDD.n597 VDD.n302 40.8219
R5161 VDD.n581 VDD.n301 40.8219
R5162 VDD.n603 VDD.n300 40.8219
R5163 VDD.n579 VDD.n299 40.8219
R5164 VDD.n609 VDD.n298 40.8219
R5165 VDD.n612 VDD.n297 40.8219
R5166 VDD.n296 VDD.n294 40.8219
R5167 VDD.n168 VDD.n167 40.8219
R5168 VDD.n166 VDD.n165 40.8219
R5169 VDD.n167 VDD.n166 40.8219
R5170 VDD.n192 VDD.n168 40.8219
R5171 VDD.n468 VDD.n467 40.8219
R5172 VDD.n591 VDD.n303 40.8219
R5173 VDD.n593 VDD.n302 40.8219
R5174 VDD.n597 VDD.n301 40.8219
R5175 VDD.n581 VDD.n300 40.8219
R5176 VDD.n603 VDD.n299 40.8219
R5177 VDD.n579 VDD.n298 40.8219
R5178 VDD.n609 VDD.n297 40.8219
R5179 VDD.n612 VDD.n296 40.8219
R5180 VDD.n313 VDD.n312 40.8219
R5181 VDD.n684 VDD.n311 40.8219
R5182 VDD.n506 VDD.n310 40.8219
R5183 VDD.n517 VDD.n309 40.8219
R5184 VDD.n675 VDD.n308 40.8219
R5185 VDD.n4651 VDD.n4650 39.5177
R5186 VDD.n5183 VDD.n5182 39.5177
R5187 VDD.n4309 VDD.n4308 39.5177
R5188 VDD.n5338 VDD.n5337 39.5177
R5189 VDD.n8605 VDD.n8604 39.5177
R5190 VDD.n8967 VDD.n8966 39.5177
R5191 VDD.n8908 VDD.n8907 39.5177
R5192 VDD.n4016 VDD.n3954 39.2068
R5193 VDD.n3379 VDD.n3376 38.7994
R5194 VDD.n3357 VDD.n3356 38.7994
R5195 VDD.n3347 VDD.n3346 38.7994
R5196 VDD.n2282 VDD.n2259 38.7994
R5197 VDD.n2277 VDD.n2258 38.7994
R5198 VDD.n2274 VDD.n2257 38.7994
R5199 VDD.n2391 VDD.n2390 38.7994
R5200 VDD.n1933 VDD.n1932 38.7994
R5201 VDD.n1867 VDD.n1843 38.7994
R5202 VDD.n1866 VDD.n1844 38.7994
R5203 VDD.n1858 VDD.n1857 38.7994
R5204 VDD.n1428 VDD.n1405 38.7994
R5205 VDD.n1423 VDD.n1404 38.7994
R5206 VDD.n1420 VDD.n1403 38.7994
R5207 VDD.n1537 VDD.n1536 38.7994
R5208 VDD.n1079 VDD.n1078 38.7994
R5209 VDD.n1013 VDD.n989 38.7994
R5210 VDD.n1012 VDD.n990 38.7994
R5211 VDD.n1004 VDD.n1003 38.7994
R5212 VDD.n573 VDD.n550 38.7994
R5213 VDD.n568 VDD.n549 38.7994
R5214 VDD.n565 VDD.n548 38.7994
R5215 VDD.n682 VDD.n681 38.7994
R5216 VDD.n224 VDD.n223 38.7994
R5217 VDD.n158 VDD.n134 38.7994
R5218 VDD.n157 VDD.n135 38.7994
R5219 VDD.n149 VDD.n148 38.7994
R5220 VDD.n2637 VDD.n2636 38.7989
R5221 VDD.n2645 VDD.n2643 38.7989
R5222 VDD.n2784 VDD.n2783 38.7989
R5223 VDD.n3379 VDD.n3378 38.7989
R5224 VDD.n3368 VDD.n3367 38.7989
R5225 VDD.n2275 VDD.n2258 38.7989
R5226 VDD.n2271 VDD.n2257 38.7989
R5227 VDD.n2282 VDD.n2281 38.7989
R5228 VDD.n2390 VDD.n2218 38.7989
R5229 VDD.n1933 VDD.n1823 38.7989
R5230 VDD.n1857 VDD.n1821 38.7989
R5231 VDD.n1856 VDD.n1844 38.7989
R5232 VDD.n1843 VDD.n1824 38.7989
R5233 VDD.n1421 VDD.n1404 38.7989
R5234 VDD.n1417 VDD.n1403 38.7989
R5235 VDD.n1428 VDD.n1427 38.7989
R5236 VDD.n1536 VDD.n1364 38.7989
R5237 VDD.n1079 VDD.n969 38.7989
R5238 VDD.n1003 VDD.n967 38.7989
R5239 VDD.n1002 VDD.n990 38.7989
R5240 VDD.n989 VDD.n970 38.7989
R5241 VDD.n566 VDD.n549 38.7989
R5242 VDD.n562 VDD.n548 38.7989
R5243 VDD.n573 VDD.n572 38.7989
R5244 VDD.n681 VDD.n509 38.7989
R5245 VDD.n224 VDD.n114 38.7989
R5246 VDD.n148 VDD.n112 38.7989
R5247 VDD.n147 VDD.n135 38.7989
R5248 VDD.n134 VDD.n115 38.7989
R5249 VDD.n2795 VDD.n2794 38.7987
R5250 VDD.n2807 VDD.n2806 38.7987
R5251 VDD.n2940 VDD.n2939 38.7987
R5252 VDD.n2951 VDD.n2950 38.7987
R5253 VDD.n2962 VDD.n2961 38.7987
R5254 VDD.n2388 VDD.n2224 38.7987
R5255 VDD.n2375 VDD.n2223 38.7987
R5256 VDD.n2388 VDD.n2387 38.7987
R5257 VDD.n2379 VDD.n2223 38.7987
R5258 VDD.n2309 VDD.n2222 38.7987
R5259 VDD.n2315 VDD.n2221 38.7987
R5260 VDD.n2324 VDD.n2220 38.7987
R5261 VDD.n2316 VDD.n2220 38.7987
R5262 VDD.n2310 VDD.n2221 38.7987
R5263 VDD.n2304 VDD.n2222 38.7987
R5264 VDD.n1534 VDD.n1370 38.7987
R5265 VDD.n1521 VDD.n1369 38.7987
R5266 VDD.n1534 VDD.n1533 38.7987
R5267 VDD.n1525 VDD.n1369 38.7987
R5268 VDD.n1455 VDD.n1368 38.7987
R5269 VDD.n1461 VDD.n1367 38.7987
R5270 VDD.n1470 VDD.n1366 38.7987
R5271 VDD.n1462 VDD.n1366 38.7987
R5272 VDD.n1456 VDD.n1367 38.7987
R5273 VDD.n1450 VDD.n1368 38.7987
R5274 VDD.n679 VDD.n515 38.7987
R5275 VDD.n666 VDD.n514 38.7987
R5276 VDD.n679 VDD.n678 38.7987
R5277 VDD.n670 VDD.n514 38.7987
R5278 VDD.n600 VDD.n513 38.7987
R5279 VDD.n606 VDD.n512 38.7987
R5280 VDD.n615 VDD.n511 38.7987
R5281 VDD.n607 VDD.n511 38.7987
R5282 VDD.n601 VDD.n512 38.7987
R5283 VDD.n595 VDD.n513 38.7987
R5284 VDD.n7619 VDD.n7618 38.777
R5285 VDD.n2373 VDD.n2372 36.539
R5286 VDD.n2365 VDD.n2238 36.539
R5287 VDD.n1519 VDD.n1518 36.539
R5288 VDD.n1511 VDD.n1384 36.539
R5289 VDD.n664 VDD.n663 36.539
R5290 VDD.n656 VDD.n529 36.539
R5291 VDD.n5287 VDD.n5286 36.2246
R5292 VDD.n54 VDD.n38 36.1417
R5293 VDD.n54 VDD.n53 36.1417
R5294 VDD.n53 VDD.n42 36.1417
R5295 VDD.n49 VDD.n42 36.1417
R5296 VDD.n19 VDD.n11 36.1417
R5297 VDD.n30 VDD.n11 36.1417
R5298 VDD.n30 VDD.n7 36.1417
R5299 VDD.n61 VDD.n7 36.1417
R5300 VDD.n905 VDD.n900 36.1417
R5301 VDD.n905 VDD.n904 36.1417
R5302 VDD.n904 VDD.n859 36.1417
R5303 VDD.n910 VDD.n859 36.1417
R5304 VDD.n877 VDD.n868 36.1417
R5305 VDD.n882 VDD.n868 36.1417
R5306 VDD.n882 VDD.n863 36.1417
R5307 VDD.n893 VDD.n863 36.1417
R5308 VDD.n1763 VDD.n1747 36.1417
R5309 VDD.n1763 VDD.n1762 36.1417
R5310 VDD.n1762 VDD.n1751 36.1417
R5311 VDD.n1758 VDD.n1751 36.1417
R5312 VDD.n1728 VDD.n1720 36.1417
R5313 VDD.n1739 VDD.n1720 36.1417
R5314 VDD.n1739 VDD.n1716 36.1417
R5315 VDD.n1770 VDD.n1716 36.1417
R5316 VDD.n2598 VDD.n2595 36.1417
R5317 VDD.n3255 VDD.n3254 35.9626
R5318 VDD.n2491 VDD.n2490 35.9626
R5319 VDD.n1637 VDD.n1636 35.9626
R5320 VDD.n782 VDD.n781 35.9626
R5321 VDD.n2814 VDD.n2813 35.2569
R5322 VDD.n2400 VDD.n2004 35.2569
R5323 VDD.n1546 VDD.n1150 35.2569
R5324 VDD.n691 VDD.n295 35.2569
R5325 VDD.n6499 VDD.n6498 34.6359
R5326 VDD.n3202 VDD.n3201 34.6159
R5327 VDD.n2530 VDD.n1810 34.6159
R5328 VDD.n1676 VDD.n956 34.6159
R5329 VDD.n821 VDD.n101 34.6159
R5330 VDD.n7119 VDD.n7116 34.3808
R5331 VDD.n5844 VDD.n5843 34.3388
R5332 VDD.n7576 VDD.n7572 34.2989
R5333 VDD.n8051 VDD.n8049 33.9026
R5334 VDD.n8564 VDD.n8560 33.8536
R5335 VDD.n8552 VDD.n8550 33.4435
R5336 VDD.n8555 VDD.n8553 33.4435
R5337 VDD.n8060 VDD.n8059 33.4435
R5338 VDD.n8130 VDD.n8129 33.4435
R5339 VDD.n8049 VDD.n8045 33.4435
R5340 VDD.n7572 VDD.n7569 33.4435
R5341 VDD.n5843 VDD.n5840 33.4435
R5342 VDD.n7116 VDD.n7112 33.4435
R5343 VDD.n2867 VDD.n2866 33.4435
R5344 VDD.n3264 VDD.n3263 33.4435
R5345 VDD.n3364 VDD.n3363 33.4435
R5346 VDD.n3354 VDD.n3353 33.4435
R5347 VDD.n3344 VDD.n3343 33.4435
R5348 VDD.n2713 VDD.n2710 33.4435
R5349 VDD.n1989 VDD.n1986 33.4435
R5350 VDD.n2500 VDD.n2499 33.4435
R5351 VDD.n1850 VDD.n1816 33.4435
R5352 VDD.n1846 VDD.n1841 33.4435
R5353 VDD.n1863 VDD.n1862 33.4435
R5354 VDD.n1849 VDD.n1848 33.4435
R5355 VDD.n1919 VDD.n1918 33.4435
R5356 VDD.n1838 VDD.n1835 33.4435
R5357 VDD.n1908 VDD.n1839 33.4435
R5358 VDD.n2071 VDD.n2069 33.4435
R5359 VDD.n2113 VDD.n2112 33.4435
R5360 VDD.n2182 VDD.n2181 33.4435
R5361 VDD.n1135 VDD.n1132 33.4435
R5362 VDD.n1646 VDD.n1645 33.4435
R5363 VDD.n996 VDD.n962 33.4435
R5364 VDD.n992 VDD.n987 33.4435
R5365 VDD.n1009 VDD.n1008 33.4435
R5366 VDD.n995 VDD.n994 33.4435
R5367 VDD.n1065 VDD.n1064 33.4435
R5368 VDD.n984 VDD.n981 33.4435
R5369 VDD.n1054 VDD.n985 33.4435
R5370 VDD.n1217 VDD.n1215 33.4435
R5371 VDD.n1259 VDD.n1258 33.4435
R5372 VDD.n1328 VDD.n1327 33.4435
R5373 VDD.n280 VDD.n277 33.4435
R5374 VDD.n791 VDD.n790 33.4435
R5375 VDD.n141 VDD.n107 33.4435
R5376 VDD.n137 VDD.n132 33.4435
R5377 VDD.n154 VDD.n153 33.4435
R5378 VDD.n140 VDD.n139 33.4435
R5379 VDD.n210 VDD.n209 33.4435
R5380 VDD.n129 VDD.n126 33.4435
R5381 VDD.n199 VDD.n130 33.4435
R5382 VDD.n362 VDD.n360 33.4435
R5383 VDD.n404 VDD.n403 33.4435
R5384 VDD.n473 VDD.n472 33.4435
R5385 VDD.n6498 VDD.n6496 33.4431
R5386 VDD.n8552 VDD.n8551 33.4431
R5387 VDD.n8555 VDD.n8554 33.4431
R5388 VDD.n8079 VDD.n8078 33.4431
R5389 VDD.n8095 VDD.n8094 33.4431
R5390 VDD.n8109 VDD.n8108 33.4431
R5391 VDD.n8123 VDD.n8122 33.4431
R5392 VDD.n7572 VDD.n7571 33.4431
R5393 VDD.n5843 VDD.n5842 33.4431
R5394 VDD.n7116 VDD.n7115 33.4431
R5395 VDD.n3337 VDD.n3336 33.4431
R5396 VDD.n3204 VDD.n3203 33.4431
R5397 VDD.n3191 VDD.n3190 33.4431
R5398 VDD.n3180 VDD.n3179 33.4431
R5399 VDD.n3119 VDD.n3118 33.4431
R5400 VDD.n3113 VDD.n3112 33.4431
R5401 VDD.n2713 VDD.n2712 33.4431
R5402 VDD.n1986 VDD.n1985 33.4431
R5403 VDD.n2499 VDD.n2498 33.4431
R5404 VDD.n1851 VDD.n1850 33.4431
R5405 VDD.n1852 VDD.n1849 33.4431
R5406 VDD.n1862 VDD.n1861 33.4431
R5407 VDD.n1847 VDD.n1846 33.4431
R5408 VDD.n1904 VDD.n1839 33.4431
R5409 VDD.n1909 VDD.n1838 33.4431
R5410 VDD.n1918 VDD.n1917 33.4431
R5411 VDD.n2112 VDD.n2111 33.4431
R5412 VDD.n2114 VDD.n2071 33.4431
R5413 VDD.n2181 VDD.n2041 33.4431
R5414 VDD.n1132 VDD.n1131 33.4431
R5415 VDD.n1645 VDD.n1644 33.4431
R5416 VDD.n997 VDD.n996 33.4431
R5417 VDD.n998 VDD.n995 33.4431
R5418 VDD.n1008 VDD.n1007 33.4431
R5419 VDD.n993 VDD.n992 33.4431
R5420 VDD.n1050 VDD.n985 33.4431
R5421 VDD.n1055 VDD.n984 33.4431
R5422 VDD.n1064 VDD.n1063 33.4431
R5423 VDD.n1258 VDD.n1257 33.4431
R5424 VDD.n1260 VDD.n1217 33.4431
R5425 VDD.n1327 VDD.n1187 33.4431
R5426 VDD.n277 VDD.n276 33.4431
R5427 VDD.n790 VDD.n789 33.4431
R5428 VDD.n142 VDD.n141 33.4431
R5429 VDD.n143 VDD.n140 33.4431
R5430 VDD.n153 VDD.n152 33.4431
R5431 VDD.n138 VDD.n137 33.4431
R5432 VDD.n195 VDD.n130 33.4431
R5433 VDD.n200 VDD.n129 33.4431
R5434 VDD.n209 VDD.n208 33.4431
R5435 VDD.n403 VDD.n402 33.4431
R5436 VDD.n405 VDD.n362 33.4431
R5437 VDD.n472 VDD.n332 33.4431
R5438 VDD.n6463 VDD.n6462 33.4428
R5439 VDD.n6452 VDD.n6451 33.4428
R5440 VDD.n6443 VDD.n6442 33.4428
R5441 VDD.n6434 VDD.n6433 33.4428
R5442 VDD.n6425 VDD.n6424 33.4428
R5443 VDD.n6384 VDD.n6383 33.4428
R5444 VDD.n6373 VDD.n6372 33.4428
R5445 VDD.n6393 VDD.n6392 33.4428
R5446 VDD.n6402 VDD.n6401 33.4428
R5447 VDD.n6411 VDD.n6410 33.4428
R5448 VDD.n6420 VDD.n6419 33.4428
R5449 VDD.n6472 VDD.n6471 33.4428
R5450 VDD.n6481 VDD.n6480 33.4428
R5451 VDD.n6490 VDD.n6489 33.4428
R5452 VDD.n2816 VDD.n2815 33.4428
R5453 VDD.n2297 VDD.n2014 33.4428
R5454 VDD.n2294 VDD.n2014 33.4428
R5455 VDD.n1443 VDD.n1160 33.4428
R5456 VDD.n1440 VDD.n1160 33.4428
R5457 VDD.n588 VDD.n305 33.4428
R5458 VDD.n585 VDD.n305 33.4428
R5459 VDD.n2858 VDD.n2857 32.9658
R5460 VDD.n2433 VDD.n1982 32.9658
R5461 VDD.n1579 VDD.n1128 32.9658
R5462 VDD.n724 VDD.n273 32.9658
R5463 VDD.n4621 VDD.n4620 32.9315
R5464 VDD.n5197 VDD.n5196 32.9315
R5465 VDD.n5257 VDD.n5256 32.9315
R5466 VDD.n8642 VDD.n8641 32.9315
R5467 VDD.n9005 VDD.n9004 32.9315
R5468 VDD.n8921 VDD.n8920 32.9315
R5469 VDD.n2714 VDD.n2713 32.6607
R5470 VDD.n2181 VDD.n2180 32.6607
R5471 VDD.n1327 VDD.n1326 32.6607
R5472 VDD.n472 VDD.n471 32.6607
R5473 VDD.n1926 VDD.n1924 30.1287
R5474 VDD.n1072 VDD.n1070 30.1287
R5475 VDD.n217 VDD.n215 30.1287
R5476 VDD.n3051 VDD.n3046 30.1181
R5477 VDD.n3403 VDD.n3399 30.1181
R5478 VDD.n3326 VDD.n3315 30.1181
R5479 VDD.n3001 VDD.n2663 30.1181
R5480 VDD.n2919 VDD.n2918 30.1181
R5481 VDD.n2280 VDD.n2267 30.1181
R5482 VDD.n1895 VDD.n1894 30.1181
R5483 VDD.n1881 VDD.n1792 30.1181
R5484 VDD.n2356 VDD.n2248 30.1181
R5485 VDD.n2348 VDD.n2347 30.1181
R5486 VDD.n1426 VDD.n1413 30.1181
R5487 VDD.n1041 VDD.n1040 30.1181
R5488 VDD.n1027 VDD.n938 30.1181
R5489 VDD.n1502 VDD.n1394 30.1181
R5490 VDD.n1494 VDD.n1493 30.1181
R5491 VDD.n571 VDD.n558 30.1181
R5492 VDD.n186 VDD.n185 30.1181
R5493 VDD.n172 VDD.n83 30.1181
R5494 VDD.n647 VDD.n539 30.1181
R5495 VDD.n639 VDD.n638 30.1181
R5496 VDD.n3173 VDD.n3172 30.0704
R5497 VDD.n3398 VDD.n3397 30.0704
R5498 VDD.n2662 VDD.n2661 30.0704
R5499 VDD.n1923 VDD.n1922 30.0704
R5500 VDD.n1893 VDD.n1892 30.0704
R5501 VDD.n2336 VDD.n2335 30.0704
R5502 VDD.n1069 VDD.n1068 30.0704
R5503 VDD.n1039 VDD.n1038 30.0704
R5504 VDD.n1482 VDD.n1481 30.0704
R5505 VDD.n214 VDD.n213 30.0704
R5506 VDD.n184 VDD.n183 30.0704
R5507 VDD.n627 VDD.n626 30.0704
R5508 VDD.n3195 VDD.n3194 30.0702
R5509 VDD.n3314 VDD.n3312 30.0702
R5510 VDD.n2346 VDD.n2345 30.0702
R5511 VDD.n1836 VDD.n1829 30.0702
R5512 VDD.n1883 VDD.n1882 30.0702
R5513 VDD.n1492 VDD.n1491 30.0702
R5514 VDD.n982 VDD.n975 30.0702
R5515 VDD.n1029 VDD.n1028 30.0702
R5516 VDD.n637 VDD.n636 30.0702
R5517 VDD.n127 VDD.n120 30.0702
R5518 VDD.n174 VDD.n173 30.0702
R5519 VDD.n4614 VDD.n4613 29.6384
R5520 VDD.n5154 VDD.n5153 29.6384
R5521 VDD.n5298 VDD.n5297 29.6384
R5522 VDD.n8662 VDD.n8661 29.6384
R5523 VDD.n8741 VDD.n8740 29.6384
R5524 VDD.n8941 VDD.n8940 29.6384
R5525 VDD.n8568 VDD.n8552 29.5303
R5526 VDD.n8568 VDD.n8555 29.5303
R5527 VDD.n8048 VDD.n8047 29.5303
R5528 VDD.n3801 VDD.n3800 29.5303
R5529 VDD.n2866 VDD.n2865 29.5303
R5530 VDD.n3263 VDD.n3262 29.5303
R5531 VDD.n3203 VDD.n3202 29.5303
R5532 VDD.n3118 VDD.n3117 29.5303
R5533 VDD.n2434 VDD.n1986 29.5303
R5534 VDD.n2499 VDD.n1954 29.5303
R5535 VDD.n1846 VDD.n1810 29.5303
R5536 VDD.n1862 VDD.n1810 29.5303
R5537 VDD.n1849 VDD.n1810 29.5303
R5538 VDD.n1850 VDD.n1810 29.5303
R5539 VDD.n1918 VDD.n1810 29.5303
R5540 VDD.n1838 VDD.n1810 29.5303
R5541 VDD.n1839 VDD.n1810 29.5303
R5542 VDD.n2072 VDD.n2071 29.5303
R5543 VDD.n2112 VDD.n2072 29.5303
R5544 VDD.n1580 VDD.n1132 29.5303
R5545 VDD.n1645 VDD.n1100 29.5303
R5546 VDD.n992 VDD.n956 29.5303
R5547 VDD.n1008 VDD.n956 29.5303
R5548 VDD.n995 VDD.n956 29.5303
R5549 VDD.n996 VDD.n956 29.5303
R5550 VDD.n1064 VDD.n956 29.5303
R5551 VDD.n984 VDD.n956 29.5303
R5552 VDD.n985 VDD.n956 29.5303
R5553 VDD.n1218 VDD.n1217 29.5303
R5554 VDD.n1258 VDD.n1218 29.5303
R5555 VDD.n725 VDD.n277 29.5303
R5556 VDD.n790 VDD.n245 29.5303
R5557 VDD.n137 VDD.n101 29.5303
R5558 VDD.n153 VDD.n101 29.5303
R5559 VDD.n140 VDD.n101 29.5303
R5560 VDD.n141 VDD.n101 29.5303
R5561 VDD.n209 VDD.n101 29.5303
R5562 VDD.n129 VDD.n101 29.5303
R5563 VDD.n130 VDD.n101 29.5303
R5564 VDD.n363 VDD.n362 29.5303
R5565 VDD.n403 VDD.n363 29.5303
R5566 VDD.n3801 VDD.n3799 29.5301
R5567 VDD.n3801 VDD.n3798 29.5301
R5568 VDD.n3801 VDD.n3797 29.5301
R5569 VDD.n3801 VDD.n3796 29.5301
R5570 VDD.n3801 VDD.n3795 29.5301
R5571 VDD.n3801 VDD.n3794 29.5301
R5572 VDD.n3801 VDD.n3793 29.5301
R5573 VDD.n3801 VDD.n3792 29.5301
R5574 VDD.n3801 VDD.n3791 29.5301
R5575 VDD.n3801 VDD.n3790 29.5301
R5576 VDD.n3801 VDD.n3789 29.5301
R5577 VDD.n3801 VDD.n3788 29.5301
R5578 VDD.n3801 VDD.n3787 29.5301
R5579 VDD.n3801 VDD.n3786 29.5301
R5580 VDD.n3801 VDD.n3785 29.5301
R5581 VDD.n3801 VDD.n3784 29.5301
R5582 VDD.n3801 VDD.n3783 29.5301
R5583 VDD.n3801 VDD.n3782 29.5301
R5584 VDD.n3801 VDD.n3781 29.5301
R5585 VDD.n3801 VDD.n3780 29.5301
R5586 VDD.n2815 VDD.n2814 29.5301
R5587 VDD.n2400 VDD.n2014 29.5301
R5588 VDD.n1546 VDD.n1160 29.5301
R5589 VDD.n691 VDD.n305 29.5301
R5590 VDD.n2553 VDD.n1787 29.4877
R5591 VDD.n2547 VDD.n1795 29.4877
R5592 VDD.n1699 VDD.n933 29.4877
R5593 VDD.n1693 VDD.n941 29.4877
R5594 VDD.n844 VDD.n78 29.4877
R5595 VDD.n838 VDD.n86 29.4877
R5596 VDD.n4240 VDD.n4239 29.4133
R5597 VDD.t19 VDD.n2244 28.8467
R5598 VDD.t154 VDD.n2285 28.8467
R5599 VDD.t104 VDD.n1796 28.8467
R5600 VDD.t8 VDD.n1390 28.8467
R5601 VDD.t148 VDD.n1431 28.8467
R5602 VDD.t149 VDD.n942 28.8467
R5603 VDD.t51 VDD.n535 28.8467
R5604 VDD.t67 VDD.n576 28.8467
R5605 VDD.t48 VDD.n87 28.8467
R5606 VDD.n3544 VDD.n3543 28.5972
R5607 VDD.n3545 VDD.n3544 28.5972
R5608 VDD.n3546 VDD.n3545 28.5972
R5609 VDD.n3547 VDD.n3546 28.5972
R5610 VDD.n3554 VDD.n3553 28.5972
R5611 VDD.n3553 VDD.n3552 28.5972
R5612 VDD.n3552 VDD.n3551 28.5972
R5613 VDD.n3551 VDD.n3550 28.5972
R5614 VDD.n3550 VDD.n3549 28.5972
R5615 VDD.n6655 VDD.n6654 28.5972
R5616 VDD.n6656 VDD.n6655 28.5972
R5617 VDD.n6657 VDD.n6656 28.5972
R5618 VDD.n6658 VDD.n6657 28.5972
R5619 VDD.n6659 VDD.n6658 28.5972
R5620 VDD.n6666 VDD.n6665 28.5972
R5621 VDD.n6665 VDD.n6664 28.5972
R5622 VDD.n6664 VDD.n6663 28.5972
R5623 VDD.n6663 VDD.n6662 28.5972
R5624 VDD.n6662 VDD.n6661 28.5972
R5625 VDD.n6661 VDD.n6660 28.5972
R5626 VDD.n8781 VDD.n8780 28.5972
R5627 VDD.n8782 VDD.n8781 28.5972
R5628 VDD.n8783 VDD.n8782 28.5972
R5629 VDD.n8784 VDD.n8783 28.5972
R5630 VDD.n8838 VDD.n8837 28.5972
R5631 VDD.n8837 VDD.n8836 28.5972
R5632 VDD.n8836 VDD.n8835 28.5972
R5633 VDD.n8785 VDD.n8784 28.1767
R5634 VDD.n58 VDD.t27 28.1564
R5635 VDD.t145 VDD.n896 28.1564
R5636 VDD.n1767 VDD.t157 28.1564
R5637 VDD.t106 VDD.n2614 28.1564
R5638 VDD.n3065 VDD.n3064 28.0793
R5639 VDD.n2119 VDD.n2068 28.0793
R5640 VDD.n1265 VDD.n1214 28.0793
R5641 VDD.n410 VDD.n359 28.0793
R5642 VDD.n2632 VDD.t118 27.6955
R5643 VDD.n2632 VDD.t120 27.6955
R5644 VDD.n2631 VDD.t123 27.6955
R5645 VDD.n2631 VDD.t122 27.6955
R5646 VDD.n1780 VDD.t18 27.6955
R5647 VDD.n1780 VDD.t20 27.6955
R5648 VDD.n1779 VDD.t36 27.6955
R5649 VDD.n1779 VDD.t105 27.6955
R5650 VDD.n926 VDD.t7 27.6955
R5651 VDD.n926 VDD.t9 27.6955
R5652 VDD.n925 VDD.t32 27.6955
R5653 VDD.n925 VDD.t150 27.6955
R5654 VDD.n71 VDD.t50 27.6955
R5655 VDD.n71 VDD.t52 27.6955
R5656 VDD.n70 VDD.t15 27.6955
R5657 VDD.n70 VDD.t49 27.6955
R5658 VDD.n2643 VDD.n2642 26.8524
R5659 VDD.n2642 VDD.n2641 26.8524
R5660 VDD.n3382 VDD.n3379 26.8524
R5661 VDD.n3367 VDD.n3366 26.8524
R5662 VDD.n2283 VDD.n2258 26.8524
R5663 VDD.n2283 VDD.n2257 26.8524
R5664 VDD.n2283 VDD.n2282 26.8524
R5665 VDD.n2390 VDD.n2389 26.8524
R5666 VDD.n1934 VDD.n1933 26.8524
R5667 VDD.n1844 VDD.n1814 26.8524
R5668 VDD.n1857 VDD.n1814 26.8524
R5669 VDD.n1843 VDD.n1814 26.8524
R5670 VDD.n1429 VDD.n1404 26.8524
R5671 VDD.n1429 VDD.n1403 26.8524
R5672 VDD.n1429 VDD.n1428 26.8524
R5673 VDD.n1536 VDD.n1535 26.8524
R5674 VDD.n1080 VDD.n1079 26.8524
R5675 VDD.n990 VDD.n960 26.8524
R5676 VDD.n1003 VDD.n960 26.8524
R5677 VDD.n989 VDD.n960 26.8524
R5678 VDD.n574 VDD.n549 26.8524
R5679 VDD.n574 VDD.n548 26.8524
R5680 VDD.n574 VDD.n573 26.8524
R5681 VDD.n681 VDD.n680 26.8524
R5682 VDD.n225 VDD.n224 26.8524
R5683 VDD.n135 VDD.n105 26.8524
R5684 VDD.n148 VDD.n105 26.8524
R5685 VDD.n134 VDD.n105 26.8524
R5686 VDD.n2806 VDD.n2805 26.8521
R5687 VDD.n2389 VDD.n2388 26.8521
R5688 VDD.n2389 VDD.n2223 26.8521
R5689 VDD.n2389 VDD.n2220 26.8521
R5690 VDD.n2389 VDD.n2221 26.8521
R5691 VDD.n2389 VDD.n2222 26.8521
R5692 VDD.n1535 VDD.n1534 26.8521
R5693 VDD.n1535 VDD.n1369 26.8521
R5694 VDD.n1535 VDD.n1366 26.8521
R5695 VDD.n1535 VDD.n1367 26.8521
R5696 VDD.n1535 VDD.n1368 26.8521
R5697 VDD.n680 VDD.n679 26.8521
R5698 VDD.n680 VDD.n514 26.8521
R5699 VDD.n680 VDD.n511 26.8521
R5700 VDD.n680 VDD.n512 26.8521
R5701 VDD.n680 VDD.n513 26.8521
R5702 VDD.n3008 VDD.n2646 26.3534
R5703 VDD.n2272 VDD.n2249 26.3534
R5704 VDD.n1418 VDD.n1395 26.3534
R5705 VDD.n563 VDD.n540 26.3534
R5706 VDD.n4613 VDD.n4612 26.3453
R5707 VDD.n5153 VDD.n5152 26.3453
R5708 VDD.n5297 VDD.n5296 26.3453
R5709 VDD.n8661 VDD.n8660 26.3453
R5710 VDD.n8740 VDD.n8739 26.3453
R5711 VDD.n8940 VDD.n8939 26.3453
R5712 VDD.n3432 VDD.n3431 25.9875
R5713 VDD.n2709 VDD.n2708 25.7394
R5714 VDD.n2184 VDD.n2183 25.7394
R5715 VDD.n1330 VDD.n1329 25.7394
R5716 VDD.n475 VDD.n474 25.7394
R5717 VDD.n7618 VDD.n7615 25.6005
R5718 VDD.n7615 VDD.n7613 25.6005
R5719 VDD.n7613 VDD.n7611 25.6005
R5720 VDD.n7611 VDD.n7609 25.6005
R5721 VDD.n7609 VDD.n7607 25.6005
R5722 VDD.n7607 VDD.n7605 25.6005
R5723 VDD.n7605 VDD.n7604 25.6005
R5724 VDD.n7604 VDD.n7603 25.6005
R5725 VDD.n7603 VDD.n7602 25.6005
R5726 VDD.n3967 VDD.n3966 25.6005
R5727 VDD.n3968 VDD.n3967 25.6005
R5728 VDD.n3456 VDD.n3455 25.6005
R5729 VDD.n3457 VDD.n3456 25.6005
R5730 VDD.n3458 VDD.n3457 25.6005
R5731 VDD.n3459 VDD.n3458 25.6005
R5732 VDD.n3460 VDD.n3459 25.6005
R5733 VDD.n3461 VDD.n3460 25.6005
R5734 VDD.n3463 VDD.n3461 25.6005
R5735 VDD.n3465 VDD.n3463 25.6005
R5736 VDD.n3467 VDD.n3465 25.6005
R5737 VDD.n3046 VDD.n3043 25.6005
R5738 VDD.n2638 VDD.n2635 25.6005
R5739 VDD.n2640 VDD.n2638 25.6005
R5740 VDD.n2646 VDD.n2640 25.6005
R5741 VDD.n3271 VDD.n3268 25.6005
R5742 VDD.n3268 VDD.n3265 25.6005
R5743 VDD.n3265 VDD.n3261 25.6005
R5744 VDD.n3261 VDD.n3259 25.6005
R5745 VDD.n2860 VDD.n2856 25.6005
R5746 VDD.n2856 VDD.n2853 25.6005
R5747 VDD.n2853 VDD.n2850 25.6005
R5748 VDD.n2850 VDD.n2847 25.6005
R5749 VDD.n2847 VDD.n2844 25.6005
R5750 VDD.n2844 VDD.n2841 25.6005
R5751 VDD.n2841 VDD.n2838 25.6005
R5752 VDD.n2838 VDD.n2835 25.6005
R5753 VDD.n2835 VDD.n2832 25.6005
R5754 VDD.n2832 VDD.n2829 25.6005
R5755 VDD.n2829 VDD.n2826 25.6005
R5756 VDD.n2826 VDD.n2823 25.6005
R5757 VDD.n2823 VDD.n2820 25.6005
R5758 VDD.n3217 VDD.n3214 25.6005
R5759 VDD.n3220 VDD.n3217 25.6005
R5760 VDD.n3223 VDD.n3220 25.6005
R5761 VDD.n3226 VDD.n3223 25.6005
R5762 VDD.n3229 VDD.n3226 25.6005
R5763 VDD.n3232 VDD.n3229 25.6005
R5764 VDD.n3235 VDD.n3232 25.6005
R5765 VDD.n3238 VDD.n3235 25.6005
R5766 VDD.n3241 VDD.n3238 25.6005
R5767 VDD.n3244 VDD.n3241 25.6005
R5768 VDD.n3247 VDD.n3244 25.6005
R5769 VDD.n3250 VDD.n3247 25.6005
R5770 VDD.n3253 VDD.n3250 25.6005
R5771 VDD.n3257 VDD.n3253 25.6005
R5772 VDD.n2874 VDD.n2871 25.6005
R5773 VDD.n2871 VDD.n2868 25.6005
R5774 VDD.n2868 VDD.n2864 25.6005
R5775 VDD.n2864 VDD.n2862 25.6005
R5776 VDD.n3399 VDD.n3394 25.6005
R5777 VDD.n3394 VDD.n3391 25.6005
R5778 VDD.n3391 VDD.n3388 25.6005
R5779 VDD.n3315 VDD.n3311 25.6005
R5780 VDD.n2663 VDD.n2657 25.6005
R5781 VDD.n2657 VDD.n2654 25.6005
R5782 VDD.n2654 VDD.n2651 25.6005
R5783 VDD.n2651 VDD.n2648 25.6005
R5784 VDD.n2280 VDD.n2279 25.6005
R5785 VDD.n2279 VDD.n2278 25.6005
R5786 VDD.n2278 VDD.n2276 25.6005
R5787 VDD.n2276 VDD.n2273 25.6005
R5788 VDD.n2273 VDD.n2272 25.6005
R5789 VDD.n2503 VDD.n2502 25.6005
R5790 VDD.n2502 VDD.n2501 25.6005
R5791 VDD.n2501 VDD.n1953 25.6005
R5792 VDD.n2496 VDD.n1953 25.6005
R5793 VDD.n2438 VDD.n2437 25.6005
R5794 VDD.n2438 VDD.n1980 25.6005
R5795 VDD.n2444 VDD.n1980 25.6005
R5796 VDD.n2445 VDD.n2444 25.6005
R5797 VDD.n2446 VDD.n2445 25.6005
R5798 VDD.n2446 VDD.n1976 25.6005
R5799 VDD.n2452 VDD.n1976 25.6005
R5800 VDD.n2453 VDD.n2452 25.6005
R5801 VDD.n2454 VDD.n2453 25.6005
R5802 VDD.n2454 VDD.n1972 25.6005
R5803 VDD.n2460 VDD.n1972 25.6005
R5804 VDD.n2461 VDD.n2460 25.6005
R5805 VDD.n2462 VDD.n2461 25.6005
R5806 VDD.n2462 VDD.n1968 25.6005
R5807 VDD.n2468 VDD.n1968 25.6005
R5808 VDD.n2469 VDD.n2468 25.6005
R5809 VDD.n2470 VDD.n2469 25.6005
R5810 VDD.n2470 VDD.n1964 25.6005
R5811 VDD.n2476 VDD.n1964 25.6005
R5812 VDD.n2477 VDD.n2476 25.6005
R5813 VDD.n2478 VDD.n2477 25.6005
R5814 VDD.n2478 VDD.n1960 25.6005
R5815 VDD.n2484 VDD.n1960 25.6005
R5816 VDD.n2485 VDD.n2484 25.6005
R5817 VDD.n2486 VDD.n2485 25.6005
R5818 VDD.n2486 VDD.n1956 25.6005
R5819 VDD.n2494 VDD.n1956 25.6005
R5820 VDD.n2495 VDD.n2494 25.6005
R5821 VDD.n2430 VDD.n2428 25.6005
R5822 VDD.n2430 VDD.n2429 25.6005
R5823 VDD.n2429 VDD.n1984 25.6005
R5824 VDD.n2436 VDD.n1984 25.6005
R5825 VDD.n1894 VDD.n1878 25.6005
R5826 VDD.n1888 VDD.n1878 25.6005
R5827 VDD.n1888 VDD.n1887 25.6005
R5828 VDD.n1887 VDD.n1880 25.6005
R5829 VDD.n1881 VDD.n1880 25.6005
R5830 VDD.n2334 VDD.n2248 25.6005
R5831 VDD.n2340 VDD.n2334 25.6005
R5832 VDD.n2341 VDD.n2340 25.6005
R5833 VDD.n2341 VDD.n2332 25.6005
R5834 VDD.n2347 VDD.n2332 25.6005
R5835 VDD.n1426 VDD.n1425 25.6005
R5836 VDD.n1425 VDD.n1424 25.6005
R5837 VDD.n1424 VDD.n1422 25.6005
R5838 VDD.n1422 VDD.n1419 25.6005
R5839 VDD.n1419 VDD.n1418 25.6005
R5840 VDD.n1649 VDD.n1648 25.6005
R5841 VDD.n1648 VDD.n1647 25.6005
R5842 VDD.n1647 VDD.n1099 25.6005
R5843 VDD.n1642 VDD.n1099 25.6005
R5844 VDD.n1584 VDD.n1583 25.6005
R5845 VDD.n1584 VDD.n1126 25.6005
R5846 VDD.n1590 VDD.n1126 25.6005
R5847 VDD.n1591 VDD.n1590 25.6005
R5848 VDD.n1592 VDD.n1591 25.6005
R5849 VDD.n1592 VDD.n1122 25.6005
R5850 VDD.n1598 VDD.n1122 25.6005
R5851 VDD.n1599 VDD.n1598 25.6005
R5852 VDD.n1600 VDD.n1599 25.6005
R5853 VDD.n1600 VDD.n1118 25.6005
R5854 VDD.n1606 VDD.n1118 25.6005
R5855 VDD.n1607 VDD.n1606 25.6005
R5856 VDD.n1608 VDD.n1607 25.6005
R5857 VDD.n1608 VDD.n1114 25.6005
R5858 VDD.n1614 VDD.n1114 25.6005
R5859 VDD.n1615 VDD.n1614 25.6005
R5860 VDD.n1616 VDD.n1615 25.6005
R5861 VDD.n1616 VDD.n1110 25.6005
R5862 VDD.n1622 VDD.n1110 25.6005
R5863 VDD.n1623 VDD.n1622 25.6005
R5864 VDD.n1624 VDD.n1623 25.6005
R5865 VDD.n1624 VDD.n1106 25.6005
R5866 VDD.n1630 VDD.n1106 25.6005
R5867 VDD.n1631 VDD.n1630 25.6005
R5868 VDD.n1632 VDD.n1631 25.6005
R5869 VDD.n1632 VDD.n1102 25.6005
R5870 VDD.n1640 VDD.n1102 25.6005
R5871 VDD.n1641 VDD.n1640 25.6005
R5872 VDD.n1576 VDD.n1574 25.6005
R5873 VDD.n1576 VDD.n1575 25.6005
R5874 VDD.n1575 VDD.n1130 25.6005
R5875 VDD.n1582 VDD.n1130 25.6005
R5876 VDD.n1040 VDD.n1024 25.6005
R5877 VDD.n1034 VDD.n1024 25.6005
R5878 VDD.n1034 VDD.n1033 25.6005
R5879 VDD.n1033 VDD.n1026 25.6005
R5880 VDD.n1027 VDD.n1026 25.6005
R5881 VDD.n1480 VDD.n1394 25.6005
R5882 VDD.n1486 VDD.n1480 25.6005
R5883 VDD.n1487 VDD.n1486 25.6005
R5884 VDD.n1487 VDD.n1478 25.6005
R5885 VDD.n1493 VDD.n1478 25.6005
R5886 VDD.n571 VDD.n570 25.6005
R5887 VDD.n570 VDD.n569 25.6005
R5888 VDD.n569 VDD.n567 25.6005
R5889 VDD.n567 VDD.n564 25.6005
R5890 VDD.n564 VDD.n563 25.6005
R5891 VDD.n794 VDD.n793 25.6005
R5892 VDD.n793 VDD.n792 25.6005
R5893 VDD.n792 VDD.n244 25.6005
R5894 VDD.n787 VDD.n244 25.6005
R5895 VDD.n729 VDD.n728 25.6005
R5896 VDD.n729 VDD.n271 25.6005
R5897 VDD.n735 VDD.n271 25.6005
R5898 VDD.n736 VDD.n735 25.6005
R5899 VDD.n737 VDD.n736 25.6005
R5900 VDD.n737 VDD.n267 25.6005
R5901 VDD.n743 VDD.n267 25.6005
R5902 VDD.n744 VDD.n743 25.6005
R5903 VDD.n745 VDD.n744 25.6005
R5904 VDD.n745 VDD.n263 25.6005
R5905 VDD.n751 VDD.n263 25.6005
R5906 VDD.n752 VDD.n751 25.6005
R5907 VDD.n753 VDD.n752 25.6005
R5908 VDD.n753 VDD.n259 25.6005
R5909 VDD.n759 VDD.n259 25.6005
R5910 VDD.n760 VDD.n759 25.6005
R5911 VDD.n761 VDD.n760 25.6005
R5912 VDD.n761 VDD.n255 25.6005
R5913 VDD.n767 VDD.n255 25.6005
R5914 VDD.n768 VDD.n767 25.6005
R5915 VDD.n769 VDD.n768 25.6005
R5916 VDD.n769 VDD.n251 25.6005
R5917 VDD.n775 VDD.n251 25.6005
R5918 VDD.n776 VDD.n775 25.6005
R5919 VDD.n777 VDD.n776 25.6005
R5920 VDD.n777 VDD.n247 25.6005
R5921 VDD.n785 VDD.n247 25.6005
R5922 VDD.n786 VDD.n785 25.6005
R5923 VDD.n721 VDD.n719 25.6005
R5924 VDD.n721 VDD.n720 25.6005
R5925 VDD.n720 VDD.n275 25.6005
R5926 VDD.n727 VDD.n275 25.6005
R5927 VDD.n185 VDD.n169 25.6005
R5928 VDD.n179 VDD.n169 25.6005
R5929 VDD.n179 VDD.n178 25.6005
R5930 VDD.n178 VDD.n171 25.6005
R5931 VDD.n172 VDD.n171 25.6005
R5932 VDD.n625 VDD.n539 25.6005
R5933 VDD.n631 VDD.n625 25.6005
R5934 VDD.n632 VDD.n631 25.6005
R5935 VDD.n632 VDD.n623 25.6005
R5936 VDD.n638 VDD.n623 25.6005
R5937 VDD.n7574 VDD.n7573 25.3507
R5938 VDD.n7130 VDD.n7129 25.3507
R5939 VDD.n3207 VDD.n3206 25.3507
R5940 VDD.n2770 VDD.n2769 25.3507
R5941 VDD.n2971 VDD.n2970 25.3507
R5942 VDD.n1903 VDD.n1902 25.3507
R5943 VDD.n2399 VDD.n2398 25.3507
R5944 VDD.n2298 VDD.n2013 25.3507
R5945 VDD.n1049 VDD.n1048 25.3507
R5946 VDD.n1545 VDD.n1544 25.3507
R5947 VDD.n1444 VDD.n1159 25.3507
R5948 VDD.n194 VDD.n193 25.3507
R5949 VDD.n690 VDD.n689 25.3507
R5950 VDD.n589 VDD.n304 25.3507
R5951 VDD.n8567 VDD.n8566 25.3505
R5952 VDD.n8549 VDD.n8548 25.3505
R5953 VDD.n7499 VDD.n7498 25.3505
R5954 VDD.n7118 VDD.n7117 25.3505
R5955 VDD.n2716 VDD.n2715 25.3505
R5956 VDD.n2725 VDD.n2724 25.3505
R5957 VDD.n2803 VDD.n2802 25.3505
R5958 VDD.n2912 VDD.n2911 25.3505
R5959 VDD.n3164 VDD.n3163 25.3505
R5960 VDD.n3170 VDD.n3169 25.3505
R5961 VDD.n3371 VDD.n3370 25.3505
R5962 VDD.n2173 VDD.n2040 25.3505
R5963 VDD.n2174 VDD.n2037 25.3505
R5964 VDD.n2377 VDD.n2016 25.3505
R5965 VDD.n2402 VDD.n2401 25.3505
R5966 VDD.n2534 VDD.n2533 25.3505
R5967 VDD.n1834 VDD.n1809 25.3505
R5968 VDD.n1873 VDD.n1872 25.3505
R5969 VDD.n1319 VDD.n1186 25.3505
R5970 VDD.n1320 VDD.n1183 25.3505
R5971 VDD.n1523 VDD.n1162 25.3505
R5972 VDD.n1548 VDD.n1547 25.3505
R5973 VDD.n1680 VDD.n1679 25.3505
R5974 VDD.n980 VDD.n955 25.3505
R5975 VDD.n1019 VDD.n1018 25.3505
R5976 VDD.n464 VDD.n331 25.3505
R5977 VDD.n465 VDD.n328 25.3505
R5978 VDD.n668 VDD.n307 25.3505
R5979 VDD.n693 VDD.n692 25.3505
R5980 VDD.n825 VDD.n824 25.3505
R5981 VDD.n125 VDD.n100 25.3505
R5982 VDD.n164 VDD.n163 25.3505
R5983 VDD.n3549 VDD.t34 24.8124
R5984 VDD.n3543 VDD.n3542 23.9713
R5985 VDD.n43 VDD.t30 23.5572
R5986 VDD.n912 VDD.t147 23.5572
R5987 VDD.n1752 VDD.t159 23.5572
R5988 VDD.n2621 VDD.t109 23.5572
R5989 VDD.n3431 VDD.n3430 23.4711
R5990 VDD.n2256 VDD.n2245 23.0774
R5991 VDD.n2352 VDD.n2283 23.0774
R5992 VDD.n1925 VDD.n1803 23.0774
R5993 VDD.n1402 VDD.n1391 23.0774
R5994 VDD.n1498 VDD.n1429 23.0774
R5995 VDD.n1071 VDD.n949 23.0774
R5996 VDD.n547 VDD.n536 23.0774
R5997 VDD.n643 VDD.n574 23.0774
R5998 VDD.n216 VDD.n94 23.0774
R5999 VDD.n4622 VDD.n4621 23.0522
R6000 VDD.n5198 VDD.n5197 23.0522
R6001 VDD.n5258 VDD.n5257 23.0522
R6002 VDD.n8643 VDD.n8642 23.0522
R6003 VDD.n9006 VDD.n9005 23.0522
R6004 VDD.n8922 VDD.n8921 23.0522
R6005 VDD.n8834 VDD.n8833 22.7097
R6006 VDD.n8780 VDD.t112 22.2891
R6007 VDD.n3377 VDD.t69 21.7954
R6008 VDD.n2237 VDD.t17 21.7954
R6009 VDD.n1931 VDD.t155 21.7954
R6010 VDD.t155 VDD.n1822 21.7954
R6011 VDD.n1383 VDD.t6 21.7954
R6012 VDD.n1077 VDD.t151 21.7954
R6013 VDD.t151 VDD.n968 21.7954
R6014 VDD.n528 VDD.t16 21.7954
R6015 VDD.n222 VDD.t47 21.7954
R6016 VDD.t47 VDD.n113 21.7954
R6017 VDD.n8764 VDD.n8763 21.468
R6018 VDD.n39 VDD.n34 21.1346
R6019 VDD.n901 VDD.n897 21.1346
R6020 VDD.n1748 VDD.n1743 21.1346
R6021 VDD.n8138 VDD.n8137 20.7186
R6022 VDD.n7631 VDD.n7630 20.7183
R6023 VDD.n7631 VDD.n7627 20.7183
R6024 VDD.n7631 VDD.n7624 20.7183
R6025 VDD.n7631 VDD.n7621 20.7183
R6026 VDD.n7631 VDD.n7620 20.7183
R6027 VDD.n3274 VDD.n3271 20.6044
R6028 VDD.n2503 VDD.n1949 20.6044
R6029 VDD.n1649 VDD.n1095 20.6044
R6030 VDD.n794 VDD.n240 20.6044
R6031 VDD.n2359 VDD.n2245 20.5133
R6032 VDD.n2286 VDD.n2283 20.5133
R6033 VDD.n2541 VDD.n1803 20.5133
R6034 VDD.n1505 VDD.n1391 20.5133
R6035 VDD.n1432 VDD.n1429 20.5133
R6036 VDD.n1687 VDD.n949 20.5133
R6037 VDD.n650 VDD.n536 20.5133
R6038 VDD.n577 VDD.n574 20.5133
R6039 VDD.n832 VDD.n94 20.5133
R6040 VDD.n4673 VDD.n4672 19.7591
R6041 VDD.n5213 VDD.n5212 19.7591
R6042 VDD.n5286 VDD.n5285 19.7591
R6043 VDD.n2877 VDD.n2874 18.7439
R6044 VDD.n2428 VDD.n2427 18.7439
R6045 VDD.n1574 VDD.n1573 18.7439
R6046 VDD.n719 VDD.n718 18.7439
R6047 VDD.n43 VDD.t116 17.8272
R6048 VDD.n912 VDD.t22 17.8272
R6049 VDD.n1752 VDD.t75 17.8272
R6050 VDD.n2621 VDD.t156 17.8272
R6051 VDD.n3803 VDD.n3801 17.8254
R6052 VDD.n49 VDD.n35 17.2489
R6053 VDD.n910 VDD.n909 17.2489
R6054 VDD.n1758 VDD.n1744 17.2489
R6055 VDD.n2619 VDD.n2618 17.2489
R6056 VDD.n3623 VDD.n3547 17.2426
R6057 VDD.n4652 VDD.n4651 16.466
R6058 VDD.n5184 VDD.n5183 16.466
R6059 VDD.n4310 VDD.n4309 16.466
R6060 VDD.n5339 VDD.n5338 16.466
R6061 VDD.n8606 VDD.n8605 16.466
R6062 VDD.n8968 VDD.n8967 16.466
R6063 VDD.n8909 VDD.n8908 16.466
R6064 VDD.n2919 VDD.n2915 15.6165
R6065 VDD.n3326 VDD.n3325 15.6165
R6066 VDD.n2350 VDD.n2348 15.6165
R6067 VDD.n2549 VDD.n1792 15.6165
R6068 VDD.n1496 VDD.n1494 15.6165
R6069 VDD.n1695 VDD.n938 15.6165
R6070 VDD.n641 VDD.n639 15.6165
R6071 VDD.n840 VDD.n83 15.6165
R6072 VDD.n3803 VDD.n3802 15.0799
R6073 VDD.n2983 VDD.t117 14.7441
R6074 VDD.n2998 VDD.t119 14.7441
R6075 VDD.n3009 VDD.t5 14.7441
R6076 VDD.n3032 VDD.t4 14.7441
R6077 VDD.n3400 VDD.t121 14.7441
R6078 VDD.t17 VDD.n2231 14.7441
R6079 VDD.n2359 VDD.t19 14.7441
R6080 VDD.n2286 VDD.t154 14.7441
R6081 VDD.t35 VDD.n1788 14.7441
R6082 VDD.n1794 VDD.t35 14.7441
R6083 VDD.n2541 VDD.t104 14.7441
R6084 VDD.t6 VDD.n1377 14.7441
R6085 VDD.n1505 VDD.t8 14.7441
R6086 VDD.n1432 VDD.t148 14.7441
R6087 VDD.t31 VDD.n934 14.7441
R6088 VDD.n940 VDD.t31 14.7441
R6089 VDD.n1687 VDD.t149 14.7441
R6090 VDD.t16 VDD.n522 14.7441
R6091 VDD.n650 VDD.t51 14.7441
R6092 VDD.n577 VDD.t67 14.7441
R6093 VDD.t14 VDD.n79 14.7441
R6094 VDD.n85 VDD.t14 14.7441
R6095 VDD.n832 VDD.t48 14.7441
R6096 VDD.n8137 VDD.n8136 14.2505
R6097 VDD.n2921 VDD.n2919 14.2085
R6098 VDD.n3328 VDD.n3326 14.2085
R6099 VDD.n2348 VDD.n2331 14.2085
R6100 VDD.n1928 VDD.n1792 14.2085
R6101 VDD.n1494 VDD.n1477 14.2085
R6102 VDD.n1074 VDD.n938 14.2085
R6103 VDD.n639 VDD.n622 14.2085
R6104 VDD.n219 VDD.n83 14.2085
R6105 VDD.n2285 VDD.n1787 14.1031
R6106 VDD.n2553 VDD.n1788 14.1031
R6107 VDD.n1795 VDD.n1794 14.1031
R6108 VDD.n2547 VDD.n1796 14.1031
R6109 VDD.n1431 VDD.n933 14.1031
R6110 VDD.n1699 VDD.n934 14.1031
R6111 VDD.n941 VDD.n940 14.1031
R6112 VDD.n1693 VDD.n942 14.1031
R6113 VDD.n576 VDD.n78 14.1031
R6114 VDD.n844 VDD.n79 14.1031
R6115 VDD.n86 VDD.n85 14.1031
R6116 VDD.n838 VDD.n87 14.1031
R6117 VDD.t68 VDD.n6659 13.8783
R6118 VDD.n8840 VDD.n8839 13.8783
R6119 VDD.n1931 VDD.n1924 13.462
R6120 VDD.n1077 VDD.n1070 13.462
R6121 VDD.n222 VDD.n215 13.462
R6122 VDD.t43 VDD.n6666 13.0372
R6123 VDD.t53 VDD.n9 12.789
R6124 VDD.n879 VDD.t23 12.789
R6125 VDD.t61 VDD.n1718 12.789
R6126 VDD.n2580 VDD.t135 12.789
R6127 VDD.n5140 VDD.n5137 12.6901
R6128 VDD.n7632 VDD.n7631 12.6672
R6129 VDD.n3433 VDD.n3432 12.1342
R6130 VDD.n5834 VDD.n5833 12.064
R6131 VDD.n2928 VDD.n2927 12.0325
R6132 VDD.n3335 VDD.n3334 12.0325
R6133 VDD.n2326 VDD.n2002 12.0325
R6134 VDD.n1939 VDD.n1938 12.0325
R6135 VDD.n1472 VDD.n1148 12.0325
R6136 VDD.n1085 VDD.n1084 12.0325
R6137 VDD.n617 VDD.n293 12.0325
R6138 VDD.n230 VDD.n229 12.0325
R6139 VDD.n3542 VDD.t10 11.8979
R6140 VDD.n3906 VDD.n3905 11.6711
R6141 VDD.n3623 VDD.n3554 11.3551
R6142 VDD.n6772 VDD.t140 11.3551
R6143 VDD.n3427 VDD.n3426 11.1178
R6144 VDD.n5238 VDD.n3762 10.8935
R6145 VDD.n3806 VDD.n3805 10.8935
R6146 VDD.n3051 VDD.n3050 10.4112
R6147 VDD.n3053 VDD.n3051 10.4112
R6148 VDD.n2267 VDD.n2242 10.4112
R6149 VDD.n2267 VDD.n2266 10.4112
R6150 VDD.n1413 VDD.n1388 10.4112
R6151 VDD.n1413 VDD.n1412 10.4112
R6152 VDD.n558 VDD.n533 10.4112
R6153 VDD.n558 VDD.n557 10.4112
R6154 VDD.n4641 VDD.n4640 9.87981
R6155 VDD.n5173 VDD.n5172 9.87981
R6156 VDD.n4294 VDD.n4293 9.87981
R6157 VDD.n5323 VDD.n5322 9.87981
R6158 VDD.n8627 VDD.n8626 9.87981
R6159 VDD.n8989 VDD.n8988 9.87981
R6160 VDD.n8899 VDD.n8898 9.87981
R6161 VDD.n6742 VDD.t141 9.67292
R6162 VDD.n8835 VDD.n8834 9.67292
R6163 VDD.n4634 VDD.n4633 9.3005
R6164 VDD.n4645 VDD.n4644 9.3005
R6165 VDD.n4658 VDD.n4657 9.3005
R6166 VDD.n4632 VDD.n4631 9.3005
R6167 VDD.n4631 VDD.n4630 9.3005
R6168 VDD.n4636 VDD.n4635 9.3005
R6169 VDD.n4643 VDD.n4642 9.3005
R6170 VDD.n4642 VDD.n4641 9.3005
R6171 VDD.n4647 VDD.n4646 9.3005
R6172 VDD.n4654 VDD.n4653 9.3005
R6173 VDD.n4653 VDD.n4652 9.3005
R6174 VDD.n4656 VDD.n4655 9.3005
R6175 VDD.n4615 VDD.n4614 9.3005
R6176 VDD.n4623 VDD.n4622 9.3005
R6177 VDD.n4713 VDD.n4712 9.3005
R6178 VDD.n4715 VDD.n4714 9.3005
R6179 VDD.n4711 VDD.n4710 9.3005
R6180 VDD.n4710 VDD.n4709 9.3005
R6181 VDD.n4699 VDD.n4698 9.3005
R6182 VDD.n4697 VDD.n4696 9.3005
R6183 VDD.n4695 VDD.n4694 9.3005
R6184 VDD.n4694 VDD.n4693 9.3005
R6185 VDD.n4723 VDD.n4722 9.3005
R6186 VDD.n4730 VDD.n4729 9.3005
R6187 VDD.n4737 VDD.n4736 9.3005
R6188 VDD.n4744 VDD.n4743 9.3005
R6189 VDD.n4751 VDD.n4750 9.3005
R6190 VDD.n4758 VDD.n4757 9.3005
R6191 VDD.n4764 VDD.n4763 9.3005
R6192 VDD.n4771 VDD.n4770 9.3005
R6193 VDD.n4778 VDD.n4777 9.3005
R6194 VDD.n4780 VDD.n4779 9.3005
R6195 VDD.n4776 VDD.n4775 9.3005
R6196 VDD.n4773 VDD.n4772 9.3005
R6197 VDD.n4769 VDD.n4768 9.3005
R6198 VDD.n4766 VDD.n4765 9.3005
R6199 VDD.n4762 VDD.n4761 9.3005
R6200 VDD.n4760 VDD.n4759 9.3005
R6201 VDD.n4756 VDD.n4755 9.3005
R6202 VDD.n4754 VDD.n4753 9.3005
R6203 VDD.n4749 VDD.n4748 9.3005
R6204 VDD.n4747 VDD.n4746 9.3005
R6205 VDD.n4742 VDD.n4741 9.3005
R6206 VDD.n4740 VDD.n4739 9.3005
R6207 VDD.n4735 VDD.n4734 9.3005
R6208 VDD.n4733 VDD.n4732 9.3005
R6209 VDD.n4728 VDD.n4727 9.3005
R6210 VDD.n4726 VDD.n4725 9.3005
R6211 VDD.n4721 VDD.n4720 9.3005
R6212 VDD.n5054 VDD.n5053 9.3005
R6213 VDD.n5056 VDD.n5055 9.3005
R6214 VDD.n5052 VDD.n5051 9.3005
R6215 VDD.n5051 VDD.n5050 9.3005
R6216 VDD.n5040 VDD.n5039 9.3005
R6217 VDD.n5038 VDD.n5037 9.3005
R6218 VDD.n5036 VDD.n5035 9.3005
R6219 VDD.n5035 VDD.n5034 9.3005
R6220 VDD.n5064 VDD.n5063 9.3005
R6221 VDD.n5071 VDD.n5070 9.3005
R6222 VDD.n5078 VDD.n5077 9.3005
R6223 VDD.n5085 VDD.n5084 9.3005
R6224 VDD.n5092 VDD.n5091 9.3005
R6225 VDD.n5099 VDD.n5098 9.3005
R6226 VDD.n5105 VDD.n5104 9.3005
R6227 VDD.n5112 VDD.n5111 9.3005
R6228 VDD.n5119 VDD.n5118 9.3005
R6229 VDD.n5121 VDD.n5120 9.3005
R6230 VDD.n5117 VDD.n5116 9.3005
R6231 VDD.n5114 VDD.n5113 9.3005
R6232 VDD.n5110 VDD.n5109 9.3005
R6233 VDD.n5107 VDD.n5106 9.3005
R6234 VDD.n5103 VDD.n5102 9.3005
R6235 VDD.n5101 VDD.n5100 9.3005
R6236 VDD.n5097 VDD.n5096 9.3005
R6237 VDD.n5095 VDD.n5094 9.3005
R6238 VDD.n5090 VDD.n5089 9.3005
R6239 VDD.n5088 VDD.n5087 9.3005
R6240 VDD.n5083 VDD.n5082 9.3005
R6241 VDD.n5081 VDD.n5080 9.3005
R6242 VDD.n5076 VDD.n5075 9.3005
R6243 VDD.n5074 VDD.n5073 9.3005
R6244 VDD.n5069 VDD.n5068 9.3005
R6245 VDD.n5067 VDD.n5066 9.3005
R6246 VDD.n5062 VDD.n5061 9.3005
R6247 VDD.n5188 VDD.n5187 9.3005
R6248 VDD.n5177 VDD.n5176 9.3005
R6249 VDD.n5166 VDD.n5165 9.3005
R6250 VDD.n5164 VDD.n5163 9.3005
R6251 VDD.n5163 VDD.n5162 9.3005
R6252 VDD.n5168 VDD.n5167 9.3005
R6253 VDD.n5175 VDD.n5174 9.3005
R6254 VDD.n5174 VDD.n5173 9.3005
R6255 VDD.n5179 VDD.n5178 9.3005
R6256 VDD.n5186 VDD.n5185 9.3005
R6257 VDD.n5185 VDD.n5184 9.3005
R6258 VDD.n5190 VDD.n5189 9.3005
R6259 VDD.n5155 VDD.n5154 9.3005
R6260 VDD.n5199 VDD.n5198 9.3005
R6261 VDD.n4470 VDD.n4469 9.3005
R6262 VDD.n4463 VDD.n4462 9.3005
R6263 VDD.n4456 VDD.n4455 9.3005
R6264 VDD.n4454 VDD.n4453 9.3005
R6265 VDD.n4459 VDD.n4458 9.3005
R6266 VDD.n4461 VDD.n4460 9.3005
R6267 VDD.n4466 VDD.n4465 9.3005
R6268 VDD.n4468 VDD.n4467 9.3005
R6269 VDD.n4540 VDD.n4539 9.3005
R6270 VDD.n4538 VDD.n4537 9.3005
R6271 VDD.n4526 VDD.n4525 9.3005
R6272 VDD.n4536 VDD.n4535 9.3005
R6273 VDD.n4529 VDD.n4528 9.3005
R6274 VDD.n4524 VDD.n4523 9.3005
R6275 VDD.n4531 VDD.n4530 9.3005
R6276 VDD.n4533 VDD.n4532 9.3005
R6277 VDD.n4446 VDD.n4445 9.3005
R6278 VDD.n4427 VDD.n4426 9.3005
R6279 VDD.n4448 VDD.n4447 9.3005
R6280 VDD.n4444 VDD.n4443 9.3005
R6281 VDD.n4443 VDD.n4442 9.3005
R6282 VDD.n4434 VDD.n4433 9.3005
R6283 VDD.n4433 VDD.n4432 9.3005
R6284 VDD.n4425 VDD.n4424 9.3005
R6285 VDD.n4516 VDD.n4515 9.3005
R6286 VDD.n4518 VDD.n4517 9.3005
R6287 VDD.n4514 VDD.n4513 9.3005
R6288 VDD.n4513 VDD.n4512 9.3005
R6289 VDD.n4420 VDD.n4419 9.3005
R6290 VDD.n4353 VDD.n4352 9.3005
R6291 VDD.n4337 VDD.n4336 9.3005
R6292 VDD.n4335 VDD.n4334 9.3005
R6293 VDD.n4333 VDD.n4332 9.3005
R6294 VDD.n4332 VDD.n4331 9.3005
R6295 VDD.n4351 VDD.n4350 9.3005
R6296 VDD.n4349 VDD.n4348 9.3005
R6297 VDD.n4348 VDD.n4347 9.3005
R6298 VDD.n4418 VDD.n4417 9.3005
R6299 VDD.n4416 VDD.n4415 9.3005
R6300 VDD.n4415 VDD.n4414 9.3005
R6301 VDD.n4362 VDD.n4361 9.3005
R6302 VDD.n4369 VDD.n4368 9.3005
R6303 VDD.n4376 VDD.n4375 9.3005
R6304 VDD.n4360 VDD.n4359 9.3005
R6305 VDD.n4365 VDD.n4364 9.3005
R6306 VDD.n4367 VDD.n4366 9.3005
R6307 VDD.n4372 VDD.n4371 9.3005
R6308 VDD.n4374 VDD.n4373 9.3005
R6309 VDD.n4287 VDD.n4286 9.3005
R6310 VDD.n4289 VDD.n4288 9.3005
R6311 VDD.n4285 VDD.n4284 9.3005
R6312 VDD.n4284 VDD.n4283 9.3005
R6313 VDD.n4311 VDD.n4310 9.3005
R6314 VDD.n4295 VDD.n4294 9.3005
R6315 VDD.n3655 VDD.n3654 9.3005
R6316 VDD.n3653 VDD.n3652 9.3005
R6317 VDD.n3652 VDD.n3651 9.3005
R6318 VDD.n3657 VDD.n3656 9.3005
R6319 VDD.n3679 VDD.n3678 9.3005
R6320 VDD.n3677 VDD.n3676 9.3005
R6321 VDD.n3665 VDD.n3664 9.3005
R6322 VDD.n3675 VDD.n3674 9.3005
R6323 VDD.n3668 VDD.n3667 9.3005
R6324 VDD.n3663 VDD.n3662 9.3005
R6325 VDD.n3670 VDD.n3669 9.3005
R6326 VDD.n3672 VDD.n3671 9.3005
R6327 VDD.n5316 VDD.n5315 9.3005
R6328 VDD.n5314 VDD.n5313 9.3005
R6329 VDD.n5313 VDD.n5312 9.3005
R6330 VDD.n5318 VDD.n5317 9.3005
R6331 VDD.n5272 VDD.n5271 9.3005
R6332 VDD.n5270 VDD.n5269 9.3005
R6333 VDD.n5269 VDD.n5268 9.3005
R6334 VDD.n5274 VDD.n5273 9.3005
R6335 VDD.n5282 VDD.n5281 9.3005
R6336 VDD.n5293 VDD.n5292 9.3005
R6337 VDD.n5304 VDD.n5303 9.3005
R6338 VDD.n5302 VDD.n5301 9.3005
R6339 VDD.n5300 VDD.n5299 9.3005
R6340 VDD.n5299 VDD.n5298 9.3005
R6341 VDD.n5291 VDD.n5290 9.3005
R6342 VDD.n5289 VDD.n5288 9.3005
R6343 VDD.n5288 VDD.n5287 9.3005
R6344 VDD.n5280 VDD.n5279 9.3005
R6345 VDD.n5259 VDD.n5258 9.3005
R6346 VDD.n5324 VDD.n5323 9.3005
R6347 VDD.n5340 VDD.n5339 9.3005
R6348 VDD.n8620 VDD.n8619 9.3005
R6349 VDD.n8618 VDD.n8617 9.3005
R6350 VDD.n8617 VDD.n8616 9.3005
R6351 VDD.n8622 VDD.n8621 9.3005
R6352 VDD.n8629 VDD.n8628 9.3005
R6353 VDD.n8628 VDD.n8627 9.3005
R6354 VDD.n8631 VDD.n8630 9.3005
R6355 VDD.n8644 VDD.n8643 9.3005
R6356 VDD.n8663 VDD.n8662 9.3005
R6357 VDD.n8633 VDD.n8632 9.3005
R6358 VDD.n8607 VDD.n8606 9.3005
R6359 VDD.n8982 VDD.n8981 9.3005
R6360 VDD.n8980 VDD.n8979 9.3005
R6361 VDD.n8979 VDD.n8978 9.3005
R6362 VDD.n8984 VDD.n8983 9.3005
R6363 VDD.n8991 VDD.n8990 9.3005
R6364 VDD.n8990 VDD.n8989 9.3005
R6365 VDD.n8993 VDD.n8992 9.3005
R6366 VDD.n9007 VDD.n9006 9.3005
R6367 VDD.n8742 VDD.n8741 9.3005
R6368 VDD.n8995 VDD.n8994 9.3005
R6369 VDD.n8969 VDD.n8968 9.3005
R6370 VDD.n8903 VDD.n8902 9.3005
R6371 VDD.n8892 VDD.n8891 9.3005
R6372 VDD.n8901 VDD.n8900 9.3005
R6373 VDD.n8900 VDD.n8899 9.3005
R6374 VDD.n8890 VDD.n8889 9.3005
R6375 VDD.n8889 VDD.n8888 9.3005
R6376 VDD.n8894 VDD.n8893 9.3005
R6377 VDD.n8905 VDD.n8904 9.3005
R6378 VDD.n8942 VDD.n8941 9.3005
R6379 VDD.n8923 VDD.n8922 9.3005
R6380 VDD.n8910 VDD.n8909 9.3005
R6381 VDD.n3910 VDD.n3909 9.3005
R6382 VDD.n3913 VDD.n3912 9.3005
R6383 VDD.n3901 VDD.n3900 9.3005
R6384 VDD.n2772 VDD.n2671 8.9605
R6385 VDD.n3166 VDD.n3063 8.9605
R6386 VDD.n2396 VDD.n2214 8.9605
R6387 VDD.n2538 VDD.n2537 8.9605
R6388 VDD.n1542 VDD.n1360 8.9605
R6389 VDD.n1684 VDD.n1683 8.9605
R6390 VDD.n687 VDD.n505 8.9605
R6391 VDD.n829 VDD.n828 8.9605
R6392 VDD.n38 VDD.n37 8.85536
R6393 VDD.n55 VDD.n54 8.85536
R6394 VDD.n53 VDD.n36 8.85536
R6395 VDD.n42 VDD.n41 8.85536
R6396 VDD.n19 VDD.n18 8.85536
R6397 VDD.n11 VDD.n10 8.85536
R6398 VDD.n10 VDD.n9 8.85536
R6399 VDD.n31 VDD.n30 8.85536
R6400 VDD.n32 VDD.n31 8.85536
R6401 VDD.n8 VDD.n7 8.85536
R6402 VDD.n33 VDD.n8 8.85536
R6403 VDD.n61 VDD.n60 8.85536
R6404 VDD.n60 VDD.n59 8.85536
R6405 VDD.n900 VDD.n899 8.85536
R6406 VDD.n906 VDD.n905 8.85536
R6407 VDD.n904 VDD.n898 8.85536
R6408 VDD.n860 VDD.n859 8.85536
R6409 VDD.n878 VDD.n877 8.85536
R6410 VDD.n869 VDD.n868 8.85536
R6411 VDD.n879 VDD.n869 8.85536
R6412 VDD.n882 VDD.n881 8.85536
R6413 VDD.n881 VDD.n880 8.85536
R6414 VDD.n863 VDD.n862 8.85536
R6415 VDD.n862 VDD.n861 8.85536
R6416 VDD.n894 VDD.n893 8.85536
R6417 VDD.n895 VDD.n894 8.85536
R6418 VDD.n1747 VDD.n1746 8.85536
R6419 VDD.n1764 VDD.n1763 8.85536
R6420 VDD.n1762 VDD.n1745 8.85536
R6421 VDD.n1751 VDD.n1750 8.85536
R6422 VDD.n1728 VDD.n1727 8.85536
R6423 VDD.n1720 VDD.n1719 8.85536
R6424 VDD.n1719 VDD.n1718 8.85536
R6425 VDD.n1740 VDD.n1739 8.85536
R6426 VDD.n1741 VDD.n1740 8.85536
R6427 VDD.n1717 VDD.n1716 8.85536
R6428 VDD.n1742 VDD.n1717 8.85536
R6429 VDD.n1770 VDD.n1769 8.85536
R6430 VDD.n1769 VDD.n1768 8.85536
R6431 VDD.n2603 VDD.n2602 8.85536
R6432 VDD.n2606 VDD.n2605 8.85536
R6433 VDD.n2609 VDD.n2608 8.85536
R6434 VDD.n2612 VDD.n2611 8.85536
R6435 VDD.n2575 VDD.n2574 8.85536
R6436 VDD.n2582 VDD.n2581 8.85536
R6437 VDD.n2581 VDD.n2580 8.85536
R6438 VDD.n2587 VDD.n2586 8.85536
R6439 VDD.n2586 VDD.n2585 8.85536
R6440 VDD.n2595 VDD.n2594 8.85536
R6441 VDD.n2594 VDD.n2593 8.85536
R6442 VDD.n2598 VDD.n2597 8.85536
R6443 VDD.n2597 VDD.n2596 8.85536
R6444 VDD.n4436 VDD.n4435 8.76429
R6445 VDD.n4341 VDD.n4340 8.76429
R6446 VDD.n2927 VDD.n2925 8.7045
R6447 VDD.n2925 VDD.n2923 8.7045
R6448 VDD.n2923 VDD.n2921 8.7045
R6449 VDD.n3319 VDD.n3317 8.7045
R6450 VDD.n3321 VDD.n3319 8.7045
R6451 VDD.n3323 VDD.n3321 8.7045
R6452 VDD.n3325 VDD.n3323 8.7045
R6453 VDD.n3330 VDD.n3328 8.7045
R6454 VDD.n3332 VDD.n3330 8.7045
R6455 VDD.n3334 VDD.n3332 8.7045
R6456 VDD.n2327 VDD.n2326 8.7045
R6457 VDD.n2328 VDD.n2327 8.7045
R6458 VDD.n2331 VDD.n2328 8.7045
R6459 VDD.n2350 VDD.n2349 8.7045
R6460 VDD.n2349 VDD.n1791 8.7045
R6461 VDD.n2551 VDD.n1791 8.7045
R6462 VDD.n2551 VDD.n2550 8.7045
R6463 VDD.n2550 VDD.n2549 8.7045
R6464 VDD.n1929 VDD.n1928 8.7045
R6465 VDD.n1929 VDD.n1819 8.7045
R6466 VDD.n1938 VDD.n1819 8.7045
R6467 VDD.n1473 VDD.n1472 8.7045
R6468 VDD.n1474 VDD.n1473 8.7045
R6469 VDD.n1477 VDD.n1474 8.7045
R6470 VDD.n1496 VDD.n1495 8.7045
R6471 VDD.n1495 VDD.n937 8.7045
R6472 VDD.n1697 VDD.n937 8.7045
R6473 VDD.n1697 VDD.n1696 8.7045
R6474 VDD.n1696 VDD.n1695 8.7045
R6475 VDD.n1075 VDD.n1074 8.7045
R6476 VDD.n1075 VDD.n965 8.7045
R6477 VDD.n1084 VDD.n965 8.7045
R6478 VDD.n618 VDD.n617 8.7045
R6479 VDD.n619 VDD.n618 8.7045
R6480 VDD.n622 VDD.n619 8.7045
R6481 VDD.n641 VDD.n640 8.7045
R6482 VDD.n640 VDD.n82 8.7045
R6483 VDD.n842 VDD.n82 8.7045
R6484 VDD.n842 VDD.n841 8.7045
R6485 VDD.n841 VDD.n840 8.7045
R6486 VDD.n220 VDD.n219 8.7045
R6487 VDD.n220 VDD.n110 8.7045
R6488 VDD.n229 VDD.n110 8.7045
R6489 VDD.n4199 VDD.n4117 8.65557
R6490 VDD.n8564 VDD.n8559 8.46493
R6491 VDD.n8869 VDD.n8868 8.45089
R6492 VDD.n3946 VDD.n3945 8.45089
R6493 VDD.n5243 VDD.n5242 8.45089
R6494 VDD.n3758 VDD.n3757 8.45089
R6495 VDD.n8817 VDD.n8816 8.45089
R6496 VDD.n8813 VDD.n8812 8.45089
R6497 VDD.n8807 VDD.n8806 8.45089
R6498 VDD.n3951 VDD.n3950 8.45089
R6499 VDD.n4073 VDD.n3953 8.45089
R6500 VDD.n3755 VDD.n3754 8.45089
R6501 VDD.n4270 VDD.n4269 8.45089
R6502 VDD.n8787 VDD.n8786 8.40959
R6503 VDD.n56 VDD.n36 8.39408
R6504 VDD.n56 VDD.n55 8.39408
R6505 VDD.n41 VDD.n35 8.39408
R6506 VDD.n907 VDD.n898 8.39408
R6507 VDD.n907 VDD.n906 8.39408
R6508 VDD.n909 VDD.n860 8.39408
R6509 VDD.n1765 VDD.n1745 8.39408
R6510 VDD.n1765 VDD.n1764 8.39408
R6511 VDD.n1750 VDD.n1744 8.39408
R6512 VDD.n37 VDD.n34 8.39405
R6513 VDD.n899 VDD.n897 8.39405
R6514 VDD.n1746 VDD.n1743 8.39405
R6515 VDD.n3971 VDD.n3970 8.06816
R6516 VDD.n4021 VDD.n4020 8.06816
R6517 VDD.n4025 VDD.n4024 8.06816
R6518 VDD.n4056 VDD.n4053 8.06816
R6519 VDD.n4052 VDD.n4049 8.06816
R6520 VDD.n4048 VDD.n4045 8.06816
R6521 VDD.n4044 VDD.n4041 8.06816
R6522 VDD.n4040 VDD.n4037 8.06816
R6523 VDD.n4215 VDD.n4214 8.06816
R6524 VDD.n4219 VDD.n4218 8.06816
R6525 VDD.n4233 VDD.n4230 8.06816
R6526 VDD.n4229 VDD.n4226 8.06816
R6527 VDD.n4084 VDD.n4083 8.06816
R6528 VDD.n4088 VDD.n4087 8.06816
R6529 VDD.n4092 VDD.n4091 8.06816
R6530 VDD.n4096 VDD.n4095 8.06816
R6531 VDD.n4100 VDD.n4099 8.06816
R6532 VDD.n4196 VDD.n4193 8.06816
R6533 VDD.n4192 VDD.n4189 8.06816
R6534 VDD.n4188 VDD.n4185 8.06816
R6535 VDD.n4184 VDD.n4181 8.06816
R6536 VDD.n4180 VDD.n4177 8.06816
R6537 VDD.n4172 VDD.n4169 8.06816
R6538 VDD.n4168 VDD.n4165 8.06816
R6539 VDD.n4164 VDD.n4161 8.06816
R6540 VDD.n4160 VDD.n4157 8.06816
R6541 VDD.n4156 VDD.n4153 8.06816
R6542 VDD.n4152 VDD.n4149 8.06816
R6543 VDD.n4148 VDD.n4145 8.06816
R6544 VDD.n4144 VDD.n4141 8.06816
R6545 VDD.n4140 VDD.n4137 8.06816
R6546 VDD.n4136 VDD.n4133 8.06816
R6547 VDD.n4132 VDD.n4129 8.06816
R6548 VDD.n4128 VDD.n4125 8.06816
R6549 VDD.n8559 VDD.n8558 8.06816
R6550 VDD.n6660 VDD.t37 7.99076
R6551 VDD.n4692 VDD.n4691 7.45411
R6552 VDD.n4708 VDD.n4707 7.45411
R6553 VDD.n5033 VDD.n5032 7.45411
R6554 VDD.n5049 VDD.n5048 7.45411
R6555 VDD.n4330 VDD.n4329 7.45411
R6556 VDD.n4346 VDD.n4345 7.45411
R6557 VDD.n4413 VDD.n4412 7.45411
R6558 VDD.n4511 VDD.n4510 7.45411
R6559 VDD.n4441 VDD.n4440 7.45411
R6560 VDD.n4431 VDD.n4430 7.45411
R6561 VDD.n3650 VDD.n3649 7.45411
R6562 VDD.n5267 VDD.n5266 7.45411
R6563 VDD.n6562 VDD.t39 7.14968
R6564 VDD.n2633 VDD.n2632 7.09014
R6565 VDD.n3040 VDD.n2631 7.09014
R6566 VDD.n1781 VDD.n1780 7.09014
R6567 VDD.n2558 VDD.n1779 7.09014
R6568 VDD.n927 VDD.n926 7.09014
R6569 VDD.n1704 VDD.n925 7.09014
R6570 VDD.n72 VDD.n71 7.09014
R6571 VDD.n849 VDD.n70 7.09014
R6572 VDD.n2707 VDD.n2704 7.07692
R6573 VDD.n2704 VDD.n2701 7.07692
R6574 VDD.n2701 VDD.n2698 7.07692
R6575 VDD.n2698 VDD.n2695 7.07692
R6576 VDD.n2695 VDD.n2692 7.07692
R6577 VDD.n2692 VDD.n2689 7.07692
R6578 VDD.n2689 VDD.n2686 7.07692
R6579 VDD.n2686 VDD.n2683 7.07692
R6580 VDD.n2683 VDD.n2680 7.07692
R6581 VDD.n2680 VDD.n2677 7.07692
R6582 VDD.n2677 VDD.n2674 7.07692
R6583 VDD.n3072 VDD.n3069 7.07692
R6584 VDD.n3075 VDD.n3072 7.07692
R6585 VDD.n3078 VDD.n3075 7.07692
R6586 VDD.n3081 VDD.n3078 7.07692
R6587 VDD.n3084 VDD.n3081 7.07692
R6588 VDD.n3087 VDD.n3084 7.07692
R6589 VDD.n3090 VDD.n3087 7.07692
R6590 VDD.n3093 VDD.n3090 7.07692
R6591 VDD.n3096 VDD.n3093 7.07692
R6592 VDD.n3099 VDD.n3096 7.07692
R6593 VDD.n3102 VDD.n3099 7.07692
R6594 VDD.n3105 VDD.n3102 7.07692
R6595 VDD.n3108 VDD.n3105 7.07692
R6596 VDD.n2171 VDD.n2042 7.07692
R6597 VDD.n2165 VDD.n2042 7.07692
R6598 VDD.n2165 VDD.n2164 7.07692
R6599 VDD.n2164 VDD.n2163 7.07692
R6600 VDD.n2163 VDD.n2046 7.07692
R6601 VDD.n2157 VDD.n2046 7.07692
R6602 VDD.n2157 VDD.n2156 7.07692
R6603 VDD.n2156 VDD.n2155 7.07692
R6604 VDD.n2155 VDD.n2050 7.07692
R6605 VDD.n2149 VDD.n2050 7.07692
R6606 VDD.n2149 VDD.n2148 7.07692
R6607 VDD.n2148 VDD.n2147 7.07692
R6608 VDD.n2147 VDD.n2054 7.07692
R6609 VDD.n2141 VDD.n2054 7.07692
R6610 VDD.n2141 VDD.n2140 7.07692
R6611 VDD.n2140 VDD.n2139 7.07692
R6612 VDD.n2139 VDD.n2058 7.07692
R6613 VDD.n2133 VDD.n2058 7.07692
R6614 VDD.n2133 VDD.n2132 7.07692
R6615 VDD.n2132 VDD.n2131 7.07692
R6616 VDD.n2131 VDD.n2062 7.07692
R6617 VDD.n2125 VDD.n2062 7.07692
R6618 VDD.n2125 VDD.n2124 7.07692
R6619 VDD.n2124 VDD.n2123 7.07692
R6620 VDD.n2123 VDD.n2066 7.07692
R6621 VDD.n1317 VDD.n1188 7.07692
R6622 VDD.n1311 VDD.n1188 7.07692
R6623 VDD.n1311 VDD.n1310 7.07692
R6624 VDD.n1310 VDD.n1309 7.07692
R6625 VDD.n1309 VDD.n1192 7.07692
R6626 VDD.n1303 VDD.n1192 7.07692
R6627 VDD.n1303 VDD.n1302 7.07692
R6628 VDD.n1302 VDD.n1301 7.07692
R6629 VDD.n1301 VDD.n1196 7.07692
R6630 VDD.n1295 VDD.n1196 7.07692
R6631 VDD.n1295 VDD.n1294 7.07692
R6632 VDD.n1294 VDD.n1293 7.07692
R6633 VDD.n1293 VDD.n1200 7.07692
R6634 VDD.n1287 VDD.n1200 7.07692
R6635 VDD.n1287 VDD.n1286 7.07692
R6636 VDD.n1286 VDD.n1285 7.07692
R6637 VDD.n1285 VDD.n1204 7.07692
R6638 VDD.n1279 VDD.n1204 7.07692
R6639 VDD.n1279 VDD.n1278 7.07692
R6640 VDD.n1278 VDD.n1277 7.07692
R6641 VDD.n1277 VDD.n1208 7.07692
R6642 VDD.n1271 VDD.n1208 7.07692
R6643 VDD.n1271 VDD.n1270 7.07692
R6644 VDD.n1270 VDD.n1269 7.07692
R6645 VDD.n1269 VDD.n1212 7.07692
R6646 VDD.n462 VDD.n333 7.07692
R6647 VDD.n456 VDD.n333 7.07692
R6648 VDD.n456 VDD.n455 7.07692
R6649 VDD.n455 VDD.n454 7.07692
R6650 VDD.n454 VDD.n337 7.07692
R6651 VDD.n448 VDD.n337 7.07692
R6652 VDD.n448 VDD.n447 7.07692
R6653 VDD.n447 VDD.n446 7.07692
R6654 VDD.n446 VDD.n341 7.07692
R6655 VDD.n440 VDD.n341 7.07692
R6656 VDD.n440 VDD.n439 7.07692
R6657 VDD.n439 VDD.n438 7.07692
R6658 VDD.n438 VDD.n345 7.07692
R6659 VDD.n432 VDD.n345 7.07692
R6660 VDD.n432 VDD.n431 7.07692
R6661 VDD.n431 VDD.n430 7.07692
R6662 VDD.n430 VDD.n349 7.07692
R6663 VDD.n424 VDD.n349 7.07692
R6664 VDD.n424 VDD.n423 7.07692
R6665 VDD.n423 VDD.n422 7.07692
R6666 VDD.n422 VDD.n353 7.07692
R6667 VDD.n416 VDD.n353 7.07692
R6668 VDD.n416 VDD.n415 7.07692
R6669 VDD.n415 VDD.n414 7.07692
R6670 VDD.n414 VDD.n357 7.07692
R6671 VDD.n2373 VDD.n2219 7.05178
R6672 VDD.n2372 VDD.n2231 7.05178
R6673 VDD.n2365 VDD.n2237 7.05178
R6674 VDD.n2244 VDD.n2238 7.05178
R6675 VDD.n1519 VDD.n1365 7.05178
R6676 VDD.n1518 VDD.n1377 7.05178
R6677 VDD.n1511 VDD.n1383 7.05178
R6678 VDD.n1390 VDD.n1384 7.05178
R6679 VDD.n664 VDD.n510 7.05178
R6680 VDD.n663 VDD.n522 7.05178
R6681 VDD.n656 VDD.n528 7.05178
R6682 VDD.n535 VDD.n529 7.05178
R6683 VDD.n4203 VDD.n4200 6.89484
R6684 VDD.n4688 VDD.n4687 6.80334
R6685 VDD.n5029 VDD.n5028 6.80334
R6686 VDD.n4326 VDD.n4325 6.80334
R6687 VDD.n3646 VDD.n3645 6.80105
R6688 VDD.n5263 VDD.n5262 6.80105
R6689 VDD.n4704 VDD.n4703 6.80104
R6690 VDD.n5045 VDD.n5044 6.80104
R6691 VDD.n4507 VDD.n4506 6.80104
R6692 VDD.n3114 VDD.n3111 6.59444
R6693 VDD.n3116 VDD.n3114 6.59444
R6694 VDD.n3120 VDD.n3116 6.59444
R6695 VDD.n3123 VDD.n3120 6.59444
R6696 VDD.n3126 VDD.n3123 6.59444
R6697 VDD.n3129 VDD.n3126 6.59444
R6698 VDD.n3132 VDD.n3129 6.59444
R6699 VDD.n3135 VDD.n3132 6.59444
R6700 VDD.n3138 VDD.n3135 6.59444
R6701 VDD.n3141 VDD.n3138 6.59444
R6702 VDD.n3144 VDD.n3141 6.59444
R6703 VDD.n3147 VDD.n3144 6.59444
R6704 VDD.n3150 VDD.n3147 6.59444
R6705 VDD.n3153 VDD.n3150 6.59444
R6706 VDD.n3156 VDD.n3153 6.59444
R6707 VDD.n3159 VDD.n3156 6.59444
R6708 VDD.n3162 VDD.n3159 6.59444
R6709 VDD.n2116 VDD.n2115 6.59444
R6710 VDD.n2115 VDD.n2070 6.59444
R6711 VDD.n2110 VDD.n2070 6.59444
R6712 VDD.n2110 VDD.n2109 6.59444
R6713 VDD.n2109 VDD.n2108 6.59444
R6714 VDD.n2108 VDD.n2074 6.59444
R6715 VDD.n2102 VDD.n2074 6.59444
R6716 VDD.n2102 VDD.n2101 6.59444
R6717 VDD.n2101 VDD.n2100 6.59444
R6718 VDD.n2100 VDD.n2079 6.59444
R6719 VDD.n2094 VDD.n2079 6.59444
R6720 VDD.n2094 VDD.n2093 6.59444
R6721 VDD.n2093 VDD.n2092 6.59444
R6722 VDD.n2092 VDD.n2083 6.59444
R6723 VDD.n2086 VDD.n2083 6.59444
R6724 VDD.n2086 VDD.n2085 6.59444
R6725 VDD.n2085 VDD.n1812 6.59444
R6726 VDD.n1262 VDD.n1261 6.59444
R6727 VDD.n1261 VDD.n1216 6.59444
R6728 VDD.n1256 VDD.n1216 6.59444
R6729 VDD.n1256 VDD.n1255 6.59444
R6730 VDD.n1255 VDD.n1254 6.59444
R6731 VDD.n1254 VDD.n1220 6.59444
R6732 VDD.n1248 VDD.n1220 6.59444
R6733 VDD.n1248 VDD.n1247 6.59444
R6734 VDD.n1247 VDD.n1246 6.59444
R6735 VDD.n1246 VDD.n1225 6.59444
R6736 VDD.n1240 VDD.n1225 6.59444
R6737 VDD.n1240 VDD.n1239 6.59444
R6738 VDD.n1239 VDD.n1238 6.59444
R6739 VDD.n1238 VDD.n1229 6.59444
R6740 VDD.n1232 VDD.n1229 6.59444
R6741 VDD.n1232 VDD.n1231 6.59444
R6742 VDD.n1231 VDD.n958 6.59444
R6743 VDD.n407 VDD.n406 6.59444
R6744 VDD.n406 VDD.n361 6.59444
R6745 VDD.n401 VDD.n361 6.59444
R6746 VDD.n401 VDD.n400 6.59444
R6747 VDD.n400 VDD.n399 6.59444
R6748 VDD.n399 VDD.n365 6.59444
R6749 VDD.n393 VDD.n365 6.59444
R6750 VDD.n393 VDD.n392 6.59444
R6751 VDD.n392 VDD.n391 6.59444
R6752 VDD.n391 VDD.n370 6.59444
R6753 VDD.n385 VDD.n370 6.59444
R6754 VDD.n385 VDD.n384 6.59444
R6755 VDD.n384 VDD.n383 6.59444
R6756 VDD.n383 VDD.n374 6.59444
R6757 VDD.n377 VDD.n374 6.59444
R6758 VDD.n377 VDD.n376 6.59444
R6759 VDD.n376 VDD.n103 6.59444
R6760 VDD.n4124 VDD.t12 6.34882
R6761 VDD.n3892 VDD.n3891 6.31321
R6762 VDD.t112 VDD.n8779 6.3086
R6763 VDD.n2913 VDD.n2910 6.17355
R6764 VDD.n2910 VDD.n2907 6.17355
R6765 VDD.n2907 VDD.n2904 6.17355
R6766 VDD.n2904 VDD.n2901 6.17355
R6767 VDD.n2901 VDD.n2898 6.17355
R6768 VDD.n2898 VDD.n2895 6.17355
R6769 VDD.n2895 VDD.n2892 6.17355
R6770 VDD.n2892 VDD.n2889 6.17355
R6771 VDD.n2889 VDD.n2886 6.17355
R6772 VDD.n2886 VDD.n2883 6.17355
R6773 VDD.n2883 VDD.n2880 6.17355
R6774 VDD.n2880 VDD.n2877 6.17355
R6775 VDD.n2404 VDD.n2403 6.17355
R6776 VDD.n2405 VDD.n2404 6.17355
R6777 VDD.n2405 VDD.n1998 6.17355
R6778 VDD.n2411 VDD.n1998 6.17355
R6779 VDD.n2412 VDD.n2411 6.17355
R6780 VDD.n2413 VDD.n2412 6.17355
R6781 VDD.n2413 VDD.n1994 6.17355
R6782 VDD.n2419 VDD.n1994 6.17355
R6783 VDD.n2420 VDD.n2419 6.17355
R6784 VDD.n2421 VDD.n2420 6.17355
R6785 VDD.n2421 VDD.n1990 6.17355
R6786 VDD.n2427 VDD.n1990 6.17355
R6787 VDD.n1550 VDD.n1549 6.17355
R6788 VDD.n1551 VDD.n1550 6.17355
R6789 VDD.n1551 VDD.n1144 6.17355
R6790 VDD.n1557 VDD.n1144 6.17355
R6791 VDD.n1558 VDD.n1557 6.17355
R6792 VDD.n1559 VDD.n1558 6.17355
R6793 VDD.n1559 VDD.n1140 6.17355
R6794 VDD.n1565 VDD.n1140 6.17355
R6795 VDD.n1566 VDD.n1565 6.17355
R6796 VDD.n1567 VDD.n1566 6.17355
R6797 VDD.n1567 VDD.n1136 6.17355
R6798 VDD.n1573 VDD.n1136 6.17355
R6799 VDD.n695 VDD.n694 6.17355
R6800 VDD.n696 VDD.n695 6.17355
R6801 VDD.n696 VDD.n289 6.17355
R6802 VDD.n702 VDD.n289 6.17355
R6803 VDD.n703 VDD.n702 6.17355
R6804 VDD.n704 VDD.n703 6.17355
R6805 VDD.n704 VDD.n285 6.17355
R6806 VDD.n710 VDD.n285 6.17355
R6807 VDD.n711 VDD.n710 6.17355
R6808 VDD.n712 VDD.n711 6.17355
R6809 VDD.n712 VDD.n281 6.17355
R6810 VDD.n718 VDD.n281 6.17355
R6811 VDD.n4017 VDD.n4016 6.08431
R6812 VDD.n4627 VDD.n4626 6.02403
R6813 VDD.n5159 VDD.n5158 6.02403
R6814 VDD.n4281 VDD.n4280 6.02403
R6815 VDD.n5309 VDD.n5308 6.02403
R6816 VDD.n8613 VDD.n8612 6.02403
R6817 VDD.n8975 VDD.n8974 6.02403
R6818 VDD.n8885 VDD.n8884 6.02403
R6819 VDD.n7490 VDD.n7489 5.96815
R6820 VDD.t80 VDD.n4173 5.95205
R6821 VDD.n2671 VDD.n2669 5.80317
R6822 VDD.n2669 VDD.n2667 5.80317
R6823 VDD.n2667 VDD.n2665 5.80317
R6824 VDD.n3050 VDD.n3048 5.80317
R6825 VDD.n3055 VDD.n3053 5.80317
R6826 VDD.n3057 VDD.n3055 5.80317
R6827 VDD.n3059 VDD.n3057 5.80317
R6828 VDD.n3061 VDD.n3059 5.80317
R6829 VDD.n3063 VDD.n3061 5.80317
R6830 VDD.n2241 VDD.n2214 5.80317
R6831 VDD.n2363 VDD.n2241 5.80317
R6832 VDD.n2363 VDD.n2362 5.80317
R6833 VDD.n2362 VDD.n2361 5.80317
R6834 VDD.n2361 VDD.n2242 5.80317
R6835 VDD.n2266 VDD.n2261 5.80317
R6836 VDD.n2262 VDD.n2261 5.80317
R6837 VDD.n2262 VDD.n1806 5.80317
R6838 VDD.n2539 VDD.n1806 5.80317
R6839 VDD.n2539 VDD.n2538 5.80317
R6840 VDD.n1387 VDD.n1360 5.80317
R6841 VDD.n1509 VDD.n1387 5.80317
R6842 VDD.n1509 VDD.n1508 5.80317
R6843 VDD.n1508 VDD.n1507 5.80317
R6844 VDD.n1507 VDD.n1388 5.80317
R6845 VDD.n1412 VDD.n1407 5.80317
R6846 VDD.n1408 VDD.n1407 5.80317
R6847 VDD.n1408 VDD.n952 5.80317
R6848 VDD.n1685 VDD.n952 5.80317
R6849 VDD.n1685 VDD.n1684 5.80317
R6850 VDD.n532 VDD.n505 5.80317
R6851 VDD.n654 VDD.n532 5.80317
R6852 VDD.n654 VDD.n653 5.80317
R6853 VDD.n653 VDD.n652 5.80317
R6854 VDD.n652 VDD.n533 5.80317
R6855 VDD.n557 VDD.n552 5.80317
R6856 VDD.n553 VDD.n552 5.80317
R6857 VDD.n553 VDD.n97 5.80317
R6858 VDD.n830 VDD.n97 5.80317
R6859 VDD.n830 VDD.n829 5.80317
R6860 VDD.n5278 VDD.n5277 5.73742
R6861 VDD.n4690 VDD.n4689 5.64756
R6862 VDD.n4706 VDD.n4705 5.64756
R6863 VDD.n5031 VDD.n5030 5.64756
R6864 VDD.n5047 VDD.n5046 5.64756
R6865 VDD.n4328 VDD.n4327 5.64756
R6866 VDD.n4344 VDD.n4343 5.64756
R6867 VDD.n4411 VDD.n4410 5.64756
R6868 VDD.n4509 VDD.n4508 5.64756
R6869 VDD.n4439 VDD.n4438 5.64756
R6870 VDD.n4429 VDD.n4428 5.64756
R6871 VDD.n3648 VDD.n3647 5.64756
R6872 VDD.n5265 VDD.n5264 5.64756
R6873 VDD.n4797 VDD.n4796 5.63005
R6874 VDD.n4829 VDD.n4828 5.63005
R6875 VDD.n4859 VDD.n4858 5.63005
R6876 VDD.n4889 VDD.n4888 5.63005
R6877 VDD.n4919 VDD.n4918 5.63005
R6878 VDD.n4949 VDD.n4948 5.63005
R6879 VDD.n5140 VDD.n5139 5.63005
R6880 VDD.n3309 VDD.n3307 5.61598
R6881 VDD.n3307 VDD.n3304 5.61598
R6882 VDD.n3304 VDD.n3301 5.61598
R6883 VDD.n3301 VDD.n3298 5.61598
R6884 VDD.n3298 VDD.n3295 5.61598
R6885 VDD.n3295 VDD.n3292 5.61598
R6886 VDD.n3292 VDD.n3289 5.61598
R6887 VDD.n3289 VDD.n3286 5.61598
R6888 VDD.n3286 VDD.n3283 5.61598
R6889 VDD.n3283 VDD.n3280 5.61598
R6890 VDD.n3280 VDD.n3277 5.61598
R6891 VDD.n3277 VDD.n3274 5.61598
R6892 VDD.n2527 VDD.n1940 5.61598
R6893 VDD.n2527 VDD.n2526 5.61598
R6894 VDD.n2526 VDD.n2525 5.61598
R6895 VDD.n2525 VDD.n1941 5.61598
R6896 VDD.n2519 VDD.n1941 5.61598
R6897 VDD.n2519 VDD.n2518 5.61598
R6898 VDD.n2518 VDD.n2517 5.61598
R6899 VDD.n2517 VDD.n1945 5.61598
R6900 VDD.n2511 VDD.n1945 5.61598
R6901 VDD.n2511 VDD.n2510 5.61598
R6902 VDD.n2510 VDD.n2509 5.61598
R6903 VDD.n2509 VDD.n1949 5.61598
R6904 VDD.n1673 VDD.n1086 5.61598
R6905 VDD.n1673 VDD.n1672 5.61598
R6906 VDD.n1672 VDD.n1671 5.61598
R6907 VDD.n1671 VDD.n1087 5.61598
R6908 VDD.n1665 VDD.n1087 5.61598
R6909 VDD.n1665 VDD.n1664 5.61598
R6910 VDD.n1664 VDD.n1663 5.61598
R6911 VDD.n1663 VDD.n1091 5.61598
R6912 VDD.n1657 VDD.n1091 5.61598
R6913 VDD.n1657 VDD.n1656 5.61598
R6914 VDD.n1656 VDD.n1655 5.61598
R6915 VDD.n1655 VDD.n1095 5.61598
R6916 VDD.n818 VDD.n231 5.61598
R6917 VDD.n818 VDD.n817 5.61598
R6918 VDD.n817 VDD.n816 5.61598
R6919 VDD.n816 VDD.n232 5.61598
R6920 VDD.n810 VDD.n232 5.61598
R6921 VDD.n810 VDD.n809 5.61598
R6922 VDD.n809 VDD.n808 5.61598
R6923 VDD.n808 VDD.n236 5.61598
R6924 VDD.n802 VDD.n236 5.61598
R6925 VDD.n802 VDD.n801 5.61598
R6926 VDD.n801 VDD.n800 5.61598
R6927 VDD.n800 VDD.n240 5.61598
R6928 VDD.n5215 VDD.n5214 5.57349
R6929 VDD.n4675 VDD.n4674 5.57349
R6930 VDD.n4811 VDD.t81 5.5395
R6931 VDD.t100 VDD.n4811 5.5395
R6932 VDD.n4812 VDD.t100 5.5395
R6933 VDD.n4812 VDD.t13 5.5395
R6934 VDD.n4845 VDD.t144 5.5395
R6935 VDD.n4845 VDD.t46 5.5395
R6936 VDD.n4875 VDD.t11 5.5395
R6937 VDD.n4875 VDD.t114 5.5395
R6938 VDD.n4905 VDD.t115 5.5395
R6939 VDD.n4905 VDD.t111 5.5395
R6940 VDD.n4935 VDD.t132 5.5395
R6941 VDD.n4935 VDD.t1 5.5395
R6942 VDD.n3851 VDD.t3 5.5395
R6943 VDD.n3851 VDD.t139 5.5395
R6944 VDD.n3818 VDD.t138 5.5395
R6945 VDD.n3818 VDD.t98 5.5395
R6946 VDD.n5137 VDD.t91 5.5395
R6947 VDD.n4380 VDD.t83 5.5395
R6948 VDD.n4380 VDD.t78 5.5395
R6949 VDD.n4473 VDD.t88 5.5395
R6950 VDD.n4543 VDD.t86 5.5395
R6951 VDD.n3682 VDD.t103 5.5395
R6952 VDD.n3682 VDD.t126 5.5395
R6953 VDD.n3725 VDD.t124 5.5395
R6954 VDD.n3725 VDD.t94 5.5395
R6955 VDD.n8682 VDD.t38 5.5395
R6956 VDD.n8682 VDD.t42 5.5395
R6957 VDD.n4104 VDD.n4103 5.42303
R6958 VDD.n915 VDD 5.2805
R6959 VDD.n2624 VDD 5.2805
R6960 VDD.n8577 VDD.t137 5.27719
R6961 VDD.n4638 VDD.n4637 5.27109
R6962 VDD.n5170 VDD.n5169 5.27109
R6963 VDD.n8624 VDD.n8623 5.27109
R6964 VDD.n8986 VDD.n8985 5.27109
R6965 VDD.n8896 VDD.n8895 5.27109
R6966 VDD.n8653 VDD.n8652 5.25364
R6967 VDD.n8732 VDD.n8731 5.25364
R6968 VDD.n8932 VDD.n8931 5.25364
R6969 VDD.n2976 VDD.n2973 5.2318
R6970 VDD.n2293 VDD.n2292 5.2318
R6971 VDD.n1439 VDD.n1438 5.2318
R6972 VDD.n584 VDD.n583 5.2318
R6973 VDD.n4237 VDD.n4222 5.15851
R6974 VDD.n3661 VDD.n3660 4.96787
R6975 VDD.n4719 VDD.n4718 4.95584
R6976 VDD.n5060 VDD.n5059 4.95584
R6977 VDD.n4358 VDD.n4357 4.95584
R6978 VDD.n4452 VDD.n4451 4.95584
R6979 VDD.n4522 VDD.n4521 4.95584
R6980 VDD.n4297 VDD.n4291 4.89462
R6981 VDD.n5326 VDD.n5320 4.89462
R6982 VDD.n4029 VDD.n4028 4.894
R6983 VDD.n8854 VDD.n8852 4.89039
R6984 VDD.n3007 VDD.n3004 4.78659
R6985 VDD.n2355 VDD.n2354 4.78659
R6986 VDD.n1501 VDD.n1500 4.78659
R6987 VDD.n646 VDD.n645 4.78659
R6988 VDD.n3956 VDD.n3955 4.7505
R6989 VDD.n3958 VDD.n3957 4.7505
R6990 VDD.n3963 VDD.n3962 4.7505
R6991 VDD.n3961 VDD.n3960 4.7505
R6992 VDD.n4701 VDD.n4700 4.73575
R6993 VDD.n4716 VDD.n4702 4.73575
R6994 VDD.n5042 VDD.n5041 4.73575
R6995 VDD.n5057 VDD.n5043 4.73575
R6996 VDD.n4339 VDD.n4338 4.73575
R6997 VDD.n4355 VDD.n4354 4.73575
R6998 VDD.n4422 VDD.n4421 4.73575
R6999 VDD.n4519 VDD.n4505 4.73575
R7000 VDD.n4449 VDD.n4423 4.73575
R7001 VDD.n4504 VDD.n4503 4.73575
R7002 VDD.n3659 VDD.n3658 4.73575
R7003 VDD.n5276 VDD.n5275 4.73575
R7004 VDD.n2719 VDD.n2717 4.73093
R7005 VDD.n2722 VDD.n2719 4.73093
R7006 VDD.n2726 VDD.n2722 4.73093
R7007 VDD.n2729 VDD.n2726 4.73093
R7008 VDD.n2732 VDD.n2729 4.73093
R7009 VDD.n2735 VDD.n2732 4.73093
R7010 VDD.n2738 VDD.n2735 4.73093
R7011 VDD.n2741 VDD.n2738 4.73093
R7012 VDD.n2744 VDD.n2741 4.73093
R7013 VDD.n2747 VDD.n2744 4.73093
R7014 VDD.n2750 VDD.n2747 4.73093
R7015 VDD.n2753 VDD.n2750 4.73093
R7016 VDD.n2756 VDD.n2753 4.73093
R7017 VDD.n2759 VDD.n2756 4.73093
R7018 VDD.n2762 VDD.n2759 4.73093
R7019 VDD.n2765 VDD.n2762 4.73093
R7020 VDD.n2768 VDD.n2765 4.73093
R7021 VDD.n2179 VDD.n2178 4.73093
R7022 VDD.n2178 VDD.n2172 4.73093
R7023 VDD.n2172 VDD.n2036 4.73093
R7024 VDD.n2187 VDD.n2036 4.73093
R7025 VDD.n2188 VDD.n2187 4.73093
R7026 VDD.n2189 VDD.n2188 4.73093
R7027 VDD.n2189 VDD.n2032 4.73093
R7028 VDD.n2195 VDD.n2032 4.73093
R7029 VDD.n2196 VDD.n2195 4.73093
R7030 VDD.n2197 VDD.n2196 4.73093
R7031 VDD.n2197 VDD.n2028 4.73093
R7032 VDD.n2203 VDD.n2028 4.73093
R7033 VDD.n2204 VDD.n2203 4.73093
R7034 VDD.n2205 VDD.n2204 4.73093
R7035 VDD.n2205 VDD.n2024 4.73093
R7036 VDD.n2212 VDD.n2024 4.73093
R7037 VDD.n2213 VDD.n2212 4.73093
R7038 VDD.n1325 VDD.n1324 4.73093
R7039 VDD.n1324 VDD.n1318 4.73093
R7040 VDD.n1318 VDD.n1182 4.73093
R7041 VDD.n1333 VDD.n1182 4.73093
R7042 VDD.n1334 VDD.n1333 4.73093
R7043 VDD.n1335 VDD.n1334 4.73093
R7044 VDD.n1335 VDD.n1178 4.73093
R7045 VDD.n1341 VDD.n1178 4.73093
R7046 VDD.n1342 VDD.n1341 4.73093
R7047 VDD.n1343 VDD.n1342 4.73093
R7048 VDD.n1343 VDD.n1174 4.73093
R7049 VDD.n1349 VDD.n1174 4.73093
R7050 VDD.n1350 VDD.n1349 4.73093
R7051 VDD.n1351 VDD.n1350 4.73093
R7052 VDD.n1351 VDD.n1170 4.73093
R7053 VDD.n1358 VDD.n1170 4.73093
R7054 VDD.n1359 VDD.n1358 4.73093
R7055 VDD.n470 VDD.n469 4.73093
R7056 VDD.n469 VDD.n463 4.73093
R7057 VDD.n463 VDD.n327 4.73093
R7058 VDD.n478 VDD.n327 4.73093
R7059 VDD.n479 VDD.n478 4.73093
R7060 VDD.n480 VDD.n479 4.73093
R7061 VDD.n480 VDD.n323 4.73093
R7062 VDD.n486 VDD.n323 4.73093
R7063 VDD.n487 VDD.n486 4.73093
R7064 VDD.n488 VDD.n487 4.73093
R7065 VDD.n488 VDD.n319 4.73093
R7066 VDD.n494 VDD.n319 4.73093
R7067 VDD.n495 VDD.n494 4.73093
R7068 VDD.n496 VDD.n495 4.73093
R7069 VDD.n496 VDD.n315 4.73093
R7070 VDD.n503 VDD.n315 4.73093
R7071 VDD.n504 VDD.n503 4.73093
R7072 VDD.n20 VDD.n19 4.6533
R7073 VDD.n877 VDD.n876 4.6533
R7074 VDD.n1729 VDD.n1728 4.6533
R7075 VDD.n2576 VDD.n2575 4.6533
R7076 VDD.n4437 VDD.n4436 4.6505
R7077 VDD.n4342 VDD.n4341 4.6505
R7078 VDD.n3435 VDD.n3425 4.6505
R7079 VDD.n6824 VDD.n6823 4.6505
R7080 VDD.n6820 VDD.n6819 4.6505
R7081 VDD.n6816 VDD.n6815 4.6505
R7082 VDD.n6812 VDD.n6811 4.6505
R7083 VDD.n6808 VDD.n6807 4.6505
R7084 VDD.n6804 VDD.n6803 4.6505
R7085 VDD.n6799 VDD.n6798 4.6505
R7086 VDD.n6794 VDD.n6793 4.6505
R7087 VDD.n6786 VDD.n6785 4.6505
R7088 VDD.n6781 VDD.n6780 4.6505
R7089 VDD.n6776 VDD.n6775 4.6505
R7090 VDD.n6771 VDD.n6770 4.6505
R7091 VDD.n6766 VDD.n6765 4.6505
R7092 VDD.n6761 VDD.n6760 4.6505
R7093 VDD.n6756 VDD.n6755 4.6505
R7094 VDD.n6751 VDD.n6750 4.6505
R7095 VDD.n6746 VDD.n6745 4.6505
R7096 VDD.n6741 VDD.n6740 4.6505
R7097 VDD.n6736 VDD.n6735 4.6505
R7098 VDD.n6731 VDD.n6730 4.6505
R7099 VDD.n6726 VDD.n6725 4.6505
R7100 VDD.n6721 VDD.n6720 4.6505
R7101 VDD.n6716 VDD.n6715 4.6505
R7102 VDD.n6711 VDD.n6710 4.6505
R7103 VDD.n6706 VDD.n6705 4.6505
R7104 VDD.n6698 VDD.n6697 4.6505
R7105 VDD.n6694 VDD.n6693 4.6505
R7106 VDD.n6690 VDD.n6689 4.6505
R7107 VDD.n6686 VDD.n6685 4.6505
R7108 VDD.n6682 VDD.n6681 4.6505
R7109 VDD.n6678 VDD.n6677 4.6505
R7110 VDD.n6674 VDD.n6673 4.6505
R7111 VDD.n6653 VDD.n6652 4.6505
R7112 VDD.n6649 VDD.n6648 4.6505
R7113 VDD.n6645 VDD.n6644 4.6505
R7114 VDD.n6641 VDD.n6640 4.6505
R7115 VDD.n6637 VDD.n6636 4.6505
R7116 VDD.n6633 VDD.n6632 4.6505
R7117 VDD.n6629 VDD.n6628 4.6505
R7118 VDD.n6624 VDD.n6623 4.6505
R7119 VDD.n6619 VDD.n6618 4.6505
R7120 VDD.n6614 VDD.n6613 4.6505
R7121 VDD.n6606 VDD.n6605 4.6505
R7122 VDD.n6601 VDD.n6600 4.6505
R7123 VDD.n6596 VDD.n6595 4.6505
R7124 VDD.n6591 VDD.n6590 4.6505
R7125 VDD.n6586 VDD.n6585 4.6505
R7126 VDD.n6581 VDD.n6580 4.6505
R7127 VDD.n6576 VDD.n6575 4.6505
R7128 VDD.n6571 VDD.n6570 4.6505
R7129 VDD.n6566 VDD.n6565 4.6505
R7130 VDD.n6561 VDD.n6560 4.6505
R7131 VDD.n6556 VDD.n6555 4.6505
R7132 VDD.n6551 VDD.n6550 4.6505
R7133 VDD.n6546 VDD.n6545 4.6505
R7134 VDD.n6541 VDD.n6540 4.6505
R7135 VDD.n6536 VDD.n6535 4.6505
R7136 VDD.n6531 VDD.n6530 4.6505
R7137 VDD.n6526 VDD.n6525 4.6505
R7138 VDD.n6520 VDD.n6519 4.6505
R7139 VDD.n6516 VDD.n6515 4.6505
R7140 VDD.n6512 VDD.n6511 4.6505
R7141 VDD.n6508 VDD.n6507 4.6505
R7142 VDD.n8058 VDD.n8057 4.6505
R7143 VDD.n8066 VDD.n8065 4.6505
R7144 VDD.n8074 VDD.n8073 4.6505
R7145 VDD.n8082 VDD.n8081 4.6505
R7146 VDD.n8090 VDD.n8089 4.6505
R7147 VDD.n8098 VDD.n8097 4.6505
R7148 VDD.n8104 VDD.n8103 4.6505
R7149 VDD.n8112 VDD.n8111 4.6505
R7150 VDD.n8118 VDD.n8117 4.6505
R7151 VDD.n8126 VDD.n8125 4.6505
R7152 VDD.n8133 VDD.n8132 4.6505
R7153 VDD.n8142 VDD.n8141 4.6505
R7154 VDD.n8147 VDD.n8146 4.6505
R7155 VDD.n8153 VDD.n8152 4.6505
R7156 VDD.n8159 VDD.n8158 4.6505
R7157 VDD.n8165 VDD.n8164 4.6505
R7158 VDD.n8171 VDD.n8170 4.6505
R7159 VDD.n8177 VDD.n8176 4.6505
R7160 VDD.n8183 VDD.n8182 4.6505
R7161 VDD.n8191 VDD.n8190 4.6505
R7162 VDD.n8197 VDD.n8196 4.6505
R7163 VDD.n8205 VDD.n8204 4.6505
R7164 VDD.n8211 VDD.n8210 4.6505
R7165 VDD.n8217 VDD.n8216 4.6505
R7166 VDD.n8223 VDD.n8222 4.6505
R7167 VDD.n8229 VDD.n8228 4.6505
R7168 VDD.n8235 VDD.n8234 4.6505
R7169 VDD.n8241 VDD.n8240 4.6505
R7170 VDD.n8247 VDD.n8246 4.6505
R7171 VDD.n8252 VDD.n8251 4.6505
R7172 VDD.n8258 VDD.n8257 4.6505
R7173 VDD.n8264 VDD.n8263 4.6505
R7174 VDD.n8270 VDD.n8269 4.6505
R7175 VDD.n8276 VDD.n8275 4.6505
R7176 VDD.n8282 VDD.n8281 4.6505
R7177 VDD.n8288 VDD.n8287 4.6505
R7178 VDD.n8296 VDD.n8295 4.6505
R7179 VDD.n8302 VDD.n8301 4.6505
R7180 VDD.n8310 VDD.n8309 4.6505
R7181 VDD.n8316 VDD.n8315 4.6505
R7182 VDD.n8322 VDD.n8321 4.6505
R7183 VDD.n8328 VDD.n8327 4.6505
R7184 VDD.n8334 VDD.n8333 4.6505
R7185 VDD.n8340 VDD.n8339 4.6505
R7186 VDD.n8346 VDD.n8345 4.6505
R7187 VDD.n8352 VDD.n8351 4.6505
R7188 VDD.n8357 VDD.n8356 4.6505
R7189 VDD.n8363 VDD.n8362 4.6505
R7190 VDD.n8369 VDD.n8368 4.6505
R7191 VDD.n8375 VDD.n8374 4.6505
R7192 VDD.n8381 VDD.n8380 4.6505
R7193 VDD.n8387 VDD.n8386 4.6505
R7194 VDD.n8393 VDD.n8392 4.6505
R7195 VDD.n8401 VDD.n8400 4.6505
R7196 VDD.n8407 VDD.n8406 4.6505
R7197 VDD.n8419 VDD.n8418 4.6505
R7198 VDD.n8429 VDD.n8428 4.6505
R7199 VDD.n8439 VDD.n8438 4.6505
R7200 VDD.n8449 VDD.n8448 4.6505
R7201 VDD.n8459 VDD.n8458 4.6505
R7202 VDD.n8468 VDD.n8467 4.6505
R7203 VDD.n8477 VDD.n8476 4.6505
R7204 VDD.n8486 VDD.n8485 4.6505
R7205 VDD.n8494 VDD.n8493 4.6505
R7206 VDD.n8503 VDD.n8502 4.6505
R7207 VDD.n8512 VDD.n8511 4.6505
R7208 VDD.n8521 VDD.n8520 4.6505
R7209 VDD.n8529 VDD.n8528 4.6505
R7210 VDD.n8537 VDD.n8536 4.6505
R7211 VDD.n8543 VDD.n8542 4.6505
R7212 VDD.n8033 VDD.n8032 4.6505
R7213 VDD.n8025 VDD.n8024 4.6505
R7214 VDD.n8017 VDD.n8016 4.6505
R7215 VDD.n8009 VDD.n8008 4.6505
R7216 VDD.n8001 VDD.n8000 4.6505
R7217 VDD.n7993 VDD.n7992 4.6505
R7218 VDD.n7985 VDD.n7984 4.6505
R7219 VDD.n7977 VDD.n7976 4.6505
R7220 VDD.n7966 VDD.n7965 4.6505
R7221 VDD.n7958 VDD.n7957 4.6505
R7222 VDD.n7947 VDD.n7946 4.6505
R7223 VDD.n7939 VDD.n7938 4.6505
R7224 VDD.n7931 VDD.n7930 4.6505
R7225 VDD.n7923 VDD.n7922 4.6505
R7226 VDD.n7915 VDD.n7914 4.6505
R7227 VDD.n7907 VDD.n7906 4.6505
R7228 VDD.n7899 VDD.n7898 4.6505
R7229 VDD.n7891 VDD.n7890 4.6505
R7230 VDD.n7883 VDD.n7882 4.6505
R7231 VDD.n7875 VDD.n7874 4.6505
R7232 VDD.n7867 VDD.n7866 4.6505
R7233 VDD.n7859 VDD.n7858 4.6505
R7234 VDD.n7851 VDD.n7850 4.6505
R7235 VDD.n7843 VDD.n7842 4.6505
R7236 VDD.n7835 VDD.n7834 4.6505
R7237 VDD.n7825 VDD.n7824 4.6505
R7238 VDD.n7819 VDD.n7818 4.6505
R7239 VDD.n7811 VDD.n7810 4.6505
R7240 VDD.n7805 VDD.n7804 4.6505
R7241 VDD.n7799 VDD.n7798 4.6505
R7242 VDD.n7791 VDD.n7790 4.6505
R7243 VDD.n7783 VDD.n7782 4.6505
R7244 VDD.n7775 VDD.n7774 4.6505
R7245 VDD.n7767 VDD.n7766 4.6505
R7246 VDD.n7759 VDD.n7758 4.6505
R7247 VDD.n7751 VDD.n7750 4.6505
R7248 VDD.n7743 VDD.n7742 4.6505
R7249 VDD.n7735 VDD.n7734 4.6505
R7250 VDD.n7727 VDD.n7726 4.6505
R7251 VDD.n7719 VDD.n7718 4.6505
R7252 VDD.n7711 VDD.n7710 4.6505
R7253 VDD.n7703 VDD.n7702 4.6505
R7254 VDD.n7692 VDD.n7691 4.6505
R7255 VDD.n7684 VDD.n7683 4.6505
R7256 VDD.n7673 VDD.n7672 4.6505
R7257 VDD.n7665 VDD.n7664 4.6505
R7258 VDD.n7657 VDD.n7656 4.6505
R7259 VDD.n7649 VDD.n7648 4.6505
R7260 VDD.n7641 VDD.n7640 4.6505
R7261 VDD.n7636 VDD.n7635 4.6505
R7262 VDD.n8044 VDD.n8043 4.6505
R7263 VDD.n7601 VDD.n7600 4.6505
R7264 VDD.n7596 VDD.n7595 4.6505
R7265 VDD.n7591 VDD.n7590 4.6505
R7266 VDD.n7586 VDD.n7585 4.6505
R7267 VDD.n7581 VDD.n7580 4.6505
R7268 VDD.n7564 VDD.n7563 4.6505
R7269 VDD.n7557 VDD.n7556 4.6505
R7270 VDD.n7552 VDD.n7551 4.6505
R7271 VDD.n7547 VDD.n7546 4.6505
R7272 VDD.n7542 VDD.n7541 4.6505
R7273 VDD.n7537 VDD.n7536 4.6505
R7274 VDD.n7531 VDD.n7530 4.6505
R7275 VDD.n7526 VDD.n7525 4.6505
R7276 VDD.n7521 VDD.n7520 4.6505
R7277 VDD.n7516 VDD.n7515 4.6505
R7278 VDD.n7511 VDD.n7510 4.6505
R7279 VDD.n7506 VDD.n7505 4.6505
R7280 VDD.n7502 VDD.n7501 4.6505
R7281 VDD.n7496 VDD.n7495 4.6505
R7282 VDD.n7492 VDD.n7491 4.6505
R7283 VDD.n7488 VDD.n7487 4.6505
R7284 VDD.n7486 VDD.n7485 4.6505
R7285 VDD.n7480 VDD.n7479 4.6505
R7286 VDD.n7476 VDD.n7475 4.6505
R7287 VDD.n7472 VDD.n7471 4.6505
R7288 VDD.n7468 VDD.n7467 4.6505
R7289 VDD.n7464 VDD.n7463 4.6505
R7290 VDD.n7460 VDD.n7459 4.6505
R7291 VDD.n7456 VDD.n7455 4.6505
R7292 VDD.n7452 VDD.n7451 4.6505
R7293 VDD.n7448 VDD.n7447 4.6505
R7294 VDD.n7445 VDD.n7444 4.6505
R7295 VDD.n7441 VDD.n7440 4.6505
R7296 VDD.n7437 VDD.n7436 4.6505
R7297 VDD.n7433 VDD.n7432 4.6505
R7298 VDD.n7429 VDD.n7428 4.6505
R7299 VDD.n7425 VDD.n7424 4.6505
R7300 VDD.n7421 VDD.n7420 4.6505
R7301 VDD.n7417 VDD.n7416 4.6505
R7302 VDD.n7411 VDD.n7410 4.6505
R7303 VDD.n7407 VDD.n7406 4.6505
R7304 VDD.n7403 VDD.n7402 4.6505
R7305 VDD.n7399 VDD.n7398 4.6505
R7306 VDD.n7395 VDD.n7394 4.6505
R7307 VDD.n7391 VDD.n7390 4.6505
R7308 VDD.n7387 VDD.n7386 4.6505
R7309 VDD.n7383 VDD.n7382 4.6505
R7310 VDD.n7379 VDD.n7378 4.6505
R7311 VDD.n7376 VDD.n7375 4.6505
R7312 VDD.n7372 VDD.n7371 4.6505
R7313 VDD.n7368 VDD.n7367 4.6505
R7314 VDD.n7364 VDD.n7363 4.6505
R7315 VDD.n7360 VDD.n7359 4.6505
R7316 VDD.n7356 VDD.n7355 4.6505
R7317 VDD.n7352 VDD.n7351 4.6505
R7318 VDD.n7348 VDD.n7347 4.6505
R7319 VDD.n7342 VDD.n7341 4.6505
R7320 VDD.n7337 VDD.n7336 4.6505
R7321 VDD.n7332 VDD.n7331 4.6505
R7322 VDD.n7327 VDD.n7326 4.6505
R7323 VDD.n7322 VDD.n7321 4.6505
R7324 VDD.n7317 VDD.n7316 4.6505
R7325 VDD.n7312 VDD.n7311 4.6505
R7326 VDD.n7307 VDD.n7306 4.6505
R7327 VDD.n7302 VDD.n7301 4.6505
R7328 VDD.n7298 VDD.n7297 4.6505
R7329 VDD.n7293 VDD.n7292 4.6505
R7330 VDD.n7288 VDD.n7287 4.6505
R7331 VDD.n7283 VDD.n7282 4.6505
R7332 VDD.n7278 VDD.n7277 4.6505
R7333 VDD.n7273 VDD.n7272 4.6505
R7334 VDD.n7268 VDD.n7267 4.6505
R7335 VDD.n7263 VDD.n7262 4.6505
R7336 VDD.n7255 VDD.n7254 4.6505
R7337 VDD.n7250 VDD.n7249 4.6505
R7338 VDD.n7245 VDD.n7244 4.6505
R7339 VDD.n7240 VDD.n7239 4.6505
R7340 VDD.n7235 VDD.n7234 4.6505
R7341 VDD.n7230 VDD.n7229 4.6505
R7342 VDD.n7225 VDD.n7224 4.6505
R7343 VDD.n7220 VDD.n7219 4.6505
R7344 VDD.n7215 VDD.n7214 4.6505
R7345 VDD.n7211 VDD.n7210 4.6505
R7346 VDD.n7206 VDD.n7205 4.6505
R7347 VDD.n7201 VDD.n7200 4.6505
R7348 VDD.n7196 VDD.n7195 4.6505
R7349 VDD.n7191 VDD.n7190 4.6505
R7350 VDD.n7186 VDD.n7185 4.6505
R7351 VDD.n7181 VDD.n7180 4.6505
R7352 VDD.n7176 VDD.n7175 4.6505
R7353 VDD.n7168 VDD.n7167 4.6505
R7354 VDD.n7163 VDD.n7162 4.6505
R7355 VDD.n7158 VDD.n7157 4.6505
R7356 VDD.n7153 VDD.n7152 4.6505
R7357 VDD.n7148 VDD.n7147 4.6505
R7358 VDD.n7143 VDD.n7142 4.6505
R7359 VDD.n7138 VDD.n7137 4.6505
R7360 VDD.n7133 VDD.n7132 4.6505
R7361 VDD.n5832 VDD.n5831 4.6505
R7362 VDD.n5827 VDD.n5826 4.6505
R7363 VDD.n5822 VDD.n5821 4.6505
R7364 VDD.n5817 VDD.n5816 4.6505
R7365 VDD.n5812 VDD.n5811 4.6505
R7366 VDD.n5807 VDD.n5806 4.6505
R7367 VDD.n5802 VDD.n5801 4.6505
R7368 VDD.n5797 VDD.n5796 4.6505
R7369 VDD.n5792 VDD.n5791 4.6505
R7370 VDD.n5787 VDD.n5786 4.6505
R7371 VDD.n5782 VDD.n5781 4.6505
R7372 VDD.n5774 VDD.n5773 4.6505
R7373 VDD.n5769 VDD.n5768 4.6505
R7374 VDD.n5764 VDD.n5763 4.6505
R7375 VDD.n5759 VDD.n5758 4.6505
R7376 VDD.n5754 VDD.n5753 4.6505
R7377 VDD.n5749 VDD.n5748 4.6505
R7378 VDD.n5744 VDD.n5743 4.6505
R7379 VDD.n5739 VDD.n5738 4.6505
R7380 VDD.n5734 VDD.n5733 4.6505
R7381 VDD.n5729 VDD.n5728 4.6505
R7382 VDD.n5724 VDD.n5723 4.6505
R7383 VDD.n5719 VDD.n5718 4.6505
R7384 VDD.n5714 VDD.n5713 4.6505
R7385 VDD.n5709 VDD.n5708 4.6505
R7386 VDD.n5704 VDD.n5703 4.6505
R7387 VDD.n5699 VDD.n5698 4.6505
R7388 VDD.n5694 VDD.n5693 4.6505
R7389 VDD.n5686 VDD.n5685 4.6505
R7390 VDD.n5681 VDD.n5680 4.6505
R7391 VDD.n5676 VDD.n5675 4.6505
R7392 VDD.n5671 VDD.n5670 4.6505
R7393 VDD.n5666 VDD.n5665 4.6505
R7394 VDD.n5661 VDD.n5660 4.6505
R7395 VDD.n5656 VDD.n5655 4.6505
R7396 VDD.n5651 VDD.n5650 4.6505
R7397 VDD.n5646 VDD.n5645 4.6505
R7398 VDD.n5641 VDD.n5640 4.6505
R7399 VDD.n5636 VDD.n5635 4.6505
R7400 VDD.n5631 VDD.n5630 4.6505
R7401 VDD.n5626 VDD.n5625 4.6505
R7402 VDD.n5621 VDD.n5620 4.6505
R7403 VDD.n5616 VDD.n5615 4.6505
R7404 VDD.n5611 VDD.n5610 4.6505
R7405 VDD.n5606 VDD.n5605 4.6505
R7406 VDD.n5598 VDD.n5597 4.6505
R7407 VDD.n5593 VDD.n5592 4.6505
R7408 VDD.n5588 VDD.n5587 4.6505
R7409 VDD.n5583 VDD.n5582 4.6505
R7410 VDD.n5578 VDD.n5577 4.6505
R7411 VDD.n5573 VDD.n5572 4.6505
R7412 VDD.n5568 VDD.n5567 4.6505
R7413 VDD.n5563 VDD.n5562 4.6505
R7414 VDD.n5558 VDD.n5557 4.6505
R7415 VDD.n5553 VDD.n5552 4.6505
R7416 VDD.n5548 VDD.n5547 4.6505
R7417 VDD.n5543 VDD.n5542 4.6505
R7418 VDD.n5538 VDD.n5537 4.6505
R7419 VDD.n5533 VDD.n5532 4.6505
R7420 VDD.n5528 VDD.n5527 4.6505
R7421 VDD.n5523 VDD.n5522 4.6505
R7422 VDD.n5518 VDD.n5517 4.6505
R7423 VDD.n5510 VDD.n5509 4.6505
R7424 VDD.n5505 VDD.n5504 4.6505
R7425 VDD.n5500 VDD.n5499 4.6505
R7426 VDD.n5495 VDD.n5494 4.6505
R7427 VDD.n5490 VDD.n5489 4.6505
R7428 VDD.n5485 VDD.n5484 4.6505
R7429 VDD.n5480 VDD.n5479 4.6505
R7430 VDD.n5475 VDD.n5474 4.6505
R7431 VDD.n5470 VDD.n5469 4.6505
R7432 VDD.n5465 VDD.n5464 4.6505
R7433 VDD.n5460 VDD.n5459 4.6505
R7434 VDD.n5455 VDD.n5454 4.6505
R7435 VDD.n6831 VDD.n6830 4.6505
R7436 VDD.n6836 VDD.n6835 4.6505
R7437 VDD.n6841 VDD.n6840 4.6505
R7438 VDD.n6846 VDD.n6845 4.6505
R7439 VDD.n6854 VDD.n6853 4.6505
R7440 VDD.n6859 VDD.n6858 4.6505
R7441 VDD.n6864 VDD.n6863 4.6505
R7442 VDD.n6869 VDD.n6868 4.6505
R7443 VDD.n6874 VDD.n6873 4.6505
R7444 VDD.n6879 VDD.n6878 4.6505
R7445 VDD.n6884 VDD.n6883 4.6505
R7446 VDD.n6889 VDD.n6888 4.6505
R7447 VDD.n6894 VDD.n6893 4.6505
R7448 VDD.n6899 VDD.n6898 4.6505
R7449 VDD.n6904 VDD.n6903 4.6505
R7450 VDD.n6909 VDD.n6908 4.6505
R7451 VDD.n6914 VDD.n6913 4.6505
R7452 VDD.n6919 VDD.n6918 4.6505
R7453 VDD.n6924 VDD.n6923 4.6505
R7454 VDD.n6929 VDD.n6928 4.6505
R7455 VDD.n6934 VDD.n6933 4.6505
R7456 VDD.n6942 VDD.n6941 4.6505
R7457 VDD.n6947 VDD.n6946 4.6505
R7458 VDD.n6952 VDD.n6951 4.6505
R7459 VDD.n6957 VDD.n6956 4.6505
R7460 VDD.n6962 VDD.n6961 4.6505
R7461 VDD.n6967 VDD.n6966 4.6505
R7462 VDD.n6972 VDD.n6971 4.6505
R7463 VDD.n6977 VDD.n6976 4.6505
R7464 VDD.n6982 VDD.n6981 4.6505
R7465 VDD.n6987 VDD.n6986 4.6505
R7466 VDD.n6992 VDD.n6991 4.6505
R7467 VDD.n6997 VDD.n6996 4.6505
R7468 VDD.n7002 VDD.n7001 4.6505
R7469 VDD.n7007 VDD.n7006 4.6505
R7470 VDD.n7012 VDD.n7011 4.6505
R7471 VDD.n7017 VDD.n7016 4.6505
R7472 VDD.n7022 VDD.n7021 4.6505
R7473 VDD.n7030 VDD.n7029 4.6505
R7474 VDD.n7035 VDD.n7034 4.6505
R7475 VDD.n7040 VDD.n7039 4.6505
R7476 VDD.n7045 VDD.n7044 4.6505
R7477 VDD.n7050 VDD.n7049 4.6505
R7478 VDD.n7055 VDD.n7054 4.6505
R7479 VDD.n7060 VDD.n7059 4.6505
R7480 VDD.n7065 VDD.n7064 4.6505
R7481 VDD.n7070 VDD.n7069 4.6505
R7482 VDD.n7075 VDD.n7074 4.6505
R7483 VDD.n7080 VDD.n7079 4.6505
R7484 VDD.n7085 VDD.n7084 4.6505
R7485 VDD.n7090 VDD.n7089 4.6505
R7486 VDD.n7095 VDD.n7094 4.6505
R7487 VDD.n7100 VDD.n7099 4.6505
R7488 VDD.n7105 VDD.n7104 4.6505
R7489 VDD.n7110 VDD.n7109 4.6505
R7490 VDD.n7125 VDD.n7124 4.6505
R7491 VDD.n6493 VDD.n6492 4.6505
R7492 VDD.n6488 VDD.n6487 4.6505
R7493 VDD.n6484 VDD.n6483 4.6505
R7494 VDD.n6479 VDD.n6478 4.6505
R7495 VDD.n6475 VDD.n6474 4.6505
R7496 VDD.n6470 VDD.n6469 4.6505
R7497 VDD.n6466 VDD.n6465 4.6505
R7498 VDD.n6459 VDD.n6458 4.6505
R7499 VDD.n6455 VDD.n6454 4.6505
R7500 VDD.n6450 VDD.n6449 4.6505
R7501 VDD.n6446 VDD.n6445 4.6505
R7502 VDD.n6441 VDD.n6440 4.6505
R7503 VDD.n6437 VDD.n6436 4.6505
R7504 VDD.n6432 VDD.n6431 4.6505
R7505 VDD.n6428 VDD.n6427 4.6505
R7506 VDD.n6423 VDD.n6422 4.6505
R7507 VDD.n6418 VDD.n6417 4.6505
R7508 VDD.n6414 VDD.n6413 4.6505
R7509 VDD.n6409 VDD.n6408 4.6505
R7510 VDD.n6405 VDD.n6404 4.6505
R7511 VDD.n6400 VDD.n6399 4.6505
R7512 VDD.n6396 VDD.n6395 4.6505
R7513 VDD.n6391 VDD.n6390 4.6505
R7514 VDD.n6387 VDD.n6386 4.6505
R7515 VDD.n6380 VDD.n6379 4.6505
R7516 VDD.n6376 VDD.n6375 4.6505
R7517 VDD.n6371 VDD.n6370 4.6505
R7518 VDD.n6366 VDD.n6365 4.6505
R7519 VDD.n6361 VDD.n6360 4.6505
R7520 VDD.n6356 VDD.n6355 4.6505
R7521 VDD.n6351 VDD.n6350 4.6505
R7522 VDD.n6346 VDD.n6345 4.6505
R7523 VDD.n6341 VDD.n6340 4.6505
R7524 VDD.n6336 VDD.n6335 4.6505
R7525 VDD.n6331 VDD.n6330 4.6505
R7526 VDD.n6326 VDD.n6325 4.6505
R7527 VDD.n6321 VDD.n6320 4.6505
R7528 VDD.n6316 VDD.n6315 4.6505
R7529 VDD.n6311 VDD.n6310 4.6505
R7530 VDD.n6306 VDD.n6305 4.6505
R7531 VDD.n6301 VDD.n6300 4.6505
R7532 VDD.n6293 VDD.n6292 4.6505
R7533 VDD.n6288 VDD.n6287 4.6505
R7534 VDD.n6283 VDD.n6282 4.6505
R7535 VDD.n6278 VDD.n6277 4.6505
R7536 VDD.n6273 VDD.n6272 4.6505
R7537 VDD.n6268 VDD.n6267 4.6505
R7538 VDD.n6263 VDD.n6262 4.6505
R7539 VDD.n6258 VDD.n6257 4.6505
R7540 VDD.n6253 VDD.n6252 4.6505
R7541 VDD.n6248 VDD.n6247 4.6505
R7542 VDD.n6243 VDD.n6242 4.6505
R7543 VDD.n6238 VDD.n6237 4.6505
R7544 VDD.n6233 VDD.n6232 4.6505
R7545 VDD.n6228 VDD.n6227 4.6505
R7546 VDD.n6223 VDD.n6222 4.6505
R7547 VDD.n6219 VDD.n6218 4.6505
R7548 VDD.n6215 VDD.n6214 4.6505
R7549 VDD.n6209 VDD.n6208 4.6505
R7550 VDD.n6205 VDD.n6204 4.6505
R7551 VDD.n6201 VDD.n6200 4.6505
R7552 VDD.n6197 VDD.n6196 4.6505
R7553 VDD.n6193 VDD.n6192 4.6505
R7554 VDD.n6189 VDD.n6188 4.6505
R7555 VDD.n6185 VDD.n6184 4.6505
R7556 VDD.n6181 VDD.n6180 4.6505
R7557 VDD.n6177 VDD.n6176 4.6505
R7558 VDD.n6173 VDD.n6172 4.6505
R7559 VDD.n6169 VDD.n6168 4.6505
R7560 VDD.n6165 VDD.n6164 4.6505
R7561 VDD.n6161 VDD.n6160 4.6505
R7562 VDD.n6157 VDD.n6156 4.6505
R7563 VDD.n6153 VDD.n6152 4.6505
R7564 VDD.n6149 VDD.n6148 4.6505
R7565 VDD.n6145 VDD.n6144 4.6505
R7566 VDD.n6139 VDD.n6138 4.6505
R7567 VDD.n6135 VDD.n6134 4.6505
R7568 VDD.n6131 VDD.n6130 4.6505
R7569 VDD.n6127 VDD.n6126 4.6505
R7570 VDD.n6123 VDD.n6122 4.6505
R7571 VDD.n6119 VDD.n6118 4.6505
R7572 VDD.n6115 VDD.n6114 4.6505
R7573 VDD.n6111 VDD.n6110 4.6505
R7574 VDD.n6107 VDD.n6106 4.6505
R7575 VDD.n6103 VDD.n6102 4.6505
R7576 VDD.n6099 VDD.n6098 4.6505
R7577 VDD.n6095 VDD.n6094 4.6505
R7578 VDD.n6091 VDD.n6090 4.6505
R7579 VDD.n6087 VDD.n6086 4.6505
R7580 VDD.n6083 VDD.n6082 4.6505
R7581 VDD.n6079 VDD.n6078 4.6505
R7582 VDD.n6075 VDD.n6074 4.6505
R7583 VDD.n6069 VDD.n6068 4.6505
R7584 VDD.n6065 VDD.n6064 4.6505
R7585 VDD.n6061 VDD.n6060 4.6505
R7586 VDD.n6057 VDD.n6056 4.6505
R7587 VDD.n6052 VDD.n6051 4.6505
R7588 VDD.n6047 VDD.n6046 4.6505
R7589 VDD.n6042 VDD.n6041 4.6505
R7590 VDD.n6037 VDD.n6036 4.6505
R7591 VDD.n6032 VDD.n6031 4.6505
R7592 VDD.n6027 VDD.n6026 4.6505
R7593 VDD.n6022 VDD.n6021 4.6505
R7594 VDD.n6017 VDD.n6016 4.6505
R7595 VDD.n6012 VDD.n6011 4.6505
R7596 VDD.n6007 VDD.n6006 4.6505
R7597 VDD.n6002 VDD.n6001 4.6505
R7598 VDD.n5997 VDD.n5996 4.6505
R7599 VDD.n5992 VDD.n5991 4.6505
R7600 VDD.n5984 VDD.n5983 4.6505
R7601 VDD.n5979 VDD.n5978 4.6505
R7602 VDD.n5974 VDD.n5973 4.6505
R7603 VDD.n5969 VDD.n5968 4.6505
R7604 VDD.n5964 VDD.n5963 4.6505
R7605 VDD.n5959 VDD.n5958 4.6505
R7606 VDD.n5954 VDD.n5953 4.6505
R7607 VDD.n5949 VDD.n5948 4.6505
R7608 VDD.n5944 VDD.n5943 4.6505
R7609 VDD.n5939 VDD.n5938 4.6505
R7610 VDD.n5934 VDD.n5933 4.6505
R7611 VDD.n5929 VDD.n5928 4.6505
R7612 VDD.n5924 VDD.n5923 4.6505
R7613 VDD.n5919 VDD.n5918 4.6505
R7614 VDD.n5914 VDD.n5913 4.6505
R7615 VDD.n5909 VDD.n5908 4.6505
R7616 VDD.n5904 VDD.n5903 4.6505
R7617 VDD.n5896 VDD.n5895 4.6505
R7618 VDD.n5891 VDD.n5890 4.6505
R7619 VDD.n5886 VDD.n5885 4.6505
R7620 VDD.n5881 VDD.n5880 4.6505
R7621 VDD.n5876 VDD.n5875 4.6505
R7622 VDD.n5871 VDD.n5870 4.6505
R7623 VDD.n5866 VDD.n5865 4.6505
R7624 VDD.n6503 VDD.n6502 4.6505
R7625 VDD.n5856 VDD.n5855 4.6505
R7626 VDD.n5851 VDD.n5850 4.6505
R7627 VDD.n5846 VDD.n5845 4.6505
R7628 VDD.n5861 VDD.n5860 4.6505
R7629 VDD.n54 VDD.n40 4.6505
R7630 VDD.n53 VDD.n52 4.6505
R7631 VDD.n51 VDD.n42 4.6505
R7632 VDD.n50 VDD.n49 4.6505
R7633 VDD.n23 VDD.n11 4.6505
R7634 VDD.n30 VDD.n29 4.6505
R7635 VDD.n14 VDD.n7 4.6505
R7636 VDD VDD.n61 4.6505
R7637 VDD.n13 VDD.n6 4.6505
R7638 VDD.n16 VDD.n13 4.6505
R7639 VDD.n22 VDD.n21 4.6505
R7640 VDD.n905 VDD.n902 4.6505
R7641 VDD.n904 VDD.n903 4.6505
R7642 VDD.n859 VDD.n858 4.6505
R7643 VDD.n911 VDD.n910 4.6505
R7644 VDD.n872 VDD.n868 4.6505
R7645 VDD.n883 VDD.n882 4.6505
R7646 VDD.n889 VDD.n863 4.6505
R7647 VDD.n893 VDD 4.6505
R7648 VDD.n892 VDD.n891 4.6505
R7649 VDD.n891 VDD.n865 4.6505
R7650 VDD.n871 VDD.n870 4.6505
R7651 VDD.n1763 VDD.n1749 4.6505
R7652 VDD.n1762 VDD.n1761 4.6505
R7653 VDD.n1760 VDD.n1751 4.6505
R7654 VDD.n1759 VDD.n1758 4.6505
R7655 VDD.n1732 VDD.n1720 4.6505
R7656 VDD.n1739 VDD.n1738 4.6505
R7657 VDD.n1723 VDD.n1716 4.6505
R7658 VDD VDD.n1770 4.6505
R7659 VDD.n1722 VDD.n1715 4.6505
R7660 VDD.n1725 VDD.n1722 4.6505
R7661 VDD.n1731 VDD.n1730 4.6505
R7662 VDD.n2607 VDD.n2606 4.6505
R7663 VDD.n2610 VDD.n2609 4.6505
R7664 VDD.n2613 VDD.n2612 4.6505
R7665 VDD.n2620 VDD.n2619 4.6505
R7666 VDD.n2583 VDD.n2582 4.6505
R7667 VDD.n2588 VDD.n2587 4.6505
R7668 VDD.n2595 VDD.n2592 4.6505
R7669 VDD VDD.n2598 4.6505
R7670 VDD.n2572 VDD.n2571 4.6505
R7671 VDD.n7131 VDD.n7127 4.58155
R7672 VDD.n4649 VDD.n4648 4.51815
R7673 VDD.n5181 VDD.n5180 4.51815
R7674 VDD.n4403 VDD.n4402 4.51815
R7675 VDD.n4496 VDD.n4495 4.51815
R7676 VDD.n4566 VDD.n4565 4.51815
R7677 VDD.n4318 VDD.n4317 4.51815
R7678 VDD.n3705 VDD.n3704 4.51815
R7679 VDD.n3748 VDD.n3747 4.51815
R7680 VDD.n5347 VDD.n5346 4.51815
R7681 VDD.n8600 VDD.n8599 4.51815
R7682 VDD.n8609 VDD.n8608 4.51815
R7683 VDD.n8678 VDD.n8677 4.51815
R7684 VDD.n8729 VDD.n8728 4.51815
R7685 VDD.n8971 VDD.n8970 4.51815
R7686 VDD.n8879 VDD.n8878 4.51815
R7687 VDD.n8912 VDD.n8911 4.51815
R7688 VDD.n4472 VDD.n4409 4.5005
R7689 VDD.n4542 VDD.n4502 4.5005
R7690 VDD.n4378 VDD.n4324 4.5005
R7691 VDD.n4556 VDD.n4555 4.5005
R7692 VDD.n4562 VDD.n4561 4.5005
R7693 VDD.n4479 VDD.n4478 4.5005
R7694 VDD.n4549 VDD.n4548 4.5005
R7695 VDD.n4393 VDD.n4392 4.5005
R7696 VDD.n4305 VDD.n4304 4.5005
R7697 VDD.n4314 VDD.n4313 4.5005
R7698 VDD.n4399 VDD.n4398 4.5005
R7699 VDD.n4386 VDD.n4385 4.5005
R7700 VDD.n4486 VDD.n4485 4.5005
R7701 VDD.n4492 VDD.n4491 4.5005
R7702 VDD.n4298 VDD.n4297 4.5005
R7703 VDD.n3681 VDD.n3644 4.5005
R7704 VDD.n5306 VDD.n5261 4.5005
R7705 VDD.n5327 VDD.n5326 4.5005
R7706 VDD.n3738 VDD.n3737 4.5005
R7707 VDD.n3744 VDD.n3743 4.5005
R7708 VDD.n3688 VDD.n3687 4.5005
R7709 VDD.n3695 VDD.n3694 4.5005
R7710 VDD.n3701 VDD.n3700 4.5005
R7711 VDD.n3731 VDD.n3730 4.5005
R7712 VDD.n5334 VDD.n5333 4.5005
R7713 VDD.n5343 VDD.n5342 4.5005
R7714 VDD.n8657 VDD.n8656 4.5005
R7715 VDD.n8705 VDD.n8704 4.5005
R7716 VDD.n8736 VDD.n8735 4.5005
R7717 VDD.n8936 VDD.n8935 4.5005
R7718 VDD.n8997 VDD.n8972 4.5005
R7719 VDD.n9001 VDD.n8965 4.5005
R7720 VDD.n9011 VDD.n9010 4.5005
R7721 VDD.n8635 VDD.n8610 4.5005
R7722 VDD.n8639 VDD.n8603 4.5005
R7723 VDD.n8648 VDD.n8647 4.5005
R7724 VDD.n8712 VDD.n8711 4.5005
R7725 VDD.n8747 VDD.n8746 4.5005
R7726 VDD.n8947 VDD.n8946 4.5005
R7727 VDD.n8927 VDD.n8926 4.5005
R7728 VDD.n8668 VDD.n8667 4.5005
R7729 VDD.n8687 VDD.n8686 4.5005
R7730 VDD.n8691 VDD.n8681 4.5005
R7731 VDD.n8696 VDD.n8695 4.5005
R7732 VDD.n8914 VDD.n8913 4.5005
R7733 VDD.n8918 VDD.n8882 4.5005
R7734 VDD.n8871 VDD.n8870 4.5005
R7735 VDD.n8809 VDD.n8808 4.5005
R7736 VDD.n3898 VDD.n3897 4.5005
R7737 VDD.n3916 VDD.n3888 4.5005
R7738 VDD.n3907 VDD.n3906 4.5005
R7739 VDD.n3925 VDD.n3924 4.5005
R7740 VDD.n3928 VDD.n3883 4.5005
R7741 VDD.n3935 VDD.n3934 4.5005
R7742 VDD.n3938 VDD.n3880 4.5005
R7743 VDD.n5124 VDD.n5027 4.5005
R7744 VDD.n3816 VDD.n3815 4.5005
R7745 VDD.n5009 VDD.n5008 4.5005
R7746 VDD.n4945 VDD.n4931 4.5005
R7747 VDD.n5207 VDD.n5156 4.5005
R7748 VDD.n5201 VDD.n5200 4.5005
R7749 VDD.n5134 VDD.n5133 4.5005
R7750 VDD.n5016 VDD.n5014 4.5005
R7751 VDD.n3843 VDD.n3840 4.5005
R7752 VDD.n3836 VDD.n3835 4.5005
R7753 VDD.n3855 VDD.n3850 4.5005
R7754 VDD.n4909 VDD.n4904 4.5005
R7755 VDD.n4939 VDD.n4934 4.5005
R7756 VDD.n4879 VDD.n4874 4.5005
R7757 VDD.n4885 VDD.n4871 4.5005
R7758 VDD.n4915 VDD.n4901 4.5005
R7759 VDD.n4855 VDD.n4841 4.5005
R7760 VDD.n4783 VDD.n4686 4.5005
R7761 VDD.n4661 VDD.n4624 4.5005
R7762 VDD.n4667 VDD.n4616 4.5005
R7763 VDD.n4825 VDD.n4809 4.5005
R7764 VDD.n4849 VDD.n4844 4.5005
R7765 VDD.n4819 VDD.n4818 4.5005
R7766 VDD.n4793 VDD.n4792 4.5005
R7767 VDD.n3434 VDD.n3433 4.48249
R7768 VDD.n4012 VDD.n4011 4.36497
R7769 VDD.n8773 VDD.n8772 4.31361
R7770 VDD.n8765 VDD.n8764 4.31361
R7771 VDD.n8788 VDD.n8787 4.31361
R7772 VDD.n5228 VDD.n3812 4.31361
R7773 VDD.n3769 VDD.n3767 4.31361
R7774 VDD.n3766 VDD.n3763 4.31361
R7775 VDD.n4254 VDD.n4253 4.31361
R7776 VDD.n4246 VDD.n4245 4.31361
R7777 VDD.n4249 VDD.n4248 4.31361
R7778 VDD.n8871 VDD.n8819 4.31327
R7779 VDD.n4632 VDD.n4625 4.23768
R7780 VDD.n5164 VDD.n5157 4.23768
R7781 VDD.n4285 VDD.n4279 4.23768
R7782 VDD.n8890 VDD.n8883 4.23768
R7783 VDD.n5314 VDD.n5307 4.23684
R7784 VDD.n8618 VDD.n8611 4.23684
R7785 VDD.n8980 VDD.n8973 4.23684
R7786 VDD.n4059 VDD.n4058 4.18565
R7787 VDD.n4199 VDD.n4198 4.18565
R7788 VDD.n3409 VDD.n3406 4.17441
R7789 VDD.n1897 VDD.n1896 4.17441
R7790 VDD.n1043 VDD.n1042 4.17441
R7791 VDD.n188 VDD.n187 4.17441
R7792 VDD.n4671 VDD.n4670 4.14168
R7793 VDD.n5211 VDD.n5210 4.14168
R7794 VDD.n4398 VDD.n4395 4.14168
R7795 VDD.n4491 VDD.n4488 4.14168
R7796 VDD.n4561 VDD.n4558 4.14168
R7797 VDD.n4313 VDD.n4307 4.14168
R7798 VDD.n3700 VDD.n3697 4.14168
R7799 VDD.n3743 VDD.n3740 4.14168
R7800 VDD.n5342 VDD.n5336 4.14168
R7801 VDD.n5288 VDD.n5284 4.14168
R7802 VDD.n8473 VDD.t85 4.10046
R7803 VDD.n6501 VDD.n6499 4.05022
R7804 VDD.n3436 VDD.n3422 4.03708
R7805 VDD.n3436 VDD.n3423 4.03708
R7806 VDD.n7580 VDD.n7579 3.94428
R7807 VDD.n8039 VDD.n8036 3.92921
R7808 VDD.n3434 VDD.n3427 3.79052
R7809 VDD.t34 VDD.n3548 3.78536
R7810 VDD.n3000 VDD.n2997 3.78485
R7811 VDD.n2357 VDD.n2247 3.78485
R7812 VDD.n2254 VDD.n2253 3.78485
R7813 VDD.n2544 VDD.n1800 3.78485
R7814 VDD.n1503 VDD.n1393 3.78485
R7815 VDD.n1400 VDD.n1399 3.78485
R7816 VDD.n1690 VDD.n946 3.78485
R7817 VDD.n648 VDD.n538 3.78485
R7818 VDD.n545 VDD.n544 3.78485
R7819 VDD.n835 VDD.n91 3.78485
R7820 VDD.n4624 VDD.n4617 3.76521
R7821 VDD.n4619 VDD.n4618 3.76521
R7822 VDD.n4686 VDD.n4683 3.76521
R7823 VDD.n4818 VDD.n4816 3.76521
R7824 VDD.n4844 VDD.n4842 3.76521
R7825 VDD.n4874 VDD.n4872 3.76521
R7826 VDD.n4904 VDD.n4902 3.76521
R7827 VDD.n4934 VDD.n4932 3.76521
R7828 VDD.n3850 VDD.n3848 3.76521
R7829 VDD.n3815 VDD.n3813 3.76521
R7830 VDD.n5027 VDD.n5024 3.76521
R7831 VDD.n5200 VDD.n5193 3.76521
R7832 VDD.n5195 VDD.n5194 3.76521
R7833 VDD.n8646 VDD.n8645 3.76521
R7834 VDD.n3433 VDD.n3429 3.76521
R7835 VDD.n9009 VDD.n9008 3.76521
R7836 VDD.n8925 VDD.n8924 3.76521
R7837 VDD.n8054 VDD.n8053 3.73911
R7838 VDD.n4011 VDD.n3974 3.70369
R7839 VDD.n39 VDD.n38 3.67828
R7840 VDD.n901 VDD.n900 3.67828
R7841 VDD.n1748 VDD.n1747 3.67828
R7842 VDD.n2604 VDD.n2603 3.67828
R7843 VDD.n2714 VDD.n2707 3.64278
R7844 VDD.n2180 VDD.n2171 3.64278
R7845 VDD.n1326 VDD.n1317 3.64278
R7846 VDD.n471 VDD.n462 3.64278
R7847 VDD.n918 VDD.n911 3.43528
R7848 VDD.n2627 VDD.n2620 3.43528
R7849 VDD.n3653 VDD.n3646 3.42768
R7850 VDD.n5270 VDD.n5263 3.42768
R7851 VDD.n4711 VDD.n4704 3.42765
R7852 VDD.n5052 VDD.n5045 3.42765
R7853 VDD.n4514 VDD.n4507 3.42765
R7854 VDD.n4695 VDD.n4688 3.42683
R7855 VDD.n5036 VDD.n5029 3.42683
R7856 VDD.n4333 VDD.n4326 3.42683
R7857 VDD.n3165 VDD.n3162 3.42221
R7858 VDD.n1812 VDD.n1807 3.42221
R7859 VDD.n958 VDD.n953 3.42221
R7860 VDD.n103 VDD.n98 3.42221
R7861 VDD.n2771 VDD.n2768 3.39504
R7862 VDD.n2397 VDD.n2213 3.39504
R7863 VDD.n1543 VDD.n1359 3.39504
R7864 VDD.n688 VDD.n504 3.39504
R7865 VDD.n4616 VDD.n4615 3.38874
R7866 VDD.n4615 VDD.n4611 3.38874
R7867 VDD.n4792 VDD.n4791 3.38874
R7868 VDD.n4809 VDD.n4808 3.38874
R7869 VDD.n4841 VDD.n4840 3.38874
R7870 VDD.n4871 VDD.n4870 3.38874
R7871 VDD.n4901 VDD.n4900 3.38874
R7872 VDD.n4931 VDD.n4930 3.38874
R7873 VDD.n3835 VDD.n3834 3.38874
R7874 VDD.n5008 VDD.n5007 3.38874
R7875 VDD.n5133 VDD.n5132 3.38874
R7876 VDD.n5156 VDD.n5155 3.38874
R7877 VDD.n5155 VDD.n5151 3.38874
R7878 VDD.n4324 VDD.n4321 3.38874
R7879 VDD.n4409 VDD.n4406 3.38874
R7880 VDD.n4502 VDD.n4499 3.38874
R7881 VDD.n3644 VDD.n3641 3.38874
R7882 VDD.n5261 VDD.n5255 3.38874
R7883 VDD.n5299 VDD.n5295 3.38874
R7884 VDD.n3770 VDD.n3766 3.33963
R7885 VDD.n3770 VDD.n3769 3.33963
R7886 VDD.n5229 VDD.n5228 3.33963
R7887 VDD.n3755 VDD.n3753 3.33963
R7888 VDD.n5243 VDD.n5241 3.33963
R7889 VDD.n4073 VDD.n4072 3.33963
R7890 VDD.n3946 VDD.n3944 3.33963
R7891 VDD.n4246 VDD.n4244 3.33963
R7892 VDD.n4630 VDD.n4629 3.2936
R7893 VDD.n5162 VDD.n5161 3.2936
R7894 VDD.n4283 VDD.n4282 3.2936
R7895 VDD.n5312 VDD.n5311 3.2936
R7896 VDD.n8616 VDD.n8615 3.2936
R7897 VDD.n8978 VDD.n8977 3.2936
R7898 VDD.n8888 VDD.n8887 3.2936
R7899 VDD.n8857 VDD.n8855 3.25377
R7900 VDD.n50 VDD.n48 3.20702
R7901 VDD.n1759 VDD.n1757 3.20702
R7902 VDD VDD.n9031 3.20632
R7903 VDD.n4030 VDD.n4029 3.17466
R7904 VDD.n4058 VDD.n4057 3.17466
R7905 VDD.n2982 VDD.n2979 3.17267
R7906 VDD.n2988 VDD.n2985 3.17267
R7907 VDD.n2994 VDD.n2991 3.17267
R7908 VDD.n2370 VDD.n2230 3.17267
R7909 VDD.n2369 VDD.n2368 3.17267
R7910 VDD.n2367 VDD.n2235 3.17267
R7911 VDD.n1516 VDD.n1376 3.17267
R7912 VDD.n1515 VDD.n1514 3.17267
R7913 VDD.n1513 VDD.n1381 3.17267
R7914 VDD.n661 VDD.n521 3.17267
R7915 VDD.n660 VDD.n659 3.17267
R7916 VDD.n658 VDD.n526 3.17267
R7917 VDD.n3965 VDD.n3959 3.16717
R7918 VDD.n3536 VDD.n3533 3.10907
R7919 VDD.n3533 VDD.n3530 3.10907
R7920 VDD.n3530 VDD.n3527 3.10907
R7921 VDD.n3527 VDD.n3524 3.10907
R7922 VDD.n3524 VDD.n3521 3.10907
R7923 VDD.n3521 VDD.n3518 3.10907
R7924 VDD.n3518 VDD.n3515 3.10907
R7925 VDD.n3515 VDD.n3512 3.10907
R7926 VDD.n3512 VDD.n3509 3.10907
R7927 VDD.n3509 VDD.n3506 3.10907
R7928 VDD.n3506 VDD.n3503 3.10907
R7929 VDD.n3503 VDD.n3500 3.10907
R7930 VDD.n3500 VDD.n3497 3.10907
R7931 VDD.n3497 VDD.n3494 3.10907
R7932 VDD.n3494 VDD.n3491 3.10907
R7933 VDD.n3491 VDD.n3488 3.10907
R7934 VDD.n3488 VDD.n3485 3.10907
R7935 VDD.n3485 VDD.n3482 3.10907
R7936 VDD.n3482 VDD.n3479 3.10907
R7937 VDD.n3479 VDD.n3477 3.10907
R7938 VDD.n3477 VDD.n3475 3.10907
R7939 VDD.n3475 VDD.n3473 3.10907
R7940 VDD.n3473 VDD.n3471 3.10907
R7941 VDD.n3471 VDD.n3469 3.10907
R7942 VDD.n21 VDD.n20 3.10102
R7943 VDD.n876 VDD.n870 3.10102
R7944 VDD.n1730 VDD.n1729 3.10102
R7945 VDD.n2576 VDD.n2573 3.10102
R7946 VDD.n13 VDD.n5 3.09792
R7947 VDD.n891 VDD.n890 3.09792
R7948 VDD.n1722 VDD.n1714 3.09792
R7949 VDD.n2571 VDD.n2570 3.09792
R7950 VDD.n4319 VDD.n4318 3.03311
R7951 VDD.n4404 VDD.n4403 3.03311
R7952 VDD.n4497 VDD.n4496 3.03311
R7953 VDD.n4567 VDD.n4566 3.03311
R7954 VDD.n3749 VDD.n3748 3.03311
R7955 VDD.n3706 VDD.n3705 3.03311
R7956 VDD.n5348 VDD.n5347 3.03311
R7957 VDD.n8651 VDD.n8600 3.03311
R7958 VDD.n8730 VDD.n8729 3.03311
R7959 VDD.n8930 VDD.n8879 3.03311
R7960 VDD.n8699 VDD.n8678 3.03311
R7961 VDD.n8818 VDD.n8817 3.03311
R7962 VDD.n8814 VDD.n8813 3.03311
R7963 VDD.n8774 VDD.n8773 3.03311
R7964 VDD.n8766 VDD.n8765 3.03311
R7965 VDD.n8789 VDD.n8788 3.03311
R7966 VDD.n3947 VDD.n3946 3.03311
R7967 VDD.n5244 VDD.n5243 3.03311
R7968 VDD.n3759 VDD.n3758 3.03311
R7969 VDD.n5228 VDD.n5227 3.03311
R7970 VDD.n3756 VDD.n3755 3.03311
R7971 VDD.n4273 VDD.n4272 3.03311
R7972 VDD.n4267 VDD.n4266 3.03311
R7973 VDD.n4271 VDD.n4270 3.03311
R7974 VDD.n4255 VDD.n4254 3.03311
R7975 VDD.n3919 VDD.n3886 3.03311
R7976 VDD.n3769 VDD.n3768 3.03311
R7977 VDD.n4250 VDD.n4249 3.03311
R7978 VDD.n4074 VDD.n4073 3.03311
R7979 VDD.n3952 VDD.n3951 3.03311
R7980 VDD.n4247 VDD.n4246 3.03311
R7981 VDD.n3766 VDD.n3765 3.03311
R7982 VDD.n4616 VDD.n4609 3.01226
R7983 VDD.n4611 VDD.n4610 3.01226
R7984 VDD.n4792 VDD.n4789 3.01226
R7985 VDD.n4809 VDD.n4806 3.01226
R7986 VDD.n4841 VDD.n4838 3.01226
R7987 VDD.n4871 VDD.n4868 3.01226
R7988 VDD.n4901 VDD.n4898 3.01226
R7989 VDD.n4931 VDD.n4928 3.01226
R7990 VDD.n3840 VDD.n3839 3.01226
R7991 VDD.n3835 VDD.n3832 3.01226
R7992 VDD.n5014 VDD.n5013 3.01226
R7993 VDD.n5008 VDD.n5005 3.01226
R7994 VDD.n5133 VDD.n5130 3.01226
R7995 VDD.n5156 VDD.n5149 3.01226
R7996 VDD.n5151 VDD.n5150 3.01226
R7997 VDD.n5295 VDD.n5294 3.01226
R7998 VDD.n8666 VDD.n8665 3.01226
R7999 VDD.n8745 VDD.n8744 3.01226
R8000 VDD.n8945 VDD.n8944 3.01226
R8001 VDD.n3924 VDD.n3923 3.01226
R8002 VDD.n3886 VDD.n3885 3.01226
R8003 VDD.n4324 VDD.n4323 2.96007
R8004 VDD.n4409 VDD.n4408 2.96007
R8005 VDD.n4502 VDD.n4501 2.96007
R8006 VDD.n3644 VDD.n3643 2.96007
R8007 VDD.n4237 VDD.n4234 2.91015
R8008 VDD.n7563 VDD.n7559 2.88677
R8009 VDD.n3890 VDD.t143 2.77
R8010 VDD.n3890 VDD.t131 2.77
R8011 VDD.n8765 VDD.n8762 2.69036
R8012 VDD.n3340 VDD.n3338 2.64609
R8013 VDD.n1853 VDD.n1818 2.64609
R8014 VDD.n999 VDD.n964 2.64609
R8015 VDD.n144 VDD.n109 2.64609
R8016 VDD.n4105 VDD.n4104 2.64563
R8017 VDD.n4198 VDD.n4197 2.64563
R8018 VDD.n4624 VDD.n4623 2.63579
R8019 VDD.n4623 VDD.n4619 2.63579
R8020 VDD.n4686 VDD.n4685 2.63579
R8021 VDD.n4818 VDD.n4817 2.63579
R8022 VDD.n4844 VDD.n4843 2.63579
R8023 VDD.n4874 VDD.n4873 2.63579
R8024 VDD.n4904 VDD.n4903 2.63579
R8025 VDD.n4934 VDD.n4933 2.63579
R8026 VDD.n3850 VDD.n3849 2.63579
R8027 VDD.n3815 VDD.n3814 2.63579
R8028 VDD.n5027 VDD.n5026 2.63579
R8029 VDD.n5200 VDD.n5199 2.63579
R8030 VDD.n5199 VDD.n5195 2.63579
R8031 VDD.n5260 VDD.n5259 2.63579
R8032 VDD.n8667 VDD.n8664 2.63579
R8033 VDD.n8711 VDD.n8709 2.63579
R8034 VDD.n3429 VDD.n3428 2.63579
R8035 VDD.n8746 VDD.n8743 2.63579
R8036 VDD.n8946 VDD.n8943 2.63579
R8037 VDD.n3934 VDD.n3933 2.63579
R8038 VDD.n2777 VDD.n2774 2.56805
R8039 VDD.n2812 VDD.n2810 2.56805
R8040 VDD.n2817 VDD.n2812 2.56805
R8041 VDD.n2972 VDD.n2969 2.56805
R8042 VDD.n2969 VDD.n2966 2.56805
R8043 VDD.n2933 VDD.n2930 2.56805
R8044 VDD.n2395 VDD.n2394 2.56805
R8045 VDD.n2295 VDD.n2228 2.56805
R8046 VDD.n2296 VDD.n2295 2.56805
R8047 VDD.n2301 VDD.n2299 2.56805
R8048 VDD.n2303 VDD.n2301 2.56805
R8049 VDD.n2322 VDD.n2320 2.56805
R8050 VDD.n1541 VDD.n1540 2.56805
R8051 VDD.n1441 VDD.n1374 2.56805
R8052 VDD.n1442 VDD.n1441 2.56805
R8053 VDD.n1447 VDD.n1445 2.56805
R8054 VDD.n1449 VDD.n1447 2.56805
R8055 VDD.n1468 VDD.n1466 2.56805
R8056 VDD.n686 VDD.n685 2.56805
R8057 VDD.n586 VDD.n519 2.56805
R8058 VDD.n587 VDD.n586 2.56805
R8059 VDD.n592 VDD.n590 2.56805
R8060 VDD.n594 VDD.n592 2.56805
R8061 VDD.n613 VDD.n611 2.56805
R8062 VDD.n8701 VDD.n8700 2.56676
R8063 VDD.n3034 VDD.n3031 2.5605
R8064 VDD.n3028 VDD.n3025 2.5605
R8065 VDD.n1798 VDD.n1784 2.5605
R8066 VDD.n2545 VDD.n1799 2.5605
R8067 VDD.n944 VDD.n930 2.5605
R8068 VDD.n1691 VDD.n945 2.5605
R8069 VDD.n89 VDD.n75 2.5605
R8070 VDD.n836 VDD.n90 2.5605
R8071 VDD.n6465 VDD.n6461 2.53157
R8072 VDD.n6386 VDD.n6382 2.53157
R8073 VDD.n6300 VDD.n6296 2.53157
R8074 VDD.n6214 VDD.n6211 2.53157
R8075 VDD.n6144 VDD.n6141 2.53157
R8076 VDD.n6074 VDD.n6071 2.53157
R8077 VDD.n5991 VDD.n5987 2.53157
R8078 VDD.n5903 VDD.n5899 2.53157
R8079 VDD.n8089 VDD.n8084 2.4386
R8080 VDD.n8204 VDD.n8199 2.4386
R8081 VDD.n8309 VDD.n8304 2.4386
R8082 VDD.n8418 VDD.n8409 2.4386
R8083 VDD.n3374 VDD.n3372 2.43651
R8084 VDD.n1871 VDD.n1826 2.43651
R8085 VDD.n1017 VDD.n972 2.43651
R8086 VDD.n162 VDD.n117 2.43651
R8087 VDD.n7485 VDD.n7484 2.42576
R8088 VDD.n7416 VDD.n7415 2.42576
R8089 VDD.n7347 VDD.n7346 2.42576
R8090 VDD.n7262 VDD.n7261 2.42576
R8091 VDD.n7175 VDD.n7174 2.42576
R8092 VDD.n914 VDD.n913 2.42534
R8093 VDD.n2623 VDD.n2622 2.42534
R8094 VDD.n6465 VDD.n6464 2.38694
R8095 VDD.n6386 VDD.n6385 2.38694
R8096 VDD.n6300 VDD.n6299 2.38694
R8097 VDD.n6214 VDD.n6213 2.38694
R8098 VDD.n6144 VDD.n6143 2.38694
R8099 VDD.n6074 VDD.n6073 2.38694
R8100 VDD.n5991 VDD.n5990 2.38694
R8101 VDD.n5903 VDD.n5902 2.38694
R8102 VDD.n5845 VDD.n5844 2.38694
R8103 VDD.n3890 VDD.n3889 2.37942
R8104 VDD.n3436 VDD.n3435 2.3755
R8105 VDD.n8571 VDD.n8570 2.37087
R8106 VDD.n25 VDD.n17 2.30684
R8107 VDD.n875 VDD.n874 2.30684
R8108 VDD.n1734 VDD.n1726 2.30684
R8109 VDD.n7124 VDD.n7123 2.30315
R8110 VDD.n7029 VDD.n7025 2.30315
R8111 VDD.n7029 VDD.n7028 2.30315
R8112 VDD.n6941 VDD.n6937 2.30315
R8113 VDD.n6941 VDD.n6940 2.30315
R8114 VDD.n6853 VDD.n6849 2.30315
R8115 VDD.n6853 VDD.n6852 2.30315
R8116 VDD.n5517 VDD.n5513 2.30315
R8117 VDD.n5517 VDD.n5516 2.30315
R8118 VDD.n5605 VDD.n5601 2.30315
R8119 VDD.n5605 VDD.n5604 2.30315
R8120 VDD.n5693 VDD.n5689 2.30315
R8121 VDD.n5693 VDD.n5692 2.30315
R8122 VDD.n5781 VDD.n5777 2.30315
R8123 VDD.n5781 VDD.n5780 2.30315
R8124 VDD.n4670 VDD.n4669 2.25932
R8125 VDD.n5210 VDD.n5209 2.25932
R8126 VDD.n4391 VDD.n4390 2.25932
R8127 VDD.n4484 VDD.n4483 2.25932
R8128 VDD.n4554 VDD.n4553 2.25932
R8129 VDD.n4303 VDD.n4302 2.25932
R8130 VDD.n3693 VDD.n3692 2.25932
R8131 VDD.n3736 VDD.n3735 2.25932
R8132 VDD.n5332 VDD.n5331 2.25932
R8133 VDD.n5284 VDD.n5283 2.25932
R8134 VDD.n8647 VDD.n8644 2.25932
R8135 VDD.n8602 VDD.n8601 2.25932
R8136 VDD.n8695 VDD.n8693 2.25932
R8137 VDD.n8680 VDD.n8679 2.25932
R8138 VDD.n9010 VDD.n9007 2.25932
R8139 VDD.n8964 VDD.n8963 2.25932
R8140 VDD.n8926 VDD.n8923 2.25932
R8141 VDD.n8881 VDD.n8880 2.25932
R8142 VDD.n3888 VDD.n3887 2.25932
R8143 VDD.n8695 VDD.n8694 2.25379
R8144 VDD.n5019 VDD.n3820 2.25051
R8145 VDD.n25 VDD.n24 2.2505
R8146 VDD.n26 VDD.n12 2.2505
R8147 VDD.n28 VDD.n27 2.2505
R8148 VDD.n15 VDD.n4 2.2505
R8149 VDD.n63 VDD.n62 2.2505
R8150 VDD.n874 VDD.n873 2.2505
R8151 VDD.n867 VDD.n866 2.2505
R8152 VDD.n885 VDD.n884 2.2505
R8153 VDD.n888 VDD.n887 2.2505
R8154 VDD.n886 VDD.n864 2.2505
R8155 VDD.n1734 VDD.n1733 2.2505
R8156 VDD.n1735 VDD.n1721 2.2505
R8157 VDD.n1737 VDD.n1736 2.2505
R8158 VDD.n1724 VDD.n1713 2.2505
R8159 VDD.n1772 VDD.n1771 2.2505
R8160 VDD.n2600 VDD.n2599 2.2505
R8161 VDD.n5019 VDD.n5018 2.24905
R8162 VDD.n6469 VDD.n6468 2.24231
R8163 VDD.n6390 VDD.n6389 2.24231
R8164 VDD.n6305 VDD.n6304 2.24231
R8165 VDD.n6218 VDD.n6217 2.24231
R8166 VDD.n6148 VDD.n6147 2.24231
R8167 VDD.n6078 VDD.n6077 2.24231
R8168 VDD.n5996 VDD.n5995 2.24231
R8169 VDD.n5908 VDD.n5907 2.24231
R8170 VDD.n5019 VDD.n5003 2.23886
R8171 VDD.n5019 VDD.n5011 2.23886
R8172 VDD.n8073 VDD.n8072 2.23542
R8173 VDD.n8190 VDD.n8189 2.23542
R8174 VDD.n8295 VDD.n8294 2.23542
R8175 VDD.n8400 VDD.n8399 2.23542
R8176 VDD.n4398 VDD.n4397 2.22452
R8177 VDD.n4491 VDD.n4490 2.22452
R8178 VDD.n4561 VDD.n4560 2.22452
R8179 VDD.n3700 VDD.n3699 2.22452
R8180 VDD.n3743 VDD.n3742 2.22452
R8181 VDD.n7976 VDD.n7975 2.21832
R8182 VDD.n7957 VDD.n7950 2.21832
R8183 VDD.n7834 VDD.n7833 2.21832
R8184 VDD.n7818 VDD.n7813 2.21832
R8185 VDD.n7702 VDD.n7701 2.21832
R8186 VDD.n7683 VDD.n7676 2.21832
R8187 VDD.n916 VDD.n915 2.19693
R8188 VDD.n2625 VDD.n2624 2.19693
R8189 VDD.n8848 VDD.n8847 2.18378
R8190 VDD.n8081 VDD.n8077 2.1677
R8191 VDD.n8196 VDD.n8193 2.1677
R8192 VDD.n8301 VDD.n8298 2.1677
R8193 VDD.n8406 VDD.n8403 2.1677
R8194 VDD.n7485 VDD.n7482 2.15629
R8195 VDD.n7479 VDD.n7478 2.15629
R8196 VDD.n7416 VDD.n7413 2.15629
R8197 VDD.n7410 VDD.n7409 2.15629
R8198 VDD.n7347 VDD.n7344 2.15629
R8199 VDD.n7341 VDD.n7340 2.15629
R8200 VDD.n7262 VDD.n7258 2.15629
R8201 VDD.n7254 VDD.n7253 2.15629
R8202 VDD.n7175 VDD.n7171 2.15629
R8203 VDD.n7167 VDD.n7166 2.15629
R8204 VDD.n4036 VDD.t142 2.11661
R8205 VDD.n4176 VDD.t80 2.11661
R8206 VDD.n4320 VDD.n4278 2.10401
R8207 VDD.n6707 VDD.t33 2.1032
R8208 VDD.n6458 VDD.n6457 2.09768
R8209 VDD.n6379 VDD.n6378 2.09768
R8210 VDD.n6292 VDD.n6291 2.09768
R8211 VDD.n6208 VDD.n6207 2.09768
R8212 VDD.n6138 VDD.n6137 2.09768
R8213 VDD.n6068 VDD.n6067 2.09768
R8214 VDD.n5983 VDD.n5982 2.09768
R8215 VDD.n5895 VDD.n5894 2.09768
R8216 VDD.n3540 VDD.n3536 2.07664
R8217 VDD.n48 VDD.n44 2.0723
R8218 VDD.n1757 VDD.n1753 2.0723
R8219 VDD.n7109 VDD.n7108 2.03225
R8220 VDD.n7034 VDD.n7033 2.03225
R8221 VDD.n7021 VDD.n7020 2.03225
R8222 VDD.n6946 VDD.n6945 2.03225
R8223 VDD.n6933 VDD.n6932 2.03225
R8224 VDD.n6858 VDD.n6857 2.03225
R8225 VDD.n6845 VDD.n6844 2.03225
R8226 VDD.n5509 VDD.n5508 2.03225
R8227 VDD.n5522 VDD.n5521 2.03225
R8228 VDD.n5597 VDD.n5596 2.03225
R8229 VDD.n5610 VDD.n5609 2.03225
R8230 VDD.n5685 VDD.n5684 2.03225
R8231 VDD.n5698 VDD.n5697 2.03225
R8232 VDD.n5773 VDD.n5772 2.03225
R8233 VDD.n5786 VDD.n5785 2.03225
R8234 VDD.n3004 VDD.n3001 2.00398
R8235 VDD.n3008 VDD.n3007 2.00398
R8236 VDD.n3406 VDD.n3403 2.00398
R8237 VDD.n2356 VDD.n2355 2.00398
R8238 VDD.n2354 VDD.n2249 2.00398
R8239 VDD.n1896 VDD.n1895 2.00398
R8240 VDD.n1502 VDD.n1501 2.00398
R8241 VDD.n1500 VDD.n1395 2.00398
R8242 VDD.n1042 VDD.n1041 2.00398
R8243 VDD.n647 VDD.n646 2.00398
R8244 VDD.n645 VDD.n540 2.00398
R8245 VDD.n187 VDD.n186 2.00398
R8246 VDD.n4016 VDD.n4015 1.98435
R8247 VDD.n3109 VDD.n3108 1.97774
R8248 VDD.n2117 VDD.n2066 1.97774
R8249 VDD.n1263 VDD.n1212 1.97774
R8250 VDD.n408 VDD.n357 1.97774
R8251 VDD.n7965 VDD.n7961 1.96486
R8252 VDD.n7965 VDD.n7964 1.96486
R8253 VDD.n7824 VDD.n7821 1.96486
R8254 VDD.n7824 VDD.n7823 1.96486
R8255 VDD.n7691 VDD.n7687 1.96486
R8256 VDD.n7691 VDD.n7690 1.96486
R8257 VDD.n8081 VDD.n8080 1.96452
R8258 VDD.n8196 VDD.n8195 1.96452
R8259 VDD.n8301 VDD.n8300 1.96452
R8260 VDD.n8406 VDD.n8405 1.96452
R8261 VDD.n2779 VDD.n2777 1.96392
R8262 VDD.n2785 VDD.n2782 1.96392
R8263 VDD.n2790 VDD.n2788 1.96392
R8264 VDD.n2796 VDD.n2793 1.96392
R8265 VDD.n2801 VDD.n2799 1.96392
R8266 VDD.n2808 VDD.n2804 1.96392
R8267 VDD.n2394 VDD.n2392 1.96392
R8268 VDD.n2225 VDD.n2216 1.96392
R8269 VDD.n2386 VDD.n2227 1.96392
R8270 VDD.n2385 VDD.n2383 1.96392
R8271 VDD.n2382 VDD.n2380 1.96392
R8272 VDD.n2378 VDD.n2376 1.96392
R8273 VDD.n1540 VDD.n1538 1.96392
R8274 VDD.n1371 VDD.n1362 1.96392
R8275 VDD.n1532 VDD.n1373 1.96392
R8276 VDD.n1531 VDD.n1529 1.96392
R8277 VDD.n1528 VDD.n1526 1.96392
R8278 VDD.n1524 VDD.n1522 1.96392
R8279 VDD.n685 VDD.n683 1.96392
R8280 VDD.n516 VDD.n507 1.96392
R8281 VDD.n677 VDD.n518 1.96392
R8282 VDD.n676 VDD.n674 1.96392
R8283 VDD.n673 VDD.n671 1.96392
R8284 VDD.n669 VDD.n667 1.96392
R8285 VDD.n6474 VDD.n6473 1.95304
R8286 VDD.n6395 VDD.n6394 1.95304
R8287 VDD.n6310 VDD.n6309 1.95304
R8288 VDD.n6222 VDD.n6221 1.95304
R8289 VDD.n6152 VDD.n6151 1.95304
R8290 VDD.n6082 VDD.n6081 1.95304
R8291 VDD.n6001 VDD.n6000 1.95304
R8292 VDD.n5913 VDD.n5912 1.95304
R8293 VDD.n3335 VDD.n3309 1.94579
R8294 VDD.n1940 VDD.n1939 1.94579
R8295 VDD.n1086 VDD.n1085 1.94579
R8296 VDD.n231 VDD.n230 1.94579
R8297 VDD.n3620 VDD.n3601 1.90031
R8298 VDD.n8056 VDD.n8054 1.8968
R8299 VDD.n8073 VDD.n8070 1.8968
R8300 VDD.n8190 VDD.n8187 1.8968
R8301 VDD.n8295 VDD.n8292 1.8968
R8302 VDD.n8400 VDD.n8397 1.8968
R8303 VDD.n2928 VDD.n2913 1.88841
R8304 VDD.n2403 VDD.n2002 1.88841
R8305 VDD.n1549 VDD.n1148 1.88841
R8306 VDD.n694 VDD.n293 1.88841
R8307 VDD.n7475 VDD.n7474 1.88682
R8308 VDD.n7420 VDD.n7419 1.88682
R8309 VDD.n7406 VDD.n7405 1.88682
R8310 VDD.n7351 VDD.n7350 1.88682
R8311 VDD.n7336 VDD.n7335 1.88682
R8312 VDD.n7267 VDD.n7266 1.88682
R8313 VDD.n7249 VDD.n7248 1.88682
R8314 VDD.n7180 VDD.n7179 1.88682
R8315 VDD.n7162 VDD.n7161 1.88682
R8316 VDD.n4653 VDD.n4649 1.88285
R8317 VDD.n5185 VDD.n5181 1.88285
R8318 VDD.n4312 VDD.n4311 1.88285
R8319 VDD.n5341 VDD.n5340 1.88285
R8320 VDD.n7495 VDD.n7494 1.88285
R8321 VDD.n8711 VDD.n8710 1.87949
R8322 VDD.n8572 VDD.n8568 1.85282
R8323 VDD.n8057 VDD.n8056 1.82907
R8324 VDD.n4811 VDD.n4810 1.81303
R8325 VDD.n5137 VDD.n5136 1.81303
R8326 VDD.n6454 VDD.n6453 1.80841
R8327 VDD.n6375 VDD.n6374 1.80841
R8328 VDD.n6287 VDD.n6286 1.80841
R8329 VDD.n6204 VDD.n6203 1.80841
R8330 VDD.n6134 VDD.n6133 1.80841
R8331 VDD.n6064 VDD.n6063 1.80841
R8332 VDD.n5978 VDD.n5977 1.80841
R8333 VDD.n5890 VDD.n5889 1.80841
R8334 VDD.n3001 VDD.n3000 1.78137
R8335 VDD.n3403 VDD.n3402 1.78137
R8336 VDD.n2357 VDD.n2356 1.78137
R8337 VDD.n1895 VDD.n1800 1.78137
R8338 VDD.n1503 VDD.n1502 1.78137
R8339 VDD.n1041 VDD.n946 1.78137
R8340 VDD.n648 VDD.n647 1.78137
R8341 VDD.n186 VDD.n91 1.78137
R8342 VDD.n7104 VDD.n7103 1.76135
R8343 VDD.n7039 VDD.n7038 1.76135
R8344 VDD.n7016 VDD.n7015 1.76135
R8345 VDD.n6951 VDD.n6950 1.76135
R8346 VDD.n6928 VDD.n6927 1.76135
R8347 VDD.n6863 VDD.n6862 1.76135
R8348 VDD.n6840 VDD.n6839 1.76135
R8349 VDD.n5504 VDD.n5503 1.76135
R8350 VDD.n5527 VDD.n5526 1.76135
R8351 VDD.n5592 VDD.n5591 1.76135
R8352 VDD.n5615 VDD.n5614 1.76135
R8353 VDD.n5680 VDD.n5679 1.76135
R8354 VDD.n5703 VDD.n5702 1.76135
R8355 VDD.n5768 VDD.n5767 1.76135
R8356 VDD.n5791 VDD.n5790 1.76135
R8357 VDD.n3111 VDD.n3109 1.74595
R8358 VDD.n2117 VDD.n2116 1.74595
R8359 VDD.n1263 VDD.n1262 1.74595
R8360 VDD.n408 VDD.n407 1.74595
R8361 VDD.t12 VDD.n4121 1.71984
R8362 VDD.n3369 VDD.n3365 1.71235
R8363 VDD.n3362 VDD.n3360 1.71235
R8364 VDD.n3358 VDD.n3355 1.71235
R8365 VDD.n3352 VDD.n3350 1.71235
R8366 VDD.n3348 VDD.n3345 1.71235
R8367 VDD.n3342 VDD.n3340 1.71235
R8368 VDD.n1870 VDD.n1869 1.71235
R8369 VDD.n1868 VDD.n1842 1.71235
R8370 VDD.n1865 VDD.n1864 1.71235
R8371 VDD.n1860 VDD.n1845 1.71235
R8372 VDD.n1859 VDD.n1855 1.71235
R8373 VDD.n1854 VDD.n1853 1.71235
R8374 VDD.n1016 VDD.n1015 1.71235
R8375 VDD.n1014 VDD.n988 1.71235
R8376 VDD.n1011 VDD.n1010 1.71235
R8377 VDD.n1006 VDD.n991 1.71235
R8378 VDD.n1005 VDD.n1001 1.71235
R8379 VDD.n1000 VDD.n999 1.71235
R8380 VDD.n161 VDD.n160 1.71235
R8381 VDD.n159 VDD.n133 1.71235
R8382 VDD.n156 VDD.n155 1.71235
R8383 VDD.n151 VDD.n136 1.71235
R8384 VDD.n150 VDD.n146 1.71235
R8385 VDD.n145 VDD.n144 1.71235
R8386 VDD.n7976 VDD.n7972 1.71139
R8387 VDD.n7957 VDD.n7956 1.71139
R8388 VDD.n7834 VDD.n7831 1.71139
R8389 VDD.n7818 VDD.n7817 1.71139
R8390 VDD.n7702 VDD.n7698 1.71139
R8391 VDD.n7683 VDD.n7682 1.71139
R8392 VDD.n5415 VDD.n5414 1.70907
R8393 VDD.n5411 VDD.n5410 1.70593
R8394 VDD.n5430 VDD.n5429 1.70592
R8395 VDD.n5417 VDD.n5373 1.70592
R8396 VDD.n5391 VDD.n5390 1.70592
R8397 VDD.n5432 VDD.n3631 1.70583
R8398 VDD.n5419 VDD.n3638 1.70583
R8399 VDD.n5401 VDD.n5400 1.70582
R8400 VDD.n5422 VDD.n3634 1.70582
R8401 VDD.n65 VDD.n3 1.7055
R8402 VDD.n920 VDD.n919 1.7055
R8403 VDD.n1774 VDD.n1712 1.7055
R8404 VDD.n2629 VDD.n2628 1.7055
R8405 VDD.n4595 VDD.n4590 1.70404
R8406 VDD.n4606 VDD.n4605 1.70006
R8407 VDD.n8089 VDD.n8088 1.69362
R8408 VDD.n8204 VDD.n8203 1.69362
R8409 VDD.n8309 VDD.n8308 1.69362
R8410 VDD.n8418 VDD.n8417 1.69362
R8411 VDD.t43 VDD.t68 1.68266
R8412 VDD.n3410 VDD.n3409 1.67007
R8413 VDD.n1898 VDD.n1897 1.67007
R8414 VDD.n1044 VDD.n1043 1.67007
R8415 VDD.n189 VDD.n188 1.67007
R8416 VDD.n6478 VDD.n6477 1.66378
R8417 VDD.n6399 VDD.n6398 1.66378
R8418 VDD.n6315 VDD.n6314 1.66378
R8419 VDD.n6227 VDD.n6226 1.66378
R8420 VDD.n6156 VDD.n6155 1.66378
R8421 VDD.n6086 VDD.n6085 1.66378
R8422 VDD.n6006 VDD.n6005 1.66378
R8423 VDD.n5918 VDD.n5917 1.66378
R8424 VDD.n2963 VDD.n2960 1.66186
R8425 VDD.n2957 VDD.n2955 1.66186
R8426 VDD.n2952 VDD.n2949 1.66186
R8427 VDD.n2946 VDD.n2944 1.66186
R8428 VDD.n2941 VDD.n2938 1.66186
R8429 VDD.n2935 VDD.n2933 1.66186
R8430 VDD.n2307 VDD.n2305 1.66186
R8431 VDD.n2308 VDD.n2291 1.66186
R8432 VDD.n2313 VDD.n2311 1.66186
R8433 VDD.n2314 VDD.n2289 1.66186
R8434 VDD.n2319 VDD.n2317 1.66186
R8435 VDD.n2323 VDD.n2322 1.66186
R8436 VDD.n1453 VDD.n1451 1.66186
R8437 VDD.n1454 VDD.n1437 1.66186
R8438 VDD.n1459 VDD.n1457 1.66186
R8439 VDD.n1460 VDD.n1435 1.66186
R8440 VDD.n1465 VDD.n1463 1.66186
R8441 VDD.n1469 VDD.n1468 1.66186
R8442 VDD.n598 VDD.n596 1.66186
R8443 VDD.n599 VDD.n582 1.66186
R8444 VDD.n604 VDD.n602 1.66186
R8445 VDD.n605 VDD.n580 1.66186
R8446 VDD.n610 VDD.n608 1.66186
R8447 VDD.n614 VDD.n613 1.66186
R8448 VDD.n4474 VDD.n4473 1.64452
R8449 VDD.n4544 VDD.n4543 1.64452
R8450 VDD.n4381 VDD.n4380 1.64447
R8451 VDD.n3683 VDD.n3682 1.64446
R8452 VDD.n3726 VDD.n3725 1.64446
R8453 VDD.n7501 VDD.n7500 1.63187
R8454 VDD.n8065 VDD.n8064 1.6259
R8455 VDD.n8182 VDD.n8181 1.6259
R8456 VDD.n8287 VDD.n8286 1.6259
R8457 VDD.n8392 VDD.n8391 1.6259
R8458 VDD.n8542 VDD.n8541 1.6259
R8459 VDD.n3629 VDD.n3436 1.62066
R8460 VDD.n7471 VDD.n7470 1.61734
R8461 VDD.n7424 VDD.n7423 1.61734
R8462 VDD.n7402 VDD.n7401 1.61734
R8463 VDD.n7355 VDD.n7354 1.61734
R8464 VDD.n7331 VDD.n7330 1.61734
R8465 VDD.n7272 VDD.n7271 1.61734
R8466 VDD.n7244 VDD.n7243 1.61734
R8467 VDD.n7185 VDD.n7184 1.61734
R8468 VDD.n7157 VDD.n7156 1.61734
R8469 VDD.n3619 VDD.n3616 1.61534
R8470 VDD.n3616 VDD.n3613 1.61534
R8471 VDD.n3613 VDD.n3610 1.61534
R8472 VDD.n3610 VDD.n3607 1.61534
R8473 VDD.n3607 VDD.n3604 1.61534
R8474 VDD.n3559 VDD.n3556 1.61534
R8475 VDD.n3562 VDD.n3559 1.61534
R8476 VDD.n3565 VDD.n3562 1.61534
R8477 VDD.n3568 VDD.n3565 1.61534
R8478 VDD.n3571 VDD.n3568 1.61534
R8479 VDD.n3575 VDD.n3571 1.61534
R8480 VDD.n3595 VDD.n3592 1.61534
R8481 VDD.n3592 VDD.n3589 1.61534
R8482 VDD.n3589 VDD.n3586 1.61534
R8483 VDD.n3586 VDD.n3583 1.61534
R8484 VDD.n3583 VDD.n3580 1.61534
R8485 VDD.n3580 VDD.n3577 1.61534
R8486 VDD.n3442 VDD.n3439 1.61534
R8487 VDD.n3445 VDD.n3442 1.61534
R8488 VDD.n3448 VDD.n3445 1.61534
R8489 VDD.n3451 VDD.n3448 1.61534
R8490 VDD.n3454 VDD.n3451 1.61534
R8491 VDD.n3012 VDD.n3011 1.61441
R8492 VDD.n2254 VDD.n2252 1.61441
R8493 VDD.n1400 VDD.n1398 1.61441
R8494 VDD.n545 VDD.n543 1.61441
R8495 VDD.n8525 VDD.t45 1.58758
R8496 VDD.n6793 VDD.n6792 1.58445
R8497 VDD.n6705 VDD.n6704 1.58445
R8498 VDD.n6613 VDD.n6612 1.58445
R8499 VDD.n6525 VDD.n6524 1.58445
R8500 VDD.n3965 VDD.n3964 1.58383
R8501 VDD.n8870 VDD.n8867 1.57731
R8502 VDD.n7124 VDD.n7120 1.55817
R8503 VDD.n8574 VDD.n8573 1.5505
R8504 VDD.n6449 VDD.n6448 1.51914
R8505 VDD.n6370 VDD.n6369 1.51914
R8506 VDD.n6282 VDD.n6281 1.51914
R8507 VDD.n6200 VDD.n6199 1.51914
R8508 VDD.n6130 VDD.n6129 1.51914
R8509 VDD.n6060 VDD.n6059 1.51914
R8510 VDD.n5973 VDD.n5972 1.51914
R8511 VDD.n5885 VDD.n5884 1.51914
R8512 VDD.n8610 VDD.n8607 1.50638
R8513 VDD.n8686 VDD.n8685 1.50638
R8514 VDD.n8972 VDD.n8969 1.50638
R8515 VDD.n8913 VDD.n8910 1.50638
R8516 VDD.n3880 VDD.n3879 1.50638
R8517 VDD.n3906 VDD.n3904 1.50638
R8518 VDD.n8683 VDD.n8682 1.50148
R8519 VDD.n3939 VDD.n3938 1.5005
R8520 VDD.n7099 VDD.n7098 1.49045
R8521 VDD.n7044 VDD.n7043 1.49045
R8522 VDD.n7011 VDD.n7010 1.49045
R8523 VDD.n6956 VDD.n6955 1.49045
R8524 VDD.n6923 VDD.n6922 1.49045
R8525 VDD.n6868 VDD.n6867 1.49045
R8526 VDD.n6835 VDD.n6834 1.49045
R8527 VDD.n5499 VDD.n5498 1.49045
R8528 VDD.n5532 VDD.n5531 1.49045
R8529 VDD.n5587 VDD.n5586 1.49045
R8530 VDD.n5620 VDD.n5619 1.49045
R8531 VDD.n5675 VDD.n5674 1.49045
R8532 VDD.n5708 VDD.n5707 1.49045
R8533 VDD.n5763 VDD.n5762 1.49045
R8534 VDD.n5796 VDD.n5795 1.49045
R8535 VDD.n4385 VDD.n4384 1.4871
R8536 VDD.n4478 VDD.n4477 1.4871
R8537 VDD.n4548 VDD.n4547 1.4871
R8538 VDD.n3687 VDD.n3686 1.4871
R8539 VDD.n3730 VDD.n3729 1.4871
R8540 VDD.n5218 VDD.n5217 1.48392
R8541 VDD.n5144 VDD.n5143 1.48392
R8542 VDD.n4923 VDD.n4922 1.48392
R8543 VDD.n4893 VDD.n4892 1.48392
R8544 VDD.n4833 VDD.n4832 1.48392
R8545 VDD.n4801 VDD.n4800 1.48392
R8546 VDD.n4678 VDD.n4677 1.48392
R8547 VDD.n4863 VDD.n4862 1.48392
R8548 VDD.n4953 VDD.n4952 1.48392
R8549 VDD.n3853 VDD.n3852 1.47597
R8550 VDD.n3820 VDD.n3819 1.47597
R8551 VDD.n4814 VDD.n4813 1.46766
R8552 VDD.n4847 VDD.n4846 1.46766
R8553 VDD.n4937 VDD.n4936 1.46766
R8554 VDD.n4877 VDD.n4876 1.46766
R8555 VDD.n4907 VDD.n4906 1.46766
R8556 VDD.n3171 VDD.n3168 1.45846
R8557 VDD.n3208 VDD.n3205 1.45846
R8558 VDD.n3211 VDD.n3208 1.45846
R8559 VDD.n2536 VDD.n1808 1.45846
R8560 VDD.n1905 VDD.n1840 1.45846
R8561 VDD.n1900 VDD.n1840 1.45846
R8562 VDD.n1682 VDD.n954 1.45846
R8563 VDD.n1051 VDD.n986 1.45846
R8564 VDD.n1046 VDD.n986 1.45846
R8565 VDD.n827 VDD.n99 1.45846
R8566 VDD.n196 VDD.n131 1.45846
R8567 VDD.n191 VDD.n131 1.45846
R8568 VDD.n7984 VDD.n7983 1.45793
R8569 VDD.n7946 VDD.n7945 1.45793
R8570 VDD.n7842 VDD.n7841 1.45793
R8571 VDD.n7810 VDD.n7809 1.45793
R8572 VDD.n7710 VDD.n7709 1.45793
R8573 VDD.n7672 VDD.n7671 1.45793
R8574 VDD.n3542 VDD.n3541 1.45532
R8575 VDD.n8097 VDD.n8096 1.42272
R8576 VDD.n8210 VDD.n8209 1.42272
R8577 VDD.n8315 VDD.n8314 1.42272
R8578 VDD.n8428 VDD.n8427 1.42272
R8579 VDD.n6785 VDD.n6784 1.41321
R8580 VDD.n6697 VDD.n6696 1.41321
R8581 VDD.n6605 VDD.n6604 1.41321
R8582 VDD.n6519 VDD.n6518 1.41321
R8583 VDD.n8859 VDD.n8850 1.41321
R8584 VDD.n8807 VDD.n8805 1.3918
R8585 VDD.n7563 VDD.n7562 1.38089
R8586 VDD.n7505 VDD.n7504 1.38089
R8587 VDD.n6483 VDD.n6482 1.37451
R8588 VDD.n6404 VDD.n6403 1.37451
R8589 VDD.n6320 VDD.n6319 1.37451
R8590 VDD.n6232 VDD.n6231 1.37451
R8591 VDD.n6160 VDD.n6159 1.37451
R8592 VDD.n6090 VDD.n6089 1.37451
R8593 VDD.n6011 VDD.n6010 1.37451
R8594 VDD.n5923 VDD.n5922 1.37451
R8595 VDD.n8176 VDD.n8175 1.355
R8596 VDD.n8281 VDD.n8280 1.355
R8597 VDD.n8386 VDD.n8385 1.355
R8598 VDD.n8536 VDD.n8535 1.355
R8599 VDD.n3385 VDD.n3382 1.35125
R8600 VDD.n1934 VDD.n1825 1.35125
R8601 VDD.n1080 VDD.n971 1.35125
R8602 VDD.n225 VDD.n116 1.35125
R8603 VDD.n7467 VDD.n7466 1.34787
R8604 VDD.n7428 VDD.n7427 1.34787
R8605 VDD.n7398 VDD.n7397 1.34787
R8606 VDD.n7359 VDD.n7358 1.34787
R8607 VDD.n7326 VDD.n7325 1.34787
R8608 VDD.n7277 VDD.n7276 1.34787
R8609 VDD.n7239 VDD.n7238 1.34787
R8610 VDD.n7190 VDD.n7189 1.34787
R8611 VDD.n7152 VDD.n7151 1.34787
R8612 VDD.n4971 VDD.n3845 1.34458
R8613 VDD.n4971 VDD.n3857 1.34227
R8614 VDD.n3038 VDD.n3037 1.33615
R8615 VDD.n2556 VDD.n2555 1.33615
R8616 VDD.n1702 VDD.n1701 1.33615
R8617 VDD.n847 VDD.n846 1.33615
R8618 VDD.n6793 VDD.n6789 1.32759
R8619 VDD.n6705 VDD.n6701 1.32759
R8620 VDD.n6613 VDD.n6609 1.32759
R8621 VDD.n6525 VDD.n6522 1.32759
R8622 VDD.n2774 VDD.n2772 1.32203
R8623 VDD.n2973 VDD.n2972 1.32203
R8624 VDD.n2396 VDD.n2395 1.32203
R8625 VDD.n2299 VDD.n2293 1.32203
R8626 VDD.n1542 VDD.n1541 1.32203
R8627 VDD.n1445 VDD.n1439 1.32203
R8628 VDD.n687 VDD.n686 1.32203
R8629 VDD.n590 VDD.n584 1.32203
R8630 VDD.n3620 VDD.n3619 1.28287
R8631 VDD.n3893 VDD.n3892 1.26837
R8632 VDD.n2717 VDD.n2714 1.25267
R8633 VDD.n2180 VDD.n2179 1.25267
R8634 VDD.n1326 VDD.n1325 1.25267
R8635 VDD.n471 VDD.n470 1.25267
R8636 VDD.n2772 VDD.n2771 1.24652
R8637 VDD.n2973 VDD.n2817 1.24652
R8638 VDD.n2397 VDD.n2396 1.24652
R8639 VDD.n2296 VDD.n2293 1.24652
R8640 VDD.n1543 VDD.n1542 1.24652
R8641 VDD.n1442 VDD.n1439 1.24652
R8642 VDD.n688 VDD.n687 1.24652
R8643 VDD.n587 VDD.n584 1.24652
R8644 VDD.n6780 VDD.n6779 1.24197
R8645 VDD.n6693 VDD.n6692 1.24197
R8646 VDD.n6600 VDD.n6599 1.24197
R8647 VDD.n6515 VDD.n6514 1.24197
R8648 VDD.n6445 VDD.n6444 1.22988
R8649 VDD.n6365 VDD.n6364 1.22988
R8650 VDD.n6277 VDD.n6276 1.22988
R8651 VDD.n6196 VDD.n6195 1.22988
R8652 VDD.n6126 VDD.n6125 1.22988
R8653 VDD.n6056 VDD.n6055 1.22988
R8654 VDD.n5968 VDD.n5967 1.22988
R8655 VDD.n5880 VDD.n5879 1.22988
R8656 VDD.n3019 VDD.n3016 1.22485
R8657 VDD.n3038 VDD.n3019 1.22485
R8658 VDD.n3037 VDD.n3034 1.22485
R8659 VDD.n3031 VDD.n3028 1.22485
R8660 VDD.n3025 VDD.n3022 1.22485
R8661 VDD.n2253 VDD.n1783 1.22485
R8662 VDD.n2556 VDD.n1783 1.22485
R8663 VDD.n2555 VDD.n1784 1.22485
R8664 VDD.n1799 VDD.n1798 1.22485
R8665 VDD.n2545 VDD.n2544 1.22485
R8666 VDD.n1399 VDD.n929 1.22485
R8667 VDD.n1702 VDD.n929 1.22485
R8668 VDD.n1701 VDD.n930 1.22485
R8669 VDD.n945 VDD.n944 1.22485
R8670 VDD.n1691 VDD.n1690 1.22485
R8671 VDD.n544 VDD.n74 1.22485
R8672 VDD.n847 VDD.n74 1.22485
R8673 VDD.n846 VDD.n75 1.22485
R8674 VDD.n90 VDD.n89 1.22485
R8675 VDD.n836 VDD.n835 1.22485
R8676 VDD.n7094 VDD.n7093 1.21955
R8677 VDD.n7049 VDD.n7048 1.21955
R8678 VDD.n7006 VDD.n7005 1.21955
R8679 VDD.n6961 VDD.n6960 1.21955
R8680 VDD.n6918 VDD.n6917 1.21955
R8681 VDD.n6873 VDD.n6872 1.21955
R8682 VDD.n6830 VDD.n6829 1.21955
R8683 VDD.n5494 VDD.n5493 1.21955
R8684 VDD.n5537 VDD.n5536 1.21955
R8685 VDD.n5582 VDD.n5581 1.21955
R8686 VDD.n5625 VDD.n5624 1.21955
R8687 VDD.n5670 VDD.n5669 1.21955
R8688 VDD.n5713 VDD.n5712 1.21955
R8689 VDD.n5758 VDD.n5757 1.21955
R8690 VDD.n5801 VDD.n5800 1.21955
R8691 VDD.n7992 VDD.n7991 1.20446
R8692 VDD.n7938 VDD.n7937 1.20446
R8693 VDD.n7850 VDD.n7849 1.20446
R8694 VDD.n7804 VDD.n7803 1.20446
R8695 VDD.n7718 VDD.n7717 1.20446
R8696 VDD.n7664 VDD.n7663 1.20446
R8697 VDD.n886 VDD.n857 1.20001
R8698 VDD.n2601 VDD.n2600 1.20001
R8699 VDD.n64 VDD.n63 1.1947
R8700 VDD.n1773 VDD.n1772 1.1947
R8701 VDD.n6798 VDD.n6797 1.15635
R8702 VDD.n6710 VDD.n6709 1.15635
R8703 VDD.n6618 VDD.n6617 1.15635
R8704 VDD.n6530 VDD.n6529 1.15635
R8705 VDD.n3629 VDD.n3628 1.15386
R8706 VDD.n8103 VDD.n8102 1.15182
R8707 VDD.n8216 VDD.n8215 1.15182
R8708 VDD.n8321 VDD.n8320 1.15182
R8709 VDD.n8438 VDD.n8437 1.15182
R8710 VDD.n8790 VDD.n8761 1.13602
R8711 VDD.n4642 VDD.n4638 1.12991
R8712 VDD.n5174 VDD.n5170 1.12991
R8713 VDD.n4296 VDD.n4295 1.12991
R8714 VDD.n5325 VDD.n5324 1.12991
R8715 VDD.n8628 VDD.n8624 1.12991
R8716 VDD.n8990 VDD.n8986 1.12991
R8717 VDD.n8900 VDD.n8896 1.12991
R8718 VDD.n7556 VDD.n7555 1.12991
R8719 VDD.n7510 VDD.n7509 1.12991
R8720 VDD.n3933 VDD.n3932 1.12991
R8721 VDD.n3923 VDD.n3922 1.12991
R8722 VDD.n3174 VDD.n3171 1.11541
R8723 VDD.n3178 VDD.n3176 1.11541
R8724 VDD.n3184 VDD.n3181 1.11541
R8725 VDD.n3189 VDD.n3186 1.11541
R8726 VDD.n3196 VDD.n3192 1.11541
R8727 VDD.n3200 VDD.n3198 1.11541
R8728 VDD.n1921 VDD.n1808 1.11541
R8729 VDD.n1920 VDD.n1833 1.11541
R8730 VDD.n1916 VDD.n1915 1.11541
R8731 VDD.n1913 VDD.n1912 1.11541
R8732 VDD.n1910 VDD.n1837 1.11541
R8733 VDD.n1907 VDD.n1906 1.11541
R8734 VDD.n1067 VDD.n954 1.11541
R8735 VDD.n1066 VDD.n979 1.11541
R8736 VDD.n1062 VDD.n1061 1.11541
R8737 VDD.n1059 VDD.n1058 1.11541
R8738 VDD.n1056 VDD.n983 1.11541
R8739 VDD.n1053 VDD.n1052 1.11541
R8740 VDD.n212 VDD.n99 1.11541
R8741 VDD.n211 VDD.n124 1.11541
R8742 VDD.n207 VDD.n206 1.11541
R8743 VDD.n204 VDD.n203 1.11541
R8744 VDD.n201 VDD.n128 1.11541
R8745 VDD.n198 VDD.n197 1.11541
R8746 VDD.n8714 VDD.n8713 1.10918
R8747 VDD.n8949 VDD.n8948 1.10899
R8748 VDD.n8672 VDD.n8669 1.10899
R8749 VDD.n48 VDD 1.09833
R8750 VDD.n1757 VDD 1.09833
R8751 VDD.n8578 VDD.n8577 1.09663
R8752 VDD.n6487 VDD.n6486 1.08525
R8753 VDD.n6408 VDD.n6407 1.08525
R8754 VDD.n6325 VDD.n6324 1.08525
R8755 VDD.n6237 VDD.n6236 1.08525
R8756 VDD.n6164 VDD.n6163 1.08525
R8757 VDD.n6094 VDD.n6093 1.08525
R8758 VDD.n6016 VDD.n6015 1.08525
R8759 VDD.n5928 VDD.n5927 1.08525
R8760 VDD.n8170 VDD.n8169 1.0841
R8761 VDD.n8275 VDD.n8274 1.0841
R8762 VDD.n8380 VDD.n8379 1.0841
R8763 VDD.n8528 VDD.n8527 1.0841
R8764 VDD.n7463 VDD.n7462 1.07839
R8765 VDD.n7432 VDD.n7431 1.07839
R8766 VDD.n7394 VDD.n7393 1.07839
R8767 VDD.n7363 VDD.n7362 1.07839
R8768 VDD.n7321 VDD.n7320 1.07839
R8769 VDD.n7282 VDD.n7281 1.07839
R8770 VDD.n7234 VDD.n7233 1.07839
R8771 VDD.n7195 VDD.n7194 1.07839
R8772 VDD.n7147 VDD.n7146 1.07839
R8773 VDD.n3601 VDD.n3600 1.07073
R8774 VDD.n6775 VDD.n6774 1.07073
R8775 VDD.n6689 VDD.n6688 1.07073
R8776 VDD.n6595 VDD.n6594 1.07073
R8777 VDD.n6511 VDD.n6510 1.07073
R8778 VDD.n8790 VDD.n8789 1.04225
R8779 VDD.n9013 VDD.n9012 1.0272
R8780 VDD.n9013 VDD.n8748 1.02649
R8781 VDD.n3626 VDD.n3454 1.02165
R8782 VDD.n4693 VDD.n4692 0.994314
R8783 VDD.n4709 VDD.n4708 0.994314
R8784 VDD.n5034 VDD.n5033 0.994314
R8785 VDD.n5050 VDD.n5049 0.994314
R8786 VDD.n4331 VDD.n4330 0.994314
R8787 VDD.n4347 VDD.n4346 0.994314
R8788 VDD.n4414 VDD.n4413 0.994314
R8789 VDD.n4512 VDD.n4511 0.994314
R8790 VDD.n4442 VDD.n4441 0.994314
R8791 VDD.n4432 VDD.n4431 0.994314
R8792 VDD.n3651 VDD.n3650 0.994314
R8793 VDD.n5268 VDD.n5267 0.994314
R8794 VDD.n6803 VDD.n6802 0.985115
R8795 VDD.n6715 VDD.n6714 0.985115
R8796 VDD.n6623 VDD.n6622 0.985115
R8797 VDD.n6535 VDD.n6534 0.985115
R8798 VDD.n8000 VDD.n7999 0.950995
R8799 VDD.n7930 VDD.n7929 0.950995
R8800 VDD.n7858 VDD.n7857 0.950995
R8801 VDD.n7798 VDD.n7797 0.950995
R8802 VDD.n7726 VDD.n7725 0.950995
R8803 VDD.n7656 VDD.n7655 0.950995
R8804 VDD.n7089 VDD.n7088 0.948648
R8805 VDD.n7054 VDD.n7053 0.948648
R8806 VDD.n7001 VDD.n7000 0.948648
R8807 VDD.n6966 VDD.n6965 0.948648
R8808 VDD.n6913 VDD.n6912 0.948648
R8809 VDD.n6878 VDD.n6877 0.948648
R8810 VDD.n5454 VDD.n5453 0.948648
R8811 VDD.n5489 VDD.n5488 0.948648
R8812 VDD.n5542 VDD.n5541 0.948648
R8813 VDD.n5577 VDD.n5576 0.948648
R8814 VDD.n5630 VDD.n5629 0.948648
R8815 VDD.n5665 VDD.n5664 0.948648
R8816 VDD.n5718 VDD.n5717 0.948648
R8817 VDD.n5753 VDD.n5752 0.948648
R8818 VDD.n5806 VDD.n5805 0.948648
R8819 VDD.n6673 VDD.n6670 0.942306
R8820 VDD.n8859 VDD.n8858 0.942306
R8821 VDD.n6440 VDD.n6439 0.940613
R8822 VDD.n6360 VDD.n6359 0.940613
R8823 VDD.n6272 VDD.n6271 0.940613
R8824 VDD.n6192 VDD.n6191 0.940613
R8825 VDD.n6122 VDD.n6121 0.940613
R8826 VDD.n6051 VDD.n6050 0.940613
R8827 VDD.n5963 VDD.n5962 0.940613
R8828 VDD.n5875 VDD.n5874 0.940613
R8829 VDD.n3372 VDD.n3369 0.934239
R8830 VDD.n3365 VDD.n3362 0.934239
R8831 VDD.n3360 VDD.n3358 0.934239
R8832 VDD.n3355 VDD.n3352 0.934239
R8833 VDD.n3350 VDD.n3348 0.934239
R8834 VDD.n3345 VDD.n3342 0.934239
R8835 VDD.n1871 VDD.n1870 0.934239
R8836 VDD.n1869 VDD.n1868 0.934239
R8837 VDD.n1865 VDD.n1842 0.934239
R8838 VDD.n1864 VDD.n1845 0.934239
R8839 VDD.n1860 VDD.n1859 0.934239
R8840 VDD.n1855 VDD.n1854 0.934239
R8841 VDD.n1017 VDD.n1016 0.934239
R8842 VDD.n1015 VDD.n1014 0.934239
R8843 VDD.n1011 VDD.n988 0.934239
R8844 VDD.n1010 VDD.n991 0.934239
R8845 VDD.n1006 VDD.n1005 0.934239
R8846 VDD.n1001 VDD.n1000 0.934239
R8847 VDD.n162 VDD.n161 0.934239
R8848 VDD.n160 VDD.n159 0.934239
R8849 VDD.n156 VDD.n133 0.934239
R8850 VDD.n155 VDD.n136 0.934239
R8851 VDD.n151 VDD.n150 0.934239
R8852 VDD.n146 VDD.n145 0.934239
R8853 VDD.n3970 VDD.n3965 0.926297
R8854 VDD.n3974 VDD.n3971 0.926297
R8855 VDD.n4015 VDD.n4012 0.926297
R8856 VDD.n4020 VDD.n4017 0.926297
R8857 VDD.n4024 VDD.n4021 0.926297
R8858 VDD.n4028 VDD.n4025 0.926297
R8859 VDD.n4033 VDD.n4030 0.926297
R8860 VDD.n4057 VDD.n4056 0.926297
R8861 VDD.n4053 VDD.n4052 0.926297
R8862 VDD.n4049 VDD.n4048 0.926297
R8863 VDD.n4045 VDD.n4044 0.926297
R8864 VDD.n4041 VDD.n4040 0.926297
R8865 VDD.n4037 VDD.n4036 0.926297
R8866 VDD.n4214 VDD.n4211 0.926297
R8867 VDD.n4218 VDD.n4215 0.926297
R8868 VDD.n4222 VDD.n4219 0.926297
R8869 VDD.n4234 VDD.n4233 0.926297
R8870 VDD.n4230 VDD.n4229 0.926297
R8871 VDD.n4226 VDD.n4225 0.926297
R8872 VDD.n4087 VDD.n4084 0.926297
R8873 VDD.n4091 VDD.n4088 0.926297
R8874 VDD.n4095 VDD.n4092 0.926297
R8875 VDD.n4099 VDD.n4096 0.926297
R8876 VDD.n4103 VDD.n4100 0.926297
R8877 VDD.n4108 VDD.n4105 0.926297
R8878 VDD.n4197 VDD.n4196 0.926297
R8879 VDD.n4193 VDD.n4192 0.926297
R8880 VDD.n4189 VDD.n4188 0.926297
R8881 VDD.n4185 VDD.n4184 0.926297
R8882 VDD.n4181 VDD.n4180 0.926297
R8883 VDD.n4177 VDD.n4176 0.926297
R8884 VDD.n4173 VDD.n4172 0.926297
R8885 VDD.n4169 VDD.n4168 0.926297
R8886 VDD.n4165 VDD.n4164 0.926297
R8887 VDD.n4161 VDD.n4160 0.926297
R8888 VDD.n4157 VDD.n4156 0.926297
R8889 VDD.n4153 VDD.n4152 0.926297
R8890 VDD.n4145 VDD.n4144 0.926297
R8891 VDD.n4141 VDD.n4140 0.926297
R8892 VDD.n4137 VDD.n4136 0.926297
R8893 VDD.n4133 VDD.n4132 0.926297
R8894 VDD.n4129 VDD.n4128 0.926297
R8895 VDD.n4125 VDD.n4124 0.926297
R8896 VDD.n4121 VDD.n4120 0.926297
R8897 VDD.n8558 VDD.n8557 0.926297
R8898 VDD.n2966 VDD.n2963 0.906695
R8899 VDD.n2960 VDD.n2957 0.906695
R8900 VDD.n2955 VDD.n2952 0.906695
R8901 VDD.n2949 VDD.n2946 0.906695
R8902 VDD.n2944 VDD.n2941 0.906695
R8903 VDD.n2938 VDD.n2935 0.906695
R8904 VDD.n2305 VDD.n2303 0.906695
R8905 VDD.n2308 VDD.n2307 0.906695
R8906 VDD.n2311 VDD.n2291 0.906695
R8907 VDD.n2314 VDD.n2313 0.906695
R8908 VDD.n2317 VDD.n2289 0.906695
R8909 VDD.n2323 VDD.n2319 0.906695
R8910 VDD.n1451 VDD.n1449 0.906695
R8911 VDD.n1454 VDD.n1453 0.906695
R8912 VDD.n1457 VDD.n1437 0.906695
R8913 VDD.n1460 VDD.n1459 0.906695
R8914 VDD.n1463 VDD.n1435 0.906695
R8915 VDD.n1469 VDD.n1465 0.906695
R8916 VDD.n596 VDD.n594 0.906695
R8917 VDD.n599 VDD.n598 0.906695
R8918 VDD.n602 VDD.n582 0.906695
R8919 VDD.n605 VDD.n604 0.906695
R8920 VDD.n608 VDD.n580 0.906695
R8921 VDD.n614 VDD.n610 0.906695
R8922 VDD.n4571 VDD.n4568 0.903353
R8923 VDD.n4585 VDD.n4320 0.903353
R8924 VDD.n3596 VDD.n3595 0.902912
R8925 VDD.n7579 VDD.n7576 0.899959
R8926 VDD.n6770 VDD.n6769 0.899497
R8927 VDD.n6685 VDD.n6684 0.899497
R8928 VDD.n6590 VDD.n6589 0.899497
R8929 VDD.n5248 VDD.n5245 0.884222
R8930 VDD.n5248 VDD.n3760 0.883499
R8931 VDD.n8111 VDD.n8110 0.880923
R8932 VDD.n8222 VDD.n8221 0.880923
R8933 VDD.n8327 VDD.n8326 0.880923
R8934 VDD.n8448 VDD.n8447 0.880923
R8935 VDD.n5844 VDD.n5839 0.880923
R8936 VDD.n7551 VDD.n7550 0.878931
R8937 VDD.n7515 VDD.n7514 0.878931
R8938 VDD.n47 VDD.n45 0.8405
R8939 VDD.n45 VDD 0.8405
R8940 VDD.n1756 VDD.n1754 0.8405
R8941 VDD.n1754 VDD 0.8405
R8942 VDD.n4257 VDD.n4256 0.825441
R8943 VDD.n7640 VDD.n7639 0.824262
R8944 VDD.n4277 VDD.n4268 0.82077
R8945 VDD.n6807 VDD.n6806 0.813878
R8946 VDD.n6720 VDD.n6719 0.813878
R8947 VDD.n6628 VDD.n6627 0.813878
R8948 VDD.n6540 VDD.n6539 0.813878
R8949 VDD.n8164 VDD.n8163 0.813198
R8950 VDD.n8269 VDD.n8268 0.813198
R8951 VDD.n8374 VDD.n8373 0.813198
R8952 VDD.n8520 VDD.n8519 0.813198
R8953 VDD.n8572 VDD.n8571 0.813198
R8954 VDD.n7459 VDD.n7458 0.808921
R8955 VDD.n7436 VDD.n7435 0.808921
R8956 VDD.n7390 VDD.n7389 0.808921
R8957 VDD.n7367 VDD.n7366 0.808921
R8958 VDD.n7316 VDD.n7315 0.808921
R8959 VDD.n7287 VDD.n7286 0.808921
R8960 VDD.n7229 VDD.n7228 0.808921
R8961 VDD.n7200 VDD.n7199 0.808921
R8962 VDD.n7142 VDD.n7141 0.808921
R8963 VDD.n6492 VDD.n6491 0.79598
R8964 VDD.n6413 VDD.n6412 0.79598
R8965 VDD.n6330 VDD.n6329 0.79598
R8966 VDD.n6242 VDD.n6241 0.79598
R8967 VDD.n6168 VDD.n6167 0.79598
R8968 VDD.n6098 VDD.n6097 0.79598
R8969 VDD.n6021 VDD.n6020 0.79598
R8970 VDD.n5933 VDD.n5932 0.79598
R8971 VDD.n5845 VDD.n5836 0.79598
R8972 VDD.n4109 VDD.n4108 0.79404
R8973 VDD.n3842 VDD.n3841 0.775778
R8974 VDD.n5018 VDD.n5017 0.775778
R8975 VDD.n40 VDD.n39 0.761777
R8976 VDD.n902 VDD.n901 0.761777
R8977 VDD.n1749 VDD.n1748 0.761777
R8978 VDD.n2607 VDD.n2604 0.761777
R8979 VDD.n7580 VDD.n7567 0.761581
R8980 VDD.n4694 VDD.n4690 0.753441
R8981 VDD.n4710 VDD.n4706 0.753441
R8982 VDD.n5035 VDD.n5031 0.753441
R8983 VDD.n5051 VDD.n5047 0.753441
R8984 VDD.n4392 VDD.n4391 0.753441
R8985 VDD.n4332 VDD.n4328 0.753441
R8986 VDD.n4348 VDD.n4344 0.753441
R8987 VDD.n4415 VDD.n4411 0.753441
R8988 VDD.n4513 VDD.n4509 0.753441
R8989 VDD.n4443 VDD.n4439 0.753441
R8990 VDD.n4433 VDD.n4429 0.753441
R8991 VDD.n4485 VDD.n4484 0.753441
R8992 VDD.n4555 VDD.n4554 0.753441
R8993 VDD.n4304 VDD.n4303 0.753441
R8994 VDD.n3694 VDD.n3693 0.753441
R8995 VDD.n3652 VDD.n3648 0.753441
R8996 VDD.n3737 VDD.n3736 0.753441
R8997 VDD.n5333 VDD.n5332 0.753441
R8998 VDD.n5269 VDD.n5265 0.753441
R8999 VDD.n8656 VDD.n8655 0.753441
R9000 VDD.n8603 VDD.n8602 0.753441
R9001 VDD.n8704 VDD.n8703 0.753441
R9002 VDD.n8681 VDD.n8680 0.753441
R9003 VDD.n8735 VDD.n8734 0.753441
R9004 VDD.n8965 VDD.n8964 0.753441
R9005 VDD.n8935 VDD.n8934 0.753441
R9006 VDD.n8882 VDD.n8881 0.753441
R9007 VDD.n3883 VDD.n3882 0.753441
R9008 VDD.n3897 VDD.n3896 0.753441
R9009 VDD.n3168 VDD.n3166 0.750919
R9010 VDD.n3410 VDD.n3385 0.750919
R9011 VDD.n2537 VDD.n2536 0.750919
R9012 VDD.n1898 VDD.n1825 0.750919
R9013 VDD.n1683 VDD.n1682 0.750919
R9014 VDD.n1044 VDD.n971 0.750919
R9015 VDD.n828 VDD.n827 0.750919
R9016 VDD.n189 VDD.n116 0.750919
R9017 VDD.n4575 VDD.n4498 0.743006
R9018 VDD.n3710 VDD.n3707 0.743006
R9019 VDD.n4580 VDD.n4405 0.742904
R9020 VDD.n6765 VDD.n6764 0.728259
R9021 VDD.n6681 VDD.n6680 0.728259
R9022 VDD.n6585 VDD.n6584 0.728259
R9023 VDD.n8850 VDD.n8848 0.728259
R9024 VDD.n4076 VDD.n3948 0.724685
R9025 VDD.n4076 VDD.n4075 0.724297
R9026 VDD.n3596 VDD.n3575 0.71293
R9027 VDD.n3166 VDD.n3165 0.708038
R9028 VDD.n2537 VDD.n1807 0.708038
R9029 VDD.n1683 VDD.n953 0.708038
R9030 VDD.n828 VDD.n98 0.708038
R9031 VDD.n3338 VDD.n3335 0.700804
R9032 VDD.n1939 VDD.n1818 0.700804
R9033 VDD.n1085 VDD.n964 0.700804
R9034 VDD.n230 VDD.n109 0.700804
R9035 VDD.n5434 VDD.n3629 0.699924
R9036 VDD.n8008 VDD.n8007 0.69753
R9037 VDD.n7922 VDD.n7921 0.69753
R9038 VDD.n7866 VDD.n7865 0.69753
R9039 VDD.n7790 VDD.n7789 0.69753
R9040 VDD.n7734 VDD.n7733 0.69753
R9041 VDD.n7648 VDD.n7647 0.69753
R9042 VDD.n4257 VDD.n4251 0.692441
R9043 VDD.n4277 VDD.n4274 0.689368
R9044 VDD.n48 VDD 0.682932
R9045 VDD.n48 VDD 0.682932
R9046 VDD.n1757 VDD 0.682932
R9047 VDD.n1757 VDD 0.682932
R9048 VDD.n8675 VDD.n8674 0.682531
R9049 VDD.n4836 VDD.n4835 0.682531
R9050 VDD.n4866 VDD.n4865 0.682531
R9051 VDD.n4896 VDD.n4895 0.682531
R9052 VDD.n4926 VDD.n4925 0.682531
R9053 VDD.n4988 VDD.n4987 0.6825
R9054 VDD.n4978 VDD.n4977 0.6825
R9055 VDD.n5369 VDD.n5365 0.6825
R9056 VDD.n2930 VDD.n2928 0.680146
R9057 VDD.n2320 VDD.n2002 0.680146
R9058 VDD.n1466 VDD.n1148 0.680146
R9059 VDD.n611 VDD.n293 0.680146
R9060 VDD.n7084 VDD.n7083 0.677749
R9061 VDD.n7059 VDD.n7058 0.677749
R9062 VDD.n6996 VDD.n6995 0.677749
R9063 VDD.n6971 VDD.n6970 0.677749
R9064 VDD.n6908 VDD.n6907 0.677749
R9065 VDD.n6883 VDD.n6882 0.677749
R9066 VDD.n5459 VDD.n5458 0.677749
R9067 VDD.n5484 VDD.n5483 0.677749
R9068 VDD.n5547 VDD.n5546 0.677749
R9069 VDD.n5572 VDD.n5571 0.677749
R9070 VDD.n5635 VDD.n5634 0.677749
R9071 VDD.n5660 VDD.n5659 0.677749
R9072 VDD.n5723 VDD.n5722 0.677749
R9073 VDD.n5748 VDD.n5747 0.677749
R9074 VDD.n5811 VDD.n5810 0.677749
R9075 VDD.t130 VDD.n4080 0.661784
R9076 VDD.n4149 VDD.t77 0.661784
R9077 VDD.n6436 VDD.n6435 0.651347
R9078 VDD.n6355 VDD.n6354 0.651347
R9079 VDD.n6267 VDD.n6266 0.651347
R9080 VDD.n6188 VDD.n6187 0.651347
R9081 VDD.n6118 VDD.n6117 0.651347
R9082 VDD.n6046 VDD.n6045 0.651347
R9083 VDD.n5958 VDD.n5957 0.651347
R9084 VDD.n5870 VDD.n5869 0.651347
R9085 VDD.n8855 VDD.n8854 0.647691
R9086 VDD.n6811 VDD.n6810 0.64264
R9087 VDD.n6725 VDD.n6724 0.64264
R9088 VDD.n6632 VDD.n6631 0.64264
R9089 VDD.n6545 VDD.n6544 0.64264
R9090 VDD.n8873 VDD.n8872 0.629701
R9091 VDD.n7546 VDD.n7545 0.627951
R9092 VDD.n7520 VDD.n7519 0.627951
R9093 VDD.n5226 VDD.n5225 0.614024
R9094 VDD.n2979 VDD.n2976 0.612674
R9095 VDD.n2985 VDD.n2982 0.612674
R9096 VDD.n2991 VDD.n2988 0.612674
R9097 VDD.n2997 VDD.n2994 0.612674
R9098 VDD.n2292 VDD.n2230 0.612674
R9099 VDD.n2370 VDD.n2369 0.612674
R9100 VDD.n2368 VDD.n2367 0.612674
R9101 VDD.n2247 VDD.n2235 0.612674
R9102 VDD.n1438 VDD.n1376 0.612674
R9103 VDD.n1516 VDD.n1515 0.612674
R9104 VDD.n1514 VDD.n1513 0.612674
R9105 VDD.n1393 VDD.n1381 0.612674
R9106 VDD.n583 VDD.n521 0.612674
R9107 VDD.n661 VDD.n660 0.612674
R9108 VDD.n659 VDD.n658 0.612674
R9109 VDD.n538 VDD.n526 0.612674
R9110 VDD.n8117 VDD.n8116 0.610024
R9111 VDD.n8228 VDD.n8227 0.610024
R9112 VDD.n8333 VDD.n8332 0.610024
R9113 VDD.n8458 VDD.n8457 0.610024
R9114 VDD.n2782 VDD.n2779 0.60463
R9115 VDD.n2788 VDD.n2785 0.60463
R9116 VDD.n2793 VDD.n2790 0.60463
R9117 VDD.n2799 VDD.n2796 0.60463
R9118 VDD.n2804 VDD.n2801 0.60463
R9119 VDD.n2810 VDD.n2808 0.60463
R9120 VDD.n2392 VDD.n2216 0.60463
R9121 VDD.n2227 VDD.n2225 0.60463
R9122 VDD.n2386 VDD.n2385 0.60463
R9123 VDD.n2383 VDD.n2382 0.60463
R9124 VDD.n2380 VDD.n2378 0.60463
R9125 VDD.n2376 VDD.n2228 0.60463
R9126 VDD.n1538 VDD.n1362 0.60463
R9127 VDD.n1373 VDD.n1371 0.60463
R9128 VDD.n1532 VDD.n1531 0.60463
R9129 VDD.n1529 VDD.n1528 0.60463
R9130 VDD.n1526 VDD.n1524 0.60463
R9131 VDD.n1522 VDD.n1374 0.60463
R9132 VDD.n683 VDD.n507 0.60463
R9133 VDD.n518 VDD.n516 0.60463
R9134 VDD.n677 VDD.n676 0.60463
R9135 VDD.n674 VDD.n673 0.60463
R9136 VDD.n671 VDD.n669 0.60463
R9137 VDD.n667 VDD.n519 0.60463
R9138 VDD.n5350 VDD.n5349 0.604026
R9139 VDD.n5364 VDD.n3750 0.603703
R9140 VDD.n3750 VDD.n3724 0.576974
R9141 VDD.n8054 VDD.n8051 0.570797
R9142 VDD.n7635 VDD.n7634 0.570797
R9143 VDD.n9018 VDD.n9017 0.568833
R9144 VDD.n6760 VDD.n6759 0.557022
R9145 VDD.n6677 VDD.n6676 0.557022
R9146 VDD.n6580 VDD.n6579 0.557022
R9147 VDD.n8858 VDD.n8857 0.557022
R9148 VDD.n46 VDD.n3 0.544383
R9149 VDD.n919 VDD.n918 0.544383
R9150 VDD.n1755 VDD.n1712 0.544383
R9151 VDD.n2628 VDD.n2627 0.544383
R9152 VDD.n8158 VDD.n8157 0.542299
R9153 VDD.n8263 VDD.n8262 0.542299
R9154 VDD.n8368 VDD.n8367 0.542299
R9155 VDD.n8511 VDD.n8510 0.542299
R9156 VDD.n7455 VDD.n7454 0.539447
R9157 VDD.n7440 VDD.n7439 0.539447
R9158 VDD.n7386 VDD.n7385 0.539447
R9159 VDD.n7371 VDD.n7370 0.539447
R9160 VDD.n7311 VDD.n7310 0.539447
R9161 VDD.n7292 VDD.n7291 0.539447
R9162 VDD.n7224 VDD.n7223 0.539447
R9163 VDD.n7205 VDD.n7204 0.539447
R9164 VDD.n7137 VDD.n7136 0.539447
R9165 VDD.n917 VDD 0.530391
R9166 VDD.n2626 VDD 0.530391
R9167 VDD.n8565 VDD.n8564 0.529527
R9168 VDD.n3625 VDD.n3540 0.522949
R9169 VDD.n3411 VDD.n3211 0.515073
R9170 VDD.n1900 VDD.n1899 0.515073
R9171 VDD.n1046 VDD.n1045 0.515073
R9172 VDD.n191 VDD.n190 0.515073
R9173 VDD.n6502 VDD.n6501 0.506715
R9174 VDD.n6417 VDD.n6416 0.506715
R9175 VDD.n6335 VDD.n6334 0.506715
R9176 VDD.n6247 VDD.n6246 0.506715
R9177 VDD.n6172 VDD.n6171 0.506715
R9178 VDD.n6102 VDD.n6101 0.506715
R9179 VDD.n6026 VDD.n6025 0.506715
R9180 VDD.n5938 VDD.n5937 0.506715
R9181 VDD.n5850 VDD.n5849 0.506715
R9182 VDD.n7576 VDD.n7575 0.502461
R9183 VDD.n916 VDD 0.497949
R9184 VDD.n2625 VDD 0.497949
R9185 VDD.n4078 VDD.n4077 0.491125
R9186 VDD.n4599 VDD.n4598 0.488891
R9187 VDD.n4079 VDD.n4078 0.488
R9188 VDD.n7585 VDD.n7584 0.484824
R9189 VDD.n4475 VDD.n4474 0.48381
R9190 VDD.n3684 VDD.n3683 0.483797
R9191 VDD.n8684 VDD.n8683 0.476817
R9192 VDD.n8064 VDD.n8061 0.474574
R9193 VDD.n8070 VDD.n8068 0.474574
R9194 VDD.n8088 VDD.n8086 0.474574
R9195 VDD.n8096 VDD.n8093 0.474574
R9196 VDD.n8102 VDD.n8100 0.474574
R9197 VDD.n8110 VDD.n8107 0.474574
R9198 VDD.n8116 VDD.n8114 0.474574
R9199 VDD.n8124 VDD.n8121 0.474574
R9200 VDD.n8131 VDD.n8128 0.474574
R9201 VDD.n8146 VDD.n8144 0.474574
R9202 VDD.n8151 VDD.n8149 0.474574
R9203 VDD.n8157 VDD.n8155 0.474574
R9204 VDD.n8163 VDD.n8161 0.474574
R9205 VDD.n8169 VDD.n8167 0.474574
R9206 VDD.n8175 VDD.n8173 0.474574
R9207 VDD.n8181 VDD.n8179 0.474574
R9208 VDD.n8187 VDD.n8185 0.474574
R9209 VDD.n8203 VDD.n8201 0.474574
R9210 VDD.n8209 VDD.n8207 0.474574
R9211 VDD.n8215 VDD.n8213 0.474574
R9212 VDD.n8221 VDD.n8219 0.474574
R9213 VDD.n8227 VDD.n8225 0.474574
R9214 VDD.n8233 VDD.n8231 0.474574
R9215 VDD.n8239 VDD.n8237 0.474574
R9216 VDD.n8251 VDD.n8249 0.474574
R9217 VDD.n8256 VDD.n8254 0.474574
R9218 VDD.n8262 VDD.n8260 0.474574
R9219 VDD.n8268 VDD.n8266 0.474574
R9220 VDD.n8274 VDD.n8272 0.474574
R9221 VDD.n8280 VDD.n8278 0.474574
R9222 VDD.n8286 VDD.n8284 0.474574
R9223 VDD.n8292 VDD.n8290 0.474574
R9224 VDD.n8308 VDD.n8306 0.474574
R9225 VDD.n8314 VDD.n8312 0.474574
R9226 VDD.n8320 VDD.n8318 0.474574
R9227 VDD.n8326 VDD.n8324 0.474574
R9228 VDD.n8332 VDD.n8330 0.474574
R9229 VDD.n8338 VDD.n8336 0.474574
R9230 VDD.n8344 VDD.n8342 0.474574
R9231 VDD.n8356 VDD.n8354 0.474574
R9232 VDD.n8361 VDD.n8359 0.474574
R9233 VDD.n8367 VDD.n8365 0.474574
R9234 VDD.n8373 VDD.n8371 0.474574
R9235 VDD.n8379 VDD.n8377 0.474574
R9236 VDD.n8385 VDD.n8383 0.474574
R9237 VDD.n8391 VDD.n8389 0.474574
R9238 VDD.n8397 VDD.n8395 0.474574
R9239 VDD.n8417 VDD.n8414 0.474574
R9240 VDD.n8427 VDD.n8424 0.474574
R9241 VDD.n8437 VDD.n8434 0.474574
R9242 VDD.n8447 VDD.n8444 0.474574
R9243 VDD.n8457 VDD.n8454 0.474574
R9244 VDD.n8466 VDD.n8463 0.474574
R9245 VDD.n8475 VDD.n8472 0.474574
R9246 VDD.n8493 VDD.n8489 0.474574
R9247 VDD.n8501 VDD.n8497 0.474574
R9248 VDD.n8510 VDD.n8506 0.474574
R9249 VDD.n8519 VDD.n8515 0.474574
R9250 VDD.n8527 VDD.n8524 0.474574
R9251 VDD.n8535 VDD.n8532 0.474574
R9252 VDD.n8541 VDD.n8539 0.474574
R9253 VDD.n3727 VDD.n3726 0.473002
R9254 VDD.n6815 VDD.n6814 0.471403
R9255 VDD.n6730 VDD.n6729 0.471403
R9256 VDD.n6636 VDD.n6635 0.471403
R9257 VDD.n6550 VDD.n6549 0.471403
R9258 VDD.n4545 VDD.n4544 0.469257
R9259 VDD.n4382 VDD.n4381 0.469245
R9260 VDD.n8800 VDD.n8799 0.461585
R9261 VDD.n5278 VDD.n5276 0.444775
R9262 VDD.n8016 VDD.n8015 0.444064
R9263 VDD.n7914 VDD.n7913 0.444064
R9264 VDD.n7874 VDD.n7873 0.444064
R9265 VDD.n7782 VDD.n7781 0.444064
R9266 VDD.n7742 VDD.n7741 0.444064
R9267 VDD.n7635 VDD.n7619 0.444064
R9268 VDD.n2630 VDD 0.435138
R9269 VDD.n6499 VDD.n6495 0.431961
R9270 VDD.n8058 VDD.n8044 0.428211
R9271 VDD.n921 VDD 0.427658
R9272 VDD.n6597 VDD.t41 0.42104
R9273 VDD.n8786 VDD.n8785 0.42104
R9274 VDD.n8862 VDD.n8840 0.42104
R9275 VDD.n8839 VDD.n8838 0.42104
R9276 VDD.n7079 VDD.n7078 0.406849
R9277 VDD.n7064 VDD.n7063 0.406849
R9278 VDD.n6991 VDD.n6990 0.406849
R9279 VDD.n6976 VDD.n6975 0.406849
R9280 VDD.n6903 VDD.n6902 0.406849
R9281 VDD.n6888 VDD.n6887 0.406849
R9282 VDD.n5464 VDD.n5463 0.406849
R9283 VDD.n5479 VDD.n5478 0.406849
R9284 VDD.n5552 VDD.n5551 0.406849
R9285 VDD.n5567 VDD.n5566 0.406849
R9286 VDD.n5640 VDD.n5639 0.406849
R9287 VDD.n5655 VDD.n5654 0.406849
R9288 VDD.n5728 VDD.n5727 0.406849
R9289 VDD.n5743 VDD.n5742 0.406849
R9290 VDD.n5816 VDD.n5815 0.406849
R9291 VDD.n5831 VDD.n5830 0.406849
R9292 VDD.n4813 VDD.n4812 0.400769
R9293 VDD.n4846 VDD.n4845 0.400769
R9294 VDD.n4936 VDD.n4935 0.400769
R9295 VDD.n4876 VDD.n4875 0.400768
R9296 VDD.n4906 VDD.n4905 0.400768
R9297 VDD.n3852 VDD.n3851 0.400768
R9298 VDD.n3819 VDD.n3818 0.400768
R9299 VDD.n4069 VDD.n4033 0.39727
R9300 VDD.n9031 VDD.n9030 0.388641
R9301 VDD.n6755 VDD.n6754 0.385784
R9302 VDD.n6673 VDD.n6672 0.385784
R9303 VDD.n6575 VDD.n6574 0.385784
R9304 VDD.n8023 VDD.n8020 0.380698
R9305 VDD.n8015 VDD.n8012 0.380698
R9306 VDD.n8007 VDD.n8004 0.380698
R9307 VDD.n7999 VDD.n7996 0.380698
R9308 VDD.n7991 VDD.n7988 0.380698
R9309 VDD.n7983 VDD.n7980 0.380698
R9310 VDD.n7972 VDD.n7969 0.380698
R9311 VDD.n7956 VDD.n7953 0.380698
R9312 VDD.n7945 VDD.n7942 0.380698
R9313 VDD.n7937 VDD.n7934 0.380698
R9314 VDD.n7929 VDD.n7926 0.380698
R9315 VDD.n7921 VDD.n7918 0.380698
R9316 VDD.n7913 VDD.n7910 0.380698
R9317 VDD.n7905 VDD.n7902 0.380698
R9318 VDD.n7881 VDD.n7878 0.380698
R9319 VDD.n7873 VDD.n7870 0.380698
R9320 VDD.n7865 VDD.n7862 0.380698
R9321 VDD.n7857 VDD.n7854 0.380698
R9322 VDD.n7849 VDD.n7846 0.380698
R9323 VDD.n7841 VDD.n7838 0.380698
R9324 VDD.n7831 VDD.n7828 0.380698
R9325 VDD.n7817 VDD.n7815 0.380698
R9326 VDD.n7809 VDD.n7807 0.380698
R9327 VDD.n7803 VDD.n7801 0.380698
R9328 VDD.n7797 VDD.n7794 0.380698
R9329 VDD.n7789 VDD.n7786 0.380698
R9330 VDD.n7781 VDD.n7778 0.380698
R9331 VDD.n7773 VDD.n7770 0.380698
R9332 VDD.n7749 VDD.n7746 0.380698
R9333 VDD.n7741 VDD.n7738 0.380698
R9334 VDD.n7733 VDD.n7730 0.380698
R9335 VDD.n7725 VDD.n7722 0.380698
R9336 VDD.n7717 VDD.n7714 0.380698
R9337 VDD.n7709 VDD.n7706 0.380698
R9338 VDD.n7698 VDD.n7695 0.380698
R9339 VDD.n7682 VDD.n7679 0.380698
R9340 VDD.n7671 VDD.n7668 0.380698
R9341 VDD.n7663 VDD.n7660 0.380698
R9342 VDD.n7655 VDD.n7652 0.380698
R9343 VDD.n7647 VDD.n7644 0.380698
R9344 VDD.n6504 VDD.n6503 0.378512
R9345 VDD.n4631 VDD.n4627 0.376971
R9346 VDD.n5163 VDD.n5159 0.376971
R9347 VDD.n4284 VDD.n4281 0.376971
R9348 VDD.n4297 VDD.n4296 0.376971
R9349 VDD.n4313 VDD.n4312 0.376971
R9350 VDD.n5313 VDD.n5309 0.376971
R9351 VDD.n5326 VDD.n5325 0.376971
R9352 VDD.n5342 VDD.n5341 0.376971
R9353 VDD.n5261 VDD.n5260 0.376971
R9354 VDD.n8664 VDD.n8663 0.376971
R9355 VDD.n8667 VDD.n8666 0.376971
R9356 VDD.n8647 VDD.n8646 0.376971
R9357 VDD.n8610 VDD.n8609 0.376971
R9358 VDD.n8617 VDD.n8613 0.376971
R9359 VDD.n8709 VDD.n8708 0.376971
R9360 VDD.n8743 VDD.n8742 0.376971
R9361 VDD.n8746 VDD.n8745 0.376971
R9362 VDD.n9010 VDD.n9009 0.376971
R9363 VDD.n8972 VDD.n8971 0.376971
R9364 VDD.n8979 VDD.n8975 0.376971
R9365 VDD.n8943 VDD.n8942 0.376971
R9366 VDD.n8946 VDD.n8945 0.376971
R9367 VDD.n8926 VDD.n8925 0.376971
R9368 VDD.n8913 VDD.n8912 0.376971
R9369 VDD.n8889 VDD.n8885 0.376971
R9370 VDD.n7541 VDD.n7540 0.376971
R9371 VDD.n7525 VDD.n7524 0.376971
R9372 VDD.n6431 VDD.n6430 0.362082
R9373 VDD.n6350 VDD.n6349 0.362082
R9374 VDD.n6262 VDD.n6261 0.362082
R9375 VDD.n6184 VDD.n6183 0.362082
R9376 VDD.n6114 VDD.n6113 0.362082
R9377 VDD.n6041 VDD.n6040 0.362082
R9378 VDD.n5953 VDD.n5952 0.362082
R9379 VDD.n5865 VDD.n5864 0.362082
R9380 VDD.n3892 VDD.n3890 0.357498
R9381 VDD.n7600 VDD.n7599 0.346446
R9382 VDD.n3176 VDD.n3174 0.343549
R9383 VDD.n3181 VDD.n3178 0.343549
R9384 VDD.n3186 VDD.n3184 0.343549
R9385 VDD.n3192 VDD.n3189 0.343549
R9386 VDD.n3198 VDD.n3196 0.343549
R9387 VDD.n3205 VDD.n3200 0.343549
R9388 VDD.n1921 VDD.n1920 0.343549
R9389 VDD.n1916 VDD.n1833 0.343549
R9390 VDD.n1915 VDD.n1913 0.343549
R9391 VDD.n1912 VDD.n1910 0.343549
R9392 VDD.n1907 VDD.n1837 0.343549
R9393 VDD.n1906 VDD.n1905 0.343549
R9394 VDD.n1067 VDD.n1066 0.343549
R9395 VDD.n1062 VDD.n979 0.343549
R9396 VDD.n1061 VDD.n1059 0.343549
R9397 VDD.n1058 VDD.n1056 0.343549
R9398 VDD.n1053 VDD.n983 0.343549
R9399 VDD.n1052 VDD.n1051 0.343549
R9400 VDD.n212 VDD.n211 0.343549
R9401 VDD.n207 VDD.n124 0.343549
R9402 VDD.n206 VDD.n204 0.343549
R9403 VDD.n203 VDD.n201 0.343549
R9404 VDD.n198 VDD.n128 0.343549
R9405 VDD.n197 VDD.n196 0.343549
R9406 VDD.n3661 VDD.n3659 0.34084
R9407 VDD.n8125 VDD.n8124 0.339124
R9408 VDD.n8234 VDD.n8233 0.339124
R9409 VDD.n8339 VDD.n8338 0.339124
R9410 VDD.n8467 VDD.n8466 0.339124
R9411 VDD.n7120 VDD.n7119 0.337342
R9412 VDD.n3762 VDD.n3761 0.33059
R9413 VDD.n5238 VDD.n3806 0.33059
R9414 VDD.n3805 VDD.n3804 0.33059
R9415 VDD.n914 VDD 0.329892
R9416 VDD.n2623 VDD 0.329892
R9417 VDD.n4583 VDD.n4582 0.324719
R9418 VDD.n4578 VDD.n4577 0.324719
R9419 VDD.n4574 VDD.n4573 0.324719
R9420 VDD.n4681 VDD.n4680 0.324719
R9421 VDD.n4804 VDD.n4803 0.324719
R9422 VDD.n5022 VDD.n5021 0.324719
R9423 VDD.n5147 VDD.n5146 0.324719
R9424 VDD.n8043 VDD.n8042 0.317332
R9425 VDD.n8032 VDD.n8028 0.317332
R9426 VDD.n7898 VDD.n7897 0.317332
R9427 VDD.n7890 VDD.n7886 0.317332
R9428 VDD.n7766 VDD.n7765 0.317332
R9429 VDD.n7758 VDD.n7754 0.317332
R9430 VDD.n7581 VDD.n7564 0.313753
R9431 VDD.n8573 VDD.n8572 0.30922
R9432 VDD.n6819 VDD.n6818 0.300166
R9433 VDD.n6735 VDD.n6734 0.300166
R9434 VDD.n6640 VDD.n6639 0.300166
R9435 VDD.n6555 VDD.n6554 0.300166
R9436 VDD.n918 VDD 0.299413
R9437 VDD.n2627 VDD 0.299413
R9438 VDD.n920 VDD.n857 0.292759
R9439 VDD.n2629 VDD.n2601 0.292759
R9440 VDD.n65 VDD.n64 0.292507
R9441 VDD.n1774 VDD.n1773 0.292507
R9442 VDD.n4950 VDD.n4949 0.278729
R9443 VDD.n4860 VDD.n4859 0.278729
R9444 VDD.n4830 VDD.n4829 0.278729
R9445 VDD.n4920 VDD.n4919 0.278729
R9446 VDD.n5141 VDD.n5140 0.278729
R9447 VDD.n4890 VDD.n4889 0.278729
R9448 VDD.n4798 VDD.n4797 0.278729
R9449 VDD.n66 VDD 0.278033
R9450 VDD.n1775 VDD 0.278033
R9451 VDD.n7133 VDD.n7125 0.27309
R9452 VDD.n8141 VDD.n8140 0.271399
R9453 VDD.n8152 VDD.n8151 0.271399
R9454 VDD.n8246 VDD.n8245 0.271399
R9455 VDD.n8257 VDD.n8256 0.271399
R9456 VDD.n8351 VDD.n8350 0.271399
R9457 VDD.n8362 VDD.n8361 0.271399
R9458 VDD.n8485 VDD.n8484 0.271399
R9459 VDD.n8502 VDD.n8501 0.271399
R9460 VDD.n7451 VDD.n7450 0.269974
R9461 VDD.n7444 VDD.n7443 0.269974
R9462 VDD.n7382 VDD.n7381 0.269974
R9463 VDD.n7375 VDD.n7374 0.269974
R9464 VDD.n7306 VDD.n7305 0.269974
R9465 VDD.n7297 VDD.n7296 0.269974
R9466 VDD.n7219 VDD.n7218 0.269974
R9467 VDD.n7210 VDD.n7209 0.269974
R9468 VDD.n7132 VDD.n7131 0.269974
R9469 VDD.n3712 VDD.n3711 0.26925
R9470 VDD.n3041 VDD.n3040 0.267107
R9471 VDD.n2559 VDD.n2558 0.267107
R9472 VDD.n1705 VDD.n1704 0.267107
R9473 VDD.n850 VDD.n849 0.267107
R9474 VDD.n4083 VDD.t130 0.265013
R9475 VDD.t77 VDD.n4148 0.265013
R9476 VDD.n52 VDD.n40 0.26137
R9477 VDD.n52 VDD.n51 0.26137
R9478 VDD.n51 VDD.n50 0.26137
R9479 VDD.n903 VDD.n902 0.26137
R9480 VDD.n903 VDD.n858 0.26137
R9481 VDD.n911 VDD.n858 0.26137
R9482 VDD.n1761 VDD.n1749 0.26137
R9483 VDD.n1761 VDD.n1760 0.26137
R9484 VDD.n1760 VDD.n1759 0.26137
R9485 VDD.n2610 VDD.n2607 0.26137
R9486 VDD.n2613 VDD.n2610 0.26137
R9487 VDD.n2620 VDD.n2613 0.26137
R9488 VDD.n3427 VDD 0.260619
R9489 VDD.n3435 VDD.n3434 0.25512
R9490 VDD.n5846 VDD.n5832 0.236946
R9491 VDD.n57 VDD.n34 0.231925
R9492 VDD.n908 VDD.n897 0.231925
R9493 VDD.n1766 VDD.n1743 0.231925
R9494 VDD.n2617 VDD.n2615 0.231925
R9495 VDD.n57 VDD.n56 0.231891
R9496 VDD.n57 VDD.n35 0.231891
R9497 VDD.n908 VDD.n907 0.231891
R9498 VDD.n909 VDD.n908 0.231891
R9499 VDD.n1766 VDD.n1765 0.231891
R9500 VDD.n1766 VDD.n1744 0.231891
R9501 VDD.n2617 VDD.n2616 0.231891
R9502 VDD.n2618 VDD.n2617 0.231891
R9503 VDD.n4717 VDD.n4701 0.229427
R9504 VDD.n4717 VDD.n4716 0.229427
R9505 VDD.n5058 VDD.n5042 0.229427
R9506 VDD.n5058 VDD.n5057 0.229427
R9507 VDD.n4356 VDD.n4339 0.229427
R9508 VDD.n4356 VDD.n4355 0.229427
R9509 VDD.n4450 VDD.n4422 0.229427
R9510 VDD.n4450 VDD.n4449 0.229427
R9511 VDD.n4520 VDD.n4504 0.229427
R9512 VDD.n4520 VDD.n4519 0.229427
R9513 VDD.n921 VDD.n920 0.223437
R9514 VDD.n2630 VDD.n2629 0.22328
R9515 VDD.n66 VDD.n65 0.222418
R9516 VDD.n1775 VDD.n1774 0.222418
R9517 VDD.n6422 VDD.n6421 0.217449
R9518 VDD.n6340 VDD.n6339 0.217449
R9519 VDD.n6252 VDD.n6251 0.217449
R9520 VDD.n6176 VDD.n6175 0.217449
R9521 VDD.n6106 VDD.n6105 0.217449
R9522 VDD.n6031 VDD.n6030 0.217449
R9523 VDD.n5943 VDD.n5942 0.217449
R9524 VDD.n5855 VDD.n5854 0.217449
R9525 VDD.n6826 VDD.n6825 0.216346
R9526 VDD.n4719 VDD.n4717 0.215848
R9527 VDD.n5060 VDD.n5058 0.215848
R9528 VDD.n4452 VDD.n4450 0.215848
R9529 VDD.n4522 VDD.n4520 0.215848
R9530 VDD.n4358 VDD.n4356 0.215848
R9531 VDD.n2633 VDD 0.215174
R9532 VDD.n1781 VDD 0.215174
R9533 VDD.n927 VDD 0.215174
R9534 VDD.n72 VDD 0.215174
R9535 VDD.n6750 VDD.n6749 0.214547
R9536 VDD.n6652 VDD.n6651 0.214547
R9537 VDD.n6570 VDD.n6569 0.214547
R9538 VDD.n7492 VDD.n7490 0.214355
R9539 VDD.n8546 VDD.n6826 0.211367
R9540 VDD.n4069 VDD.n4059 0.211364
R9541 VDD.n4242 VDD.n4199 0.211364
R9542 VDD.n8717 VDD.n8716 0.210656
R9543 VDD.n4674 VDD.n4671 0.210461
R9544 VDD.n5214 VDD.n5211 0.210461
R9545 VDD.n7590 VDD.n7589 0.208068
R9546 VDD.n9028 VDD.n5446 0.204334
R9547 VDD.n8141 VDD.n8135 0.203675
R9548 VDD.n8246 VDD.n8243 0.203675
R9549 VDD.n8351 VDD.n8348 0.203675
R9550 VDD.n8485 VDD.n8480 0.203675
R9551 VDD.n4956 VDD.n4955 0.202844
R9552 VDD.n3411 VDD.n3410 0.193465
R9553 VDD.n1899 VDD.n1898 0.193465
R9554 VDD.n1045 VDD.n1044 0.193465
R9555 VDD.n190 VDD.n189 0.193465
R9556 VDD.n4762 VDD.n4760 0.190717
R9557 VDD.n5103 VDD.n5101 0.190717
R9558 VDD.n4349 VDD.n4342 0.190717
R9559 VDD.n4444 VDD.n4437 0.190717
R9560 VDD.n4437 VDD.n4434 0.190717
R9561 VDD.n8024 VDD.n8023 0.190599
R9562 VDD.n7906 VDD.n7905 0.190599
R9563 VDD.n7882 VDD.n7881 0.190599
R9564 VDD.n7774 VDD.n7773 0.190599
R9565 VDD.n7750 VDD.n7749 0.190599
R9566 VDD.n3912 VDD.n3911 0.189124
R9567 VDD.n8808 VDD.n8807 0.186007
R9568 VDD.n3886 VDD.n3884 0.178063
R9569 VDD.n64 VDD 0.174685
R9570 VDD.n1773 VDD 0.174685
R9571 VDD VDD.n857 0.174507
R9572 VDD VDD.n2601 0.174507
R9573 VDD.n47 VDD 0.167831
R9574 VDD.n1756 VDD 0.167831
R9575 VDD.n3012 VDD.n3008 0.167457
R9576 VDD.n2252 VDD.n2249 0.167457
R9577 VDD.n1398 VDD.n1395 0.167457
R9578 VDD.n543 VDD.n540 0.167457
R9579 VDD.n3882 VDD.n3881 0.166946
R9580 VDD.n4721 VDD.n4719 0.164777
R9581 VDD.n5062 VDD.n5060 0.164777
R9582 VDD.n4454 VDD.n4452 0.164777
R9583 VDD.n4524 VDD.n4522 0.164777
R9584 VDD.n4360 VDD.n4358 0.164777
R9585 VDD.n5280 VDD.n5278 0.164777
R9586 VDD.n4796 VDD.n4795 0.161367
R9587 VDD.n4725 VDD.n4724 0.161367
R9588 VDD.n4828 VDD.n4827 0.161367
R9589 VDD.n4858 VDD.n4857 0.161367
R9590 VDD.n4888 VDD.n4887 0.161367
R9591 VDD.n4918 VDD.n4917 0.161367
R9592 VDD.n4948 VDD.n4947 0.161367
R9593 VDD.n3839 VDD.n3838 0.161367
R9594 VDD.n5013 VDD.n5012 0.161367
R9595 VDD.n5139 VDD.n5138 0.161367
R9596 VDD.n5066 VDD.n5065 0.161367
R9597 VDD.n4364 VDD.n4363 0.161367
R9598 VDD.n4458 VDD.n4457 0.161367
R9599 VDD.n4528 VDD.n4527 0.161367
R9600 VDD.n3667 VDD.n3666 0.161367
R9601 VDD.n4701 VDD.n4699 0.15935
R9602 VDD.n4716 VDD.n4715 0.15935
R9603 VDD.n5042 VDD.n5040 0.15935
R9604 VDD.n5057 VDD.n5056 0.15935
R9605 VDD.n4339 VDD.n4337 0.15935
R9606 VDD.n4355 VDD.n4353 0.15935
R9607 VDD.n4422 VDD.n4420 0.15935
R9608 VDD.n4449 VDD.n4448 0.15935
R9609 VDD.n4519 VDD.n4518 0.15935
R9610 VDD.n3659 VDD.n3657 0.15935
R9611 VDD.n5276 VDD.n5274 0.15935
R9612 VDD.n8575 VDD.n8574 0.157987
R9613 VDD.n4791 VDD.n4790 0.150167
R9614 VDD.n4732 VDD.n4731 0.150167
R9615 VDD.n4808 VDD.n4807 0.150167
R9616 VDD.n4840 VDD.n4839 0.150167
R9617 VDD.n4870 VDD.n4869 0.150167
R9618 VDD.n4900 VDD.n4899 0.150167
R9619 VDD.n4930 VDD.n4929 0.150167
R9620 VDD.n3834 VDD.n3833 0.150167
R9621 VDD.n5007 VDD.n5006 0.150167
R9622 VDD.n5132 VDD.n5131 0.150167
R9623 VDD.n5073 VDD.n5072 0.150167
R9624 VDD.n4371 VDD.n4370 0.150167
R9625 VDD.n4465 VDD.n4464 0.150167
R9626 VDD.n4535 VDD.n4534 0.150167
R9627 VDD.n3674 VDD.n3673 0.150167
R9628 VDD.n3420 VDD 0.145785
R9629 VDD.n2564 VDD 0.145785
R9630 VDD.n1710 VDD 0.145785
R9631 VDD.n855 VDD 0.145785
R9632 VDD.n4654 VDD.n4647 0.144522
R9633 VDD.n4643 VDD.n4636 0.144522
R9634 VDD.n4776 VDD.n4773 0.144522
R9635 VDD.n4769 VDD.n4766 0.144522
R9636 VDD.n4756 VDD.n4754 0.144522
R9637 VDD.n4749 VDD.n4747 0.144522
R9638 VDD.n4742 VDD.n4740 0.144522
R9639 VDD.n4735 VDD.n4733 0.144522
R9640 VDD.n4728 VDD.n4726 0.144522
R9641 VDD.n5117 VDD.n5114 0.144522
R9642 VDD.n5110 VDD.n5107 0.144522
R9643 VDD.n5097 VDD.n5095 0.144522
R9644 VDD.n5090 VDD.n5088 0.144522
R9645 VDD.n5083 VDD.n5081 0.144522
R9646 VDD.n5076 VDD.n5074 0.144522
R9647 VDD.n5069 VDD.n5067 0.144522
R9648 VDD.n5186 VDD.n5179 0.144522
R9649 VDD.n5175 VDD.n5168 0.144522
R9650 VDD.n4468 VDD.n4466 0.144522
R9651 VDD.n4461 VDD.n4459 0.144522
R9652 VDD.n4538 VDD.n4536 0.144522
R9653 VDD.n4531 VDD.n4529 0.144522
R9654 VDD.n4374 VDD.n4372 0.144522
R9655 VDD.n4367 VDD.n4365 0.144522
R9656 VDD.n3677 VDD.n3675 0.144522
R9657 VDD.n3670 VDD.n3668 0.144522
R9658 VDD.n5302 VDD.n5300 0.144522
R9659 VDD.n5291 VDD.n5289 0.144522
R9660 VDD.n8629 VDD.n8622 0.144522
R9661 VDD.n8991 VDD.n8984 0.144522
R9662 VDD.n8901 VDD.n8894 0.144522
R9663 VDD.n3663 VDD.n3661 0.141804
R9664 VDD.n4685 VDD.n4684 0.138912
R9665 VDD.n4739 VDD.n4738 0.138912
R9666 VDD.n5026 VDD.n5025 0.138912
R9667 VDD.n5080 VDD.n5079 0.138912
R9668 VDD.n7074 VDD.n7073 0.13595
R9669 VDD.n7069 VDD.n7068 0.13595
R9670 VDD.n6986 VDD.n6985 0.13595
R9671 VDD.n6981 VDD.n6980 0.13595
R9672 VDD.n6898 VDD.n6897 0.13595
R9673 VDD.n6893 VDD.n6892 0.13595
R9674 VDD.n5469 VDD.n5468 0.13595
R9675 VDD.n5474 VDD.n5473 0.13595
R9676 VDD.n5557 VDD.n5556 0.13595
R9677 VDD.n5562 VDD.n5561 0.13595
R9678 VDD.n5645 VDD.n5644 0.13595
R9679 VDD.n5650 VDD.n5649 0.13595
R9680 VDD.n5733 VDD.n5732 0.13595
R9681 VDD.n5738 VDD.n5737 0.13595
R9682 VDD.n5821 VDD.n5820 0.13595
R9683 VDD.n5826 VDD.n5825 0.13595
R9684 VDD.n3013 VDD.n2633 0.134558
R9685 VDD.n1782 VDD.n1781 0.134558
R9686 VDD.n928 VDD.n927 0.134558
R9687 VDD.n73 VDD.n72 0.134558
R9688 VDD.n4242 VDD.n4109 0.132757
R9689 VDD.n6823 VDD.n6822 0.128928
R9690 VDD.n6740 VDD.n6739 0.128928
R9691 VDD.n6644 VDD.n6643 0.128928
R9692 VDD.n6560 VDD.n6559 0.128928
R9693 VDD.n4775 VDD.n4774 0.127599
R9694 VDD.n4746 VDD.n4745 0.127599
R9695 VDD.n5116 VDD.n5115 0.127599
R9696 VDD.n5087 VDD.n5086 0.127599
R9697 VDD.n9027 VDD.n9026 0.1274
R9698 VDD.n7536 VDD.n7535 0.12599
R9699 VDD.n7530 VDD.n7529 0.12599
R9700 VDD.n9028 VDD.n9027 0.122353
R9701 VDD.n9029 VDD.n9028 0.119879
R9702 VDD.n5435 VDD.n5434 0.117099
R9703 VDD.n4768 VDD.n4767 0.116231
R9704 VDD.n4753 VDD.n4752 0.116231
R9705 VDD.n5109 VDD.n5108 0.116231
R9706 VDD.n5094 VDD.n5093 0.116231
R9707 VDD.n3422 VDD 0.116103
R9708 VDD.n3423 VDD 0.116103
R9709 VDD.n5395 VDD.n5394 0.110519
R9710 VDD.n4607 VDD.n4606 0.109875
R9711 VDD.n4588 VDD.n4587 0.109094
R9712 VDD.n8044 VDD.n8033 0.108934
R9713 VDD.n8033 VDD.n8025 0.108934
R9714 VDD.n8025 VDD.n8017 0.108934
R9715 VDD.n8017 VDD.n8009 0.108934
R9716 VDD.n8009 VDD.n8001 0.108934
R9717 VDD.n8001 VDD.n7993 0.108934
R9718 VDD.n7993 VDD.n7985 0.108934
R9719 VDD.n7985 VDD.n7977 0.108934
R9720 VDD.n7977 VDD.n7966 0.108934
R9721 VDD.n7966 VDD.n7958 0.108934
R9722 VDD.n7958 VDD.n7947 0.108934
R9723 VDD.n7947 VDD.n7939 0.108934
R9724 VDD.n7939 VDD.n7931 0.108934
R9725 VDD.n7931 VDD.n7923 0.108934
R9726 VDD.n7923 VDD.n7915 0.108934
R9727 VDD.n7915 VDD.n7907 0.108934
R9728 VDD.n7907 VDD.n7899 0.108934
R9729 VDD.n7899 VDD.n7891 0.108934
R9730 VDD.n7891 VDD.n7883 0.108934
R9731 VDD.n7883 VDD.n7875 0.108934
R9732 VDD.n7875 VDD.n7867 0.108934
R9733 VDD.n7867 VDD.n7859 0.108934
R9734 VDD.n7859 VDD.n7851 0.108934
R9735 VDD.n7851 VDD.n7843 0.108934
R9736 VDD.n7843 VDD.n7835 0.108934
R9737 VDD.n7835 VDD.n7825 0.108934
R9738 VDD.n7825 VDD.n7819 0.108934
R9739 VDD.n7819 VDD.n7811 0.108934
R9740 VDD.n7811 VDD.n7805 0.108934
R9741 VDD.n7805 VDD.n7799 0.108934
R9742 VDD.n7799 VDD.n7791 0.108934
R9743 VDD.n7791 VDD.n7783 0.108934
R9744 VDD.n7783 VDD.n7775 0.108934
R9745 VDD.n7775 VDD.n7767 0.108934
R9746 VDD.n7767 VDD.n7759 0.108934
R9747 VDD.n7759 VDD.n7751 0.108934
R9748 VDD.n7751 VDD.n7743 0.108934
R9749 VDD.n7743 VDD.n7735 0.108934
R9750 VDD.n7735 VDD.n7727 0.108934
R9751 VDD.n7727 VDD.n7719 0.108934
R9752 VDD.n7719 VDD.n7711 0.108934
R9753 VDD.n7711 VDD.n7703 0.108934
R9754 VDD.n7703 VDD.n7692 0.108934
R9755 VDD.n7692 VDD.n7684 0.108934
R9756 VDD.n7684 VDD.n7673 0.108934
R9757 VDD.n7673 VDD.n7665 0.108934
R9758 VDD.n7665 VDD.n7657 0.108934
R9759 VDD.n7657 VDD.n7649 0.108934
R9760 VDD.n7649 VDD.n7641 0.108934
R9761 VDD.n7641 VDD.n7636 0.108934
R9762 VDD.n7636 VDD.n7601 0.108934
R9763 VDD.n7601 VDD.n7596 0.108934
R9764 VDD.n7596 VDD.n7591 0.108934
R9765 VDD.n7591 VDD.n7586 0.108934
R9766 VDD.n7586 VDD.n7581 0.108934
R9767 VDD.n7564 VDD.n7557 0.108934
R9768 VDD.n7557 VDD.n7552 0.108934
R9769 VDD.n7552 VDD.n7547 0.108934
R9770 VDD.n7547 VDD.n7542 0.108934
R9771 VDD.n7542 VDD.n7537 0.108934
R9772 VDD.n7537 VDD.n7531 0.108934
R9773 VDD.n7531 VDD.n7526 0.108934
R9774 VDD.n7526 VDD.n7521 0.108934
R9775 VDD.n7521 VDD.n7516 0.108934
R9776 VDD.n7516 VDD.n7511 0.108934
R9777 VDD.n7511 VDD.n7506 0.108934
R9778 VDD.n7506 VDD.n7502 0.108934
R9779 VDD.n7502 VDD.n7496 0.108934
R9780 VDD.n7496 VDD.n7492 0.108934
R9781 VDD.n7490 VDD.n7488 0.108934
R9782 VDD.n7488 VDD.n7486 0.108934
R9783 VDD.n7486 VDD.n7480 0.108934
R9784 VDD.n7480 VDD.n7476 0.108934
R9785 VDD.n7476 VDD.n7472 0.108934
R9786 VDD.n7472 VDD.n7468 0.108934
R9787 VDD.n7468 VDD.n7464 0.108934
R9788 VDD.n7464 VDD.n7460 0.108934
R9789 VDD.n7460 VDD.n7456 0.108934
R9790 VDD.n7456 VDD.n7452 0.108934
R9791 VDD.n7452 VDD.n7448 0.108934
R9792 VDD.n7448 VDD.n7445 0.108934
R9793 VDD.n7445 VDD.n7441 0.108934
R9794 VDD.n7441 VDD.n7437 0.108934
R9795 VDD.n7437 VDD.n7433 0.108934
R9796 VDD.n7433 VDD.n7429 0.108934
R9797 VDD.n7429 VDD.n7425 0.108934
R9798 VDD.n7425 VDD.n7421 0.108934
R9799 VDD.n7421 VDD.n7417 0.108934
R9800 VDD.n7417 VDD.n7411 0.108934
R9801 VDD.n7411 VDD.n7407 0.108934
R9802 VDD.n7407 VDD.n7403 0.108934
R9803 VDD.n7403 VDD.n7399 0.108934
R9804 VDD.n7399 VDD.n7395 0.108934
R9805 VDD.n7395 VDD.n7391 0.108934
R9806 VDD.n7391 VDD.n7387 0.108934
R9807 VDD.n7387 VDD.n7383 0.108934
R9808 VDD.n7383 VDD.n7379 0.108934
R9809 VDD.n7379 VDD.n7376 0.108934
R9810 VDD.n7376 VDD.n7372 0.108934
R9811 VDD.n7372 VDD.n7368 0.108934
R9812 VDD.n7368 VDD.n7364 0.108934
R9813 VDD.n7364 VDD.n7360 0.108934
R9814 VDD.n7360 VDD.n7356 0.108934
R9815 VDD.n7356 VDD.n7352 0.108934
R9816 VDD.n7352 VDD.n7348 0.108934
R9817 VDD.n7348 VDD.n7342 0.108934
R9818 VDD.n7342 VDD.n7337 0.108934
R9819 VDD.n7337 VDD.n7332 0.108934
R9820 VDD.n7332 VDD.n7327 0.108934
R9821 VDD.n7327 VDD.n7322 0.108934
R9822 VDD.n7322 VDD.n7317 0.108934
R9823 VDD.n7317 VDD.n7312 0.108934
R9824 VDD.n7312 VDD.n7307 0.108934
R9825 VDD.n7307 VDD.n7302 0.108934
R9826 VDD.n7302 VDD.n7298 0.108934
R9827 VDD.n7298 VDD.n7293 0.108934
R9828 VDD.n7293 VDD.n7288 0.108934
R9829 VDD.n7288 VDD.n7283 0.108934
R9830 VDD.n7283 VDD.n7278 0.108934
R9831 VDD.n7278 VDD.n7273 0.108934
R9832 VDD.n7273 VDD.n7268 0.108934
R9833 VDD.n7268 VDD.n7263 0.108934
R9834 VDD.n7263 VDD.n7255 0.108934
R9835 VDD.n7255 VDD.n7250 0.108934
R9836 VDD.n7250 VDD.n7245 0.108934
R9837 VDD.n7245 VDD.n7240 0.108934
R9838 VDD.n7240 VDD.n7235 0.108934
R9839 VDD.n7235 VDD.n7230 0.108934
R9840 VDD.n7230 VDD.n7225 0.108934
R9841 VDD.n7225 VDD.n7220 0.108934
R9842 VDD.n7220 VDD.n7215 0.108934
R9843 VDD.n7215 VDD.n7211 0.108934
R9844 VDD.n7211 VDD.n7206 0.108934
R9845 VDD.n7206 VDD.n7201 0.108934
R9846 VDD.n7201 VDD.n7196 0.108934
R9847 VDD.n7196 VDD.n7191 0.108934
R9848 VDD.n7191 VDD.n7186 0.108934
R9849 VDD.n7186 VDD.n7181 0.108934
R9850 VDD.n7181 VDD.n7176 0.108934
R9851 VDD.n7176 VDD.n7168 0.108934
R9852 VDD.n7168 VDD.n7163 0.108934
R9853 VDD.n7163 VDD.n7158 0.108934
R9854 VDD.n7158 VDD.n7153 0.108934
R9855 VDD.n7153 VDD.n7148 0.108934
R9856 VDD.n7148 VDD.n7143 0.108934
R9857 VDD.n7143 VDD.n7138 0.108934
R9858 VDD.n7138 VDD.n7133 0.108934
R9859 VDD.n7125 VDD.n7110 0.108934
R9860 VDD.n7110 VDD.n7105 0.108934
R9861 VDD.n7105 VDD.n7100 0.108934
R9862 VDD.n7100 VDD.n7095 0.108934
R9863 VDD.n7095 VDD.n7090 0.108934
R9864 VDD.n7090 VDD.n7085 0.108934
R9865 VDD.n7085 VDD.n7080 0.108934
R9866 VDD.n7080 VDD.n7075 0.108934
R9867 VDD.n7075 VDD.n7070 0.108934
R9868 VDD.n7070 VDD.n7065 0.108934
R9869 VDD.n7065 VDD.n7060 0.108934
R9870 VDD.n7060 VDD.n7055 0.108934
R9871 VDD.n7055 VDD.n7050 0.108934
R9872 VDD.n7050 VDD.n7045 0.108934
R9873 VDD.n7045 VDD.n7040 0.108934
R9874 VDD.n7040 VDD.n7035 0.108934
R9875 VDD.n7035 VDD.n7030 0.108934
R9876 VDD.n7030 VDD.n7022 0.108934
R9877 VDD.n7022 VDD.n7017 0.108934
R9878 VDD.n7017 VDD.n7012 0.108934
R9879 VDD.n7012 VDD.n7007 0.108934
R9880 VDD.n7007 VDD.n7002 0.108934
R9881 VDD.n7002 VDD.n6997 0.108934
R9882 VDD.n6997 VDD.n6992 0.108934
R9883 VDD.n6992 VDD.n6987 0.108934
R9884 VDD.n6987 VDD.n6982 0.108934
R9885 VDD.n6982 VDD.n6977 0.108934
R9886 VDD.n6977 VDD.n6972 0.108934
R9887 VDD.n6972 VDD.n6967 0.108934
R9888 VDD.n6967 VDD.n6962 0.108934
R9889 VDD.n6962 VDD.n6957 0.108934
R9890 VDD.n6957 VDD.n6952 0.108934
R9891 VDD.n6952 VDD.n6947 0.108934
R9892 VDD.n6947 VDD.n6942 0.108934
R9893 VDD.n6942 VDD.n6934 0.108934
R9894 VDD.n6934 VDD.n6929 0.108934
R9895 VDD.n6929 VDD.n6924 0.108934
R9896 VDD.n6924 VDD.n6919 0.108934
R9897 VDD.n6919 VDD.n6914 0.108934
R9898 VDD.n6914 VDD.n6909 0.108934
R9899 VDD.n6909 VDD.n6904 0.108934
R9900 VDD.n6904 VDD.n6899 0.108934
R9901 VDD.n6899 VDD.n6894 0.108934
R9902 VDD.n6894 VDD.n6889 0.108934
R9903 VDD.n6889 VDD.n6884 0.108934
R9904 VDD.n6884 VDD.n6879 0.108934
R9905 VDD.n6879 VDD.n6874 0.108934
R9906 VDD.n6874 VDD.n6869 0.108934
R9907 VDD.n6869 VDD.n6864 0.108934
R9908 VDD.n6864 VDD.n6859 0.108934
R9909 VDD.n6859 VDD.n6854 0.108934
R9910 VDD.n6854 VDD.n6846 0.108934
R9911 VDD.n6846 VDD.n6841 0.108934
R9912 VDD.n6841 VDD.n6836 0.108934
R9913 VDD.n6836 VDD.n6831 0.108934
R9914 VDD.n5460 VDD.n5455 0.108934
R9915 VDD.n5465 VDD.n5460 0.108934
R9916 VDD.n5470 VDD.n5465 0.108934
R9917 VDD.n5475 VDD.n5470 0.108934
R9918 VDD.n5480 VDD.n5475 0.108934
R9919 VDD.n5485 VDD.n5480 0.108934
R9920 VDD.n5490 VDD.n5485 0.108934
R9921 VDD.n5495 VDD.n5490 0.108934
R9922 VDD.n5500 VDD.n5495 0.108934
R9923 VDD.n5505 VDD.n5500 0.108934
R9924 VDD.n5510 VDD.n5505 0.108934
R9925 VDD.n5518 VDD.n5510 0.108934
R9926 VDD.n5523 VDD.n5518 0.108934
R9927 VDD.n5528 VDD.n5523 0.108934
R9928 VDD.n5533 VDD.n5528 0.108934
R9929 VDD.n5538 VDD.n5533 0.108934
R9930 VDD.n5543 VDD.n5538 0.108934
R9931 VDD.n5548 VDD.n5543 0.108934
R9932 VDD.n5553 VDD.n5548 0.108934
R9933 VDD.n5558 VDD.n5553 0.108934
R9934 VDD.n5563 VDD.n5558 0.108934
R9935 VDD.n5568 VDD.n5563 0.108934
R9936 VDD.n5573 VDD.n5568 0.108934
R9937 VDD.n5578 VDD.n5573 0.108934
R9938 VDD.n5583 VDD.n5578 0.108934
R9939 VDD.n5588 VDD.n5583 0.108934
R9940 VDD.n5593 VDD.n5588 0.108934
R9941 VDD.n5598 VDD.n5593 0.108934
R9942 VDD.n5606 VDD.n5598 0.108934
R9943 VDD.n5611 VDD.n5606 0.108934
R9944 VDD.n5616 VDD.n5611 0.108934
R9945 VDD.n5621 VDD.n5616 0.108934
R9946 VDD.n5626 VDD.n5621 0.108934
R9947 VDD.n5631 VDD.n5626 0.108934
R9948 VDD.n5636 VDD.n5631 0.108934
R9949 VDD.n5641 VDD.n5636 0.108934
R9950 VDD.n5646 VDD.n5641 0.108934
R9951 VDD.n5651 VDD.n5646 0.108934
R9952 VDD.n5656 VDD.n5651 0.108934
R9953 VDD.n5661 VDD.n5656 0.108934
R9954 VDD.n5666 VDD.n5661 0.108934
R9955 VDD.n5671 VDD.n5666 0.108934
R9956 VDD.n5676 VDD.n5671 0.108934
R9957 VDD.n5681 VDD.n5676 0.108934
R9958 VDD.n5686 VDD.n5681 0.108934
R9959 VDD.n5694 VDD.n5686 0.108934
R9960 VDD.n5699 VDD.n5694 0.108934
R9961 VDD.n5704 VDD.n5699 0.108934
R9962 VDD.n5709 VDD.n5704 0.108934
R9963 VDD.n5714 VDD.n5709 0.108934
R9964 VDD.n5719 VDD.n5714 0.108934
R9965 VDD.n5724 VDD.n5719 0.108934
R9966 VDD.n5729 VDD.n5724 0.108934
R9967 VDD.n5734 VDD.n5729 0.108934
R9968 VDD.n5739 VDD.n5734 0.108934
R9969 VDD.n5744 VDD.n5739 0.108934
R9970 VDD.n5749 VDD.n5744 0.108934
R9971 VDD.n5754 VDD.n5749 0.108934
R9972 VDD.n5759 VDD.n5754 0.108934
R9973 VDD.n5764 VDD.n5759 0.108934
R9974 VDD.n5769 VDD.n5764 0.108934
R9975 VDD.n5774 VDD.n5769 0.108934
R9976 VDD.n5782 VDD.n5774 0.108934
R9977 VDD.n5787 VDD.n5782 0.108934
R9978 VDD.n5792 VDD.n5787 0.108934
R9979 VDD.n5797 VDD.n5792 0.108934
R9980 VDD.n5802 VDD.n5797 0.108934
R9981 VDD.n5807 VDD.n5802 0.108934
R9982 VDD.n5812 VDD.n5807 0.108934
R9983 VDD.n5817 VDD.n5812 0.108934
R9984 VDD.n5822 VDD.n5817 0.108934
R9985 VDD.n5827 VDD.n5822 0.108934
R9986 VDD.n5832 VDD.n5827 0.108934
R9987 VDD.n6503 VDD.n6493 0.108934
R9988 VDD.n6493 VDD.n6488 0.108934
R9989 VDD.n6488 VDD.n6484 0.108934
R9990 VDD.n6484 VDD.n6479 0.108934
R9991 VDD.n6479 VDD.n6475 0.108934
R9992 VDD.n6475 VDD.n6470 0.108934
R9993 VDD.n6470 VDD.n6466 0.108934
R9994 VDD.n6466 VDD.n6459 0.108934
R9995 VDD.n6459 VDD.n6455 0.108934
R9996 VDD.n6455 VDD.n6450 0.108934
R9997 VDD.n6450 VDD.n6446 0.108934
R9998 VDD.n6446 VDD.n6441 0.108934
R9999 VDD.n6441 VDD.n6437 0.108934
R10000 VDD.n6437 VDD.n6432 0.108934
R10001 VDD.n6432 VDD.n6428 0.108934
R10002 VDD.n6428 VDD.n6423 0.108934
R10003 VDD.n6423 VDD.n6418 0.108934
R10004 VDD.n6418 VDD.n6414 0.108934
R10005 VDD.n6414 VDD.n6409 0.108934
R10006 VDD.n6409 VDD.n6405 0.108934
R10007 VDD.n6405 VDD.n6400 0.108934
R10008 VDD.n6400 VDD.n6396 0.108934
R10009 VDD.n6396 VDD.n6391 0.108934
R10010 VDD.n6391 VDD.n6387 0.108934
R10011 VDD.n6387 VDD.n6380 0.108934
R10012 VDD.n6380 VDD.n6376 0.108934
R10013 VDD.n6376 VDD.n6371 0.108934
R10014 VDD.n6371 VDD.n6366 0.108934
R10015 VDD.n6366 VDD.n6361 0.108934
R10016 VDD.n6361 VDD.n6356 0.108934
R10017 VDD.n6356 VDD.n6351 0.108934
R10018 VDD.n6351 VDD.n6346 0.108934
R10019 VDD.n6346 VDD.n6341 0.108934
R10020 VDD.n6341 VDD.n6336 0.108934
R10021 VDD.n6336 VDD.n6331 0.108934
R10022 VDD.n6331 VDD.n6326 0.108934
R10023 VDD.n6326 VDD.n6321 0.108934
R10024 VDD.n6321 VDD.n6316 0.108934
R10025 VDD.n6316 VDD.n6311 0.108934
R10026 VDD.n6311 VDD.n6306 0.108934
R10027 VDD.n6306 VDD.n6301 0.108934
R10028 VDD.n6301 VDD.n6293 0.108934
R10029 VDD.n6293 VDD.n6288 0.108934
R10030 VDD.n6288 VDD.n6283 0.108934
R10031 VDD.n6283 VDD.n6278 0.108934
R10032 VDD.n6278 VDD.n6273 0.108934
R10033 VDD.n6273 VDD.n6268 0.108934
R10034 VDD.n6268 VDD.n6263 0.108934
R10035 VDD.n6263 VDD.n6258 0.108934
R10036 VDD.n6258 VDD.n6253 0.108934
R10037 VDD.n6253 VDD.n6248 0.108934
R10038 VDD.n6248 VDD.n6243 0.108934
R10039 VDD.n6243 VDD.n6238 0.108934
R10040 VDD.n6238 VDD.n6233 0.108934
R10041 VDD.n6233 VDD.n6228 0.108934
R10042 VDD.n6228 VDD.n6223 0.108934
R10043 VDD.n6223 VDD.n6219 0.108934
R10044 VDD.n6219 VDD.n6215 0.108934
R10045 VDD.n6215 VDD.n6209 0.108934
R10046 VDD.n6209 VDD.n6205 0.108934
R10047 VDD.n6205 VDD.n6201 0.108934
R10048 VDD.n6201 VDD.n6197 0.108934
R10049 VDD.n6197 VDD.n6193 0.108934
R10050 VDD.n6193 VDD.n6189 0.108934
R10051 VDD.n6189 VDD.n6185 0.108934
R10052 VDD.n6185 VDD.n6181 0.108934
R10053 VDD.n6181 VDD.n6177 0.108934
R10054 VDD.n6177 VDD.n6173 0.108934
R10055 VDD.n6173 VDD.n6169 0.108934
R10056 VDD.n6169 VDD.n6165 0.108934
R10057 VDD.n6165 VDD.n6161 0.108934
R10058 VDD.n6161 VDD.n6157 0.108934
R10059 VDD.n6157 VDD.n6153 0.108934
R10060 VDD.n6153 VDD.n6149 0.108934
R10061 VDD.n6149 VDD.n6145 0.108934
R10062 VDD.n6145 VDD.n6139 0.108934
R10063 VDD.n6139 VDD.n6135 0.108934
R10064 VDD.n6135 VDD.n6131 0.108934
R10065 VDD.n6131 VDD.n6127 0.108934
R10066 VDD.n6127 VDD.n6123 0.108934
R10067 VDD.n6123 VDD.n6119 0.108934
R10068 VDD.n6119 VDD.n6115 0.108934
R10069 VDD.n6115 VDD.n6111 0.108934
R10070 VDD.n6111 VDD.n6107 0.108934
R10071 VDD.n6107 VDD.n6103 0.108934
R10072 VDD.n6103 VDD.n6099 0.108934
R10073 VDD.n6099 VDD.n6095 0.108934
R10074 VDD.n6095 VDD.n6091 0.108934
R10075 VDD.n6091 VDD.n6087 0.108934
R10076 VDD.n6087 VDD.n6083 0.108934
R10077 VDD.n6083 VDD.n6079 0.108934
R10078 VDD.n6079 VDD.n6075 0.108934
R10079 VDD.n6075 VDD.n6069 0.108934
R10080 VDD.n6069 VDD.n6065 0.108934
R10081 VDD.n6065 VDD.n6061 0.108934
R10082 VDD.n6061 VDD.n6057 0.108934
R10083 VDD.n6057 VDD.n6052 0.108934
R10084 VDD.n6052 VDD.n6047 0.108934
R10085 VDD.n6047 VDD.n6042 0.108934
R10086 VDD.n6042 VDD.n6037 0.108934
R10087 VDD.n6037 VDD.n6032 0.108934
R10088 VDD.n6032 VDD.n6027 0.108934
R10089 VDD.n6027 VDD.n6022 0.108934
R10090 VDD.n6022 VDD.n6017 0.108934
R10091 VDD.n6017 VDD.n6012 0.108934
R10092 VDD.n6012 VDD.n6007 0.108934
R10093 VDD.n6007 VDD.n6002 0.108934
R10094 VDD.n6002 VDD.n5997 0.108934
R10095 VDD.n5997 VDD.n5992 0.108934
R10096 VDD.n5992 VDD.n5984 0.108934
R10097 VDD.n5984 VDD.n5979 0.108934
R10098 VDD.n5979 VDD.n5974 0.108934
R10099 VDD.n5974 VDD.n5969 0.108934
R10100 VDD.n5969 VDD.n5964 0.108934
R10101 VDD.n5964 VDD.n5959 0.108934
R10102 VDD.n5959 VDD.n5954 0.108934
R10103 VDD.n5954 VDD.n5949 0.108934
R10104 VDD.n5949 VDD.n5944 0.108934
R10105 VDD.n5944 VDD.n5939 0.108934
R10106 VDD.n5939 VDD.n5934 0.108934
R10107 VDD.n5934 VDD.n5929 0.108934
R10108 VDD.n5929 VDD.n5924 0.108934
R10109 VDD.n5924 VDD.n5919 0.108934
R10110 VDD.n5919 VDD.n5914 0.108934
R10111 VDD.n5914 VDD.n5909 0.108934
R10112 VDD.n5909 VDD.n5904 0.108934
R10113 VDD.n5904 VDD.n5896 0.108934
R10114 VDD.n5896 VDD.n5891 0.108934
R10115 VDD.n5891 VDD.n5886 0.108934
R10116 VDD.n5886 VDD.n5881 0.108934
R10117 VDD.n5881 VDD.n5876 0.108934
R10118 VDD.n5876 VDD.n5871 0.108934
R10119 VDD.n5871 VDD.n5866 0.108934
R10120 VDD.n5866 VDD.n5861 0.108934
R10121 VDD.n5861 VDD.n5856 0.108934
R10122 VDD.n5856 VDD.n5851 0.108934
R10123 VDD.n5851 VDD.n5846 0.108934
R10124 VDD.n6825 VDD.n6824 0.108934
R10125 VDD.n6824 VDD.n6820 0.108934
R10126 VDD.n6820 VDD.n6816 0.108934
R10127 VDD.n6816 VDD.n6812 0.108934
R10128 VDD.n6812 VDD.n6808 0.108934
R10129 VDD.n6808 VDD.n6804 0.108934
R10130 VDD.n6804 VDD.n6799 0.108934
R10131 VDD.n6799 VDD.n6794 0.108934
R10132 VDD.n6794 VDD.n6786 0.108934
R10133 VDD.n6786 VDD.n6781 0.108934
R10134 VDD.n6781 VDD.n6776 0.108934
R10135 VDD.n6776 VDD.n6771 0.108934
R10136 VDD.n6771 VDD.n6766 0.108934
R10137 VDD.n6766 VDD.n6761 0.108934
R10138 VDD.n6761 VDD.n6756 0.108934
R10139 VDD.n6756 VDD.n6751 0.108934
R10140 VDD.n6751 VDD.n6746 0.108934
R10141 VDD.n6746 VDD.n6741 0.108934
R10142 VDD.n6741 VDD.n6736 0.108934
R10143 VDD.n6736 VDD.n6731 0.108934
R10144 VDD.n6731 VDD.n6726 0.108934
R10145 VDD.n6726 VDD.n6721 0.108934
R10146 VDD.n6721 VDD.n6716 0.108934
R10147 VDD.n6716 VDD.n6711 0.108934
R10148 VDD.n6711 VDD.n6706 0.108934
R10149 VDD.n6706 VDD.n6698 0.108934
R10150 VDD.n6698 VDD.n6694 0.108934
R10151 VDD.n6694 VDD.n6690 0.108934
R10152 VDD.n6690 VDD.n6686 0.108934
R10153 VDD.n6686 VDD.n6682 0.108934
R10154 VDD.n6682 VDD.n6678 0.108934
R10155 VDD.n6678 VDD.n6674 0.108934
R10156 VDD.n6674 VDD.n6653 0.108934
R10157 VDD.n6653 VDD.n6649 0.108934
R10158 VDD.n6649 VDD.n6645 0.108934
R10159 VDD.n6645 VDD.n6641 0.108934
R10160 VDD.n6641 VDD.n6637 0.108934
R10161 VDD.n6637 VDD.n6633 0.108934
R10162 VDD.n6633 VDD.n6629 0.108934
R10163 VDD.n6629 VDD.n6624 0.108934
R10164 VDD.n6624 VDD.n6619 0.108934
R10165 VDD.n6619 VDD.n6614 0.108934
R10166 VDD.n6614 VDD.n6606 0.108934
R10167 VDD.n6606 VDD.n6601 0.108934
R10168 VDD.n6601 VDD.n6596 0.108934
R10169 VDD.n6596 VDD.n6591 0.108934
R10170 VDD.n6591 VDD.n6586 0.108934
R10171 VDD.n6586 VDD.n6581 0.108934
R10172 VDD.n6581 VDD.n6576 0.108934
R10173 VDD.n6576 VDD.n6571 0.108934
R10174 VDD.n6571 VDD.n6566 0.108934
R10175 VDD.n6566 VDD.n6561 0.108934
R10176 VDD.n6561 VDD.n6556 0.108934
R10177 VDD.n6556 VDD.n6551 0.108934
R10178 VDD.n6551 VDD.n6546 0.108934
R10179 VDD.n6546 VDD.n6541 0.108934
R10180 VDD.n6541 VDD.n6536 0.108934
R10181 VDD.n6536 VDD.n6531 0.108934
R10182 VDD.n6531 VDD.n6526 0.108934
R10183 VDD.n6526 VDD.n6520 0.108934
R10184 VDD.n6520 VDD.n6516 0.108934
R10185 VDD.n6516 VDD.n6512 0.108934
R10186 VDD.n6512 VDD.n6508 0.108934
R10187 VDD.n6508 VDD.n6506 0.108934
R10188 VDD.n6506 VDD.n6505 0.108934
R10189 VDD.n6505 VDD.n6504 0.108934
R10190 VDD.n8066 VDD.n8058 0.108934
R10191 VDD.n8074 VDD.n8066 0.108934
R10192 VDD.n8082 VDD.n8074 0.108934
R10193 VDD.n8090 VDD.n8082 0.108934
R10194 VDD.n8098 VDD.n8090 0.108934
R10195 VDD.n8104 VDD.n8098 0.108934
R10196 VDD.n8112 VDD.n8104 0.108934
R10197 VDD.n8118 VDD.n8112 0.108934
R10198 VDD.n8126 VDD.n8118 0.108934
R10199 VDD.n8133 VDD.n8126 0.108934
R10200 VDD.n8142 VDD.n8133 0.108934
R10201 VDD.n8147 VDD.n8142 0.108934
R10202 VDD.n8153 VDD.n8147 0.108934
R10203 VDD.n8159 VDD.n8153 0.108934
R10204 VDD.n8165 VDD.n8159 0.108934
R10205 VDD.n8171 VDD.n8165 0.108934
R10206 VDD.n8177 VDD.n8171 0.108934
R10207 VDD.n8183 VDD.n8177 0.108934
R10208 VDD.n8191 VDD.n8183 0.108934
R10209 VDD.n8197 VDD.n8191 0.108934
R10210 VDD.n8205 VDD.n8197 0.108934
R10211 VDD.n8211 VDD.n8205 0.108934
R10212 VDD.n8217 VDD.n8211 0.108934
R10213 VDD.n8223 VDD.n8217 0.108934
R10214 VDD.n8229 VDD.n8223 0.108934
R10215 VDD.n8235 VDD.n8229 0.108934
R10216 VDD.n8241 VDD.n8235 0.108934
R10217 VDD.n8247 VDD.n8241 0.108934
R10218 VDD.n8252 VDD.n8247 0.108934
R10219 VDD.n8258 VDD.n8252 0.108934
R10220 VDD.n8264 VDD.n8258 0.108934
R10221 VDD.n8270 VDD.n8264 0.108934
R10222 VDD.n8276 VDD.n8270 0.108934
R10223 VDD.n8282 VDD.n8276 0.108934
R10224 VDD.n8288 VDD.n8282 0.108934
R10225 VDD.n8296 VDD.n8288 0.108934
R10226 VDD.n8302 VDD.n8296 0.108934
R10227 VDD.n8310 VDD.n8302 0.108934
R10228 VDD.n8316 VDD.n8310 0.108934
R10229 VDD.n8322 VDD.n8316 0.108934
R10230 VDD.n8328 VDD.n8322 0.108934
R10231 VDD.n8334 VDD.n8328 0.108934
R10232 VDD.n8340 VDD.n8334 0.108934
R10233 VDD.n8346 VDD.n8340 0.108934
R10234 VDD.n8352 VDD.n8346 0.108934
R10235 VDD.n8357 VDD.n8352 0.108934
R10236 VDD.n8363 VDD.n8357 0.108934
R10237 VDD.n8369 VDD.n8363 0.108934
R10238 VDD.n8375 VDD.n8369 0.108934
R10239 VDD.n8381 VDD.n8375 0.108934
R10240 VDD.n8387 VDD.n8381 0.108934
R10241 VDD.n8393 VDD.n8387 0.108934
R10242 VDD.n8401 VDD.n8393 0.108934
R10243 VDD.n8407 VDD.n8401 0.108934
R10244 VDD.n8419 VDD.n8407 0.108934
R10245 VDD.n8429 VDD.n8419 0.108934
R10246 VDD.n8439 VDD.n8429 0.108934
R10247 VDD.n8449 VDD.n8439 0.108934
R10248 VDD.n8459 VDD.n8449 0.108934
R10249 VDD.n8468 VDD.n8459 0.108934
R10250 VDD.n8477 VDD.n8468 0.108934
R10251 VDD.n8486 VDD.n8477 0.108934
R10252 VDD.n8494 VDD.n8486 0.108934
R10253 VDD.n8503 VDD.n8494 0.108934
R10254 VDD.n8512 VDD.n8503 0.108934
R10255 VDD.n8521 VDD.n8512 0.108934
R10256 VDD.n8529 VDD.n8521 0.108934
R10257 VDD.n8537 VDD.n8529 0.108934
R10258 VDD.n8543 VDD.n8537 0.108934
R10259 VDD.n8544 VDD.n8543 0.108934
R10260 VDD.n8545 VDD.n8544 0.108934
R10261 VDD.n3760 VDD.n3759 0.10877
R10262 VDD.n3382 VDD.n3374 0.107703
R10263 VDD.n1934 VDD.n1826 0.107703
R10264 VDD.n1080 VDD.n972 0.107703
R10265 VDD.n225 VDD.n117 0.107703
R10266 VDD.n4659 VDD.n4658 0.0995999
R10267 VDD.n4781 VDD.n4780 0.0995999
R10268 VDD.n5122 VDD.n5121 0.0995999
R10269 VDD.n5191 VDD.n5190 0.0995999
R10270 VDD.n4256 VDD.n4255 0.0980399
R10271 VDD.n8870 VDD.n8869 0.0932536
R10272 VDD.n2563 VDD.n2562 0.0926226
R10273 VDD.n1709 VDD.n1708 0.0926226
R10274 VDD.n854 VDD.n853 0.0926226
R10275 VDD.n45 VDD 0.0926053
R10276 VDD.n1754 VDD 0.0926053
R10277 VDD.n4251 VDD.n4250 0.0923441
R10278 VDD.n4075 VDD.n3952 0.0897616
R10279 VDD.n8952 VDD.n8951 0.0895625
R10280 VDD.n9030 VDD 0.0872245
R10281 VDD.n5251 VDD.n5250 0.0856562
R10282 VDD.n3865 VDD.n3864 0.0825312
R10283 VDD.n3862 VDD.n3861 0.0825312
R10284 VDD.n2564 VDD.n2563 0.0745132
R10285 VDD.n1710 VDD.n1709 0.0745132
R10286 VDD.n855 VDD.n854 0.0745132
R10287 VDD.n5221 VDD 0.0739375
R10288 VDD.n3857 VDD.n3847 0.0736942
R10289 VDD.n4274 VDD.n4271 0.0736373
R10290 VDD.n6427 VDD.n6426 0.0728164
R10291 VDD.n6345 VDD.n6344 0.0728164
R10292 VDD.n6257 VDD.n6256 0.0728164
R10293 VDD.n6180 VDD.n6179 0.0728164
R10294 VDD.n6110 VDD.n6109 0.0728164
R10295 VDD.n6036 VDD.n6035 0.0728164
R10296 VDD.n5948 VDD.n5947 0.0728164
R10297 VDD.n5860 VDD.n5859 0.0728164
R10298 VDD.n3626 VDD.n3625 0.071743
R10299 VDD.n4268 VDD.n4267 0.0711193
R10300 VDD.n4568 VDD.n4567 0.0707228
R10301 VDD.n4320 VDD.n4319 0.0707228
R10302 VDD.n4274 VDD.n4273 0.0703248
R10303 VDD.n7595 VDD.n7594 0.0696892
R10304 VDD.n4290 VDD.n4289 0.0692474
R10305 VDD.n3040 VDD.n3039 0.0688877
R10306 VDD.n2558 VDD.n2557 0.0688877
R10307 VDD.n1704 VDD.n1703 0.0688877
R10308 VDD.n849 VDD.n848 0.0688877
R10309 VDD.n8132 VDD.n8131 0.0682249
R10310 VDD.n8240 VDD.n8239 0.0682249
R10311 VDD.n8345 VDD.n8344 0.0682249
R10312 VDD.n8476 VDD.n8475 0.0682249
R10313 VDD.n5319 VDD.n5318 0.0679494
R10314 VDD.n8876 VDD 0.0645625
R10315 VDD.n3039 VDD.n3013 0.0643587
R10316 VDD.n2557 VDD.n1782 0.0643587
R10317 VDD.n1703 VDD.n928 0.0643587
R10318 VDD.n848 VDD.n73 0.0643587
R10319 VDD.n8043 VDD.n8039 0.0638663
R10320 VDD.n8032 VDD.n8031 0.0638663
R10321 VDD.n7898 VDD.n7894 0.0638663
R10322 VDD.n7890 VDD.n7889 0.0638663
R10323 VDD.n7766 VDD.n7762 0.0638663
R10324 VDD.n7758 VDD.n7757 0.0638663
R10325 VDD.n5227 VDD.n5226 0.0636644
R10326 VDD.n4832 VDD.n4826 0.0631347
R10327 VDD.n4922 VDD.n4916 0.0631347
R10328 VDD.n5217 VDD.n5208 0.0631347
R10329 VDD.n5143 VDD.n5135 0.0631347
R10330 VDD.n4892 VDD.n4886 0.0631347
R10331 VDD.n4677 VDD.n4668 0.0631347
R10332 VDD.n4800 VDD.n4794 0.0631347
R10333 VDD.n4862 VDD.n4856 0.0627929
R10334 VDD.n4952 VDD.n4946 0.0627929
R10335 VDD.n8640 VDD.n8639 0.0608156
R10336 VDD.n46 VDD 0.060807
R10337 VDD.n1755 VDD 0.060807
R10338 VDD.n4492 VDD.n4487 0.0604712
R10339 VDD.n4399 VDD.n4394 0.0604712
R10340 VDD.n4314 VDD.n4306 0.0604712
R10341 VDD.n3701 VDD.n3696 0.0604712
R10342 VDD.n9031 VDD 0.0596514
R10343 VDD.n4405 VDD.n4404 0.0595872
R10344 VDD.n8927 VDD.n8919 0.0595049
R10345 VDD.n8696 VDD.n8692 0.0591683
R10346 VDD.n4498 VDD.n4497 0.0591603
R10347 VDD.n3707 VDD.n3706 0.0591603
R10348 VDD.n8872 VDD.n8818 0.0589865
R10349 VDD.n5343 VDD.n5335 0.0586853
R10350 VDD.n3845 VDD.n3837 0.0581563
R10351 VDD.n26 VDD.n25 0.056838
R10352 VDD.n27 VDD.n26 0.056838
R10353 VDD.n27 VDD.n4 0.056838
R10354 VDD.n63 VDD.n4 0.056838
R10355 VDD.n874 VDD.n866 0.056838
R10356 VDD.n885 VDD.n866 0.056838
R10357 VDD.n887 VDD.n885 0.056838
R10358 VDD.n887 VDD.n886 0.056838
R10359 VDD.n1735 VDD.n1734 0.056838
R10360 VDD.n1736 VDD.n1735 0.056838
R10361 VDD.n1736 VDD.n1713 0.056838
R10362 VDD.n1772 VDD.n1713 0.056838
R10363 VDD.n2567 VDD.n2566 0.056838
R10364 VDD.n2568 VDD.n2567 0.056838
R10365 VDD.n2569 VDD.n2568 0.056838
R10366 VDD.n2600 VDD.n2569 0.056838
R10367 VDD VDD.n8875 0.05675
R10368 VDD.n3765 VDD.n3764 0.0566413
R10369 VDD.n4665 VDD.n4664 0.0565323
R10370 VDD.n4787 VDD.n4786 0.0565323
R10371 VDD.n4823 VDD.n4822 0.0565323
R10372 VDD.n4853 VDD.n4852 0.0565323
R10373 VDD.n4883 VDD.n4882 0.0565323
R10374 VDD.n4913 VDD.n4912 0.0565323
R10375 VDD.n4943 VDD.n4942 0.0565323
R10376 VDD.n5003 VDD.n5002 0.0565323
R10377 VDD.n5128 VDD.n5127 0.0565323
R10378 VDD.n5205 VDD.n5204 0.0565323
R10379 VDD.n3750 VDD.n3749 0.0561943
R10380 VDD.n5349 VDD.n5348 0.0558794
R10381 VDD.n8634 VDD.n8633 0.0547109
R10382 VDD.n8996 VDD.n8995 0.0547109
R10383 VDD.n8906 VDD.n8905 0.0547109
R10384 VDD VDD.n3421 0.0526991
R10385 VDD.n4251 VDD.n4247 0.0521995
R10386 VDD.n4075 VDD.n4074 0.0521189
R10387 VDD VDD.n1711 0.0517913
R10388 VDD.n8546 VDD.n8545 0.0517048
R10389 VDD.n3948 VDD.n3947 0.0513458
R10390 VDD.n3902 VDD.n3901 0.0493281
R10391 VDD.n4664 VDD.n4663 0.0487198
R10392 VDD.n4786 VDD.n4785 0.0487198
R10393 VDD.n4822 VDD.n4821 0.0487198
R10394 VDD.n4852 VDD.n4851 0.0487198
R10395 VDD.n4882 VDD.n4881 0.0487198
R10396 VDD.n4912 VDD.n4911 0.0487198
R10397 VDD.n4942 VDD.n4941 0.0487198
R10398 VDD.n5127 VDD.n5126 0.0487198
R10399 VDD.n5204 VDD.n5203 0.0487198
R10400 VDD VDD.n856 0.0482611
R10401 VDD VDD.n2565 0.0482611
R10402 VDD.n3845 VDD.n3844 0.0479088
R10403 VDD.n5421 VDD.n5420 0.0472468
R10404 VDD.n9012 VDD.n9001 0.0462851
R10405 VDD.n22 VDD.n17 0.0461081
R10406 VDD.n875 VDD.n871 0.0461081
R10407 VDD.n1731 VDD.n1726 0.0461081
R10408 VDD.n2578 VDD.n2577 0.0461081
R10409 VDD.n4562 VDD.n4557 0.0459877
R10410 VDD.n8669 VDD.n8651 0.0459833
R10411 VDD.n8948 VDD.n8930 0.0459833
R10412 VDD.n3744 VDD.n3739 0.0457021
R10413 VDD.n8713 VDD.n8699 0.0456006
R10414 VDD.n8748 VDD.n8730 0.0455549
R10415 VDD.n8748 VDD.n8747 0.0454465
R10416 VDD.n3939 VDD.n3875 0.0454219
R10417 VDD.n3872 VDD.n3871 0.0454219
R10418 VDD.n3868 VDD.n3867 0.0454219
R10419 VDD.n8713 VDD.n8712 0.0454042
R10420 VDD.n3739 VDD.n3738 0.0453096
R10421 VDD.n4557 VDD.n4556 0.045025
R10422 VDD.n8669 VDD.n8668 0.0450203
R10423 VDD.n8948 VDD.n8947 0.0450203
R10424 VDD.n5011 VDD.n5010 0.0448136
R10425 VDD.n9012 VDD.n9011 0.0447244
R10426 VDD.n8815 VDD.n8814 0.044241
R10427 VDD.n4636 VDD.n4634 0.0439783
R10428 VDD.n4766 VDD.n4764 0.0439783
R10429 VDD.n4758 VDD.n4756 0.0439783
R10430 VDD.n5107 VDD.n5105 0.0439783
R10431 VDD.n5099 VDD.n5097 0.0439783
R10432 VDD.n5168 VDD.n5166 0.0439783
R10433 VDD.n4289 VDD.n4287 0.0439783
R10434 VDD.n5318 VDD.n5316 0.0439783
R10435 VDD.n8622 VDD.n8620 0.0439783
R10436 VDD.n8984 VDD.n8982 0.0439783
R10437 VDD.n8894 VDD.n8892 0.0439783
R10438 VDD.n8818 VDD.n8815 0.0439172
R10439 VDD.n23 VDD.n12 0.0435743
R10440 VDD.n872 VDD.n867 0.0435743
R10441 VDD.n1732 VDD.n1721 0.0435743
R10442 VDD.n2584 VDD.n2583 0.0435743
R10443 VDD.n3714 VDD.n3713 0.0434688
R10444 VDD.n3715 VDD.n3714 0.0434688
R10445 VDD.n3716 VDD.n3715 0.0434688
R10446 VDD.n3719 VDD.n3718 0.0434688
R10447 VDD.n3720 VDD.n3719 0.0434688
R10448 VDD.n3721 VDD.n3720 0.0434688
R10449 VDD.n3722 VDD.n3721 0.0434688
R10450 VDD.n5361 VDD.n5360 0.0434688
R10451 VDD.n5360 VDD.n5359 0.0434688
R10452 VDD.n5359 VDD.n5358 0.0434688
R10453 VDD.n5356 VDD.n5355 0.0434688
R10454 VDD.n5355 VDD.n5354 0.0434688
R10455 VDD.n5354 VDD.n5353 0.0434688
R10456 VDD.n8719 VDD.n8718 0.0434688
R10457 VDD.n8720 VDD.n8719 0.0434688
R10458 VDD.n8721 VDD.n8720 0.0434688
R10459 VDD.n8722 VDD.n8721 0.0434688
R10460 VDD.n8725 VDD.n8724 0.0434688
R10461 VDD.n8726 VDD.n8725 0.0434688
R10462 VDD.n8727 VDD.n8726 0.0434688
R10463 VDD.n9017 VDD.n8727 0.0434688
R10464 VDD.n9017 VDD.n9016 0.0434688
R10465 VDD.n8960 VDD.n8959 0.0434688
R10466 VDD.n8959 VDD.n8958 0.0434688
R10467 VDD.n8958 VDD.n8957 0.0434688
R10468 VDD.n8955 VDD.n8954 0.0434688
R10469 VDD.n8954 VDD.n8953 0.0434688
R10470 VDD.n3920 VDD.n3919 0.0434688
R10471 VDD.n3869 VDD.n3868 0.0434688
R10472 VDD.n4958 VDD.n4957 0.0434688
R10473 VDD.n4959 VDD.n4958 0.0434688
R10474 VDD.n4960 VDD.n4959 0.0434688
R10475 VDD.n4961 VDD.n4960 0.0434688
R10476 VDD.n4964 VDD.n4963 0.0434688
R10477 VDD.n4965 VDD.n4964 0.0434688
R10478 VDD.n4966 VDD.n4965 0.0434688
R10479 VDD.n4967 VDD.n4966 0.0434688
R10480 VDD.n4968 VDD.n4967 0.0434688
R10481 VDD.n4977 VDD.n4974 0.0434688
R10482 VDD.n4977 VDD.n4976 0.0434688
R10483 VDD.n4976 VDD.n4975 0.0434688
R10484 VDD.n3822 VDD.n3821 0.0434688
R10485 VDD.n3823 VDD.n3822 0.0434688
R10486 VDD.n4988 VDD.n3823 0.0434688
R10487 VDD.n4989 VDD.n4988 0.0434688
R10488 VDD.n4990 VDD.n4989 0.0434688
R10489 VDD.n4991 VDD.n4990 0.0434688
R10490 VDD.n4992 VDD.n4991 0.0434688
R10491 VDD.n4993 VDD.n4992 0.0434688
R10492 VDD.n4994 VDD.n4993 0.0434688
R10493 VDD.n4995 VDD.n4994 0.0434688
R10494 VDD.n3600 VDD.n3599 0.0433094
R10495 VDD.n6745 VDD.n6744 0.0433094
R10496 VDD.n6648 VDD.n6647 0.0433094
R10497 VDD.n6565 VDD.n6564 0.0433094
R10498 VDD.n4862 VDD.n4861 0.0430273
R10499 VDD.n4952 VDD.n4951 0.0430273
R10500 VDD.n4549 VDD.n4545 0.0429751
R10501 VDD.n4386 VDD.n4382 0.0429751
R10502 VDD.n8635 VDD.n8634 0.042958
R10503 VDD.n8687 VDD.n8684 0.042958
R10504 VDD.n8997 VDD.n8996 0.042958
R10505 VDD.n8914 VDD.n8906 0.042958
R10506 VDD.n5003 VDD.n5000 0.0428604
R10507 VDD.n4677 VDD.n4676 0.0426869
R10508 VDD.n4800 VDD.n4799 0.0426869
R10509 VDD.n4832 VDD.n4831 0.0426869
R10510 VDD.n4892 VDD.n4891 0.0426869
R10511 VDD.n4922 VDD.n4921 0.0426869
R10512 VDD.n5143 VDD.n5142 0.0426869
R10513 VDD.n5217 VDD.n5216 0.0426869
R10514 VDD.n4323 VDD.n4322 0.0420568
R10515 VDD.n4408 VDD.n4407 0.0420568
R10516 VDD.n4501 VDD.n4500 0.0420568
R10517 VDD.n3643 VDD.n3642 0.0420568
R10518 VDD.n3925 VDD.n3921 0.0415156
R10519 VDD.n3914 VDD.n3913 0.0415156
R10520 VDD.n3871 VDD.n3870 0.0415156
R10521 VDD.n4699 VDD.n4697 0.0412609
R10522 VDD.n4715 VDD.n4713 0.0412609
R10523 VDD.n5040 VDD.n5038 0.0412609
R10524 VDD.n5056 VDD.n5054 0.0412609
R10525 VDD.n4337 VDD.n4335 0.0412609
R10526 VDD.n4353 VDD.n4351 0.0412609
R10527 VDD.n4420 VDD.n4418 0.0412609
R10528 VDD.n4448 VDD.n4446 0.0412609
R10529 VDD.n4427 VDD.n4425 0.0412609
R10530 VDD.n4518 VDD.n4516 0.0412609
R10531 VDD.n3657 VDD.n3655 0.0412609
R10532 VDD.n5274 VDD.n5272 0.0412609
R10533 VDD VDD.n917 0.0412609
R10534 VDD VDD.n2626 0.0412609
R10535 VDD.n3717 VDD.n3716 0.041125
R10536 VDD.n8956 VDD.n8955 0.041125
R10537 VDD VDD.n5220 0.041125
R10538 VDD.n3723 VDD.n3722 0.0403437
R10539 VDD.n8961 VDD.n8960 0.0403437
R10540 VDD.n4974 VDD.n4973 0.0403437
R10541 VDD.n3731 VDD.n3727 0.0398734
R10542 VDD.n3873 VDD.n3872 0.0395625
R10543 VDD.n4647 VDD.n4645 0.0385435
R10544 VDD.n4773 VDD.n4771 0.0385435
R10545 VDD.n4751 VDD.n4749 0.0385435
R10546 VDD.n5114 VDD.n5112 0.0385435
R10547 VDD.n5092 VDD.n5090 0.0385435
R10548 VDD.n5179 VDD.n5177 0.0385435
R10549 VDD.n8633 VDD.n8631 0.0385435
R10550 VDD.n8995 VDD.n8993 0.0385435
R10551 VDD.n8905 VDD.n8903 0.0385435
R10552 VDD.n29 VDD.n12 0.0385068
R10553 VDD.n62 VDD 0.0385068
R10554 VDD.n6 VDD 0.0385068
R10555 VDD.n883 VDD.n867 0.0385068
R10556 VDD VDD.n864 0.0385068
R10557 VDD.n892 VDD 0.0385068
R10558 VDD.n1738 VDD.n1721 0.0385068
R10559 VDD.n1771 VDD 0.0385068
R10560 VDD.n1715 VDD 0.0385068
R10561 VDD.n2588 VDD.n2584 0.0385068
R10562 VDD.n2599 VDD 0.0385068
R10563 VDD.n2572 VDD 0.0385068
R10564 VDD.n8814 VDD.n8811 0.0380981
R10565 VDD.n8654 VDD.n8653 0.0380882
R10566 VDD.n8702 VDD.n8701 0.0380882
R10567 VDD.n8733 VDD.n8732 0.0380882
R10568 VDD.n8933 VDD.n8932 0.0380882
R10569 VDD.n4957 VDD.n4956 0.038
R10570 VDD.n4996 VDD.n4995 0.038
R10571 VDD.n3935 VDD.n3931 0.0376094
R10572 VDD.n3875 VDD.n3874 0.0376094
R10573 VDD.n3419 VDD.n3417 0.0364779
R10574 VDD.n922 VDD.n1 0.0358522
R10575 VDD.n3930 VDD.n3929 0.0356562
R10576 VDD.n3760 VDD.n3756 0.035222
R10577 VDD.n5349 VDD.n5306 0.0351381
R10578 VDD.n8811 VDD.n8810 0.0345604
R10579 VDD.n48 VDD.n47 0.0343645
R10580 VDD.n1757 VDD.n1756 0.0343645
R10581 VDD.n9027 VDD.n8578 0.034112
R10582 VDD.n5245 VDD.n5244 0.0338623
R10583 VDD.n3916 VDD.n3915 0.0337031
R10584 VDD.n3867 VDD.n3866 0.0337031
R10585 VDD.n67 VDD.n2 0.033419
R10586 VDD.n1776 VDD.n0 0.033419
R10587 VDD.n4658 VDD.n4656 0.0331087
R10588 VDD.n4780 VDD.n4778 0.0331087
R10589 VDD.n4744 VDD.n4742 0.0331087
R10590 VDD.n5121 VDD.n5119 0.0331087
R10591 VDD.n5085 VDD.n5083 0.0331087
R10592 VDD.n5190 VDD.n5188 0.0331087
R10593 VDD.n5011 VDD.n5004 0.0330948
R10594 VDD.n3857 VDD.n3856 0.0322427
R10595 VDD.n5335 VDD.n5334 0.0319008
R10596 VDD.n3940 VDD.n3939 0.03175
R10597 VDD.n8692 VDD.n8691 0.0314198
R10598 VDD.n4498 VDD.n4472 0.0312849
R10599 VDD.n3707 VDD.n3681 0.0312849
R10600 VDD.n5327 VDD.n5319 0.0311134
R10601 VDD.n8919 VDD.n8918 0.0310804
R10602 VDD.n4405 VDD.n4378 0.0308558
R10603 VDD.n4726 VDD.n4723 0.0303913
R10604 VDD.n5067 VDD.n5064 0.0303913
R10605 VDD.n4459 VDD.n4456 0.0303913
R10606 VDD.n4529 VDD.n4526 0.0303913
R10607 VDD.n4365 VDD.n4362 0.0303913
R10608 VDD.n3668 VDD.n3665 0.0303913
R10609 VDD.n5289 VDD.n5282 0.0303913
R10610 VDD.n4397 VDD.n4396 0.0303633
R10611 VDD.n4490 VDD.n4489 0.0303633
R10612 VDD.n4560 VDD.n4559 0.0303633
R10613 VDD.n3699 VDD.n3698 0.0303633
R10614 VDD.n3742 VDD.n3741 0.0303633
R10615 VDD.n3713 VDD.n3712 0.0301875
R10616 VDD.n8718 VDD.n8717 0.0301875
R10617 VDD.n8953 VDD.n8952 0.0301875
R10618 VDD.n4394 VDD.n4393 0.0301368
R10619 VDD.n4306 VDD.n4305 0.0301368
R10620 VDD.n4487 VDD.n4486 0.0301368
R10621 VDD.n3696 VDD.n3695 0.0301368
R10622 VDD.n8753 VDD.n8752 0.0299811
R10623 VDD.n8768 VDD.n8767 0.0299811
R10624 VDD.n8658 VDD.n8657 0.0297969
R10625 VDD.n8706 VDD.n8705 0.0297969
R10626 VDD.n8737 VDD.n8736 0.0297969
R10627 VDD.n8937 VDD.n8936 0.0297969
R10628 VDD.n3901 VDD.n3899 0.0297969
R10629 VDD.n8648 VDD.n8640 0.0297952
R10630 VDD.n4479 VDD.n4475 0.0291557
R10631 VDD.n4298 VDD.n4290 0.0291557
R10632 VDD.n3688 VDD.n3684 0.0291557
R10633 VDD.n8795 VDD.n8794 0.0288019
R10634 VDD.n8770 VDD.n8769 0.0288019
R10635 VDD.n8776 VDD.n8775 0.0288019
R10636 VDD.n3421 VDD.n3419 0.0285752
R10637 VDD.n8872 VDD.n8871 0.0282045
R10638 VDD VDD.n3 0.0281786
R10639 VDD.n919 VDD 0.0281786
R10640 VDD VDD.n1712 0.0281786
R10641 VDD.n2628 VDD 0.0281786
R10642 VDD.n1711 VDD.n1 0.028087
R10643 VDD.n4660 VDD.n4659 0.0278438
R10644 VDD.n4782 VDD.n4781 0.0278438
R10645 VDD.n4815 VDD.n4814 0.0278438
R10646 VDD.n4848 VDD.n4847 0.0278438
R10647 VDD.n4878 VDD.n4877 0.0278438
R10648 VDD.n4908 VDD.n4907 0.0278438
R10649 VDD.n4938 VDD.n4937 0.0278438
R10650 VDD.n5123 VDD.n5122 0.0278438
R10651 VDD.n5192 VDD.n5191 0.0278438
R10652 VDD.n4737 VDD.n4735 0.0276739
R10653 VDD.n5078 VDD.n5076 0.0276739
R10654 VDD.n8778 VDD.n8777 0.0276226
R10655 VDD.n28 VDD.n16 0.027527
R10656 VDD.n16 VDD.n15 0.027527
R10657 VDD.n884 VDD.n865 0.027527
R10658 VDD.n888 VDD.n865 0.027527
R10659 VDD.n1737 VDD.n1725 0.027527
R10660 VDD.n1725 VDD.n1724 0.027527
R10661 VDD.n2590 VDD.n2589 0.027527
R10662 VDD.n2591 VDD.n2590 0.027527
R10663 VDD.n5449 VDD.n5448 0.0273817
R10664 VDD.n5450 VDD.n5447 0.0273817
R10665 VDD.n8723 VDD.n8722 0.0270625
R10666 VDD.n8791 VDD.n8790 0.0264434
R10667 VDD.n8789 VDD.n8778 0.0264434
R10668 VDD.n856 VDD.n2 0.0261883
R10669 VDD.n2565 VDD.n0 0.0261883
R10670 VDD.n3938 VDD.n3937 0.0258906
R10671 VDD.n3910 VDD.n3908 0.0258906
R10672 VDD.n3907 VDD.n3903 0.0258906
R10673 VDD.n3903 VDD.n3902 0.0258906
R10674 VDD.n3864 VDD.n3863 0.0258906
R10675 VDD.n3863 VDD.n3862 0.0258906
R10676 VDD.n8790 VDD.n8756 0.0252642
R10677 VDD.n8789 VDD.n8770 0.0252642
R10678 VDD.n4733 VDD.n4730 0.0249565
R10679 VDD.n5074 VDD.n5071 0.0249565
R10680 VDD.n4471 VDD.n4470 0.0249565
R10681 VDD.n4466 VDD.n4463 0.0249565
R10682 VDD.n4541 VDD.n4540 0.0249565
R10683 VDD.n4536 VDD.n4533 0.0249565
R10684 VDD.n4377 VDD.n4376 0.0249565
R10685 VDD.n4372 VDD.n4369 0.0249565
R10686 VDD.n3680 VDD.n3679 0.0249565
R10687 VDD.n3675 VDD.n3672 0.0249565
R10688 VDD.n5305 VDD.n5304 0.0249565
R10689 VDD.n5300 VDD.n5293 0.0249565
R10690 VDD.n4963 VDD.n4962 0.0247187
R10691 VDD.n62 VDD.n5 0.024466
R10692 VDD.n890 VDD.n864 0.024466
R10693 VDD.n1771 VDD.n1714 0.024466
R10694 VDD.n2599 VDD.n2570 0.024466
R10695 VDD.n4497 VDD.n4494 0.0239375
R10696 VDD.n4567 VDD.n4564 0.0239375
R10697 VDD.n4404 VDD.n4401 0.0239375
R10698 VDD.n4319 VDD.n4316 0.0239375
R10699 VDD.n3706 VDD.n3703 0.0239375
R10700 VDD.n3749 VDD.n3746 0.0239375
R10701 VDD.n5348 VDD.n5345 0.0239375
R10702 VDD.n8651 VDD.n8650 0.0239375
R10703 VDD.n8699 VDD.n8698 0.0239375
R10704 VDD.n8930 VDD.n8929 0.0239375
R10705 VDD.n3878 VDD.n3877 0.0239375
R10706 VDD.n3928 VDD.n3927 0.0239375
R10707 VDD VDD.n45 0.0235263
R10708 VDD VDD.n1754 0.0235263
R10709 VDD.n5357 VDD.n5356 0.0231563
R10710 VDD.n5253 VDD.n5252 0.022375
R10711 VDD.n4730 VDD.n4728 0.0222391
R10712 VDD.n5071 VDD.n5069 0.0222391
R10713 VDD.n4470 VDD.n4468 0.0222391
R10714 VDD.n4463 VDD.n4461 0.0222391
R10715 VDD.n4540 VDD.n4538 0.0222391
R10716 VDD.n4533 VDD.n4531 0.0222391
R10717 VDD.n4376 VDD.n4374 0.0222391
R10718 VDD.n4369 VDD.n4367 0.0222391
R10719 VDD.n3679 VDD.n3677 0.0222391
R10720 VDD.n3672 VDD.n3670 0.0222391
R10721 VDD.n5304 VDD.n5302 0.0222391
R10722 VDD.n5293 VDD.n5291 0.0222391
R10723 VDD.n4481 VDD.n4480 0.0219844
R10724 VDD.n4551 VDD.n4550 0.0219844
R10725 VDD.n4388 VDD.n4387 0.0219844
R10726 VDD.n4300 VDD.n4299 0.0219844
R10727 VDD.n3690 VDD.n3689 0.0219844
R10728 VDD.n3733 VDD.n3732 0.0219844
R10729 VDD.n5329 VDD.n5328 0.0219844
R10730 VDD.n8637 VDD.n8636 0.0219844
R10731 VDD.n8689 VDD.n8688 0.0219844
R10732 VDD.n8999 VDD.n8998 0.0219844
R10733 VDD.n8916 VDD.n8915 0.0219844
R10734 VDD.n3894 VDD.n3893 0.0219844
R10735 VDD.n8755 VDD.n8754 0.0217264
R10736 VDD.n8793 VDD.n8792 0.0217264
R10737 VDD.n8774 VDD.n8771 0.0217264
R10738 VDD.n14 VDD.n5 0.0215953
R10739 VDD.n890 VDD.n889 0.0215953
R10740 VDD.n1723 VDD.n1714 0.0215953
R10741 VDD.n2592 VDD.n2570 0.0215953
R10742 VDD.n9029 VDD.n5445 0.0211408
R10743 VDD.n5434 VDD.n5433 0.0210308
R10744 VDD.n5358 VDD.n5357 0.0208125
R10745 VDD.n3854 VDD.n3853 0.0205059
R10746 VDD.n3820 VDD.n3817 0.0205059
R10747 VDD.n3417 VDD.n2630 0.0202566
R10748 VDD.n3856 VDD.n3855 0.0200312
R10749 VDD.n3877 VDD.n3876 0.0200312
R10750 VDD.n3941 VDD.n3940 0.0200312
R10751 VDD.n922 VDD.n921 0.019913
R10752 VDD.n4596 VDD.n4595 0.0198977
R10753 VDD.n4603 VDD.n4602 0.0197278
R10754 VDD.n4568 VDD.n4542 0.0196275
R10755 VDD.n4740 VDD.n4737 0.0195217
R10756 VDD.n5081 VDD.n5078 0.0195217
R10757 VDD.n8873 VDD.n8801 0.0193679
R10758 VDD.n4962 VDD.n4961 0.01925
R10759 VDD.n4384 VDD.n4383 0.0186403
R10760 VDD.n4477 VDD.n4476 0.0186403
R10761 VDD.n4547 VDD.n4546 0.0186403
R10762 VDD.n3686 VDD.n3685 0.0186403
R10763 VDD.n3729 VDD.n3728 0.0186403
R10764 VDD.n4663 VDD.n4662 0.0185773
R10765 VDD.n4851 VDD.n4850 0.0185773
R10766 VDD.n4881 VDD.n4880 0.0185773
R10767 VDD.n4941 VDD.n4940 0.0185773
R10768 VDD.n67 VDD.n66 0.0185769
R10769 VDD.n1776 VDD.n1775 0.0185769
R10770 VDD.n8804 VDD.n8803 0.0181887
R10771 VDD.n3918 VDD.n3917 0.0180781
R10772 VDD.n3915 VDD.n3914 0.0180781
R10773 VDD.n3898 VDD.n3895 0.0180781
R10774 VDD.n3866 VDD.n3865 0.0180781
R10775 VDD.n3861 VDD.n3860 0.0180781
R10776 VDD.n4575 VDD.n4574 0.0176875
R10777 VDD.n3711 VDD.n3710 0.0176875
R10778 VDD.n8873 VDD.n8802 0.0176875
R10779 VDD.n4077 VDD.n4076 0.0176875
R10780 VDD.n4590 VDD.n4589 0.0169062
R10781 VDD.n8724 VDD.n8723 0.0169062
R10782 VDD.n4076 VDD.n3949 0.0169062
R10783 VDD.n4257 VDD.n4079 0.0169062
R10784 VDD.n4472 VDD.n4471 0.0168893
R10785 VDD.n4542 VDD.n4541 0.0168893
R10786 VDD.n4378 VDD.n4377 0.0168893
R10787 VDD.n3681 VDD.n3680 0.0168893
R10788 VDD.n5306 VDD.n5305 0.0168893
R10789 VDD.n4723 VDD.n4721 0.0168043
R10790 VDD.n5064 VDD.n5062 0.0168043
R10791 VDD.n4456 VDD.n4454 0.0168043
R10792 VDD.n4526 VDD.n4524 0.0168043
R10793 VDD.n4362 VDD.n4360 0.0168043
R10794 VDD.n3665 VDD.n3663 0.0168043
R10795 VDD.n5282 VDD.n5280 0.0168043
R10796 VDD.n29 VDD.n28 0.0165473
R10797 VDD.n884 VDD.n883 0.0165473
R10798 VDD.n1738 VDD.n1737 0.0165473
R10799 VDD.n2589 VDD.n2588 0.0165473
R10800 VDD.n4676 VDD.n4675 0.016125
R10801 VDD.n4668 VDD.n4667 0.016125
R10802 VDD.n4799 VDD.n4798 0.016125
R10803 VDD.n4794 VDD.n4793 0.016125
R10804 VDD.n4785 VDD.n4784 0.016125
R10805 VDD.n4831 VDD.n4830 0.016125
R10806 VDD.n4826 VDD.n4825 0.016125
R10807 VDD.n4821 VDD.n4820 0.016125
R10808 VDD.n4861 VDD.n4860 0.016125
R10809 VDD.n4856 VDD.n4855 0.016125
R10810 VDD.n4891 VDD.n4890 0.016125
R10811 VDD.n4886 VDD.n4885 0.016125
R10812 VDD.n4921 VDD.n4920 0.016125
R10813 VDD.n4916 VDD.n4915 0.016125
R10814 VDD.n4911 VDD.n4910 0.016125
R10815 VDD.n4951 VDD.n4950 0.016125
R10816 VDD.n4946 VDD.n4945 0.016125
R10817 VDD.n3844 VDD.n3843 0.016125
R10818 VDD.n3837 VDD.n3836 0.016125
R10819 VDD.n5016 VDD.n5015 0.016125
R10820 VDD.n5010 VDD.n5009 0.016125
R10821 VDD.n5142 VDD.n5141 0.016125
R10822 VDD.n5135 VDD.n5134 0.016125
R10823 VDD.n5126 VDD.n5125 0.016125
R10824 VDD.n5216 VDD.n5215 0.016125
R10825 VDD.n5208 VDD.n5207 0.016125
R10826 VDD.n5203 VDD.n5202 0.016125
R10827 VDD.n5350 VDD.n5254 0.016125
R10828 VDD.n3926 VDD.n3925 0.016125
R10829 VDD.n3919 VDD.n3918 0.016125
R10830 VDD.n4078 VDD.n3941 0.016125
R10831 VDD.n4260 VDD.n4259 0.016125
R10832 VDD.n20 VDD.n17 0.0157415
R10833 VDD.n876 VDD.n875 0.0157415
R10834 VDD.n1729 VDD.n1726 0.0157415
R10835 VDD.n2577 VDD.n2576 0.0157415
R10836 VDD.n9013 VDD.n8962 0.0145625
R10837 VDD.n4972 VDD.n4971 0.0145625
R10838 VDD.n3638 VDD.n3635 0.0143978
R10839 VDD.n3638 VDD.n3637 0.0143978
R10840 VDD.n3637 VDD.n3636 0.0143978
R10841 VDD.n5373 VDD.n3640 0.0143978
R10842 VDD.n5373 VDD.n5372 0.0143978
R10843 VDD.n5372 VDD.n5371 0.0143978
R10844 VDD.n5371 VDD.n5370 0.0143978
R10845 VDD.n5370 VDD.n5369 0.0143978
R10846 VDD.n5367 VDD.n5366 0.0143978
R10847 VDD.n5404 VDD.n5403 0.0143978
R10848 VDD.n5407 VDD.n5406 0.0143978
R10849 VDD.n5408 VDD.n5407 0.0143978
R10850 VDD.n5410 VDD.n5408 0.0143978
R10851 VDD.n8583 VDD.n8582 0.0143978
R10852 VDD.n8584 VDD.n8583 0.0143978
R10853 VDD.n9025 VDD.n9024 0.0143978
R10854 VDD.n9022 VDD.n9021 0.0143978
R10855 VDD.n9021 VDD.n9020 0.0143978
R10856 VDD.n9020 VDD.n9019 0.0143978
R10857 VDD.n9019 VDD.n9018 0.0143978
R10858 VDD.n9018 VDD.n8598 0.0143978
R10859 VDD.n8596 VDD.n8595 0.0143978
R10860 VDD.n8595 VDD.n8594 0.0143978
R10861 VDD.n8594 VDD.n8593 0.0143978
R10862 VDD.n8593 VDD.n8592 0.0143978
R10863 VDD.n8590 VDD.n8589 0.0143978
R10864 VDD.n8589 VDD.n8588 0.0143978
R10865 VDD.n5390 VDD.n5384 0.0143978
R10866 VDD.n5390 VDD.n5389 0.0143978
R10867 VDD.n5389 VDD.n5388 0.0143978
R10868 VDD.n5388 VDD.n5387 0.0143978
R10869 VDD.n3825 VDD.n3824 0.0143978
R10870 VDD.n3826 VDD.n3825 0.0143978
R10871 VDD.n3827 VDD.n3826 0.0143978
R10872 VDD.n3828 VDD.n3827 0.0143978
R10873 VDD.n3831 VDD.n3830 0.0143978
R10874 VDD.n4978 VDD.n3831 0.0143978
R10875 VDD.n4979 VDD.n4978 0.0143978
R10876 VDD.n4980 VDD.n4979 0.0143978
R10877 VDD.n4981 VDD.n4980 0.0143978
R10878 VDD.n4982 VDD.n4981 0.0143978
R10879 VDD.n4983 VDD.n4982 0.0143978
R10880 VDD.n4987 VDD.n4983 0.0143978
R10881 VDD.n4987 VDD.n4986 0.0143978
R10882 VDD.n4986 VDD.n4985 0.0143978
R10883 VDD.n4985 VDD.n4984 0.0143978
R10884 VDD.n4984 VDD.n3631 0.0143978
R10885 VDD.n3631 VDD.n3630 0.0143978
R10886 VDD.n5429 VDD.n5428 0.0143978
R10887 VDD.n4661 VDD.n4660 0.0141719
R10888 VDD.n4783 VDD.n4782 0.0141719
R10889 VDD.n4819 VDD.n4815 0.0141719
R10890 VDD.n4849 VDD.n4848 0.0141719
R10891 VDD.n4879 VDD.n4878 0.0141719
R10892 VDD.n4909 VDD.n4908 0.0141719
R10893 VDD.n4939 VDD.n4938 0.0141719
R10894 VDD.n3855 VDD.n3854 0.0141719
R10895 VDD.n3817 VDD.n3816 0.0141719
R10896 VDD.n5124 VDD.n5123 0.0141719
R10897 VDD.n5201 VDD.n5192 0.0141719
R10898 VDD.n8668 VDD.n8659 0.0141719
R10899 VDD.n8712 VDD.n8707 0.0141719
R10900 VDD.n8747 VDD.n8738 0.0141719
R10901 VDD.n8947 VDD.n8938 0.0141719
R10902 VDD.n3936 VDD.n3935 0.0141719
R10903 VDD.n4656 VDD.n4654 0.014087
R10904 VDD.n4778 VDD.n4776 0.014087
R10905 VDD.n4747 VDD.n4744 0.014087
R10906 VDD.n5119 VDD.n5117 0.014087
R10907 VDD.n5088 VDD.n5085 0.014087
R10908 VDD.n5188 VDD.n5186 0.014087
R10909 VDD.n9026 VDD.n8584 0.0138925
R10910 VDD.n5365 VDD.n5364 0.0137813
R10911 VDD.n8591 VDD.n8590 0.0136398
R10912 VDD.n5362 VDD.n5361 0.013
R10913 VDD.n9016 VDD.n9015 0.013
R10914 VDD.n4969 VDD.n4968 0.013
R10915 VDD.n4605 VDD.n4601 0.0128788
R10916 VDD.n4594 VDD.n4593 0.0128788
R10917 VDD.n4593 VDD.n4592 0.0128788
R10918 VDD.n4605 VDD.n4604 0.0128788
R10919 VDD.n4788 VDD.n4787 0.0127111
R10920 VDD.n4824 VDD.n4823 0.0127111
R10921 VDD.n4914 VDD.n4913 0.0127111
R10922 VDD.n5129 VDD.n5128 0.0127111
R10923 VDD.n5206 VDD.n5205 0.0127111
R10924 VDD.n5384 VDD.n5383 0.012629
R10925 VDD.n8798 VDD.n8797 0.0122925
R10926 VDD.n8801 VDD.n8800 0.0122925
R10927 VDD.n8810 VDD.n8809 0.0122925
R10928 VDD.n4667 VDD.n4666 0.0122188
R10929 VDD.n4855 VDD.n4854 0.0122188
R10930 VDD.n4885 VDD.n4884 0.0122188
R10931 VDD.n4945 VDD.n4944 0.0122188
R10932 VDD.n4482 VDD.n4481 0.0122188
R10933 VDD.n4493 VDD.n4492 0.0122188
R10934 VDD.n4552 VDD.n4551 0.0122188
R10935 VDD.n4563 VDD.n4562 0.0122188
R10936 VDD.n4389 VDD.n4388 0.0122188
R10937 VDD.n4400 VDD.n4399 0.0122188
R10938 VDD.n4301 VDD.n4300 0.0122188
R10939 VDD.n4315 VDD.n4314 0.0122188
R10940 VDD.n3691 VDD.n3690 0.0122188
R10941 VDD.n3702 VDD.n3701 0.0122188
R10942 VDD.n3734 VDD.n3733 0.0122188
R10943 VDD.n3745 VDD.n3744 0.0122188
R10944 VDD.n5330 VDD.n5329 0.0122188
R10945 VDD.n5344 VDD.n5343 0.0122188
R10946 VDD.n8649 VDD.n8648 0.0122188
R10947 VDD.n8638 VDD.n8637 0.0122188
R10948 VDD.n8697 VDD.n8696 0.0122188
R10949 VDD.n8690 VDD.n8689 0.0122188
R10950 VDD.n9011 VDD.n9003 0.0122188
R10951 VDD.n9000 VDD.n8999 0.0122188
R10952 VDD.n8928 VDD.n8927 0.0122188
R10953 VDD.n8917 VDD.n8916 0.0122188
R10954 VDD.n3931 VDD.n3930 0.0122188
R10955 VDD.n3917 VDD.n3916 0.0122188
R10956 VDD.n3895 VDD.n3894 0.0122188
R10957 VDD.n3874 VDD.n3873 0.0122188
R10958 VDD.n24 VDD.n23 0.0114797
R10959 VDD.n15 VDD.n14 0.0114797
R10960 VDD.n873 VDD.n872 0.0114797
R10961 VDD.n889 VDD.n888 0.0114797
R10962 VDD.n1733 VDD.n1732 0.0114797
R10963 VDD.n1724 VDD.n1723 0.0114797
R10964 VDD.n2583 VDD.n2579 0.0114797
R10965 VDD.n2592 VDD.n2591 0.0114797
R10966 VDD.n5353 VDD.n5352 0.0114375
R10967 VDD.n2560 VDD.n1777 0.0111838
R10968 VDD.n1706 VDD.n923 0.0111838
R10969 VDD.n851 VDD.n68 0.0111838
R10970 VDD.n8750 VDD.n8749 0.0111132
R10971 VDD.n8799 VDD.n8798 0.0111132
R10972 VDD.n5019 VDD.n4998 0.0106562
R10973 VDD.n5020 VDD.n5019 0.0106562
R10974 VDD.n4494 VDD.n4493 0.0102656
R10975 VDD.n4564 VDD.n4563 0.0102656
R10976 VDD.n4401 VDD.n4400 0.0102656
R10977 VDD.n4316 VDD.n4315 0.0102656
R10978 VDD.n3703 VDD.n3702 0.0102656
R10979 VDD.n3746 VDD.n3745 0.0102656
R10980 VDD.n5345 VDD.n5344 0.0102656
R10981 VDD.n8650 VDD.n8649 0.0102656
R10982 VDD.n8698 VDD.n8697 0.0102656
R10983 VDD.n9003 VDD.n9002 0.0102656
R10984 VDD.n8929 VDD.n8928 0.0102656
R10985 VDD.n5368 VDD.n5367 0.0101021
R10986 VDD.n8582 VDD.n8581 0.0101021
R10987 VDD.n8588 VDD.n8587 0.0101021
R10988 VDD.n3415 VDD.n3414 0.0100583
R10989 VDD.n2562 VDD.n2561 0.0100583
R10990 VDD.n1708 VDD.n1707 0.0100583
R10991 VDD.n853 VDD.n852 0.0100583
R10992 VDD.n8751 VDD.n8750 0.00993396
R10993 VDD.n8797 VDD.n8796 0.00993396
R10994 VDD.n8598 VDD.n8597 0.00984946
R10995 VDD.n3829 VDD.n3828 0.00984946
R10996 VDD.n4585 VDD.n4584 0.00957737
R10997 VDD.n4579 VDD.n4578 0.00957737
R10998 VDD.n4570 VDD.n4569 0.00957737
R10999 VDD.n4584 VDD.n4583 0.00957737
R11000 VDD.n4580 VDD.n4579 0.00957737
R11001 VDD.n4571 VDD.n4570 0.00957737
R11002 VDD.n5363 VDD.n5362 0.00957737
R11003 VDD.n5247 VDD.n5246 0.00957737
R11004 VDD.n5364 VDD.n5363 0.00957737
R11005 VDD.n5248 VDD.n5247 0.00957737
R11006 VDD.n8674 VDD.n8673 0.00957737
R11007 VDD.n8716 VDD.n8715 0.00957737
R11008 VDD.n8877 VDD.n8876 0.00957737
R11009 VDD.n8673 VDD.n8672 0.00957737
R11010 VDD.n8715 VDD.n8714 0.00957737
R11011 VDD.n8949 VDD.n8877 0.00957737
R11012 VDD.n4679 VDD.n4678 0.00957737
R11013 VDD.n4802 VDD.n4801 0.00957737
R11014 VDD.n4835 VDD.n4834 0.00957737
R11015 VDD.n4865 VDD.n4864 0.00957737
R11016 VDD.n4894 VDD.n4893 0.00957737
R11017 VDD.n4925 VDD.n4924 0.00957737
R11018 VDD.n4955 VDD.n4954 0.00957737
R11019 VDD.n5145 VDD.n5144 0.00957737
R11020 VDD.n5220 VDD.n5219 0.00957737
R11021 VDD.n5224 VDD.n5223 0.00957737
R11022 VDD.n5219 VDD.n5218 0.00957737
R11023 VDD.n4954 VDD.n4953 0.00957737
R11024 VDD.n4924 VDD.n4923 0.00957737
R11025 VDD.n4864 VDD.n4863 0.00957737
R11026 VDD.n4895 VDD.n4894 0.00957737
R11027 VDD.n4834 VDD.n4833 0.00957737
R11028 VDD.n4680 VDD.n4679 0.00957737
R11029 VDD.n4803 VDD.n4802 0.00957737
R11030 VDD.n5146 VDD.n5145 0.00957737
R11031 VDD.n5225 VDD.n5224 0.00957737
R11032 VDD.n4277 VDD.n4261 0.00955797
R11033 VDD.n4258 VDD.n3859 0.00955797
R11034 VDD.n5410 VDD.n5409 0.00934409
R11035 VDD.n47 VDD.n46 0.00927193
R11036 VDD.n1756 VDD.n1755 0.00927193
R11037 VDD.n5225 VDD.n5222 0.00923422
R11038 VDD.n4277 VDD.n4264 0.0091882
R11039 VDD.n4587 VDD.n4586 0.0091882
R11040 VDD.n4581 VDD.n4580 0.0091882
R11041 VDD.n4576 VDD.n4575 0.0091882
R11042 VDD.n4572 VDD.n4571 0.0091882
R11043 VDD.n4586 VDD.n4585 0.0091882
R11044 VDD.n4573 VDD.n4572 0.0091882
R11045 VDD.n4577 VDD.n4576 0.0091882
R11046 VDD.n4582 VDD.n4581 0.0091882
R11047 VDD.n4264 VDD.n4263 0.0091882
R11048 VDD.n3710 VDD.n3709 0.0091882
R11049 VDD.n5351 VDD.n5350 0.0091882
R11050 VDD.n5250 VDD.n5249 0.0091882
R11051 VDD.n5352 VDD.n5351 0.0091882
R11052 VDD.n5249 VDD.n5248 0.0091882
R11053 VDD.n3709 VDD.n3708 0.0091882
R11054 VDD.n8671 VDD.n8670 0.0091882
R11055 VDD.n8676 VDD.n8675 0.0091882
R11056 VDD.n9015 VDD.n9014 0.0091882
R11057 VDD.n8951 VDD.n8950 0.0091882
R11058 VDD.n8875 VDD.n8874 0.0091882
R11059 VDD.n9014 VDD.n9013 0.0091882
R11060 VDD.n8672 VDD.n8671 0.0091882
R11061 VDD.n8950 VDD.n8949 0.0091882
R11062 VDD.n8714 VDD.n8676 0.0091882
R11063 VDD.n8874 VDD.n8873 0.0091882
R11064 VDD.n4678 VDD.n4608 0.0091882
R11065 VDD.n4801 VDD.n4682 0.0091882
R11066 VDD.n4805 VDD.n4804 0.0091882
R11067 VDD.n4837 VDD.n4836 0.0091882
R11068 VDD.n4893 VDD.n4867 0.0091882
R11069 VDD.n4923 VDD.n4897 0.0091882
R11070 VDD.n4927 VDD.n4926 0.0091882
R11071 VDD.n4970 VDD.n4969 0.0091882
R11072 VDD.n5144 VDD.n5023 0.0091882
R11073 VDD.n5148 VDD.n5147 0.0091882
R11074 VDD.n4953 VDD.n4927 0.0091882
R11075 VDD.n5023 VDD.n5022 0.0091882
R11076 VDD.n5218 VDD.n5148 0.0091882
R11077 VDD.n4971 VDD.n4970 0.0091882
R11078 VDD.n4897 VDD.n4896 0.0091882
R11079 VDD.n4867 VDD.n4866 0.0091882
R11080 VDD.n4863 VDD.n4837 0.0091882
R11081 VDD.n4608 VDD.n4607 0.0091882
R11082 VDD.n4682 VDD.n4681 0.0091882
R11083 VDD.n4833 VDD.n4805 0.0091882
R11084 VDD.n5222 VDD.n5221 0.00914234
R11085 VDD.n9024 VDD.n9023 0.0090914
R11086 VDD.n24 VDD.n22 0.00894595
R11087 VDD.n873 VDD.n871 0.00894595
R11088 VDD.n1733 VDD.n1731 0.00894595
R11089 VDD.n2579 VDD.n2578 0.00894595
R11090 VDD.n917 VDD.n914 0.00887321
R11091 VDD.n917 VDD.n916 0.00887321
R11092 VDD.n2626 VDD.n2623 0.00887321
R11093 VDD.n2626 VDD.n2625 0.00887321
R11094 VDD.n4600 VDD.n4599 0.00867391
R11095 VDD.n4645 VDD.n4643 0.00865217
R11096 VDD.n4771 VDD.n4769 0.00865217
R11097 VDD.n4754 VDD.n4751 0.00865217
R11098 VDD.n5112 VDD.n5110 0.00865217
R11099 VDD.n5095 VDD.n5092 0.00865217
R11100 VDD.n5177 VDD.n5175 0.00865217
R11101 VDD.n8631 VDD.n8629 0.00865217
R11102 VDD.n8993 VDD.n8991 0.00865217
R11103 VDD.n8903 VDD.n8901 0.00865217
R11104 VDD.n4258 VDD.n3858 0.00865217
R11105 VDD.n5386 VDD.n5385 0.00833333
R11106 VDD.n4480 VDD.n4479 0.0083125
R11107 VDD.n4550 VDD.n4549 0.0083125
R11108 VDD.n4387 VDD.n4386 0.0083125
R11109 VDD.n4299 VDD.n4298 0.0083125
R11110 VDD.n3689 VDD.n3688 0.0083125
R11111 VDD.n3732 VDD.n3731 0.0083125
R11112 VDD.n5328 VDD.n5327 0.0083125
R11113 VDD.n8636 VDD.n8635 0.0083125
R11114 VDD.n8688 VDD.n8687 0.0083125
R11115 VDD.n8998 VDD.n8997 0.0083125
R11116 VDD.n8915 VDD.n8914 0.0083125
R11117 VDD.n3938 VDD.n3878 0.0083125
R11118 VDD.n3913 VDD.n3910 0.0083125
R11119 VDD.n3908 VDD.n3907 0.0083125
R11120 VDD.n8759 VDD.n5446 0.0081375
R11121 VDD.n5397 VDD.n5396 0.00808064
R11122 VDD.n2560 VDD.n2559 0.00794532
R11123 VDD.n1706 VDD.n1705 0.00794532
R11124 VDD.n851 VDD.n850 0.00794532
R11125 VDD.n5406 VDD.n5405 0.00782796
R11126 VDD.n4277 VDD.n4276 0.00774638
R11127 VDD.n8756 VDD.n8755 0.00757547
R11128 VDD.n5021 VDD.n5020 0.00753125
R11129 VDD.n5405 VDD.n5404 0.00706989
R11130 VDD.n8761 VDD.n8757 0.00694587
R11131 VDD.n5207 VDD.n5206 0.00685176
R11132 VDD.n5134 VDD.n5129 0.00685176
R11133 VDD.n4915 VDD.n4914 0.00685176
R11134 VDD.n4825 VDD.n4824 0.00685176
R11135 VDD.n4793 VDD.n4788 0.00685176
R11136 VDD.n5382 VDD.n5381 0.0068172
R11137 VDD.n4604 VDD.n4603 0.00678574
R11138 VDD.n5252 VDD.n5251 0.00675
R11139 VDD.n4998 VDD.n4997 0.00675
R11140 VDD.n4595 VDD.n4594 0.00661507
R11141 VDD.n5387 VDD.n5386 0.00656452
R11142 VDD.n8792 VDD.n8791 0.00639623
R11143 VDD.n3414 VDD.n3412 0.00638768
R11144 VDD.n2561 VDD.n1778 0.00638768
R11145 VDD.n1707 VDD.n924 0.00638768
R11146 VDD.n852 VDD.n69 0.00638768
R11147 VDD.n4666 VDD.n4665 0.00635938
R11148 VDD.n4854 VDD.n4853 0.00635938
R11149 VDD.n4884 VDD.n4883 0.00635938
R11150 VDD.n4944 VDD.n4943 0.00635938
R11151 VDD.n3847 VDD.n3846 0.00635938
R11152 VDD.n5002 VDD.n5001 0.00635938
R11153 VDD.n5000 VDD.n4999 0.00635938
R11154 VDD.n4267 VDD.n4265 0.00635938
R11155 VDD.n3937 VDD.n3936 0.00635938
R11156 VDD.n3927 VDD.n3926 0.00635938
R11157 VDD.n4697 VDD.n4695 0.00593478
R11158 VDD.n4713 VDD.n4711 0.00593478
R11159 VDD.n5038 VDD.n5036 0.00593478
R11160 VDD.n5054 VDD.n5052 0.00593478
R11161 VDD.n4335 VDD.n4333 0.00593478
R11162 VDD.n4351 VDD.n4349 0.00593478
R11163 VDD.n4418 VDD.n4416 0.00593478
R11164 VDD.n4446 VDD.n4444 0.00593478
R11165 VDD.n4434 VDD.n4427 0.00593478
R11166 VDD.n4516 VDD.n4514 0.00593478
R11167 VDD.n3655 VDD.n3653 0.00593478
R11168 VDD.n5272 VDD.n5270 0.00593478
R11169 VDD.n9023 VDD.n9022 0.00580645
R11170 VDD.n4598 VDD.n4597 0.0056087
R11171 VDD.n4589 VDD.n4588 0.0051875
R11172 VDD.n4606 VDD.n4260 0.0051875
R11173 VDD.n8597 VDD.n8596 0.00504839
R11174 VDD.n3830 VDD.n3829 0.00504839
R11175 VDD.n4597 VDD.n4596 0.00492754
R11176 VDD.n5018 VDD.n5016 0.00490286
R11177 VDD.n3843 VDD.n3842 0.00490286
R11178 VDD.n5414 VDD.n5413 0.0047957
R11179 VDD.n5369 VDD.n5368 0.0047957
R11180 VDD.n5400 VDD.n5398 0.0047957
R11181 VDD.n8581 VDD.n8580 0.0047957
R11182 VDD.n8587 VDD.n8586 0.0047957
R11183 VDD.n8759 VDD.n8758 0.00449057
R11184 VDD.n4784 VDD.n4783 0.00440625
R11185 VDD.n4820 VDD.n4819 0.00440625
R11186 VDD.n4910 VDD.n4909 0.00440625
R11187 VDD.n5125 VDD.n5124 0.00440625
R11188 VDD.n5202 VDD.n5201 0.00440625
R11189 VDD.n4486 VDD.n4482 0.00440625
R11190 VDD.n4556 VDD.n4552 0.00440625
R11191 VDD.n4393 VDD.n4389 0.00440625
R11192 VDD.n4305 VDD.n4301 0.00440625
R11193 VDD.n4263 VDD.n4262 0.00440625
R11194 VDD.n3695 VDD.n3691 0.00440625
R11195 VDD.n3738 VDD.n3734 0.00440625
R11196 VDD.n5334 VDD.n5330 0.00440625
R11197 VDD.n8657 VDD.n8654 0.00440625
R11198 VDD.n8639 VDD.n8638 0.00440625
R11199 VDD.n8705 VDD.n8702 0.00440625
R11200 VDD.n8691 VDD.n8690 0.00440625
R11201 VDD.n8736 VDD.n8733 0.00440625
R11202 VDD.n9001 VDD.n9000 0.00440625
R11203 VDD.n8936 VDD.n8933 0.00440625
R11204 VDD.n8918 VDD.n8917 0.00440625
R11205 VDD.n3929 VDD.n3928 0.00440625
R11206 VDD.n3921 VDD.n3920 0.00440625
R11207 VDD.n3899 VDD.n3898 0.00440625
R11208 VDD.n3870 VDD.n3869 0.00440625
R11209 VDD.n4255 VDD.n4252 0.00433093
R11210 VDD.n5400 VDD.n5399 0.00429032
R11211 VDD.n8580 VDD.n8579 0.00429032
R11212 VDD.n8586 VDD.n8585 0.00429032
R11213 VDD.n8761 VDD.n8760 0.00397228
R11214 VDD.n5365 VDD.n3723 0.003625
R11215 VDD.n8962 VDD.n8961 0.003625
R11216 VDD.n4973 VDD.n4972 0.003625
R11217 VDD.n4997 VDD.n4996 0.003625
R11218 VDD.n4634 VDD.n4632 0.00321739
R11219 VDD.n4764 VDD.n4762 0.00321739
R11220 VDD.n4760 VDD.n4758 0.00321739
R11221 VDD.n5105 VDD.n5103 0.00321739
R11222 VDD.n5101 VDD.n5099 0.00321739
R11223 VDD.n5166 VDD.n5164 0.00321739
R11224 VDD.n4287 VDD.n4285 0.00321739
R11225 VDD.n5316 VDD.n5314 0.00321739
R11226 VDD.n8620 VDD.n8618 0.00321739
R11227 VDD.n8982 VDD.n8980 0.00321739
R11228 VDD.n8892 VDD.n8890 0.00321739
R11229 VDD VDD.n6 0.00303378
R11230 VDD VDD.n892 0.00303378
R11231 VDD VDD.n1715 0.00303378
R11232 VDD VDD.n2572 0.00303378
R11233 VDD.n4662 VDD.n4661 0.00295228
R11234 VDD.n4850 VDD.n4849 0.00295228
R11235 VDD.n4880 VDD.n4879 0.00295228
R11236 VDD.n4940 VDD.n4939 0.00295228
R11237 VDD.n8794 VDD.n8793 0.00285849
R11238 VDD.n8777 VDD.n8776 0.00285849
R11239 VDD.n8809 VDD.n8804 0.00285849
R11240 VDD.n3718 VDD.n3717 0.00284375
R11241 VDD.n8957 VDD.n8956 0.00284375
R11242 VDD.n5440 VDD.n5439 0.00278115
R11243 VDD.n5441 VDD.n5440 0.00278115
R11244 VDD.n5379 VDD.n5378 0.00262546
R11245 VDD.n5380 VDD.n5379 0.00262546
R11246 VDD.n5398 VDD.n5397 0.00252151
R11247 VDD.n8574 VDD.n8546 0.00251613
R11248 VDD.n8659 VDD.n8658 0.00245312
R11249 VDD.n8707 VDD.n8706 0.00245312
R11250 VDD.n8738 VDD.n8737 0.00245312
R11251 VDD.n8938 VDD.n8937 0.00245312
R11252 VDD.n8865 VDD.n8864 0.00244542
R11253 VDD.n5426 VDD.n5425 0.00243946
R11254 VDD.n5415 VDD.n5412 0.00243946
R11255 VDD.n5416 VDD.n5415 0.00243946
R11256 VDD.n5427 VDD.n5426 0.00243946
R11257 VDD.n5383 VDD.n5382 0.00226882
R11258 VDD.n3634 VDD.n3632 0.00226882
R11259 VDD.n4592 VDD.n4591 0.0022029
R11260 VDD.n8827 VDD.n8826 0.00207156
R11261 VDD.n8830 VDD.n8829 0.00207156
R11262 VDD.n3943 VDD.n3942 0.00207156
R11263 VDD.n4071 VDD.n4070 0.00207156
R11264 VDD.n3752 VDD.n3751 0.00207156
R11265 VDD.n5240 VDD.n5239 0.00207156
R11266 VDD.n4203 VDD.n4202 0.00207156
R11267 VDD.n5254 VDD.n5253 0.0020625
R11268 VDD.n8821 VDD.n8820 0.00194557
R11269 VDD.n8862 VDD.n8821 0.00194557
R11270 VDD.n8845 VDD.n8844 0.00194557
R11271 VDD.n8862 VDD.n8845 0.00194557
R11272 VDD.n8826 VDD.n8825 0.00194557
R11273 VDD.n8829 VDD.n8828 0.00194557
R11274 VDD.n8864 VDD.n8863 0.00194557
R11275 VDD.n3944 VDD.n3943 0.00194557
R11276 VDD.n4072 VDD.n4071 0.00194557
R11277 VDD.n3753 VDD.n3752 0.00194557
R11278 VDD.n5241 VDD.n5240 0.00194557
R11279 VDD.n5230 VDD.n5229 0.00194557
R11280 VDD.n5238 VDD.n5230 0.00194557
R11281 VDD.n3771 VDD.n3770 0.00194557
R11282 VDD.n5238 VDD.n3771 0.00194557
R11283 VDD.n4202 VDD.n4201 0.00194557
R11284 VDD.n4210 VDD.n4209 0.00194557
R11285 VDD.n4242 VDD.n4210 0.00194557
R11286 VDD.n4244 VDD.n4243 0.00194557
R11287 VDD.n4243 VDD.n4242 0.00194557
R11288 VDD.n4111 VDD.n4110 0.00194557
R11289 VDD.n4242 VDD.n4111 0.00194557
R11290 VDD.n4601 VDD.n4600 0.00186232
R11291 VDD.n3634 VDD.n3633 0.00176344
R11292 VDD.n3622 VDD.n3597 0.00175186
R11293 VDD.n8752 VDD.n8751 0.00167925
R11294 VDD.n8754 VDD.n8753 0.00167925
R11295 VDD.n8796 VDD.n8795 0.00167925
R11296 VDD.n8767 VDD.n8766 0.00167925
R11297 VDD.n8769 VDD.n8768 0.00167925
R11298 VDD.n8775 VDD.n8774 0.00167925
R11299 VDD.n5437 VDD.n5436 0.00145036
R11300 VDD.n5436 VDD.n5435 0.00145036
R11301 VDD.n5445 VDD.n5444 0.00143078
R11302 VDD.n5444 VDD.n5443 0.00143078
R11303 VDD.n5394 VDD.n5393 0.00141098
R11304 VDD.n5393 VDD.n5392 0.00141098
R11305 VDD.n4276 VDD.n4275 0.0014058
R11306 VDD.n5375 VDD.n5374 0.00139311
R11307 VDD.n5376 VDD.n5375 0.00139311
R11308 VDD.n8862 VDD.n8827 0.00137395
R11309 VDD.n8862 VDD.n8830 0.00137395
R11310 VDD.n4070 VDD.n4069 0.00137395
R11311 VDD.n5239 VDD.n5238 0.00137395
R11312 VDD.n4242 VDD.n4203 0.00137395
R11313 VDD.n5422 VDD.n5421 0.00136393
R11314 VDD.n5402 VDD.n5401 0.00136393
R11315 VDD.n5423 VDD.n5422 0.00136393
R11316 VDD.n5401 VDD.n5395 0.00136393
R11317 VDD.n5432 VDD.n5431 0.00134811
R11318 VDD.n5419 VDD.n5418 0.00134811
R11319 VDD.n5420 VDD.n5419 0.00134811
R11320 VDD.n5433 VDD.n5432 0.00134811
R11321 VDD.n4590 VDD.n4277 0.00128125
R11322 VDD.n4258 VDD.n4257 0.00128125
R11323 VDD.n4259 VDD.n4258 0.00128125
R11324 VDD.n3640 VDD.n3639 0.00125806
R11325 VDD.n8592 VDD.n8591 0.00125806
R11326 VDD.n5443 VDD.n5442 0.00119582
R11327 VDD.n5442 VDD.n5441 0.00119582
R11328 VDD.n5378 VDD.n5377 0.0011787
R11329 VDD.n5377 VDD.n5376 0.0011787
R11330 VDD.n8576 VDD.n8575 0.00117707
R11331 VDD.n5439 VDD.n5438 0.00117624
R11332 VDD.n5438 VDD.n5437 0.00117624
R11333 VDD.n5392 VDD.n5391 0.00116083
R11334 VDD.n5391 VDD.n5380 0.00116083
R11335 VDD.n5431 VDD.n5430 0.00115824
R11336 VDD.n5417 VDD.n5416 0.00115824
R11337 VDD.n5418 VDD.n5417 0.00115824
R11338 VDD.n5430 VDD.n5427 0.00115824
R11339 VDD.n5424 VDD.n5423 0.00114242
R11340 VDD.n5412 VDD.n5411 0.00114242
R11341 VDD.n5411 VDD.n5402 0.00114242
R11342 VDD.n5425 VDD.n5424 0.00114242
R11343 VDD.n9030 VDD.n9029 0.00112121
R11344 VDD.n5237 VDD.n5232 0.00105433
R11345 VDD.n4208 VDD.n4207 0.00104275
R11346 VDD.n3622 VDD.n3621 0.00104275
R11347 VDD.n5237 VDD.n5236 0.00104275
R11348 VDD.n8862 VDD.n8861 0.00103737
R11349 VDD.n3623 VDD.n3622 0.00103651
R11350 VDD.n4208 VDD.n4205 0.00101611
R11351 VDD.n8824 VDD.n8823 0.00101576
R11352 VDD.n3779 VDD.n3778 0.00101522
R11353 VDD.n8843 VDD.n8842 0.00100772
R11354 VDD.n8861 VDD.n8860 0.00100538
R11355 VDD.n9026 VDD.n9025 0.00100538
R11356 VDD.n4116 VDD.n4113 0.00100409
R11357 VDD.n3776 VDD.n3773 0.00100409
R11358 VDD.n8866 VDD.n8865 0.00100372
R11359 VDD.n4064 VDD.n4063 0.00100292
R11360 VDD.n4064 VDD.n4061 0.00100251
R11361 VDD.n3776 VDD.n3775 0.00100251
R11362 VDD.n4116 VDD.n4115 0.00100251
R11363 VDD.n8862 VDD.n8824 0.00100095
R11364 VDD.n5238 VDD.n3779 0.00100089
R11365 VDD.n8862 VDD.n8843 0.00100024
R11366 VDD.n3628 VDD.n3627 0.00100002
R11367 VDD.n3412 VDD.n3041 0.00100001
R11368 VDD.n2559 VDD.n1778 0.00100001
R11369 VDD.n1705 VDD.n924 0.00100001
R11370 VDD.n850 VDD.n69 0.00100001
R11371 VDD.n853 VDD.n68 0.001
R11372 VDD.n1708 VDD.n923 0.001
R11373 VDD.n2562 VDD.n1777 0.001
R11374 VDD.n3416 VDD.n3415 0.001
R11375 VDD.n8865 VDD.n8862 0.001
R11376 VDD.n4069 VDD.n4064 0.001
R11377 VDD.n5238 VDD.n3776 0.001
R11378 VDD.n5238 VDD.n5237 0.001
R11379 VDD.n4242 VDD.n4208 0.001
R11380 VDD.n4242 VDD.n4116 0.001
R11381 VDD.n8577 VDD.n5450 0.000855023
R11382 VDD.n8577 VDD.n8576 0.000855023
R11383 VDD.n5450 VDD.n5449 0.000855004
R11384 VDD.n8760 VDD.n8759 0.00079375
R11385 VDD.n5232 VDD.n5231 0.000554326
R11386 VDD.n8832 VDD.n8831 0.000542748
R11387 VDD.n8862 VDD.n8832 0.000542748
R11388 VDD.n8860 VDD.n8859 0.000542748
R11389 VDD.n3621 VDD.n3620 0.000542748
R11390 VDD.n3625 VDD.n3624 0.000542748
R11391 VDD.n3624 VDD.n3623 0.000542748
R11392 VDD.n5236 VDD.n5235 0.000542748
R11393 VDD.n3811 VDD.n3810 0.000542748
R11394 VDD.n5238 VDD.n3811 0.000542748
R11395 VDD.n4207 VDD.n4206 0.000542748
R11396 VDD.n4066 VDD.n4065 0.000542748
R11397 VDD.n4069 VDD.n4066 0.000542748
R11398 VDD.n4069 VDD.n4068 0.000523923
R11399 VDD.n4242 VDD.n4241 0.000523923
R11400 VDD.n4241 VDD.n4240 0.000523923
R11401 VDD.n4068 VDD.n4067 0.000523923
R11402 VDD.n8823 VDD.n8822 0.000516711
R11403 VDD.n3778 VDD.n3777 0.000516107
R11404 VDD.n4205 VDD.n4204 0.000516107
R11405 VDD.n8842 VDD.n8841 0.000507966
R11406 VDD.n3773 VDD.n3772 0.000504095
R11407 VDD.n4113 VDD.n4112 0.000504095
R11408 VDD.n8867 VDD.n8866 0.000503718
R11409 VDD.n4063 VDD.n4062 0.000502918
R11410 VDD.n4237 VDD.n4236 0.000502851
R11411 VDD.n4236 VDD.n4235 0.000502851
R11412 VDD.n4061 VDD.n4060 0.000502515
R11413 VDD.n3775 VDD.n3774 0.000502515
R11414 VDD.n4115 VDD.n4114 0.000502515
R11415 VDD.n3597 VDD.n3596 0.000501859
R11416 VDD.n4239 VDD.n4238 0.000501425
R11417 VDD.n4238 VDD.n4237 0.000501425
R11418 VDD.n3412 VDD.n3411 0.000500887
R11419 VDD.n1899 VDD.n1778 0.000500887
R11420 VDD.n1045 VDD.n924 0.000500887
R11421 VDD.n190 VDD.n69 0.000500887
R11422 VDD.n3414 VDD.n3413 0.000500755
R11423 VDD.n2561 VDD.n2560 0.000500755
R11424 VDD.n1707 VDD.n1706 0.000500755
R11425 VDD.n852 VDD.n851 0.000500755
R11426 VDD.n6668 VDD.n6667 0.000500648
R11427 VDD.t43 VDD.n6668 0.000500648
R11428 VDD.n6670 VDD.n6669 0.000500648
R11429 VDD.n6669 VDD.t43 0.000500648
R11430 VDD.n856 VDD.n855 0.0005006
R11431 VDD.n1711 VDD.n1710 0.0005006
R11432 VDD.n2565 VDD.n2564 0.0005006
R11433 VDD.n3421 VDD.n3420 0.0005006
R11434 VDD.n5234 VDD.n5233 0.000500389
R11435 VDD.n3809 VDD.n3808 0.000500389
R11436 VDD.n3808 VDD.n3807 0.000500389
R11437 VDD.n3013 VDD.n3012 0.000500314
R11438 VDD.n2252 VDD.n1782 0.000500314
R11439 VDD.n1398 VDD.n928 0.000500314
R11440 VDD.n543 VDD.n73 0.000500314
R11441 VDD.n68 VDD.n67 0.000500314
R11442 VDD.n923 VDD.n922 0.000500314
R11443 VDD.n1777 VDD.n1776 0.000500314
R11444 VDD.n3417 VDD.n3416 0.000500314
R11445 VDD.n854 VDD.n2 0.000500311
R11446 VDD.n1709 VDD.n1 0.000500311
R11447 VDD.n2563 VDD.n0 0.000500311
R11448 VDD.n3419 VDD.n3418 0.000500311
R11449 VDD.n3039 VDD.n3038 0.000500201
R11450 VDD.n2557 VDD.n2556 0.000500201
R11451 VDD.n1703 VDD.n1702 0.000500201
R11452 VDD.n848 VDD.n847 0.000500201
R11453 VDD.n3627 VDD.n3626 0.000500031
R11454 VSS.n474 VSS.t46 1049.46
R11455 VSS.n300 VSS.t24 1045.16
R11456 VSS.t55 VSS.t57 984.947
R11457 VSS.t27 VSS.t53 984.947
R11458 VSS.t39 VSS.t36 671.51
R11459 VSS.t36 VSS.t12 671.51
R11460 VSS.t16 VSS.t6 671.51
R11461 VSS.t17 VSS.t16 671.51
R11462 VSS.t15 VSS.t17 671.51
R11463 VSS.t62 VSS.t61 671.51
R11464 VSS.t61 VSS.t8 671.51
R11465 VSS.t8 VSS.t10 671.51
R11466 VSS.t4 VSS.t2 671.51
R11467 VSS.t19 VSS.t4 671.51
R11468 VSS.t32 VSS.t19 671.51
R11469 VSS.n1379 VSS.t39 561.547
R11470 VSS.n731 VSS.t32 561.547
R11471 VSS.n485 VSS.t55 492.474
R11472 VSS.n485 VSS.t27 492.474
R11473 VSS.n1386 VSS.n1385 417.392
R11474 VSS.n1373 VSS.n1372 357.288
R11475 VSS.n1370 VSS.t14 335.755
R11476 VSS.n1370 VSS.t62 335.755
R11477 VSS.n1385 VSS.n1382 291.457
R11478 VSS.n994 VSS.t0 197.935
R11479 VSS.n487 VSS.n482 142.119
R11480 VSS.n495 VSS.n487 142.119
R11481 VSS.n986 VSS.t66 96.7682
R11482 VSS.n1435 VSS.t50 68.2323
R11483 VSS.n747 VSS.t34 68.2319
R11484 VSS.n338 VSS.t45 60.2505
R11485 VSS.n63 VSS.t26 60.2505
R11486 VSS.n176 VSS.t23 60.2505
R11487 VSS.n1840 VSS.t43 60.2505
R11488 VSS.n1726 VSS.t51 60.2505
R11489 VSS.n1865 VSS.t29 60.2505
R11490 VSS.n1951 VSS.t21 60.2505
R11491 VSS.n895 VSS.t41 60.2505
R11492 VSS.n786 VSS.t31 60.2505
R11493 VSS.n1522 VSS.t48 60.2505
R11494 VSS.n1506 VSS.t18 60.2505
R11495 VSS.n1252 VSS.t35 60.2505
R11496 VSS.n1236 VSS.t38 60.2505
R11497 VSS.n1383 VSS.t15 57.1814
R11498 VSS.n1380 VSS.n1379 48.3844
R11499 VSS.n977 VSS.n976 48.3844
R11500 VSS.n422 VSS.t47 35.3798
R11501 VSS.n261 VSS.t25 35.3798
R11502 VSS.t52 VSS.n1787 35.3798
R11503 VSS.t40 VSS.n1203 35.3798
R11504 VSS.n416 VSS.n415 31.4488
R11505 VSS.n423 VSS.n422 31.4488
R11506 VSS.n255 VSS.n254 31.4488
R11507 VSS.n262 VSS.n261 31.4488
R11508 VSS.n751 VSS.n750 31.4488
R11509 VSS.n1439 VSS.n1438 31.4488
R11510 VSS.n307 VSS.n303 30.0212
R11511 VSS.n298 VSS.n297 30.0212
R11512 VSS.n405 VSS.n404 27.5177
R11513 VSS.n434 VSS.n433 27.5177
R11514 VSS.n244 VSS.n243 27.5177
R11515 VSS.n273 VSS.n272 27.5177
R11516 VSS.n550 VSS.n549 27.5177
R11517 VSS.n761 VSS.n760 27.5177
R11518 VSS.n1450 VSS.n1449 27.5177
R11519 VSS.n1106 VSS.n1105 27.5177
R11520 VSS.n733 VSS.n732 26.5914
R11521 VSS.n394 VSS.n393 23.5867
R11522 VSS.n447 VSS.n446 23.5867
R11523 VSS.n233 VSS.n232 23.5867
R11524 VSS.n286 VSS.n285 23.5867
R11525 VSS.n575 VSS.n574 23.5867
R11526 VSS.n774 VSS.n773 23.5867
R11527 VSS.n1461 VSS.n1460 23.5867
R11528 VSS.n1117 VSS.n1116 23.5867
R11529 VSS.n1354 VSS.n1353 23.4593
R11530 VSS.n362 VSS.n361 21.6212
R11531 VSS.n201 VSS.n200 21.6212
R11532 VSS.n810 VSS.n809 21.6212
R11533 VSS.n1423 VSS.n1422 21.6212
R11534 VSS.n1077 VSS.n1076 21.6212
R11535 VSS.n383 VSS.n382 19.6557
R11536 VSS.n328 VSS.n327 19.6557
R11537 VSS.n222 VSS.n221 19.6557
R11538 VSS.n167 VSS.n166 19.6557
R11539 VSS.n830 VSS.n829 19.6557
R11540 VSS.n1474 VSS.n1473 19.6557
R11541 VSS.n1130 VSS.n1129 19.6557
R11542 VSS.n373 VSS.n372 17.6902
R11543 VSS.n313 VSS.n312 17.6902
R11544 VSS.n212 VSS.n211 17.6902
R11545 VSS.n155 VSS.n154 17.6902
R11546 VSS.n821 VSS.n820 17.6902
R11547 VSS.n1412 VSS.n1411 17.6902
R11548 VSS.n1069 VSS.n1068 17.6902
R11549 VSS.n372 VSS.n371 15.7246
R11550 VSS.n312 VSS.n311 15.7246
R11551 VSS.n211 VSS.n210 15.7246
R11552 VSS.n154 VSS.n153 15.7246
R11553 VSS.n820 VSS.n819 15.7246
R11554 VSS.n1411 VSS.n1410 15.7246
R11555 VSS.n1068 VSS.n1067 15.7246
R11556 VSS.n384 VSS.n383 13.7591
R11557 VSS.n329 VSS.n328 13.7591
R11558 VSS.n223 VSS.n222 13.7591
R11559 VSS.n168 VSS.n167 13.7591
R11560 VSS.n831 VSS.n830 13.7591
R11561 VSS.n1475 VSS.n1474 13.7591
R11562 VSS.n1131 VSS.n1130 13.7591
R11563 VSS.n146 VSS.n143 12.0077
R11564 VSS.n361 VSS.n360 11.7936
R11565 VSS.n303 VSS.n302 11.7936
R11566 VSS.n200 VSS.n199 11.7936
R11567 VSS.n297 VSS.n296 11.7936
R11568 VSS.n809 VSS.n808 11.7936
R11569 VSS.n1422 VSS.n1421 11.7936
R11570 VSS.n1076 VSS.n1075 11.7936
R11571 VSS.n395 VSS.n394 9.82809
R11572 VSS.n448 VSS.n447 9.82809
R11573 VSS.n234 VSS.n233 9.82809
R11574 VSS.n287 VSS.n286 9.82809
R11575 VSS.n576 VSS.n575 9.82809
R11576 VSS.n775 VSS.n774 9.82809
R11577 VSS.n1462 VSS.n1461 9.82809
R11578 VSS.n1118 VSS.n1117 9.82809
R11579 VSS.n348 VSS.n347 9.3005
R11580 VSS.n350 VSS.n349 9.3005
R11581 VSS.n346 VSS.n345 9.3005
R11582 VSS.n345 VSS.n344 9.3005
R11583 VSS.n439 VSS.n438 9.3005
R11584 VSS.n428 VSS.n427 9.3005
R11585 VSS.n412 VSS.n411 9.3005
R11586 VSS.n401 VSS.n400 9.3005
R11587 VSS.n390 VSS.n389 9.3005
R11588 VSS.n379 VSS.n378 9.3005
R11589 VSS.n368 VSS.n367 9.3005
R11590 VSS.n357 VSS.n356 9.3005
R11591 VSS.n355 VSS.n354 9.3005
R11592 VSS.n364 VSS.n363 9.3005
R11593 VSS.n363 VSS.n362 9.3005
R11594 VSS.n366 VSS.n365 9.3005
R11595 VSS.n375 VSS.n374 9.3005
R11596 VSS.n374 VSS.n373 9.3005
R11597 VSS.n377 VSS.n376 9.3005
R11598 VSS.n386 VSS.n385 9.3005
R11599 VSS.n385 VSS.n384 9.3005
R11600 VSS.n388 VSS.n387 9.3005
R11601 VSS.n397 VSS.n396 9.3005
R11602 VSS.n396 VSS.n395 9.3005
R11603 VSS.n399 VSS.n398 9.3005
R11604 VSS.n408 VSS.n407 9.3005
R11605 VSS.n407 VSS.n406 9.3005
R11606 VSS.n410 VSS.n409 9.3005
R11607 VSS.n419 VSS.n418 9.3005
R11608 VSS.n418 VSS.n417 9.3005
R11609 VSS.n426 VSS.n425 9.3005
R11610 VSS.n425 VSS.n424 9.3005
R11611 VSS.n430 VSS.n429 9.3005
R11612 VSS.n437 VSS.n436 9.3005
R11613 VSS.n436 VSS.n435 9.3005
R11614 VSS.n441 VSS.n440 9.3005
R11615 VSS.n449 VSS.n448 9.3005
R11616 VSS.n330 VSS.n329 9.3005
R11617 VSS.n314 VSS.n313 9.3005
R11618 VSS.n73 VSS.n72 9.3005
R11619 VSS.n75 VSS.n74 9.3005
R11620 VSS.n71 VSS.n70 9.3005
R11621 VSS.n70 VSS.n69 9.3005
R11622 VSS.n131 VSS.n130 9.3005
R11623 VSS.n124 VSS.n123 9.3005
R11624 VSS.n118 VSS.n117 9.3005
R11625 VSS.n111 VSS.n110 9.3005
R11626 VSS.n104 VSS.n103 9.3005
R11627 VSS.n97 VSS.n96 9.3005
R11628 VSS.n90 VSS.n89 9.3005
R11629 VSS.n83 VSS.n82 9.3005
R11630 VSS.n81 VSS.n80 9.3005
R11631 VSS.n86 VSS.n85 9.3005
R11632 VSS.n88 VSS.n87 9.3005
R11633 VSS.n93 VSS.n92 9.3005
R11634 VSS.n95 VSS.n94 9.3005
R11635 VSS.n100 VSS.n99 9.3005
R11636 VSS.n102 VSS.n101 9.3005
R11637 VSS.n107 VSS.n106 9.3005
R11638 VSS.n109 VSS.n108 9.3005
R11639 VSS.n114 VSS.n113 9.3005
R11640 VSS.n116 VSS.n115 9.3005
R11641 VSS.n120 VSS.n119 9.3005
R11642 VSS.n122 VSS.n121 9.3005
R11643 VSS.n126 VSS.n125 9.3005
R11644 VSS.n129 VSS.n128 9.3005
R11645 VSS.n133 VSS.n132 9.3005
R11646 VSS.n186 VSS.n185 9.3005
R11647 VSS.n188 VSS.n187 9.3005
R11648 VSS.n184 VSS.n183 9.3005
R11649 VSS.n183 VSS.n182 9.3005
R11650 VSS.n278 VSS.n277 9.3005
R11651 VSS.n267 VSS.n266 9.3005
R11652 VSS.n251 VSS.n250 9.3005
R11653 VSS.n240 VSS.n239 9.3005
R11654 VSS.n229 VSS.n228 9.3005
R11655 VSS.n218 VSS.n217 9.3005
R11656 VSS.n207 VSS.n206 9.3005
R11657 VSS.n196 VSS.n195 9.3005
R11658 VSS.n194 VSS.n193 9.3005
R11659 VSS.n203 VSS.n202 9.3005
R11660 VSS.n202 VSS.n201 9.3005
R11661 VSS.n205 VSS.n204 9.3005
R11662 VSS.n214 VSS.n213 9.3005
R11663 VSS.n213 VSS.n212 9.3005
R11664 VSS.n216 VSS.n215 9.3005
R11665 VSS.n225 VSS.n224 9.3005
R11666 VSS.n224 VSS.n223 9.3005
R11667 VSS.n227 VSS.n226 9.3005
R11668 VSS.n236 VSS.n235 9.3005
R11669 VSS.n235 VSS.n234 9.3005
R11670 VSS.n238 VSS.n237 9.3005
R11671 VSS.n247 VSS.n246 9.3005
R11672 VSS.n246 VSS.n245 9.3005
R11673 VSS.n249 VSS.n248 9.3005
R11674 VSS.n258 VSS.n257 9.3005
R11675 VSS.n257 VSS.n256 9.3005
R11676 VSS.n265 VSS.n264 9.3005
R11677 VSS.n264 VSS.n263 9.3005
R11678 VSS.n269 VSS.n268 9.3005
R11679 VSS.n276 VSS.n275 9.3005
R11680 VSS.n275 VSS.n274 9.3005
R11681 VSS.n280 VSS.n279 9.3005
R11682 VSS.n156 VSS.n155 9.3005
R11683 VSS.n288 VSS.n287 9.3005
R11684 VSS.n169 VSS.n168 9.3005
R11685 VSS.n1971 VSS.n1970 9.3005
R11686 VSS.n1978 VSS.n1977 9.3005
R11687 VSS.n1985 VSS.n1984 9.3005
R11688 VSS.n1983 VSS.n1982 9.3005
R11689 VSS.n1981 VSS.n1980 9.3005
R11690 VSS.n1976 VSS.n1975 9.3005
R11691 VSS.n1974 VSS.n1973 9.3005
R11692 VSS.n1969 VSS.n1968 9.3005
R11693 VSS.n1889 VSS.n1888 9.3005
R11694 VSS.n1893 VSS.n1892 9.3005
R11695 VSS.n1891 VSS.n1890 9.3005
R11696 VSS.n1896 VSS.n1895 9.3005
R11697 VSS.n1898 VSS.n1897 9.3005
R11698 VSS.n1900 VSS.n1899 9.3005
R11699 VSS.n1886 VSS.n1885 9.3005
R11700 VSS.n1884 VSS.n1883 9.3005
R11701 VSS.n1876 VSS.n1875 9.3005
R11702 VSS.n1857 VSS.n1856 9.3005
R11703 VSS.n1961 VSS.n1960 9.3005
R11704 VSS.n1963 VSS.n1962 9.3005
R11705 VSS.n1959 VSS.n1958 9.3005
R11706 VSS.n1958 VSS.n1957 9.3005
R11707 VSS.n1878 VSS.n1877 9.3005
R11708 VSS.n1874 VSS.n1873 9.3005
R11709 VSS.n1873 VSS.n1872 9.3005
R11710 VSS.n1864 VSS.n1863 9.3005
R11711 VSS.n1863 VSS.n1862 9.3005
R11712 VSS.n1948 VSS.n1947 9.3005
R11713 VSS.n1738 VSS.n1737 9.3005
R11714 VSS.n1736 VSS.n1735 9.3005
R11715 VSS.n1734 VSS.n1733 9.3005
R11716 VSS.n1733 VSS.n1732 9.3005
R11717 VSS.n1752 VSS.n1751 9.3005
R11718 VSS.n1748 VSS.n1747 9.3005
R11719 VSS.n1747 VSS.n1746 9.3005
R11720 VSS.n1750 VSS.n1749 9.3005
R11721 VSS.n1849 VSS.n1848 9.3005
R11722 VSS.n1848 VSS.n1847 9.3005
R11723 VSS.n1853 VSS.n1852 9.3005
R11724 VSS.n1851 VSS.n1850 9.3005
R11725 VSS.n1760 VSS.n1759 9.3005
R11726 VSS.n1767 VSS.n1766 9.3005
R11727 VSS.n1774 VSS.n1773 9.3005
R11728 VSS.n1772 VSS.n1771 9.3005
R11729 VSS.n1770 VSS.n1769 9.3005
R11730 VSS.n1765 VSS.n1764 9.3005
R11731 VSS.n1763 VSS.n1762 9.3005
R11732 VSS.n1758 VSS.n1757 9.3005
R11733 VSS.n562 VSS.n561 9.3005
R11734 VSS.n561 VSS.n560 9.3005
R11735 VSS.n564 VSS.n563 9.3005
R11736 VSS.n577 VSS.n576 9.3005
R11737 VSS.n566 VSS.n565 9.3005
R11738 VSS.n552 VSS.n551 9.3005
R11739 VSS.n903 VSS.n902 9.3005
R11740 VSS.n902 VSS.n901 9.3005
R11741 VSS.n907 VSS.n906 9.3005
R11742 VSS.n905 VSS.n904 9.3005
R11743 VSS.n914 VSS.n913 9.3005
R11744 VSS.n921 VSS.n920 9.3005
R11745 VSS.n928 VSS.n927 9.3005
R11746 VSS.n926 VSS.n925 9.3005
R11747 VSS.n924 VSS.n923 9.3005
R11748 VSS.n919 VSS.n918 9.3005
R11749 VSS.n917 VSS.n916 9.3005
R11750 VSS.n912 VSS.n911 9.3005
R11751 VSS.n756 VSS.n755 9.3005
R11752 VSS.n754 VSS.n753 9.3005
R11753 VSS.n753 VSS.n752 9.3005
R11754 VSS.n794 VSS.n793 9.3005
R11755 VSS.n793 VSS.n792 9.3005
R11756 VSS.n798 VSS.n797 9.3005
R11757 VSS.n796 VSS.n795 9.3005
R11758 VSS.n805 VSS.n804 9.3005
R11759 VSS.n816 VSS.n815 9.3005
R11760 VSS.n827 VSS.n826 9.3005
R11761 VSS.n832 VSS.n831 9.3005
R11762 VSS.n825 VSS.n824 9.3005
R11763 VSS.n823 VSS.n822 9.3005
R11764 VSS.n822 VSS.n821 9.3005
R11765 VSS.n814 VSS.n813 9.3005
R11766 VSS.n812 VSS.n811 9.3005
R11767 VSS.n811 VSS.n810 9.3005
R11768 VSS.n803 VSS.n802 9.3005
R11769 VSS.n758 VSS.n757 9.3005
R11770 VSS.n763 VSS.n762 9.3005
R11771 VSS.n776 VSS.n775 9.3005
R11772 VSS.n1518 VSS.n1517 9.3005
R11773 VSS.n1516 VSS.n1515 9.3005
R11774 VSS.n1514 VSS.n1513 9.3005
R11775 VSS.n1513 VSS.n1512 9.3005
R11776 VSS.n1534 VSS.n1533 9.3005
R11777 VSS.n1530 VSS.n1529 9.3005
R11778 VSS.n1529 VSS.n1528 9.3005
R11779 VSS.n1532 VSS.n1531 9.3005
R11780 VSS.n1542 VSS.n1541 9.3005
R11781 VSS.n1549 VSS.n1548 9.3005
R11782 VSS.n1556 VSS.n1555 9.3005
R11783 VSS.n1563 VSS.n1562 9.3005
R11784 VSS.n1570 VSS.n1569 9.3005
R11785 VSS.n1577 VSS.n1576 9.3005
R11786 VSS.n1583 VSS.n1582 9.3005
R11787 VSS.n1590 VSS.n1589 9.3005
R11788 VSS.n1597 VSS.n1596 9.3005
R11789 VSS.n1599 VSS.n1598 9.3005
R11790 VSS.n1595 VSS.n1594 9.3005
R11791 VSS.n1592 VSS.n1591 9.3005
R11792 VSS.n1588 VSS.n1587 9.3005
R11793 VSS.n1585 VSS.n1584 9.3005
R11794 VSS.n1581 VSS.n1580 9.3005
R11795 VSS.n1579 VSS.n1578 9.3005
R11796 VSS.n1575 VSS.n1574 9.3005
R11797 VSS.n1573 VSS.n1572 9.3005
R11798 VSS.n1568 VSS.n1567 9.3005
R11799 VSS.n1566 VSS.n1565 9.3005
R11800 VSS.n1561 VSS.n1560 9.3005
R11801 VSS.n1559 VSS.n1558 9.3005
R11802 VSS.n1554 VSS.n1553 9.3005
R11803 VSS.n1552 VSS.n1551 9.3005
R11804 VSS.n1547 VSS.n1546 9.3005
R11805 VSS.n1545 VSS.n1544 9.3005
R11806 VSS.n1540 VSS.n1539 9.3005
R11807 VSS.n1602 VSS.n1601 9.3005
R11808 VSS.n1444 VSS.n1443 9.3005
R11809 VSS.n1455 VSS.n1454 9.3005
R11810 VSS.n1442 VSS.n1441 9.3005
R11811 VSS.n1441 VSS.n1440 9.3005
R11812 VSS.n1446 VSS.n1445 9.3005
R11813 VSS.n1453 VSS.n1452 9.3005
R11814 VSS.n1452 VSS.n1451 9.3005
R11815 VSS.n1457 VSS.n1456 9.3005
R11816 VSS.n1464 VSS.n1463 9.3005
R11817 VSS.n1463 VSS.n1462 9.3005
R11818 VSS.n1468 VSS.n1467 9.3005
R11819 VSS.n1466 VSS.n1465 9.3005
R11820 VSS.n1424 VSS.n1423 9.3005
R11821 VSS.n1413 VSS.n1412 9.3005
R11822 VSS.n1476 VSS.n1475 9.3005
R11823 VSS.n1471 VSS.n1470 9.3005
R11824 VSS.n1100 VSS.n1099 9.3005
R11825 VSS.n1111 VSS.n1110 9.3005
R11826 VSS.n1098 VSS.n1097 9.3005
R11827 VSS.n1097 VSS.n1096 9.3005
R11828 VSS.n1102 VSS.n1101 9.3005
R11829 VSS.n1109 VSS.n1108 9.3005
R11830 VSS.n1108 VSS.n1107 9.3005
R11831 VSS.n1113 VSS.n1112 9.3005
R11832 VSS.n1120 VSS.n1119 9.3005
R11833 VSS.n1119 VSS.n1118 9.3005
R11834 VSS.n1124 VSS.n1123 9.3005
R11835 VSS.n1122 VSS.n1121 9.3005
R11836 VSS.n1070 VSS.n1069 9.3005
R11837 VSS.n1078 VSS.n1077 9.3005
R11838 VSS.n1132 VSS.n1131 9.3005
R11839 VSS.n1127 VSS.n1126 9.3005
R11840 VSS.n1248 VSS.n1247 9.3005
R11841 VSS.n1246 VSS.n1245 9.3005
R11842 VSS.n1244 VSS.n1243 9.3005
R11843 VSS.n1243 VSS.n1242 9.3005
R11844 VSS.n1264 VSS.n1263 9.3005
R11845 VSS.n1260 VSS.n1259 9.3005
R11846 VSS.n1259 VSS.n1258 9.3005
R11847 VSS.n1262 VSS.n1261 9.3005
R11848 VSS.n1272 VSS.n1271 9.3005
R11849 VSS.n1279 VSS.n1278 9.3005
R11850 VSS.n1286 VSS.n1285 9.3005
R11851 VSS.n1293 VSS.n1292 9.3005
R11852 VSS.n1300 VSS.n1299 9.3005
R11853 VSS.n1307 VSS.n1306 9.3005
R11854 VSS.n1313 VSS.n1312 9.3005
R11855 VSS.n1320 VSS.n1319 9.3005
R11856 VSS.n1327 VSS.n1326 9.3005
R11857 VSS.n1329 VSS.n1328 9.3005
R11858 VSS.n1325 VSS.n1324 9.3005
R11859 VSS.n1322 VSS.n1321 9.3005
R11860 VSS.n1318 VSS.n1317 9.3005
R11861 VSS.n1315 VSS.n1314 9.3005
R11862 VSS.n1311 VSS.n1310 9.3005
R11863 VSS.n1309 VSS.n1308 9.3005
R11864 VSS.n1305 VSS.n1304 9.3005
R11865 VSS.n1303 VSS.n1302 9.3005
R11866 VSS.n1298 VSS.n1297 9.3005
R11867 VSS.n1296 VSS.n1295 9.3005
R11868 VSS.n1291 VSS.n1290 9.3005
R11869 VSS.n1289 VSS.n1288 9.3005
R11870 VSS.n1284 VSS.n1283 9.3005
R11871 VSS.n1282 VSS.n1281 9.3005
R11872 VSS.n1277 VSS.n1276 9.3005
R11873 VSS.n1275 VSS.n1274 9.3005
R11874 VSS.n1270 VSS.n1269 9.3005
R11875 VSS.n1332 VSS.n1331 9.3005
R11876 VSS.n1035 VSS.n1034 9.3005
R11877 VSS.n1355 VSS.n1354 9.3005
R11878 VSS.n1365 VSS.n1362 9.19092
R11879 VSS.n967 VSS.n964 9.19092
R11880 VSS.n1866 VSS.n1865 8.76429
R11881 VSS.n1841 VSS.n1840 8.76429
R11882 VSS.n1357 VSS.n1356 8.44701
R11883 VSS.n343 VSS.n342 8.21641
R11884 VSS.n68 VSS.n67 8.21641
R11885 VSS.n181 VSS.n180 8.21641
R11886 VSS.n1731 VSS.n1730 8.21641
R11887 VSS.n1956 VSS.n1955 8.21641
R11888 VSS.n1871 VSS.n1870 8.21641
R11889 VSS.n1861 VSS.n1860 8.21641
R11890 VSS.n1745 VSS.n1744 8.21641
R11891 VSS.n1846 VSS.n1845 8.21641
R11892 VSS.n900 VSS.n899 8.21641
R11893 VSS.n791 VSS.n790 8.21641
R11894 VSS.n1511 VSS.n1510 8.21641
R11895 VSS.n1527 VSS.n1526 8.21641
R11896 VSS.n1241 VSS.n1240 8.21641
R11897 VSS.n1257 VSS.n1256 8.21641
R11898 VSS.n1361 VSS.n1358 7.69718
R11899 VSS.n957 VSS.n735 7.69718
R11900 VSS.n963 VSS.n958 7.69718
R11901 VSS.n1377 VSS.n1355 7.3129
R11902 VSS.n1727 VSS.n1726 6.92242
R11903 VSS.n1507 VSS.n1506 6.92242
R11904 VSS.n1237 VSS.n1236 6.92242
R11905 VSS.n64 VSS.n63 6.92012
R11906 VSS.n177 VSS.n176 6.92012
R11907 VSS.n1952 VSS.n1951 6.92012
R11908 VSS.n1523 VSS.n1522 6.92012
R11909 VSS.n1253 VSS.n1252 6.92012
R11910 VSS.n339 VSS.n338 6.92011
R11911 VSS.n896 VSS.n895 6.92007
R11912 VSS.n787 VSS.n786 6.92007
R11913 VSS.n972 VSS.n971 6.81049
R11914 VSS.n1400 VSS.n1399 6.81049
R11915 VSS.n734 VSS.n733 6.81049
R11916 VSS.n1417 VSS.n1416 6.55106
R11917 VSS.n1082 VSS.n1081 6.55006
R11918 VSS.n801 VSS.n800 6.43466
R11919 VSS.n353 VSS.n352 6.43466
R11920 VSS.n192 VSS.n191 6.43466
R11921 VSS.n414 VSS.n413 6.02403
R11922 VSS.n421 VSS.n420 6.02403
R11923 VSS.n253 VSS.n252 6.02403
R11924 VSS.n260 VSS.n259 6.02403
R11925 VSS.n558 VSS.n557 6.02403
R11926 VSS.n749 VSS.n748 6.02403
R11927 VSS.n1437 VSS.n1436 6.02403
R11928 VSS.n1094 VSS.n1093 6.02403
R11929 VSS.n406 VSS.n405 5.89705
R11930 VSS.n435 VSS.n434 5.89705
R11931 VSS.n245 VSS.n244 5.89705
R11932 VSS.n274 VSS.n273 5.89705
R11933 VSS.n551 VSS.n550 5.89705
R11934 VSS.n762 VSS.n761 5.89705
R11935 VSS.n1451 VSS.n1450 5.89705
R11936 VSS.n1107 VSS.n1106 5.89705
R11937 VSS.n341 VSS.n340 5.64756
R11938 VSS.n66 VSS.n65 5.64756
R11939 VSS.n179 VSS.n178 5.64756
R11940 VSS.n1729 VSS.n1728 5.64756
R11941 VSS.n1954 VSS.n1953 5.64756
R11942 VSS.n1869 VSS.n1868 5.64756
R11943 VSS.n1859 VSS.n1858 5.64756
R11944 VSS.n1743 VSS.n1742 5.64756
R11945 VSS.n1844 VSS.n1843 5.64756
R11946 VSS.n898 VSS.n897 5.64756
R11947 VSS.n789 VSS.n788 5.64756
R11948 VSS.n1509 VSS.n1508 5.64756
R11949 VSS.n1525 VSS.n1524 5.64756
R11950 VSS.n1239 VSS.n1238 5.64756
R11951 VSS.n1255 VSS.n1254 5.64756
R11952 VSS.n41 VSS.n40 5.61038
R11953 VSS.n146 VSS.n145 5.61038
R11954 VSS.n1143 VSS.n1142 5.39982
R11955 VSS.n1635 VSS.n1634 5.39151
R11956 VSS.n1488 VSS.n1487 5.39151
R11957 VSS.n1218 VSS.n1217 5.39151
R11958 VSS.n634 VSS.n633 5.39051
R11959 VSS.n659 VSS.n658 5.39051
R11960 VSS.n684 VSS.n683 5.39051
R11961 VSS.n709 VSS.n708 5.39051
R11962 VSS.n1193 VSS.n1192 5.39051
R11963 VSS.n1060 VSS.n1059 5.38802
R11964 VSS.n308 VSS.n307 5.3711
R11965 VSS.n299 VSS.n298 5.3711
R11966 VSS.n910 VSS.n909 5.28653
R11967 VSS.n79 VSS.n78 5.28613
R11968 VSS.n1756 VSS.n1755 5.2751
R11969 VSS.n1967 VSS.n1966 5.2751
R11970 VSS.n1882 VSS.n1881 5.2751
R11971 VSS.n1538 VSS.n1537 5.27461
R11972 VSS.n1268 VSS.n1267 5.27461
R11973 VSS.n403 VSS.n402 5.27109
R11974 VSS.n432 VSS.n431 5.27109
R11975 VSS.n242 VSS.n241 5.27109
R11976 VSS.n271 VSS.n270 5.27109
R11977 VSS.n1448 VSS.n1447 5.27109
R11978 VSS.n1104 VSS.n1103 5.27109
R11979 VSS.n646 VSS.n645 5.13412
R11980 VSS.n671 VSS.n670 5.13412
R11981 VSS.n1647 VSS.n1646 5.13412
R11982 VSS.n696 VSS.n695 5.13412
R11983 VSS.n723 VSS.n722 5.13412
R11984 VSS.n1208 VSS.n1207 5.13412
R11985 VSS.n988 VSS.n985 4.83275
R11986 VSS.n351 VSS.n337 4.76425
R11987 VSS.n77 VSS.n76 4.76425
R11988 VSS.n190 VSS.n189 4.76425
R11989 VSS.n1740 VSS.n1739 4.76425
R11990 VSS.n1964 VSS.n1950 4.76425
R11991 VSS.n1879 VSS.n1855 4.76425
R11992 VSS.n1949 VSS.n1946 4.76425
R11993 VSS.n1753 VSS.n1741 4.76425
R11994 VSS.n1854 VSS.n1839 4.76425
R11995 VSS.n908 VSS.n894 4.76425
R11996 VSS.n799 VSS.n785 4.76425
R11997 VSS.n1520 VSS.n1519 4.76425
R11998 VSS.n1535 VSS.n1521 4.76425
R11999 VSS.n1250 VSS.n1249 4.76425
R12000 VSS.n1265 VSS.n1251 4.76425
R12001 VSS.n754 VSS.n747 4.68469
R12002 VSS.n562 VSS.n556 4.68392
R12003 VSS.n1442 VSS.n1435 4.68392
R12004 VSS.n1098 VSS.n1092 4.68392
R12005 VSS.n1867 VSS.n1866 4.6505
R12006 VSS.n1842 VSS.n1841 4.6505
R12007 VSS.n36 VSS.n35 4.51815
R12008 VSS.n392 VSS.n391 4.51815
R12009 VSS.n445 VSS.n444 4.51815
R12010 VSS.n451 VSS.n450 4.51815
R12011 VSS.n139 VSS.n138 4.51815
R12012 VSS.n231 VSS.n230 4.51815
R12013 VSS.n284 VSS.n283 4.51815
R12014 VSS.n290 VSS.n289 4.51815
R12015 VSS.n555 VSS.n554 4.51815
R12016 VSS.n766 VSS.n765 4.51815
R12017 VSS.n1459 VSS.n1458 4.51815
R12018 VSS.n1115 VSS.n1114 4.51815
R12019 VSS.n37 VSS.n36 4.5005
R12020 VSS.n452 VSS.n451 4.5005
R12021 VSS.n140 VSS.n139 4.5005
R12022 VSS.n291 VSS.n290 4.5005
R12023 VSS.n50 VSS.n46 4.5005
R12024 VSS.n59 VSS.n58 4.5005
R12025 VSS.n172 VSS.n171 4.5005
R12026 VSS.n320 VSS.n316 4.5005
R12027 VSS.n333 VSS.n332 4.5005
R12028 VSS.n17 VSS.n13 4.5005
R12029 VSS.n26 VSS.n25 4.5005
R12030 VSS.n159 VSS.n158 4.5005
R12031 VSS.n1991 VSS.n1990 4.5005
R12032 VSS.n1906 VSS.n1905 4.5005
R12033 VSS.n1780 VSS.n1779 4.5005
R12034 VSS.n934 VSS.n933 4.5005
R12035 VSS.n836 VSS.n835 4.5005
R12036 VSS.n848 VSS.n844 4.5005
R12037 VSS.n852 VSS.n841 4.5005
R12038 VSS.n858 VSS.n857 4.5005
R12039 VSS.n864 VSS.n863 4.5005
R12040 VSS.n879 VSS.n878 4.5005
R12041 VSS.n883 VSS.n872 4.5005
R12042 VSS.n889 VSS.n888 4.5005
R12043 VSS.n892 VSS.n869 4.5005
R12044 VSS.n767 VSS.n766 4.5005
R12045 VSS.n771 VSS.n746 4.5005
R12046 VSS.n780 VSS.n779 4.5005
R12047 VSS.n783 VSS.n743 4.5005
R12048 VSS.n1062 VSS.n1058 4.5005
R12049 VSS.n1050 VSS.n1049 4.5005
R12050 VSS.n1040 VSS.n1039 4.5005
R12051 VSS.n1029 VSS.n1028 4.5005
R12052 VSS.n1024 VSS.n1023 4.5005
R12053 VSS.n1155 VSS.n1153 4.5005
R12054 VSS.n1162 VSS.n1161 4.5005
R12055 VSS.n1224 VSS.n1223 4.5005
R12056 VSS.n1234 VSS.n1233 4.5005
R12057 VSS.n1135 VSS.n1134 4.5005
R12058 VSS.n1084 VSS.n1080 4.5005
R12059 VSS.n1479 VSS.n1478 4.5005
R12060 VSS.n1494 VSS.n1493 4.5005
R12061 VSS.n1504 VSS.n1503 4.5005
R12062 VSS.n711 VSS.n707 4.5005
R12063 VSS.n686 VSS.n682 4.5005
R12064 VSS.n692 VSS.n678 4.5005
R12065 VSS.n1433 VSS.n1415 4.5005
R12066 VSS.n1427 VSS.n1426 4.5005
R12067 VSS.n717 VSS.n703 4.5005
R12068 VSS.n1643 VSS.n1629 4.5005
R12069 VSS.n661 VSS.n657 4.5005
R12070 VSS.n1637 VSS.n1633 4.5005
R12071 VSS.n1195 VSS.n1191 4.5005
R12072 VSS.n1201 VSS.n1187 4.5005
R12073 VSS.n1090 VSS.n1072 4.5005
R12074 VSS.n1145 VSS.n1141 4.5005
R12075 VSS.n636 VSS.n632 4.5005
R12076 VSS.n642 VSS.n628 4.5005
R12077 VSS.n667 VSS.n653 4.5005
R12078 VSS.n1608 VSS.n1607 4.5005
R12079 VSS.n1338 VSS.n1337 4.5005
R12080 VSS.n568 VSS.n555 4.5005
R12081 VSS.n572 VSS.n548 4.5005
R12082 VSS.n581 VSS.n580 4.5005
R12083 VSS.n587 VSS.n586 4.5005
R12084 VSS.n1932 VSS.n1909 4.5005
R12085 VSS.n2004 VSS.n2003 4.5005
R12086 VSS.n2008 VSS.n1997 4.5005
R12087 VSS.n2014 VSS.n2013 4.5005
R12088 VSS.n2017 VSS.n1994 4.5005
R12089 VSS.n1807 VSS.n1783 4.5005
R12090 VSS.n1804 VSS.n1803 4.5005
R12091 VSS.n1794 VSS.n1793 4.5005
R12092 VSS.n1798 VSS.n1786 4.5005
R12093 VSS.n1929 VSS.n1928 4.5005
R12094 VSS.n1919 VSS.n1918 4.5005
R12095 VSS.n1923 VSS.n1912 4.5005
R12096 VSS.n363 VSS.n359 4.14168
R12097 VSS.n306 VSS.n305 4.14168
R12098 VSS.n202 VSS.n198 4.14168
R12099 VSS.n295 VSS.n294 4.14168
R12100 VSS.n1783 VSS.n1782 4.14168
R12101 VSS.n1994 VSS.n1993 4.14168
R12102 VSS.n1909 VSS.n1908 4.14168
R12103 VSS.n586 VSS.n585 4.14168
R12104 VSS.n869 VSS.n868 4.14168
R12105 VSS.n863 VSS.n862 4.14168
R12106 VSS.n811 VSS.n807 4.14168
R12107 VSS.n743 VSS.n742 4.14168
R12108 VSS.n632 VSS.n630 4.14168
R12109 VSS.n657 VSS.n655 4.14168
R12110 VSS.n1633 VSS.n1631 4.14168
R12111 VSS.n682 VSS.n680 4.14168
R12112 VSS.n707 VSS.n705 4.14168
R12113 VSS.n1493 VSS.n1491 4.14168
R12114 VSS.n1424 VSS.n1420 4.14168
R12115 VSS.n1426 VSS.n1424 4.14168
R12116 VSS.n1078 VSS.n1074 4.14168
R12117 VSS.n1080 VSS.n1078 4.14168
R12118 VSS.n1223 VSS.n1221 4.14168
R12119 VSS.n1191 VSS.n1189 4.14168
R12120 VSS.n1141 VSS.n1139 4.14168
R12121 VSS.n1039 VSS.n1037 4.14168
R12122 VSS.n1058 VSS.n1056 4.14168
R12123 VSS.n25 VSS.n24 3.76521
R12124 VSS.n381 VSS.n380 3.76521
R12125 VSS.n326 VSS.n325 3.76521
R12126 VSS.n332 VSS.n331 3.76521
R12127 VSS.n58 VSS.n57 3.76521
R12128 VSS.n220 VSS.n219 3.76521
R12129 VSS.n165 VSS.n164 3.76521
R12130 VSS.n171 VSS.n170 3.76521
R12131 VSS.n1803 VSS.n1802 3.76521
R12132 VSS.n2013 VSS.n2012 3.76521
R12133 VSS.n1928 VSS.n1927 3.76521
R12134 VSS.n580 VSS.n579 3.76521
R12135 VSS.n888 VSS.n887 3.76521
R12136 VSS.n857 VSS.n856 3.76521
R12137 VSS.n779 VSS.n778 3.76521
R12138 VSS.n1601 VSS.n1600 3.76521
R12139 VSS.n1607 VSS.n1605 3.76521
R12140 VSS.n1470 VSS.n1469 3.76521
R12141 VSS.n1478 VSS.n1476 3.76521
R12142 VSS.n1126 VSS.n1125 3.76521
R12143 VSS.n1134 VSS.n1132 3.76521
R12144 VSS.n1331 VSS.n1330 3.76521
R12145 VSS.n1337 VSS.n1335 3.76521
R12146 VSS.n1014 VSS.n1012 3.49117
R12147 VSS.n903 VSS.n896 3.47842
R12148 VSS.n794 VSS.n787 3.47842
R12149 VSS.n1959 VSS.n1952 3.47756
R12150 VSS.n71 VSS.n64 3.47756
R12151 VSS.n184 VSS.n177 3.47756
R12152 VSS.n1530 VSS.n1523 3.47756
R12153 VSS.n1260 VSS.n1253 3.47756
R12154 VSS.n346 VSS.n339 3.47753
R12155 VSS.n1734 VSS.n1727 3.4767
R12156 VSS.n1514 VSS.n1507 3.4767
R12157 VSS.n1244 VSS.n1237 3.4767
R12158 VSS.n997 VSS.n993 3.41629
R12159 VSS.n13 VSS.n11 3.38874
R12160 VSS.n374 VSS.n370 3.38874
R12161 VSS.n314 VSS.n310 3.38874
R12162 VSS.n316 VSS.n314 3.38874
R12163 VSS.n46 VSS.n44 3.38874
R12164 VSS.n213 VSS.n209 3.38874
R12165 VSS.n156 VSS.n152 3.38874
R12166 VSS.n158 VSS.n156 3.38874
R12167 VSS.n822 VSS.n818 3.38874
R12168 VSS.n628 VSS.n626 3.38874
R12169 VSS.n653 VSS.n651 3.38874
R12170 VSS.n1629 VSS.n1627 3.38874
R12171 VSS.n678 VSS.n676 3.38874
R12172 VSS.n703 VSS.n701 3.38874
R12173 VSS.n1503 VSS.n1501 3.38874
R12174 VSS.n1413 VSS.n1409 3.38874
R12175 VSS.n1415 VSS.n1413 3.38874
R12176 VSS.n1070 VSS.n1066 3.38874
R12177 VSS.n1072 VSS.n1070 3.38874
R12178 VSS.n1233 VSS.n1231 3.38874
R12179 VSS.n1187 VSS.n1185 3.38874
R12180 VSS.n1153 VSS.n1151 3.38874
R12181 VSS.n1049 VSS.n1047 3.38874
R12182 VSS.n955 VSS.n738 3.33963
R12183 VSS.n955 VSS.n954 3.33963
R12184 VSS.n961 VSS.n960 3.33963
R12185 VSS.n1398 VSS.n734 3.33963
R12186 VSS.n1400 VSS.n1398 3.33963
R12187 VSS.n973 VSS.n972 3.33963
R12188 VSS.n30 VSS.t58 3.3065
R12189 VSS.n30 VSS.t56 3.3065
R12190 VSS.n143 VSS.t28 3.3065
R12191 VSS.n143 VSS.t54 3.3065
R12192 VSS.n1788 VSS.t52 3.3065
R12193 VSS.n1998 VSS.t22 3.3065
R12194 VSS.n1913 VSS.t44 3.3065
R12195 VSS.n1913 VSS.t30 3.3065
R12196 VSS.n873 VSS.t42 3.3065
R12197 VSS.n873 VSS.t60 3.3065
R12198 VSS.n845 VSS.t59 3.3065
R12199 VSS.n845 VSS.t33 3.3065
R12200 VSS.n644 VSS.t63 3.3065
R12201 VSS.n644 VSS.t68 3.3065
R12202 VSS.n669 VSS.t69 3.3065
R12203 VSS.n669 VSS.t65 3.3065
R12204 VSS.n1645 VSS.t70 3.3065
R12205 VSS.n1645 VSS.t9 3.3065
R12206 VSS.n694 VSS.t11 3.3065
R12207 VSS.n694 VSS.t3 3.3065
R12208 VSS.n721 VSS.t5 3.3065
R12209 VSS.n721 VSS.t20 3.3065
R12210 VSS.t20 VSS.n720 3.3065
R12211 VSS.n720 VSS.t49 3.3065
R12212 VSS.n1205 VSS.t40 3.3065
R12213 VSS.t37 VSS.n1205 3.3065
R12214 VSS.n1206 VSS.t37 3.3065
R12215 VSS.n1206 VSS.t13 3.3065
R12216 VSS.n1157 VSS.t7 3.3065
R12217 VSS.n1157 VSS.t64 3.3065
R12218 VSS.n1013 VSS.t67 3.3065
R12219 VSS.n1013 VSS.t1 3.3065
R12220 VSS.n1779 VSS.n1777 3.22952
R12221 VSS.n1990 VSS.n1988 3.22952
R12222 VSS.n1905 VSS.n1903 3.22952
R12223 VSS.n933 VSS.n931 3.22952
R12224 VSS.n734 VSS.n730 3.03311
R12225 VSS.n738 VSS.n737 3.03311
R12226 VSS.n972 VSS.n970 3.03311
R12227 VSS.n1401 VSS.n1400 3.03311
R12228 VSS.n960 VSS.n959 3.03311
R12229 VSS.n954 VSS.n953 3.03311
R12230 VSS.n592 VSS.n591 3.03311
R12231 VSS.n594 VSS.n593 3.03311
R12232 VSS.n597 VSS.n596 3.03311
R12233 VSS.n13 VSS.n12 3.01226
R12234 VSS.n370 VSS.n369 3.01226
R12235 VSS.n310 VSS.n309 3.01226
R12236 VSS.n316 VSS.n315 3.01226
R12237 VSS.n46 VSS.n45 3.01226
R12238 VSS.n209 VSS.n208 3.01226
R12239 VSS.n152 VSS.n151 3.01226
R12240 VSS.n158 VSS.n157 3.01226
R12241 VSS.n1779 VSS.n1778 3.01226
R12242 VSS.n1990 VSS.n1989 3.01226
R12243 VSS.n1905 VSS.n1904 3.01226
R12244 VSS.n933 VSS.n932 3.01226
R12245 VSS.n818 VSS.n817 3.01226
R12246 VSS.n835 VSS.n834 3.01226
R12247 VSS.n628 VSS.n627 3.01226
R12248 VSS.n653 VSS.n652 3.01226
R12249 VSS.n1629 VSS.n1628 3.01226
R12250 VSS.n678 VSS.n677 3.01226
R12251 VSS.n703 VSS.n702 3.01226
R12252 VSS.n1503 VSS.n1502 3.01226
R12253 VSS.n1409 VSS.n1408 3.01226
R12254 VSS.n1415 VSS.n1414 3.01226
R12255 VSS.n1066 VSS.n1065 3.01226
R12256 VSS.n1072 VSS.n1071 3.01226
R12257 VSS.n1233 VSS.n1232 3.01226
R12258 VSS.n1187 VSS.n1186 3.01226
R12259 VSS.n1153 VSS.n1152 3.01226
R12260 VSS.n1049 VSS.n1048 3.01226
R12261 VSS.n25 VSS.n23 2.63579
R12262 VSS.n385 VSS.n381 2.63579
R12263 VSS.n330 VSS.n326 2.63579
R12264 VSS.n332 VSS.n330 2.63579
R12265 VSS.n58 VSS.n56 2.63579
R12266 VSS.n224 VSS.n220 2.63579
R12267 VSS.n169 VSS.n165 2.63579
R12268 VSS.n171 VSS.n169 2.63579
R12269 VSS.n833 VSS.n832 2.63579
R12270 VSS.n1607 VSS.n1606 2.63579
R12271 VSS.n1478 VSS.n1477 2.63579
R12272 VSS.n1134 VSS.n1133 2.63579
R12273 VSS.n1337 VSS.n1336 2.63579
R12274 VSS.n1161 VSS.n1160 2.63579
R12275 VSS.n1023 VSS.n1019 2.63579
R12276 VSS.n1803 VSS.n1801 2.529
R12277 VSS.n2013 VSS.n2011 2.529
R12278 VSS.n1928 VSS.n1926 2.529
R12279 VSS.n888 VSS.n886 2.529
R12280 VSS.n857 VSS.n855 2.529
R12281 VSS.n590 VSS.n589 2.35698
R12282 VSS.n359 VSS.n358 2.25932
R12283 VSS.n305 VSS.n304 2.25932
R12284 VSS.n198 VSS.n197 2.25932
R12285 VSS.n294 VSS.n293 2.25932
R12286 VSS.n1785 VSS.n1784 2.25932
R12287 VSS.n1996 VSS.n1995 2.25932
R12288 VSS.n1911 VSS.n1910 2.25932
R12289 VSS.n547 VSS.n546 2.25932
R12290 VSS.n871 VSS.n870 2.25932
R12291 VSS.n840 VSS.n839 2.25932
R12292 VSS.n807 VSS.n806 2.25932
R12293 VSS.n745 VSS.n744 2.25932
R12294 VSS.n632 VSS.n631 2.25932
R12295 VSS.n657 VSS.n656 2.25932
R12296 VSS.n1633 VSS.n1632 2.25932
R12297 VSS.n682 VSS.n681 2.25932
R12298 VSS.n707 VSS.n706 2.25932
R12299 VSS.n1493 VSS.n1492 2.25932
R12300 VSS.n1420 VSS.n1419 2.25932
R12301 VSS.n1426 VSS.n1425 2.25932
R12302 VSS.n1074 VSS.n1073 2.25932
R12303 VSS.n1080 VSS.n1079 2.25932
R12304 VSS.n1223 VSS.n1222 2.25932
R12305 VSS.n1191 VSS.n1190 2.25932
R12306 VSS.n1141 VSS.n1140 2.25932
R12307 VSS.n1039 VSS.n1038 2.25932
R12308 VSS.n1058 VSS.n1057 2.25932
R12309 VSS.n496 VSS.n495 2.24394
R12310 VSS.n1034 VSS.n1033 2.24086
R12311 VSS.n417 VSS.n416 1.96602
R12312 VSS.n424 VSS.n423 1.96602
R12313 VSS.n256 VSS.n255 1.96602
R12314 VSS.n263 VSS.n262 1.96602
R12315 VSS.n560 VSS.n559 1.96602
R12316 VSS.n752 VSS.n751 1.96602
R12317 VSS.n1440 VSS.n1439 1.96602
R12318 VSS.n1096 VSS.n1095 1.96602
R12319 VSS.n36 VSS.n34 1.88285
R12320 VSS.n396 VSS.n392 1.88285
R12321 VSS.n449 VSS.n445 1.88285
R12322 VSS.n451 VSS.n449 1.88285
R12323 VSS.n139 VSS.n137 1.88285
R12324 VSS.n235 VSS.n231 1.88285
R12325 VSS.n288 VSS.n284 1.88285
R12326 VSS.n290 VSS.n288 1.88285
R12327 VSS.n578 VSS.n577 1.88285
R12328 VSS.n777 VSS.n776 1.88285
R12329 VSS.n1463 VSS.n1459 1.88285
R12330 VSS.n1119 VSS.n1115 1.88285
R12331 VSS.n1023 VSS.n1022 1.88285
R12332 VSS.n1793 VSS.n1792 1.82308
R12333 VSS.n2003 VSS.n2002 1.82308
R12334 VSS.n1918 VSS.n1917 1.82308
R12335 VSS.n878 VSS.n877 1.82308
R12336 VSS.n844 VSS.n843 1.82308
R12337 VSS.n1714 VSS.n1713 1.71198
R12338 VSS.n497 VSS.n496 1.70717
R12339 VSS.n1710 VSS.n1709 1.70597
R12340 VSS.n1716 VSS.n1691 1.70596
R12341 VSS.n1835 VSS.n617 1.70596
R12342 VSS.n1718 VSS.n621 1.70592
R12343 VSS.n2030 VSS.n2029 1.70592
R12344 VSS.n1696 VSS.n1695 1.70592
R12345 VSS.n2043 VSS.n538 1.7059
R12346 VSS.n2045 VSS.n8 1.70578
R12347 VSS.n1833 VSS.n1832 1.70567
R12348 VSS.n2041 VSS.n2040 1.70511
R12349 VSS.n1349 VSS.n1064 1.6655
R12350 VSS.n1014 VSS.n1013 1.60574
R12351 VSS.n720 VSS.n719 1.60111
R12352 VSS.n1205 VSS.n1204 1.60111
R12353 VSS.n143 VSS.n142 1.60111
R12354 VSS.n993 VSS.n988 1.59802
R12355 VSS.n32 VSS.n31 1.52198
R12356 VSS.n515 VSS.n42 1.51434
R12357 VSS.n506 VSS.n147 1.51434
R12358 VSS.n502 VSS.n299 1.51434
R12359 VSS.n466 VSS.n308 1.51289
R12360 VSS.n1028 VSS.n1027 1.50638
R12361 VSS.n1482 VSS.n1481 1.48392
R12362 VSS.n1616 VSS.n726 1.48392
R12363 VSS.n1621 VSS.n699 1.48392
R12364 VSS.n1212 VSS.n1211 1.48392
R12365 VSS.n1346 VSS.n1137 1.48392
R12366 VSS.n1661 VSS.n649 1.48392
R12367 VSS.n1656 VSS.n674 1.48392
R12368 VSS.n1341 VSS.n1340 1.48392
R12369 VSS.n1611 VSS.n1610 1.48392
R12370 VSS.n1651 VSS.n1650 1.48392
R12371 VSS.n1914 VSS.n1913 1.46886
R12372 VSS.n874 VSS.n873 1.46886
R12373 VSS.n1789 VSS.n1788 1.46879
R12374 VSS.n1999 VSS.n1998 1.46879
R12375 VSS.n846 VSS.n845 1.46878
R12376 VSS.n732 VSS.n731 1.46668
R12377 VSS.n1396 VSS.n977 1.46668
R12378 VSS.n976 VSS.n975 1.46668
R12379 VSS.n646 VSS.n644 1.41292
R12380 VSS.n671 VSS.n669 1.41292
R12381 VSS.n1647 VSS.n1645 1.41292
R12382 VSS.n696 VSS.n694 1.41292
R12383 VSS.n723 VSS.n721 1.41292
R12384 VSS.n1208 VSS.n1206 1.41292
R12385 VSS.n1165 VSS.n1164 1.34465
R12386 VSS.n1165 VSS.n1148 1.34235
R12387 VSS.n1823 VSS.n1822 1.13717
R12388 VSS.n1830 VSS.n1829 1.13717
R12389 VSS.n2026 VSS.n2025 1.13717
R12390 VSS.n1941 VSS.n1940 1.13717
R12391 VSS.n1816 VSS.n1815 1.13717
R12392 VSS.n615 VSS.n614 1.13717
R12393 VSS.n515 VSS.n38 1.13083
R12394 VSS.n506 VSS.n141 1.13027
R12395 VSS.n502 VSS.n292 1.13027
R12396 VSS.n466 VSS.n453 1.13002
R12397 VSS.n407 VSS.n403 1.12991
R12398 VSS.n436 VSS.n432 1.12991
R12399 VSS.n246 VSS.n242 1.12991
R12400 VSS.n275 VSS.n271 1.12991
R12401 VSS.n553 VSS.n552 1.12991
R12402 VSS.n764 VSS.n763 1.12991
R12403 VSS.n1452 VSS.n1448 1.12991
R12404 VSS.n1108 VSS.n1104 1.12991
R12405 VSS.n1021 VSS.n1020 1.12991
R12406 VSS.n1063 VSS.n1062 1.1255
R12407 VSS.n344 VSS.n343 1.09595
R12408 VSS.n69 VSS.n68 1.09595
R12409 VSS.n182 VSS.n181 1.09595
R12410 VSS.n1732 VSS.n1731 1.09595
R12411 VSS.n1957 VSS.n1956 1.09595
R12412 VSS.n1872 VSS.n1871 1.09595
R12413 VSS.n1862 VSS.n1861 1.09595
R12414 VSS.n1746 VSS.n1745 1.09595
R12415 VSS.n1847 VSS.n1846 1.09595
R12416 VSS.n901 VSS.n900 1.09595
R12417 VSS.n792 VSS.n791 1.09595
R12418 VSS.n1512 VSS.n1511 1.09595
R12419 VSS.n1528 VSS.n1527 1.09595
R12420 VSS.n1242 VSS.n1241 1.09595
R12421 VSS.n1258 VSS.n1257 1.09595
R12422 VSS.n1158 VSS.n1157 1.0555
R12423 VSS.n942 VSS.n866 0.903813
R12424 VSS.n2021 VSS.n2019 0.903813
R12425 VSS.n605 VSS.n590 0.903541
R12426 VSS.n938 VSS.n935 0.90354
R12427 VSS.n947 VSS.n837 0.90354
R12428 VSS.n472 VSS.n471 0.787987
R12429 VSS.n345 VSS.n341 0.753441
R12430 VSS.n70 VSS.n66 0.753441
R12431 VSS.n183 VSS.n179 0.753441
R12432 VSS.n1733 VSS.n1729 0.753441
R12433 VSS.n1958 VSS.n1954 0.753441
R12434 VSS.n1873 VSS.n1869 0.753441
R12435 VSS.n1863 VSS.n1859 0.753441
R12436 VSS.n1747 VSS.n1743 0.753441
R12437 VSS.n1848 VSS.n1844 0.753441
R12438 VSS.n580 VSS.n578 0.753441
R12439 VSS.n555 VSS.n553 0.753441
R12440 VSS.n902 VSS.n898 0.753441
R12441 VSS.n835 VSS.n833 0.753441
R12442 VSS.n779 VSS.n777 0.753441
R12443 VSS.n766 VSS.n764 0.753441
R12444 VSS.n793 VSS.n789 0.753441
R12445 VSS.n1513 VSS.n1509 0.753441
R12446 VSS.n1529 VSS.n1525 0.753441
R12447 VSS.n1243 VSS.n1239 0.753441
R12448 VSS.n1259 VSS.n1255 0.753441
R12449 VSS.n1022 VSS.n1021 0.753441
R12450 VSS.n1403 VSS.n1402 0.720975
R12451 VSS.n952 VSS.n951 0.720975
R12452 VSS.n1376 VSS.n1357 0.720717
R12453 VSS.n1940 VSS.n1934 0.707257
R12454 VSS.n1815 VSS.n1809 0.707257
R12455 VSS.n504 VSS.n503 0.682531
R12456 VSS.n940 VSS.n939 0.682531
R12457 VSS.n1659 VSS.n1658 0.682531
R12458 VSS.n1654 VSS.n1653 0.682531
R12459 VSS.n1624 VSS.n1623 0.682531
R12460 VSS.n1619 VSS.n1618 0.682531
R12461 VSS.n1682 VSS.n1679 0.6825
R12462 VSS.n1159 VSS.n1158 0.640088
R12463 VSS.n601 VSS.n598 0.614024
R12464 VSS.n866 VSS.n838 0.594417
R12465 VSS.n875 VSS.n874 0.575661
R12466 VSS.n2000 VSS.n1999 0.575335
R12467 VSS.n1790 VSS.n1789 0.574421
R12468 VSS.n1915 VSS.n1914 0.574409
R12469 VSS.n524 VSS.n523 0.568833
R12470 VSS.n847 VSS.n846 0.561441
R12471 VSS.n508 VSS.n507 0.534875
R12472 VSS.n1378 VSS.n1352 0.496624
R12473 VSS.n40 VSS.n39 0.461175
R12474 VSS.n145 VSS.n144 0.461175
R12475 VSS.n1762 VSS.n1761 0.461175
R12476 VSS.n1973 VSS.n1972 0.461175
R12477 VSS.n1888 VSS.n1887 0.461175
R12478 VSS.n916 VSS.n915 0.461175
R12479 VSS.n630 VSS.n629 0.461175
R12480 VSS.n655 VSS.n654 0.461175
R12481 VSS.n1631 VSS.n1630 0.461175
R12482 VSS.n680 VSS.n679 0.461175
R12483 VSS.n705 VSS.n704 0.461175
R12484 VSS.n1544 VSS.n1543 0.461175
R12485 VSS.n1491 VSS.n1490 0.461175
R12486 VSS.n1274 VSS.n1273 0.461175
R12487 VSS.n1221 VSS.n1220 0.461175
R12488 VSS.n1189 VSS.n1188 0.461175
R12489 VSS.n1139 VSS.n1138 0.461175
R12490 VSS.n1056 VSS.n1055 0.461175
R12491 VSS.n85 VSS.n84 0.460679
R12492 VSS.n1352 VSS.n1351 0.430441
R12493 VSS.n11 VSS.n10 0.430121
R12494 VSS.n44 VSS.n43 0.430121
R12495 VSS.n1769 VSS.n1768 0.430121
R12496 VSS.n1980 VSS.n1979 0.430121
R12497 VSS.n1895 VSS.n1894 0.430121
R12498 VSS.n923 VSS.n922 0.430121
R12499 VSS.n626 VSS.n625 0.430121
R12500 VSS.n651 VSS.n650 0.430121
R12501 VSS.n1627 VSS.n1626 0.430121
R12502 VSS.n676 VSS.n675 0.430121
R12503 VSS.n701 VSS.n700 0.430121
R12504 VSS.n1551 VSS.n1550 0.430121
R12505 VSS.n1501 VSS.n1500 0.430121
R12506 VSS.n1281 VSS.n1280 0.430121
R12507 VSS.n1231 VSS.n1230 0.430121
R12508 VSS.n1185 VSS.n1184 0.430121
R12509 VSS.n1151 VSS.n1150 0.430121
R12510 VSS.n1047 VSS.n1046 0.430121
R12511 VSS.n92 VSS.n91 0.429625
R12512 VSS.n353 VSS.n351 0.420318
R12513 VSS.n192 VSS.n190 0.420318
R12514 VSS.n801 VSS.n799 0.420318
R12515 VSS.n23 VSS.n22 0.398603
R12516 VSS.n56 VSS.n55 0.398603
R12517 VSS.n1558 VSS.n1557 0.398603
R12518 VSS.n1288 VSS.n1287 0.398603
R12519 VSS.n99 VSS.n98 0.398108
R12520 VSS.n469 VSS.n468 0.382531
R12521 VSS.n31 VSS.n30 0.378264
R12522 VSS.n418 VSS.n414 0.376971
R12523 VSS.n425 VSS.n421 0.376971
R12524 VSS.n257 VSS.n253 0.376971
R12525 VSS.n264 VSS.n260 0.376971
R12526 VSS.n1783 VSS.n1781 0.376971
R12527 VSS.n1786 VSS.n1785 0.376971
R12528 VSS.n1994 VSS.n1992 0.376971
R12529 VSS.n1997 VSS.n1996 0.376971
R12530 VSS.n1909 VSS.n1907 0.376971
R12531 VSS.n1912 VSS.n1911 0.376971
R12532 VSS.n586 VSS.n584 0.376971
R12533 VSS.n548 VSS.n547 0.376971
R12534 VSS.n561 VSS.n558 0.376971
R12535 VSS.n869 VSS.n867 0.376971
R12536 VSS.n872 VSS.n871 0.376971
R12537 VSS.n863 VSS.n861 0.376971
R12538 VSS.n841 VSS.n840 0.376971
R12539 VSS.n743 VSS.n741 0.376971
R12540 VSS.n746 VSS.n745 0.376971
R12541 VSS.n753 VSS.n749 0.376971
R12542 VSS.n1441 VSS.n1437 0.376971
R12543 VSS.n1097 VSS.n1094 0.376971
R12544 VSS.n137 VSS.n136 0.366615
R12545 VSS.n1565 VSS.n1564 0.366615
R12546 VSS.n1295 VSS.n1294 0.366615
R12547 VSS.n106 VSS.n105 0.366119
R12548 VSS.n1594 VSS.n1593 0.366119
R12549 VSS.n1324 VSS.n1323 0.366119
R12550 VSS.n307 VSS.n306 0.337513
R12551 VSS.n298 VSS.n295 0.337513
R12552 VSS.n128 VSS.n127 0.334147
R12553 VSS.n1572 VSS.n1571 0.334147
R12554 VSS.n1302 VSS.n1301 0.334147
R12555 VSS.n113 VSS.n112 0.333652
R12556 VSS.n1587 VSS.n1586 0.333652
R12557 VSS.n1317 VSS.n1316 0.333652
R12558 VSS.n945 VSS.n944 0.324719
R12559 VSS.n1344 VSS.n1343 0.324719
R12560 VSS.n1215 VSS.n1214 0.324719
R12561 VSS.n1614 VSS.n1613 0.324719
R12562 VSS.n1485 VSS.n1484 0.324719
R12563 VSS.n79 VSS.n77 0.316384
R12564 VSS.n910 VSS.n908 0.316384
R12565 VSS VSS.n499 0.313
R12566 VSS.n1349 VSS.n1348 0.298156
R12567 VSS.n42 VSS.n41 0.297854
R12568 VSS.n147 VSS.n146 0.297854
R12569 VSS.n672 VSS.n671 0.251319
R12570 VSS.n724 VSS.n723 0.251319
R12571 VSS.n1209 VSS.n1208 0.251319
R12572 VSS.n1648 VSS.n1647 0.251319
R12573 VSS.n697 VSS.n696 0.251319
R12574 VSS.n647 VSS.n646 0.251319
R12575 VSS.n2024 VSS.n2023 0.234094
R12576 VSS.n1015 VSS.n1014 0.23152
R12577 VSS.n1754 VSS.n1740 0.229427
R12578 VSS.n1754 VSS.n1753 0.229427
R12579 VSS.n1880 VSS.n1854 0.229427
R12580 VSS.n1880 VSS.n1879 0.229427
R12581 VSS.n1965 VSS.n1949 0.229427
R12582 VSS.n1965 VSS.n1964 0.229427
R12583 VSS.n1536 VSS.n1520 0.229427
R12584 VSS.n1536 VSS.n1535 0.229427
R12585 VSS.n1266 VSS.n1250 0.229427
R12586 VSS.n1266 VSS.n1265 0.229427
R12587 VSS.n1967 VSS.n1965 0.191391
R12588 VSS.n1882 VSS.n1880 0.191391
R12589 VSS.n1756 VSS.n1754 0.191391
R12590 VSS.n1538 VSS.n1536 0.191391
R12591 VSS.n1268 VSS.n1266 0.191391
R12592 VSS.n426 VSS.n419 0.190717
R12593 VSS.n122 VSS.n120 0.190717
R12594 VSS.n265 VSS.n258 0.190717
R12595 VSS.n1849 VSS.n1842 0.190717
R12596 VSS.n1874 VSS.n1867 0.190717
R12597 VSS.n1867 VSS.n1864 0.190717
R12598 VSS.n1581 VSS.n1579 0.190717
R12599 VSS.n1311 VSS.n1309 0.190717
R12600 VSS.n355 VSS.n353 0.164777
R12601 VSS.n194 VSS.n192 0.164777
R12602 VSS.n1969 VSS.n1967 0.164777
R12603 VSS.n1884 VSS.n1882 0.164777
R12604 VSS.n1758 VSS.n1756 0.164777
R12605 VSS.n803 VSS.n801 0.164777
R12606 VSS.n1540 VSS.n1538 0.164777
R12607 VSS.n1270 VSS.n1268 0.164777
R12608 VSS.n351 VSS.n350 0.15935
R12609 VSS.n77 VSS.n75 0.15935
R12610 VSS.n190 VSS.n188 0.15935
R12611 VSS.n1740 VSS.n1738 0.15935
R12612 VSS.n1753 VSS.n1752 0.15935
R12613 VSS.n1854 VSS.n1853 0.15935
R12614 VSS.n1879 VSS.n1878 0.15935
R12615 VSS.n1949 VSS.n1948 0.15935
R12616 VSS.n1964 VSS.n1963 0.15935
R12617 VSS.n908 VSS.n907 0.15935
R12618 VSS.n799 VSS.n798 0.15935
R12619 VSS.n1520 VSS.n1518 0.15935
R12620 VSS.n1535 VSS.n1534 0.15935
R12621 VSS.n1250 VSS.n1248 0.15935
R12622 VSS.n1265 VSS.n1264 0.15935
R12623 VSS.n1182 VSS.n1181 0.15675
R12624 VSS.n2032 VSS.n2031 0.149462
R12625 VSS.n366 VSS.n364 0.144522
R12626 VSS.n377 VSS.n375 0.144522
R12627 VSS.n388 VSS.n386 0.144522
R12628 VSS.n399 VSS.n397 0.144522
R12629 VSS.n410 VSS.n408 0.144522
R12630 VSS.n437 VSS.n430 0.144522
R12631 VSS.n88 VSS.n86 0.144522
R12632 VSS.n95 VSS.n93 0.144522
R12633 VSS.n102 VSS.n100 0.144522
R12634 VSS.n109 VSS.n107 0.144522
R12635 VSS.n116 VSS.n114 0.144522
R12636 VSS.n129 VSS.n126 0.144522
R12637 VSS.n205 VSS.n203 0.144522
R12638 VSS.n216 VSS.n214 0.144522
R12639 VSS.n227 VSS.n225 0.144522
R12640 VSS.n238 VSS.n236 0.144522
R12641 VSS.n249 VSS.n247 0.144522
R12642 VSS.n276 VSS.n269 0.144522
R12643 VSS.n1976 VSS.n1974 0.144522
R12644 VSS.n1983 VSS.n1981 0.144522
R12645 VSS.n1891 VSS.n1889 0.144522
R12646 VSS.n1898 VSS.n1896 0.144522
R12647 VSS.n1765 VSS.n1763 0.144522
R12648 VSS.n1772 VSS.n1770 0.144522
R12649 VSS.n919 VSS.n917 0.144522
R12650 VSS.n926 VSS.n924 0.144522
R12651 VSS.n814 VSS.n812 0.144522
R12652 VSS.n825 VSS.n823 0.144522
R12653 VSS.n1547 VSS.n1545 0.144522
R12654 VSS.n1554 VSS.n1552 0.144522
R12655 VSS.n1561 VSS.n1559 0.144522
R12656 VSS.n1568 VSS.n1566 0.144522
R12657 VSS.n1575 VSS.n1573 0.144522
R12658 VSS.n1588 VSS.n1585 0.144522
R12659 VSS.n1595 VSS.n1592 0.144522
R12660 VSS.n1453 VSS.n1446 0.144522
R12661 VSS.n1464 VSS.n1457 0.144522
R12662 VSS.n1109 VSS.n1102 0.144522
R12663 VSS.n1120 VSS.n1113 0.144522
R12664 VSS.n1277 VSS.n1275 0.144522
R12665 VSS.n1284 VSS.n1282 0.144522
R12666 VSS.n1291 VSS.n1289 0.144522
R12667 VSS.n1298 VSS.n1296 0.144522
R12668 VSS.n1305 VSS.n1303 0.144522
R12669 VSS.n1318 VSS.n1315 0.144522
R12670 VSS.n1325 VSS.n1322 0.144522
R12671 VSS.n81 VSS.n79 0.141804
R12672 VSS.n912 VSS.n910 0.141804
R12673 VSS.n1777 VSS.n1776 0.125448
R12674 VSS.n1988 VSS.n1987 0.125448
R12675 VSS.n1903 VSS.n1902 0.125448
R12676 VSS.n931 VSS.n930 0.125448
R12677 VSS.n1605 VSS.n1604 0.125448
R12678 VSS.n1335 VSS.n1334 0.125448
R12679 VSS.n1602 VSS.n1599 0.122443
R12680 VSS.n1471 VSS.n1468 0.122443
R12681 VSS.n1127 VSS.n1124 0.122443
R12682 VSS.n1332 VSS.n1329 0.122443
R12683 VSS VSS.n2046 0.11659
R12684 VSS.n949 VSS.n948 0.113781
R12685 VSS.n603 VSS.n602 0.113781
R12686 VSS.n442 VSS.n441 0.106563
R12687 VSS.n134 VSS.n133 0.106563
R12688 VSS.n281 VSS.n280 0.106563
R12689 VSS.n1801 VSS.n1800 0.0902327
R12690 VSS.n2011 VSS.n2010 0.0902327
R12691 VSS.n1926 VSS.n1925 0.0902327
R12692 VSS.n886 VSS.n885 0.0902327
R12693 VSS.n855 VSS.n854 0.0902327
R12694 VSS.n597 VSS.n595 0.0861908
R12695 VSS.n598 VSS.n597 0.0777426
R12696 VSS.n1148 VSS.n1147 0.07529
R12697 VSS.n935 VSS.n893 0.0699908
R12698 VSS.n837 VSS.n784 0.0699908
R12699 VSS.n590 VSS.n588 0.0699908
R12700 VSS.n2019 VSS.n2018 0.0695895
R12701 VSS.n866 VSS.n865 0.0695894
R12702 VSS.n953 VSS.n952 0.0683603
R12703 VSS.n1402 VSS.n1401 0.0683603
R12704 VSS.n759 VSS.n758 0.0679423
R12705 VSS.n567 VSS.n566 0.0676044
R12706 VSS.n500 VSS 0.066125
R12707 VSS VSS.n1405 0.066125
R12708 VSS.n1934 VSS.n1933 0.0638939
R12709 VSS.n1809 VSS.n1808 0.0638939
R12710 VSS.n598 VSS.n592 0.0636644
R12711 VSS.n16 VSS.n15 0.0618569
R12712 VSS.n49 VSS.n48 0.0618569
R12713 VSS.n150 VSS.n149 0.0618569
R12714 VSS.n319 VSS.n318 0.0615154
R12715 VSS.n674 VSS.n668 0.0611815
R12716 VSS.n726 VSS.n718 0.0611815
R12717 VSS.n1481 VSS.n1434 0.0611815
R12718 VSS.n1137 VSS.n1091 0.0611815
R12719 VSS.n1211 VSS.n1202 0.0611815
R12720 VSS.n699 VSS.n693 0.0611815
R12721 VSS.n649 VSS.n643 0.0611815
R12722 VSS.n1650 VSS.n1644 0.0608398
R12723 VSS.n1610 VSS.n1505 0.0608398
R12724 VSS.n1340 VSS.n1235 0.0608398
R12725 VSS.n573 VSS.n572 0.0604712
R12726 VSS.n640 VSS.n639 0.0584854
R12727 VSS.n665 VSS.n664 0.0584854
R12728 VSS.n1641 VSS.n1640 0.0584854
R12729 VSS.n690 VSS.n689 0.0584854
R12730 VSS.n715 VSS.n714 0.0584854
R12731 VSS.n1498 VSS.n1497 0.0584854
R12732 VSS.n1431 VSS.n1430 0.0584854
R12733 VSS.n1088 VSS.n1087 0.0584854
R12734 VSS.n1228 VSS.n1227 0.0584854
R12735 VSS.n1199 VSS.n1198 0.0584854
R12736 VSS.n737 VSS.n736 0.0566413
R12737 VSS.n730 VSS.n729 0.0566413
R12738 VSS.n595 VSS.n594 0.0566413
R12739 VSS.n20 VSS.n19 0.0565323
R12740 VSS.n323 VSS.n322 0.0565323
R12741 VSS.n53 VSS.n52 0.0565323
R12742 VSS.n162 VSS.n161 0.0565323
R12743 VSS.n1164 VSS.n1156 0.0558464
R12744 VSS.n1792 VSS.n1791 0.0547459
R12745 VSS.n2002 VSS.n2001 0.0547459
R12746 VSS.n1917 VSS.n1916 0.0547459
R12747 VSS.n877 VSS.n876 0.0547459
R12748 VSS.n843 VSS.n842 0.0547459
R12749 VSS.n1004 VSS.n1003 0.053
R12750 VSS.n29 VSS.n28 0.0526261
R12751 VSS.n28 VSS.n27 0.0526261
R12752 VSS.n336 VSS.n335 0.0526261
R12753 VSS.n335 VSS.n334 0.0526261
R12754 VSS.n62 VSS.n61 0.0526261
R12755 VSS.n61 VSS.n60 0.0526261
R12756 VSS.n175 VSS.n174 0.0526261
R12757 VSS.n174 VSS.n173 0.0526261
R12758 VSS.n1164 VSS.n1163 0.0502162
R12759 VSS.n1664 VSS.n1663 0.0497188
R12760 VSS.n1035 VSS.n1032 0.0493281
R12761 VSS.n1044 VSS.n1043 0.0493281
R12762 VSS.n1053 VSS.n1052 0.0493281
R12763 VSS.n1406 VSS 0.0489375
R12764 VSS.n21 VSS.n20 0.0487198
R12765 VSS.n324 VSS.n323 0.0487198
R12766 VSS.n54 VSS.n53 0.0487198
R12767 VSS.n163 VSS.n162 0.0487198
R12768 VSS.n608 VSS.n607 0.0481562
R12769 VSS.n639 VSS.n638 0.0467667
R12770 VSS.n664 VSS.n663 0.0467667
R12771 VSS.n1640 VSS.n1639 0.0467667
R12772 VSS.n689 VSS.n688 0.0467667
R12773 VSS.n714 VSS.n713 0.0467667
R12774 VSS.n1497 VSS.n1496 0.0467667
R12775 VSS.n1430 VSS.n1429 0.0467667
R12776 VSS.n1087 VSS.n1086 0.0467667
R12777 VSS.n1227 VSS.n1226 0.0467667
R12778 VSS.n1198 VSS.n1197 0.0467667
R12779 VSS.n1799 VSS.n1798 0.0464244
R12780 VSS.n1924 VSS.n1923 0.0464244
R12781 VSS.n853 VSS.n852 0.0461141
R12782 VSS.n884 VSS.n883 0.0461141
R12783 VSS.n772 VSS.n771 0.0461141
R12784 VSS.n2009 VSS.n2008 0.045605
R12785 VSS.n2014 VSS.n2009 0.0454086
R12786 VSS.n1650 VSS.n1649 0.0449804
R12787 VSS.n1610 VSS.n1609 0.0449804
R12788 VSS.n1340 VSS.n1339 0.0449804
R12789 VSS.n889 VSS.n884 0.0448907
R12790 VSS.n858 VSS.n853 0.0448907
R12791 VSS.n780 VSS.n772 0.0448907
R12792 VSS.n649 VSS.n648 0.04464
R12793 VSS.n674 VSS.n673 0.04464
R12794 VSS.n699 VSS.n698 0.04464
R12795 VSS.n726 VSS.n725 0.04464
R12796 VSS.n1481 VSS.n1480 0.04464
R12797 VSS.n1137 VSS.n1136 0.04464
R12798 VSS.n1211 VSS.n1210 0.04464
R12799 VSS.n1929 VSS.n1924 0.0445792
R12800 VSS.n1804 VSS.n1799 0.0445792
R12801 VSS.n318 VSS.n317 0.0443642
R12802 VSS.n15 VSS.n14 0.0440244
R12803 VSS.n48 VSS.n47 0.0440244
R12804 VSS.n149 VSS.n148 0.0440244
R12805 VSS.n412 VSS.n410 0.0439783
R12806 VSS.n430 VSS.n428 0.0439783
R12807 VSS.n118 VSS.n116 0.0439783
R12808 VSS.n126 VSS.n124 0.0439783
R12809 VSS.n251 VSS.n249 0.0439783
R12810 VSS.n269 VSS.n267 0.0439783
R12811 VSS.n566 VSS.n564 0.0439783
R12812 VSS.n758 VSS.n756 0.0439783
R12813 VSS.n1577 VSS.n1575 0.0439783
R12814 VSS.n1585 VSS.n1583 0.0439783
R12815 VSS.n1446 VSS.n1444 0.0439783
R12816 VSS.n1102 VSS.n1100 0.0439783
R12817 VSS.n1307 VSS.n1305 0.0439783
R12818 VSS.n1315 VSS.n1313 0.0439783
R12819 VSS.n462 VSS.n461 0.0434688
R12820 VSS.n461 VSS.n460 0.0434688
R12821 VSS.n460 VSS.n459 0.0434688
R12822 VSS.n459 VSS.n458 0.0434688
R12823 VSS.n458 VSS.n457 0.0434688
R12824 VSS.n457 VSS.n456 0.0434688
R12825 VSS.n454 VSS.n9 0.0434688
R12826 VSS.n523 VSS.n9 0.0434688
R12827 VSS.n523 VSS.n522 0.0434688
R12828 VSS.n522 VSS.n521 0.0434688
R12829 VSS.n521 VSS.n520 0.0434688
R12830 VSS.n520 VSS.n519 0.0434688
R12831 VSS.n519 VSS.n518 0.0434688
R12832 VSS.n512 VSS.n511 0.0434688
R12833 VSS.n1180 VSS.n1179 0.0434688
R12834 VSS.n1179 VSS.n1178 0.0434688
R12835 VSS.n1178 VSS.n1177 0.0434688
R12836 VSS.n1177 VSS.n1176 0.0434688
R12837 VSS.n1174 VSS.n1173 0.0434688
R12838 VSS.n1173 VSS.n1172 0.0434688
R12839 VSS.n1172 VSS.n1171 0.0434688
R12840 VSS.n1171 VSS.n1170 0.0434688
R12841 VSS.n1170 VSS.n1169 0.0434688
R12842 VSS.n1169 VSS.n1168 0.0434688
R12843 VSS.n1679 VSS.n1678 0.0434688
R12844 VSS.n1678 VSS.n1677 0.0434688
R12845 VSS.n1677 VSS.n1676 0.0434688
R12846 VSS.n1676 VSS.n1675 0.0434688
R12847 VSS.n1675 VSS.n1674 0.0434688
R12848 VSS.n1674 VSS.n1673 0.0434688
R12849 VSS.n1671 VSS.n1670 0.0434688
R12850 VSS.n1670 VSS.n1669 0.0434688
R12851 VSS.n1669 VSS.n1668 0.0434688
R12852 VSS.n1668 VSS.n1667 0.0434688
R12853 VSS.n1667 VSS.n1666 0.0434688
R12854 VSS.n1666 VSS.n1665 0.0434688
R12855 VSS.n610 VSS.n609 0.0434688
R12856 VSS.n611 VSS.n610 0.0434688
R12857 VSS.n613 VSS.n612 0.0434688
R12858 VSS.n1820 VSS.n1819 0.0434688
R12859 VSS.n1828 VSS.n1827 0.0434688
R12860 VSS.n1945 VSS.n1944 0.0434688
R12861 VSS.n1176 VSS.n1175 0.0426875
R12862 VSS.n848 VSS.n847 0.0419945
R12863 VSS.n1936 VSS.n1935 0.0419063
R12864 VSS.n1024 VSS.n1018 0.0415156
R12865 VSS.n350 VSS.n348 0.0412609
R12866 VSS.n75 VSS.n73 0.0412609
R12867 VSS.n188 VSS.n186 0.0412609
R12868 VSS.n1738 VSS.n1736 0.0412609
R12869 VSS.n1752 VSS.n1750 0.0412609
R12870 VSS.n1853 VSS.n1851 0.0412609
R12871 VSS.n1878 VSS.n1876 0.0412609
R12872 VSS.n1963 VSS.n1961 0.0412609
R12873 VSS.n907 VSS.n905 0.0412609
R12874 VSS.n798 VSS.n796 0.0412609
R12875 VSS.n1518 VSS.n1516 0.0412609
R12876 VSS.n1534 VSS.n1532 0.0412609
R12877 VSS.n1248 VSS.n1246 0.0412609
R12878 VSS.n1264 VSS.n1262 0.0412609
R12879 VSS.n1822 VSS.n1821 0.041125
R12880 VSS.n401 VSS.n399 0.0385435
R12881 VSS.n441 VSS.n439 0.0385435
R12882 VSS.n111 VSS.n109 0.0385435
R12883 VSS.n133 VSS.n131 0.0385435
R12884 VSS.n240 VSS.n238 0.0385435
R12885 VSS.n280 VSS.n278 0.0385435
R12886 VSS.n1570 VSS.n1568 0.0385435
R12887 VSS.n1592 VSS.n1590 0.0385435
R12888 VSS.n1457 VSS.n1455 0.0385435
R12889 VSS.n1113 VSS.n1111 0.0385435
R12890 VSS.n1300 VSS.n1298 0.0385435
R12891 VSS.n1322 VSS.n1320 0.0385435
R12892 VSS.n1181 VSS.n1180 0.038
R12893 VSS.n1665 VSS.n1664 0.038
R12894 VSS.n510 VSS.n509 0.0372187
R12895 VSS.n1679 VSS.n624 0.0372187
R12896 VSS.n1017 VSS.n1016 0.0356562
R12897 VSS.n1052 VSS.n1051 0.0356562
R12898 VSS.n614 VSS.n613 0.0356562
R12899 VSS.n1829 VSS.n1828 0.0356562
R12900 VSS.n609 VSS.n608 0.034875
R12901 VSS.n2025 VSS.n2024 0.034875
R12902 VSS.n1673 VSS.n1672 0.0340938
R12903 VSS.n390 VSS.n388 0.0331087
R12904 VSS.n104 VSS.n102 0.0331087
R12905 VSS.n229 VSS.n227 0.0331087
R12906 VSS.n1563 VSS.n1561 0.0331087
R12907 VSS.n1599 VSS.n1597 0.0331087
R12908 VSS.n1468 VSS.n1466 0.0331087
R12909 VSS.n1124 VSS.n1122 0.0331087
R12910 VSS.n1293 VSS.n1291 0.0331087
R12911 VSS.n1329 VSS.n1327 0.0331087
R12912 VSS.n513 VSS.n512 0.0325312
R12913 VSS.n1061 VSS.n1060 0.03175
R12914 VSS.n1007 VSS.n1006 0.03175
R12915 VSS.n1011 VSS.n1010 0.03175
R12916 VSS.n464 VSS.n463 0.0309688
R12917 VSS.n456 VSS.n455 0.0309688
R12918 VSS.n1148 VSS.n1146 0.0306452
R12919 VSS.n1794 VSS.n1790 0.0304205
R12920 VSS.n1919 VSS.n1915 0.0304205
R12921 VSS.n364 VSS.n357 0.0303913
R12922 VSS.n86 VSS.n83 0.0303913
R12923 VSS.n203 VSS.n196 0.0303913
R12924 VSS.n1974 VSS.n1971 0.0303913
R12925 VSS.n1889 VSS.n1886 0.0303913
R12926 VSS.n1763 VSS.n1760 0.0303913
R12927 VSS.n917 VSS.n914 0.0303913
R12928 VSS.n812 VSS.n805 0.0303913
R12929 VSS.n1545 VSS.n1542 0.0303913
R12930 VSS.n1275 VSS.n1272 0.0303913
R12931 VSS.n463 VSS.n462 0.0301875
R12932 VSS.n509 VSS.n508 0.0301875
R12933 VSS.n581 VSS.n573 0.0301368
R12934 VSS.n635 VSS.n634 0.0297969
R12935 VSS.n660 VSS.n659 0.0297969
R12936 VSS.n1636 VSS.n1635 0.0297969
R12937 VSS.n685 VSS.n684 0.0297969
R12938 VSS.n710 VSS.n709 0.0297969
R12939 VSS.n1489 VSS.n1488 0.0297969
R12940 VSS.n1418 VSS.n1417 0.0297969
R12941 VSS.n1083 VSS.n1082 0.0297969
R12942 VSS.n1219 VSS.n1218 0.0297969
R12943 VSS.n1194 VSS.n1193 0.0297969
R12944 VSS.n1001 VSS.n1000 0.02925
R12945 VSS.n568 VSS.n567 0.0288505
R12946 VSS.n2004 VSS.n2000 0.0288505
R12947 VSS.n879 VSS.n875 0.0285117
R12948 VSS.n767 VSS.n759 0.0285117
R12949 VSS.n1064 VSS.n1063 0.028
R12950 VSS.n1043 VSS.n1042 0.0278438
R12951 VSS.n1811 VSS.n1810 0.0278438
R12952 VSS.n379 VSS.n377 0.0276739
R12953 VSS.n97 VSS.n95 0.0276739
R12954 VSS.n218 VSS.n216 0.0276739
R12955 VSS.n1556 VSS.n1554 0.0276739
R12956 VSS.n1286 VSS.n1284 0.0276739
R12957 VSS.n1000 VSS.n999 0.02675
R12958 VSS.n1063 VSS.n1011 0.02675
R12959 VSS.n1029 VSS.n1026 0.0258906
R12960 VSS.n1934 VSS.n1906 0.0250149
R12961 VSS.n1809 VSS.n1780 0.0250149
R12962 VSS.n375 VSS.n368 0.0249565
R12963 VSS.n93 VSS.n90 0.0249565
R12964 VSS.n214 VSS.n207 0.0249565
R12965 VSS.n1981 VSS.n1978 0.0249565
R12966 VSS.n1985 VSS.n1983 0.0249565
R12967 VSS.n1896 VSS.n1893 0.0249565
R12968 VSS.n1900 VSS.n1898 0.0249565
R12969 VSS.n1770 VSS.n1767 0.0249565
R12970 VSS.n1774 VSS.n1772 0.0249565
R12971 VSS.n924 VSS.n921 0.0249565
R12972 VSS.n928 VSS.n926 0.0249565
R12973 VSS.n823 VSS.n816 0.0249565
R12974 VSS.n827 VSS.n825 0.0249565
R12975 VSS.n1552 VSS.n1549 0.0249565
R12976 VSS.n1282 VSS.n1279 0.0249565
R12977 VSS.n33 VSS.n32 0.0239375
R12978 VSS.n443 VSS.n442 0.0239375
R12979 VSS.n135 VSS.n134 0.0239375
R12980 VSS.n282 VSS.n281 0.0239375
R12981 VSS.n1031 VSS.n1030 0.0239375
R12982 VSS.n1350 VSS.n997 0.0232776
R12983 VSS.n1010 VSS.n1009 0.023
R12984 VSS.n1144 VSS.n1143 0.022459
R12985 VSS.n1720 VSS.n1719 0.0223109
R12986 VSS.n368 VSS.n366 0.0222391
R12987 VSS.n90 VSS.n88 0.0222391
R12988 VSS.n207 VSS.n205 0.0222391
R12989 VSS.n1978 VSS.n1976 0.0222391
R12990 VSS.n1986 VSS.n1985 0.0222391
R12991 VSS.n1893 VSS.n1891 0.0222391
R12992 VSS.n1901 VSS.n1900 0.0222391
R12993 VSS.n1767 VSS.n1765 0.0222391
R12994 VSS.n1775 VSS.n1774 0.0222391
R12995 VSS.n921 VSS.n919 0.0222391
R12996 VSS.n929 VSS.n928 0.0222391
R12997 VSS.n816 VSS.n814 0.0222391
R12998 VSS.n828 VSS.n827 0.0222391
R12999 VSS.n1549 VSS.n1547 0.0222391
R13000 VSS.n1279 VSS.n1277 0.0222391
R13001 VSS.n2017 VSS.n2016 0.0219844
R13002 VSS.n2006 VSS.n2005 0.0219844
R13003 VSS.n1932 VSS.n1931 0.0219844
R13004 VSS.n1921 VSS.n1920 0.0219844
R13005 VSS.n1807 VSS.n1806 0.0219844
R13006 VSS.n1796 VSS.n1795 0.0219844
R13007 VSS.n587 VSS.n583 0.0219844
R13008 VSS.n570 VSS.n569 0.0219844
R13009 VSS.n892 VSS.n891 0.0219844
R13010 VSS.n881 VSS.n880 0.0219844
R13011 VSS.n864 VSS.n860 0.0219844
R13012 VSS.n850 VSS.n849 0.0219844
R13013 VSS.n783 VSS.n782 0.0219844
R13014 VSS.n769 VSS.n768 0.0219844
R13015 VSS.n1146 VSS.n1145 0.0219844
R13016 VSS.n1040 VSS.n1036 0.0219844
R13017 VSS.n1062 VSS.n1054 0.0219844
R13018 VSS.n1008 VSS.n1007 0.02175
R13019 VSS.n518 VSS.n517 0.0208125
R13020 VSS.n638 VSS.n637 0.0205304
R13021 VSS.n1639 VSS.n1638 0.0205304
R13022 VSS.n688 VSS.n687 0.0205304
R13023 VSS.n1496 VSS.n1495 0.0205304
R13024 VSS.n1226 VSS.n1225 0.0205304
R13025 VSS.n1197 VSS.n1196 0.0205304
R13026 VSS.n1002 VSS.n1001 0.0205
R13027 VSS.n453 VSS.n336 0.0204768
R13028 VSS.n141 VSS.n62 0.0204759
R13029 VSS.n292 VSS.n175 0.0204759
R13030 VSS.n38 VSS.n29 0.020474
R13031 VSS.n26 VSS.n21 0.0200312
R13032 VSS.n333 VSS.n324 0.0200312
R13033 VSS.n59 VSS.n54 0.0200312
R13034 VSS.n172 VSS.n163 0.0200312
R13035 VSS.n1608 VSS.n1603 0.0200312
R13036 VSS.n1479 VSS.n1472 0.0200312
R13037 VSS.n1135 VSS.n1128 0.0200312
R13038 VSS.n1338 VSS.n1333 0.0200312
R13039 VSS.n1032 VSS.n1031 0.0200312
R13040 VSS.n1054 VSS.n1053 0.0200312
R13041 VSS.n386 VSS.n379 0.0195217
R13042 VSS.n100 VSS.n97 0.0195217
R13043 VSS.n225 VSS.n218 0.0195217
R13044 VSS.n1559 VSS.n1556 0.0195217
R13045 VSS.n1289 VSS.n1286 0.0195217
R13046 VSS.n2019 VSS.n1991 0.0188525
R13047 VSS.n1991 VSS.n1986 0.0188424
R13048 VSS.n1906 VSS.n1901 0.0188424
R13049 VSS.n1780 VSS.n1775 0.0188424
R13050 VSS.n934 VSS.n929 0.0188424
R13051 VSS.n836 VSS.n828 0.0188424
R13052 VSS.n935 VSS.n934 0.0184465
R13053 VSS.n837 VSS.n836 0.0184465
R13054 VSS.n643 VSS.n642 0.0180781
R13055 VSS.n668 VSS.n667 0.0180781
R13056 VSS.n663 VSS.n662 0.0180781
R13057 VSS.n1644 VSS.n1643 0.0180781
R13058 VSS.n693 VSS.n692 0.0180781
R13059 VSS.n718 VSS.n717 0.0180781
R13060 VSS.n713 VSS.n712 0.0180781
R13061 VSS.n1505 VSS.n1504 0.0180781
R13062 VSS.n1434 VSS.n1433 0.0180781
R13063 VSS.n1429 VSS.n1428 0.0180781
R13064 VSS.n1091 VSS.n1090 0.0180781
R13065 VSS.n1086 VSS.n1085 0.0180781
R13066 VSS.n1235 VSS.n1234 0.0180781
R13067 VSS.n1202 VSS.n1201 0.0180781
R13068 VSS.n1156 VSS.n1155 0.0180781
R13069 VSS.n1050 VSS.n1045 0.0180781
R13070 VSS.n1006 VSS.n1005 0.018
R13071 VSS.n939 VSS.n938 0.0176875
R13072 VSS.n948 VSS.n947 0.0176875
R13073 VSS.n602 VSS.n601 0.0176875
R13074 VSS.n2021 VSS.n2020 0.0176875
R13075 VSS.n507 VSS.n506 0.0169062
R13076 VSS.n503 VSS.n502 0.0169062
R13077 VSS.n357 VSS.n355 0.0168043
R13078 VSS.n83 VSS.n81 0.0168043
R13079 VSS.n196 VSS.n194 0.0168043
R13080 VSS.n1971 VSS.n1969 0.0168043
R13081 VSS.n1886 VSS.n1884 0.0168043
R13082 VSS.n1760 VSS.n1758 0.0168043
R13083 VSS.n914 VSS.n912 0.0168043
R13084 VSS.n805 VSS.n803 0.0168043
R13085 VSS.n1542 VSS.n1540 0.0168043
R13086 VSS.n1272 VSS.n1270 0.0168043
R13087 VSS.n17 VSS.n16 0.016125
R13088 VSS.n320 VSS.n319 0.016125
R13089 VSS.n50 VSS.n49 0.016125
R13090 VSS.n159 VSS.n150 0.016125
R13091 VSS.n1045 VSS.n1044 0.016125
R13092 VSS.n1051 VSS.n1050 0.016125
R13093 VSS.n1168 VSS.n1167 0.016125
R13094 VSS.n1812 VSS.n1811 0.016125
R13095 VSS.n1005 VSS.n1004 0.0155
R13096 VSS.n1940 VSS.n1937 0.0153437
R13097 VSS.n8 VSS.n7 0.0143978
R13098 VSS.n7 VSS.n6 0.0143978
R13099 VSS.n6 VSS.n5 0.0143978
R13100 VSS.n5 VSS.n4 0.0143978
R13101 VSS.n4 VSS.n3 0.0143978
R13102 VSS.n1 VSS.n0 0.0143978
R13103 VSS.n525 VSS.n524 0.0143978
R13104 VSS.n526 VSS.n525 0.0143978
R13105 VSS.n527 VSS.n526 0.0143978
R13106 VSS.n528 VSS.n527 0.0143978
R13107 VSS.n529 VSS.n528 0.0143978
R13108 VSS.n532 VSS.n531 0.0143978
R13109 VSS.n538 VSS.n532 0.0143978
R13110 VSS.n621 VSS.n618 0.0143978
R13111 VSS.n621 VSS.n620 0.0143978
R13112 VSS.n620 VSS.n619 0.0143978
R13113 VSS.n1691 VSS.n1690 0.0143978
R13114 VSS.n1690 VSS.n1689 0.0143978
R13115 VSS.n1689 VSS.n1688 0.0143978
R13116 VSS.n1688 VSS.n1687 0.0143978
R13117 VSS.n1687 VSS.n1686 0.0143978
R13118 VSS.n1686 VSS.n1685 0.0143978
R13119 VSS.n1683 VSS.n1682 0.0143978
R13120 VSS.n1682 VSS.n1681 0.0143978
R13121 VSS.n1681 VSS.n1680 0.0143978
R13122 VSS.n1699 VSS.n1698 0.0143978
R13123 VSS.n1700 VSS.n1699 0.0143978
R13124 VSS.n1701 VSS.n1700 0.0143978
R13125 VSS.n1704 VSS.n1703 0.0143978
R13126 VSS.n1705 VSS.n1704 0.0143978
R13127 VSS.n1706 VSS.n1705 0.0143978
R13128 VSS.n1707 VSS.n1706 0.0143978
R13129 VSS.n1709 VSS.n1707 0.0143978
R13130 VSS.n1709 VSS.n1708 0.0143978
R13131 VSS.n617 VSS.n542 0.0143978
R13132 VSS.n617 VSS.n616 0.0143978
R13133 VSS.n545 VSS.n544 0.0143978
R13134 VSS.n544 VSS.n543 0.0143978
R13135 VSS.n1818 VSS.n1817 0.0143978
R13136 VSS.n1832 VSS.n1831 0.0143978
R13137 VSS.n1825 VSS.n1824 0.0143978
R13138 VSS.n1838 VSS.n1837 0.0143978
R13139 VSS.n1943 VSS.n1942 0.0143978
R13140 VSS.n27 VSS.n26 0.0141719
R13141 VSS.n334 VSS.n333 0.0141719
R13142 VSS.n60 VSS.n59 0.0141719
R13143 VSS.n173 VSS.n172 0.0141719
R13144 VSS.n2015 VSS.n2014 0.0141719
R13145 VSS.n1930 VSS.n1929 0.0141719
R13146 VSS.n1805 VSS.n1804 0.0141719
R13147 VSS.n582 VSS.n581 0.0141719
R13148 VSS.n890 VSS.n889 0.0141719
R13149 VSS.n859 VSS.n858 0.0141719
R13150 VSS.n781 VSS.n780 0.0141719
R13151 VSS.n648 VSS.n647 0.0141719
R13152 VSS.n673 VSS.n672 0.0141719
R13153 VSS.n1649 VSS.n1648 0.0141719
R13154 VSS.n698 VSS.n697 0.0141719
R13155 VSS.n725 VSS.n724 0.0141719
R13156 VSS.n1603 VSS.n1602 0.0141719
R13157 VSS.n1609 VSS.n1608 0.0141719
R13158 VSS.n1472 VSS.n1471 0.0141719
R13159 VSS.n1480 VSS.n1479 0.0141719
R13160 VSS.n1128 VSS.n1127 0.0141719
R13161 VSS.n1136 VSS.n1135 0.0141719
R13162 VSS.n1333 VSS.n1332 0.0141719
R13163 VSS.n1339 VSS.n1338 0.0141719
R13164 VSS.n1210 VSS.n1209 0.0141719
R13165 VSS.n1163 VSS.n1162 0.0141719
R13166 VSS.n1025 VSS.n1024 0.0141719
R13167 VSS.n623 VSS.n622 0.0141452
R13168 VSS.n1817 VSS.n1816 0.0141452
R13169 VSS.n397 VSS.n390 0.014087
R13170 VSS.n107 VSS.n104 0.014087
R13171 VSS.n236 VSS.n229 0.014087
R13172 VSS.n1566 VSS.n1563 0.014087
R13173 VSS.n1597 VSS.n1595 0.014087
R13174 VSS.n1466 VSS.n1464 0.014087
R13175 VSS.n1122 VSS.n1120 0.014087
R13176 VSS.n1296 VSS.n1293 0.014087
R13177 VSS.n1327 VSS.n1325 0.014087
R13178 VSS.n1832 VSS.n1823 0.0136398
R13179 VSS.n455 VSS.n454 0.013
R13180 VSS.n1003 VSS.n1002 0.013
R13181 VSS.n517 VSS.n516 0.012435
R13182 VSS.n501 VSS.n500 0.0124292
R13183 VSS.n505 VSS.n504 0.0124292
R13184 VSS.n530 VSS.n529 0.0123763
R13185 VSS.n537 VSS.n536 0.0123763
R13186 VSS.n2007 VSS.n2006 0.0122188
R13187 VSS.n1922 VSS.n1921 0.0122188
R13188 VSS.n1797 VSS.n1796 0.0122188
R13189 VSS.n571 VSS.n570 0.0122188
R13190 VSS.n882 VSS.n881 0.0122188
R13191 VSS.n851 VSS.n850 0.0122188
R13192 VSS.n770 VSS.n769 0.0122188
R13193 VSS.n642 VSS.n641 0.0122188
R13194 VSS.n636 VSS.n635 0.0122188
R13195 VSS.n661 VSS.n660 0.0122188
R13196 VSS.n1643 VSS.n1642 0.0122188
R13197 VSS.n1637 VSS.n1636 0.0122188
R13198 VSS.n692 VSS.n691 0.0122188
R13199 VSS.n686 VSS.n685 0.0122188
R13200 VSS.n711 VSS.n710 0.0122188
R13201 VSS.n1504 VSS.n1499 0.0122188
R13202 VSS.n1494 VSS.n1489 0.0122188
R13203 VSS.n1427 VSS.n1418 0.0122188
R13204 VSS.n1084 VSS.n1083 0.0122188
R13205 VSS.n1234 VSS.n1229 0.0122188
R13206 VSS.n1224 VSS.n1219 0.0122188
R13207 VSS.n1201 VSS.n1200 0.0122188
R13208 VSS.n1195 VSS.n1194 0.0122188
R13209 VSS.n1145 VSS.n1144 0.0122188
R13210 VSS.n1036 VSS.n1035 0.0122188
R13211 VSS.n1041 VSS.n1040 0.0122188
R13212 VSS.n1042 VSS.n1041 0.0122188
R13213 VSS.n1062 VSS.n1061 0.0122188
R13214 VSS.n950 VSS.n949 0.0118907
R13215 VSS.n1405 VSS.n1404 0.0118907
R13216 VSS.n600 VSS.n599 0.0118907
R13217 VSS.n615 VSS.n545 0.011871
R13218 VSS.n1830 VSS.n1825 0.011871
R13219 VSS.n542 VSS.n541 0.0116183
R13220 VSS.n2027 VSS.n2026 0.0116183
R13221 VSS.n514 VSS.n513 0.0114375
R13222 VSS.n1165 VSS.n1149 0.0114375
R13223 VSS.n1702 VSS.n1701 0.0113656
R13224 VSS.n1685 VSS.n1684 0.0108602
R13225 VSS.n666 VSS.n665 0.010758
R13226 VSS.n716 VSS.n715 0.010758
R13227 VSS.n1432 VSS.n1431 0.010758
R13228 VSS.n1089 VSS.n1088 0.010758
R13229 VSS.n322 VSS.n321 0.0107521
R13230 VSS.n52 VSS.n51 0.0107521
R13231 VSS.n161 VSS.n160 0.0107521
R13232 VSS.n1009 VSS.n1008 0.0105
R13233 VSS.n1382 VSS.n1378 0.0104225
R13234 VSS.n3 VSS.n2 0.0103548
R13235 VSS.n37 VSS.n33 0.0102656
R13236 VSS.n452 VSS.n443 0.0102656
R13237 VSS.n140 VSS.n135 0.0102656
R13238 VSS.n291 VSS.n282 0.0102656
R13239 VSS.n2016 VSS.n2015 0.0102656
R13240 VSS.n2005 VSS.n2004 0.0102656
R13241 VSS.n1931 VSS.n1930 0.0102656
R13242 VSS.n1920 VSS.n1919 0.0102656
R13243 VSS.n1806 VSS.n1805 0.0102656
R13244 VSS.n1795 VSS.n1794 0.0102656
R13245 VSS.n583 VSS.n582 0.0102656
R13246 VSS.n569 VSS.n568 0.0102656
R13247 VSS.n891 VSS.n890 0.0102656
R13248 VSS.n880 VSS.n879 0.0102656
R13249 VSS.n860 VSS.n859 0.0102656
R13250 VSS.n849 VSS.n848 0.0102656
R13251 VSS.n782 VSS.n781 0.0102656
R13252 VSS.n768 VSS.n767 0.0102656
R13253 VSS.n2040 VSS.n2039 0.0101021
R13254 VSS.n536 VSS.n535 0.0101021
R13255 VSS.n1672 VSS.n1671 0.009875
R13256 VSS.n18 VSS.n17 0.00987154
R13257 VSS.n19 VSS.n18 0.00967578
R13258 VSS.n951 VSS.n740 0.00962927
R13259 VSS.n1403 VSS.n728 0.00962927
R13260 VSS.n1942 VSS.n1941 0.00959677
R13261 VSS.n465 VSS.n464 0.00957737
R13262 VSS.n466 VSS.n465 0.00957737
R13263 VSS.n944 VSS.n943 0.00957737
R13264 VSS.n943 VSS.n942 0.00957737
R13265 VSS.n1345 VSS.n1344 0.00957737
R13266 VSS.n1341 VSS.n1216 0.00957737
R13267 VSS.n1183 VSS.n1182 0.00957737
R13268 VSS.n1661 VSS.n1660 0.00957737
R13269 VSS.n1655 VSS.n1654 0.00957737
R13270 VSS.n1625 VSS.n1624 0.00957737
R13271 VSS.n1621 VSS.n1620 0.00957737
R13272 VSS.n1615 VSS.n1614 0.00957737
R13273 VSS.n1611 VSS.n1486 0.00957737
R13274 VSS.n1407 VSS.n1406 0.00957737
R13275 VSS.n1212 VSS.n1183 0.00957737
R13276 VSS.n1216 VSS.n1215 0.00957737
R13277 VSS.n1346 VSS.n1345 0.00957737
R13278 VSS.n1482 VSS.n1407 0.00957737
R13279 VSS.n1486 VSS.n1485 0.00957737
R13280 VSS.n1616 VSS.n1615 0.00957737
R13281 VSS.n1651 VSS.n1625 0.00957737
R13282 VSS.n1620 VSS.n1619 0.00957737
R13283 VSS.n1656 VSS.n1655 0.00957737
R13284 VSS.n1660 VSS.n1659 0.00957737
R13285 VSS.n607 VSS.n606 0.00957737
R13286 VSS.n1815 VSS.n1814 0.00957737
R13287 VSS.n1940 VSS.n1939 0.00957737
R13288 VSS.n606 VSS.n605 0.00957737
R13289 VSS.n1939 VSS.n1938 0.00957737
R13290 VSS.n1814 VSS.n1813 0.00957737
R13291 VSS.n740 VSS.n739 0.00952566
R13292 VSS.n728 VSS.n727 0.00952566
R13293 VSS.n468 VSS.n467 0.0091882
R13294 VSS.n467 VSS.n466 0.0091882
R13295 VSS.n938 VSS.n937 0.0091882
R13296 VSS.n941 VSS.n940 0.0091882
R13297 VSS.n947 VSS.n946 0.0091882
R13298 VSS.n946 VSS.n945 0.0091882
R13299 VSS.n942 VSS.n941 0.0091882
R13300 VSS.n937 VSS.n936 0.0091882
R13301 VSS.n1347 VSS.n1346 0.0091882
R13302 VSS.n1342 VSS.n1341 0.0091882
R13303 VSS.n1214 VSS.n1213 0.0091882
R13304 VSS.n1166 VSS.n1165 0.0091882
R13305 VSS.n1662 VSS.n1661 0.0091882
R13306 VSS.n1657 VSS.n1656 0.0091882
R13307 VSS.n1653 VSS.n1652 0.0091882
R13308 VSS.n1622 VSS.n1621 0.0091882
R13309 VSS.n1617 VSS.n1616 0.0091882
R13310 VSS.n1612 VSS.n1611 0.0091882
R13311 VSS.n1484 VSS.n1483 0.0091882
R13312 VSS.n1343 VSS.n1342 0.0091882
R13313 VSS.n1348 VSS.n1347 0.0091882
R13314 VSS.n1613 VSS.n1612 0.0091882
R13315 VSS.n1618 VSS.n1617 0.0091882
R13316 VSS.n1623 VSS.n1622 0.0091882
R13317 VSS.n1483 VSS.n1482 0.0091882
R13318 VSS.n1652 VSS.n1651 0.0091882
R13319 VSS.n1658 VSS.n1657 0.0091882
R13320 VSS.n1213 VSS.n1212 0.0091882
R13321 VSS.n1167 VSS.n1166 0.0091882
R13322 VSS.n1663 VSS.n1662 0.0091882
R13323 VSS.n605 VSS.n604 0.0091882
R13324 VSS.n2022 VSS.n2021 0.0091882
R13325 VSS.n604 VSS.n603 0.0091882
R13326 VSS.n2023 VSS.n2022 0.0091882
R13327 VSS.n321 VSS.n320 0.00879896
R13328 VSS.n51 VSS.n50 0.00879896
R13329 VSS.n160 VSS.n159 0.00879896
R13330 VSS.n408 VSS.n401 0.00865217
R13331 VSS.n439 VSS.n437 0.00865217
R13332 VSS.n114 VSS.n111 0.00865217
R13333 VSS.n131 VSS.n129 0.00865217
R13334 VSS.n247 VSS.n240 0.00865217
R13335 VSS.n278 VSS.n276 0.00865217
R13336 VSS.n1573 VSS.n1570 0.00865217
R13337 VSS.n1590 VSS.n1588 0.00865217
R13338 VSS.n1455 VSS.n1453 0.00865217
R13339 VSS.n1111 VSS.n1109 0.00865217
R13340 VSS.n1303 VSS.n1300 0.00865217
R13341 VSS.n1320 VSS.n1318 0.00865217
R13342 VSS.n1018 VSS.n1017 0.0083125
R13343 VSS.n1030 VSS.n1029 0.0083125
R13344 VSS.n614 VSS.n611 0.0083125
R13345 VSS.n1829 VSS.n1826 0.0083125
R13346 VSS.n1155 VSS.n1154 0.00765694
R13347 VSS.n1433 VSS.n1432 0.00685176
R13348 VSS.n717 VSS.n716 0.00685176
R13349 VSS.n1090 VSS.n1089 0.00685176
R13350 VSS.n667 VSS.n666 0.00685176
R13351 VSS.n1695 VSS.n1694 0.0068172
R13352 VSS.n515 VSS.n514 0.00675
R13353 VSS.n511 VSS.n510 0.00675
R13354 VSS.n1149 VSS.n624 0.00675
R13355 VSS.n506 VSS.n505 0.00671462
R13356 VSS.n502 VSS.n501 0.00671462
R13357 VSS.n2029 VSS.n2028 0.00656452
R13358 VSS.n951 VSS.n950 0.00647588
R13359 VSS.n1404 VSS.n1403 0.00647588
R13360 VSS.n601 VSS.n600 0.00647588
R13361 VSS.n1026 VSS.n1025 0.00635938
R13362 VSS.n348 VSS.n346 0.00593478
R13363 VSS.n73 VSS.n71 0.00593478
R13364 VSS.n186 VSS.n184 0.00593478
R13365 VSS.n1736 VSS.n1734 0.00593478
R13366 VSS.n1750 VSS.n1748 0.00593478
R13367 VSS.n1851 VSS.n1849 0.00593478
R13368 VSS.n1876 VSS.n1874 0.00593478
R13369 VSS.n1864 VSS.n1857 0.00593478
R13370 VSS.n1961 VSS.n1959 0.00593478
R13371 VSS.n905 VSS.n903 0.00593478
R13372 VSS.n796 VSS.n794 0.00593478
R13373 VSS.n1516 VSS.n1514 0.00593478
R13374 VSS.n1532 VSS.n1530 0.00593478
R13375 VSS.n1246 VSS.n1244 0.00593478
R13376 VSS.n1262 VSS.n1260 0.00593478
R13377 VSS.n516 VSS.n515 0.00592961
R13378 VSS.n540 VSS.n539 0.00580645
R13379 VSS.n999 VSS.n998 0.0055
R13380 VSS.n1941 VSS.n1838 0.00530108
R13381 VSS.n974 VSS.n973 0.00507113
R13382 VSS.n1396 VSS.n974 0.00507113
R13383 VSS.n1398 VSS.n1397 0.00507113
R13384 VSS.n1397 VSS.n1396 0.00507113
R13385 VSS.n962 VSS.n961 0.00507113
R13386 VSS.n956 VSS.n955 0.00507113
R13387 VSS.n1367 VSS.n1366 0.00507113
R13388 VSS.n1376 VSS.n1367 0.00507113
R13389 VSS.n1360 VSS.n1359 0.00507113
R13390 VSS.n38 VSS.n37 0.00492302
R13391 VSS.n141 VSS.n140 0.00492108
R13392 VSS.n292 VSS.n291 0.00492108
R13393 VSS.n453 VSS.n452 0.00492021
R13394 VSS.n1162 VSS.n1159 0.00490286
R13395 VSS.n2040 VSS.n2038 0.0047957
R13396 VSS.n535 VSS.n534 0.0047957
R13397 VSS.n963 VSS.n962 0.00478282
R13398 VSS.n957 VSS.n956 0.00478282
R13399 VSS.n1361 VSS.n1360 0.00478282
R13400 VSS.n2 VSS.n1 0.00454301
R13401 VSS.n641 VSS.n640 0.00440625
R13402 VSS.n662 VSS.n661 0.00440625
R13403 VSS.n1642 VSS.n1641 0.00440625
R13404 VSS.n691 VSS.n690 0.00440625
R13405 VSS.n712 VSS.n711 0.00440625
R13406 VSS.n1499 VSS.n1498 0.00440625
R13407 VSS.n1428 VSS.n1427 0.00440625
R13408 VSS.n1085 VSS.n1084 0.00440625
R13409 VSS.n1229 VSS.n1228 0.00440625
R13410 VSS.n1200 VSS.n1199 0.00440625
R13411 VSS.n1016 VSS.n1015 0.00440625
R13412 VSS.n2038 VSS.n2037 0.00429032
R13413 VSS.n534 VSS.n533 0.00429032
R13414 VSS.n1684 VSS.n1683 0.00403763
R13415 VSS.n1703 VSS.n1702 0.00353226
R13416 VSS.n541 VSS.n540 0.00327957
R13417 VSS.n419 VSS.n412 0.00321739
R13418 VSS.n428 VSS.n426 0.00321739
R13419 VSS.n120 VSS.n118 0.00321739
R13420 VSS.n124 VSS.n122 0.00321739
R13421 VSS.n258 VSS.n251 0.00321739
R13422 VSS.n267 VSS.n265 0.00321739
R13423 VSS.n564 VSS.n562 0.00321739
R13424 VSS.n756 VSS.n754 0.00321739
R13425 VSS.n1579 VSS.n1577 0.00321739
R13426 VSS.n1583 VSS.n1581 0.00321739
R13427 VSS.n1444 VSS.n1442 0.00321739
R13428 VSS.n1100 VSS.n1098 0.00321739
R13429 VSS.n1309 VSS.n1307 0.00321739
R13430 VSS.n1313 VSS.n1311 0.00321739
R13431 VSS.n616 VSS.n615 0.00302688
R13432 VSS.n1831 VSS.n1830 0.00302688
R13433 VSS.n637 VSS.n636 0.00295228
R13434 VSS.n1638 VSS.n1637 0.00295228
R13435 VSS.n687 VSS.n686 0.00295228
R13436 VSS.n1495 VSS.n1494 0.00295228
R13437 VSS.n1225 VSS.n1224 0.00295228
R13438 VSS.n1196 VSS.n1195 0.00295228
R13439 VSS.n1822 VSS.n1820 0.00284375
R13440 VSS.n2025 VSS.n1945 0.00284375
R13441 VSS.n2041 VSS.n2036 0.00278115
R13442 VSS.n2042 VSS.n2041 0.00278115
R13443 VSS.n499 VSS.n498 0.00269167
R13444 VSS.n531 VSS.n530 0.00252151
R13445 VSS.n538 VSS.n537 0.00252151
R13446 VSS.n2029 VSS.n2027 0.00252151
R13447 VSS.n2018 VSS.n2017 0.00245312
R13448 VSS.n2008 VSS.n2007 0.00245312
R13449 VSS.n1933 VSS.n1932 0.00245312
R13450 VSS.n1923 VSS.n1922 0.00245312
R13451 VSS.n1808 VSS.n1807 0.00245312
R13452 VSS.n1798 VSS.n1797 0.00245312
R13453 VSS.n588 VSS.n587 0.00245312
R13454 VSS.n572 VSS.n571 0.00245312
R13455 VSS.n893 VSS.n892 0.00245312
R13456 VSS.n883 VSS.n882 0.00245312
R13457 VSS.n865 VSS.n864 0.00245312
R13458 VSS.n852 VSS.n851 0.00245312
R13459 VSS.n784 VSS.n783 0.00245312
R13460 VSS.n771 VSS.n770 0.00245312
R13461 VSS.n1713 VSS.n1712 0.00226882
R13462 VSS.n1695 VSS.n1693 0.00226882
R13463 VSS.n1937 VSS.n1936 0.0020625
R13464 VSS.n1396 VSS.n963 0.00178792
R13465 VSS.n1396 VSS.n957 0.00178792
R13466 VSS.n1376 VSS.n1361 0.00178792
R13467 VSS.n1834 VSS.n1833 0.00166815
R13468 VSS.n1714 VSS.n1711 0.00166815
R13469 VSS.n1715 VSS.n1714 0.00166815
R13470 VSS.n1833 VSS.n1724 0.00166815
R13471 VSS.n301 VSS.n300 0.00149427
R13472 VSS.n2033 VSS.n2032 0.00145036
R13473 VSS.n2034 VSS.n2033 0.00145036
R13474 VSS.n2045 VSS.n2044 0.00143078
R13475 VSS.n2046 VSS.n2045 0.00143078
R13476 VSS.n498 VSS.n497 0.00130794
R13477 VSS.n1175 VSS.n1174 0.00128125
R13478 VSS.n1815 VSS.n1812 0.00128125
R13479 VSS.n1823 VSS.n1818 0.00125806
R13480 VSS.n2026 VSS.n1943 0.00125806
R13481 VSS.n2043 VSS.n2042 0.00119582
R13482 VSS.n2044 VSS.n2043 0.00119582
R13483 VSS.n2036 VSS.n2035 0.00117624
R13484 VSS.n2035 VSS.n2034 0.00117624
R13485 VSS.n1390 VSS.n1389 0.00117024
R13486 VSS.n1721 VSS.n1720 0.0011689
R13487 VSS.n1697 VSS.n1696 0.0011689
R13488 VSS.n1722 VSS.n1721 0.0011689
R13489 VSS.n1696 VSS.n1692 0.0011689
R13490 VSS.n2031 VSS.n2030 0.00116156
R13491 VSS.n1718 VSS.n1717 0.00116156
R13492 VSS.n2030 VSS.n1836 0.00116156
R13493 VSS.n1719 VSS.n1718 0.00116156
R13494 VSS.n982 VSS.n979 0.00113518
R13495 VSS.n1375 VSS.n1374 0.00113518
R13496 VSS.n1395 VSS.n1394 0.00113518
R13497 VSS.n1390 VSS.n1387 0.00113518
R13498 VSS.n1835 VSS.n1834 0.00107344
R13499 VSS.n1716 VSS.n1715 0.00107344
R13500 VSS.n1836 VSS.n1835 0.00107344
R13501 VSS.n1717 VSS.n1716 0.00107344
R13502 VSS.n1723 VSS.n1722 0.00106609
R13503 VSS.n1711 VSS.n1710 0.00106609
R13504 VSS.n1710 VSS.n1697 0.00106609
R13505 VSS.n1724 VSS.n1723 0.00106609
R13506 VSS.n1395 VSS.n1392 0.00105224
R13507 VSS.n1375 VSS.n1369 0.00105224
R13508 VSS.n967 VSS.n966 0.00100786
R13509 VSS.n1365 VSS.n1364 0.00100786
R13510 VSS.n982 VSS.n981 0.00100398
R13511 VSS.n492 VSS.n491 0.00100166
R13512 VSS.n479 VSS.n478 0.00100166
R13513 VSS.n492 VSS.n489 0.00100102
R13514 VSS.n479 VSS.n476 0.00100102
R13515 VSS.n480 VSS.n474 0.00100018
R13516 VSS.n1396 VSS.n967 0.00100009
R13517 VSS.n1376 VSS.n1365 0.00100009
R13518 VSS.n997 VSS.n996 0.00100007
R13519 VSS.n470 VSS.n469 0.00100006
R13520 VSS.n1351 VSS.n1350 0.00100002
R13521 VSS.n472 VSS.n470 0.00100001
R13522 VSS.n1396 VSS.n1390 0.001
R13523 VSS.n493 VSS.n492 0.001
R13524 VSS.n474 VSS.n473 0.001
R13525 VSS.n480 VSS.n479 0.001
R13526 VSS.n983 VSS.n982 0.001
R13527 VSS.n1376 VSS.n1375 0.001
R13528 VSS.n1396 VSS.n1395 0.001
R13529 VSS.n1691 VSS.n623 0.000752688
R13530 VSS.n1816 VSS.n1725 0.000752688
R13531 VSS.n1389 VSS.n1388 0.000670243
R13532 VSS.n979 VSS.n978 0.000635176
R13533 VSS.n1374 VSS.n1373 0.000635176
R13534 VSS.n1394 VSS.n1393 0.000635176
R13535 VSS.n1387 VSS.n1386 0.000635176
R13536 VSS.n984 VSS.n983 0.000635176
R13537 VSS.n985 VSS.n984 0.000635176
R13538 VSS.n1382 VSS.n1381 0.000631513
R13539 VSS.n1381 VSS.n1380 0.000631513
R13540 VSS.n1392 VSS.n1391 0.000552238
R13541 VSS.n1369 VSS.n1368 0.000552238
R13542 VSS.n969 VSS.n968 0.000512877
R13543 VSS.n1396 VSS.n969 0.000512877
R13544 VSS.n988 VSS.n987 0.00051244
R13545 VSS.n987 VSS.n986 0.00051244
R13546 VSS.n1378 VSS.n1377 0.000511972
R13547 VSS.n1377 VSS.n1376 0.000511972
R13548 VSS.n990 VSS.n989 0.000509014
R13549 VSS.n991 VSS.n990 0.000509014
R13550 VSS.n966 VSS.n965 0.000507954
R13551 VSS.n1364 VSS.n1363 0.000507954
R13552 VSS.n495 VSS.n494 0.000505303
R13553 VSS.n494 VSS.n493 0.000505303
R13554 VSS.n482 VSS.n481 0.000505303
R13555 VSS.n481 VSS.n480 0.000505303
R13556 VSS.n981 VSS.n980 0.000503977
R13557 VSS.n487 VSS.n486 0.000503145
R13558 VSS.n486 VSS.n485 0.000503145
R13559 VSS.n485 VSS.n484 0.000503145
R13560 VSS.n484 VSS.n483 0.000503145
R13561 VSS.n491 VSS.n490 0.000501661
R13562 VSS.n478 VSS.n477 0.000501661
R13563 VSS.n1372 VSS.n1371 0.000501229
R13564 VSS.n1371 VSS.n1370 0.000501229
R13565 VSS.n1385 VSS.n1384 0.000501048
R13566 VSS.n1384 VSS.n1383 0.000501048
R13567 VSS.n489 VSS.n488 0.000501025
R13568 VSS.n476 VSS.n475 0.000501025
R13569 VSS.n992 VSS.n991 0.000500725
R13570 VSS.n993 VSS.n992 0.000500725
R13571 VSS.n996 VSS.n995 0.000500479
R13572 VSS.n995 VSS.n994 0.000500479
R13573 VSS.n497 VSS.n301 0.000500181
R13574 VSS.n473 VSS.n472 0.000500181
R13575 VSS.n1350 VSS.n1349 0.000500106
R13576 a_2151_4783.n51 a_2151_4783.t8 60.2505
R13577 a_2151_4783.n72 a_2151_4783.t9 60.2505
R13578 a_2151_4783.n94 a_2151_4783.t2 60.2505
R13579 a_2151_4783.n39 a_2151_4783.t0 60.2505
R13580 a_2151_4783.n5 a_2151_4783.n60 9.3005
R13581 a_2151_4783.n7 a_2151_4783.n64 9.3005
R13582 a_2151_4783.n8 a_2151_4783.n82 9.3005
R13583 a_2151_4783.n10 a_2151_4783.n86 9.3005
R13584 a_2151_4783.n11 a_2151_4783.n104 9.3005
R13585 a_2151_4783.n12 a_2151_4783.n48 9.3005
R13586 a_2151_4783.n12 a_2151_4783.n47 9.3005
R13587 a_2151_4783.n12 a_2151_4783.n46 9.3005
R13588 a_2151_4783.n46 a_2151_4783.n45 9.3005
R13589 a_2151_4783.n11 a_2151_4783.n103 9.3005
R13590 a_2151_4783.n11 a_2151_4783.n102 9.3005
R13591 a_2151_4783.n102 a_2151_4783.n101 9.3005
R13592 a_2151_4783.n10 a_2151_4783.n87 9.3005
R13593 a_2151_4783.n10 a_2151_4783.n93 9.3005
R13594 a_2151_4783.n93 a_2151_4783.n92 9.3005
R13595 a_2151_4783.n8 a_2151_4783.n81 9.3005
R13596 a_2151_4783.n8 a_2151_4783.n80 9.3005
R13597 a_2151_4783.n80 a_2151_4783.n79 9.3005
R13598 a_2151_4783.n7 a_2151_4783.n65 9.3005
R13599 a_2151_4783.n7 a_2151_4783.n71 9.3005
R13600 a_2151_4783.n71 a_2151_4783.n70 9.3005
R13601 a_2151_4783.n5 a_2151_4783.n58 9.3005
R13602 a_2151_4783.n58 a_2151_4783.n57 9.3005
R13603 a_2151_4783.n5 a_2151_4783.n59 9.3005
R13604 a_2151_4783.n0 a_2151_4783.n109 9.3005
R13605 a_2151_4783.n95 a_2151_4783.n94 8.76429
R13606 a_2151_4783.n73 a_2151_4783.n72 8.76429
R13607 a_2151_4783.n44 a_2151_4783.n43 7.45411
R13608 a_2151_4783.n100 a_2151_4783.n99 7.45411
R13609 a_2151_4783.n91 a_2151_4783.n90 7.45411
R13610 a_2151_4783.n78 a_2151_4783.n77 7.45411
R13611 a_2151_4783.n69 a_2151_4783.n68 7.45411
R13612 a_2151_4783.n56 a_2151_4783.n55 7.45411
R13613 a_2151_4783.n40 a_2151_4783.n39 6.80334
R13614 a_2151_4783.n52 a_2151_4783.n51 6.80105
R13615 a_2151_4783.n111 a_2151_4783.n110 6.31679
R13616 a_2151_4783.n42 a_2151_4783.n41 5.64756
R13617 a_2151_4783.n98 a_2151_4783.n97 5.64756
R13618 a_2151_4783.n89 a_2151_4783.n88 5.64756
R13619 a_2151_4783.n76 a_2151_4783.n75 5.64756
R13620 a_2151_4783.n67 a_2151_4783.n66 5.64756
R13621 a_2151_4783.n54 a_2151_4783.n53 5.64756
R13622 a_2151_4783.n112 a_2151_4783.t1 5.5395
R13623 a_2151_4783.t3 a_2151_4783.n112 5.5395
R13624 a_2151_4783.n0 a_2151_4783.n108 4.95534
R13625 a_2151_4783.n50 a_2151_4783.n49 4.73575
R13626 a_2151_4783.n106 a_2151_4783.n105 4.73575
R13627 a_2151_4783.n9 a_2151_4783.n85 4.73575
R13628 a_2151_4783.n84 a_2151_4783.n83 4.73575
R13629 a_2151_4783.n6 a_2151_4783.n63 4.73575
R13630 a_2151_4783.n62 a_2151_4783.n61 4.73575
R13631 a_2151_4783.n1 a_2151_4783.n13 4.6673
R13632 a_2151_4783.n96 a_2151_4783.n95 4.6505
R13633 a_2151_4783.n74 a_2151_4783.n73 4.6505
R13634 a_2151_4783.n4 a_2151_4783.n31 4.5005
R13635 a_2151_4783.n4 a_2151_4783.n28 4.5005
R13636 a_2151_4783.n2 a_2151_4783.n20 4.5005
R13637 a_2151_4783.n2 a_2151_4783.n23 4.5005
R13638 a_2151_4783.n0 a_2151_4783.n38 4.5005
R13639 a_2151_4783.n1 a_2151_4783.n36 4.5005
R13640 a_2151_4783.n1 a_2151_4783.n15 4.5005
R13641 a_2151_4783.n28 a_2151_4783.n27 4.14168
R13642 a_2151_4783.n23 a_2151_4783.n22 4.14168
R13643 a_2151_4783.n15 a_2151_4783.n14 3.76521
R13644 a_2151_4783.n5 a_2151_4783.n52 3.42768
R13645 a_2151_4783.n12 a_2151_4783.n40 3.42683
R13646 a_2151_4783.n38 a_2151_4783.n37 3.38874
R13647 a_2151_4783.n32 a_2151_4783.t4 3.3065
R13648 a_2151_4783.n32 a_2151_4783.t7 3.3065
R13649 a_2151_4783.n16 a_2151_4783.t6 3.3065
R13650 a_2151_4783.n16 a_2151_4783.t5 3.3065
R13651 a_2151_4783.n36 a_2151_4783.n35 3.01226
R13652 a_2151_4783.n30 a_2151_4783.n29 2.25932
R13653 a_2151_4783.n19 a_2151_4783.n18 2.25932
R13654 a_2151_4783.n111 a_2151_4783.n1 1.50789
R13655 a_2151_4783.n17 a_2151_4783.n16 1.46878
R13656 a_2151_4783.n45 a_2151_4783.n44 0.994314
R13657 a_2151_4783.n101 a_2151_4783.n100 0.994314
R13658 a_2151_4783.n92 a_2151_4783.n91 0.994314
R13659 a_2151_4783.n79 a_2151_4783.n78 0.994314
R13660 a_2151_4783.n70 a_2151_4783.n69 0.994314
R13661 a_2151_4783.n57 a_2151_4783.n56 0.994314
R13662 a_2151_4783.n34 a_2151_4783.n25 0.920917
R13663 a_2151_4783.n46 a_2151_4783.n42 0.753441
R13664 a_2151_4783.n102 a_2151_4783.n98 0.753441
R13665 a_2151_4783.n93 a_2151_4783.n89 0.753441
R13666 a_2151_4783.n80 a_2151_4783.n76 0.753441
R13667 a_2151_4783.n71 a_2151_4783.n67 0.753441
R13668 a_2151_4783.n58 a_2151_4783.n54 0.753441
R13669 a_2151_4783.n13 a_2151_4783.n2 0.70141
R13670 a_2151_4783.n13 a_2151_4783.n34 0.700686
R13671 a_2151_4783.n2 a_2151_4783.n24 0.604067
R13672 a_2151_4783.n25 a_2151_4783.n33 0.594011
R13673 a_2151_4783.n4 a_2151_4783.n32 2.11687
R13674 a_2151_4783.n3 a_2151_4783.n17 0.555028
R13675 a_2151_4783.n9 a_2151_4783.n84 0.458354
R13676 a_2151_4783.n6 a_2151_4783.n62 0.458354
R13677 a_2151_4783.n1 a_2151_4783.n0 0.452411
R13678 a_2151_4783.n112 a_2151_4783.n111 0.400755
R13679 a_2151_4783.n28 a_2151_4783.n26 0.376971
R13680 a_2151_4783.n31 a_2151_4783.n30 0.376971
R13681 a_2151_4783.n23 a_2151_4783.n21 0.376971
R13682 a_2151_4783.n20 a_2151_4783.n19 0.376971
R13683 a_2151_4783.n2 a_2151_4783.n3 0.29091
R13684 a_2151_4783.n107 a_2151_4783.n50 0.229427
R13685 a_2151_4783.n107 a_2151_4783.n106 0.229427
R13686 a_2151_4783.n0 a_2151_4783.n107 0.215848
R13687 a_2151_4783.n25 a_2151_4783.n4 0.206871
R13688 a_2151_4783.n50 a_2151_4783.n12 0.205546
R13689 a_2151_4783.n106 a_2151_4783.n11 0.205546
R13690 a_2151_4783.n10 a_2151_4783.n9 0.205546
R13691 a_2151_4783.n84 a_2151_4783.n8 0.205546
R13692 a_2151_4783.n7 a_2151_4783.n6 0.205546
R13693 a_2151_4783.n62 a_2151_4783.n5 0.205546
R13694 a_2151_4783.n11 a_2151_4783.n96 0.190717
R13695 a_2151_4783.n96 a_2151_4783.n10 0.190717
R13696 a_2151_4783.n8 a_2151_4783.n74 0.190717
R13697 a_2151_4783.n74 a_2151_4783.n7 0.190717
R13698 a_2551_4880.n67 a_2551_4880.t4 60.2505
R13699 a_2551_4880.n46 a_2551_4880.t7 60.2505
R13700 a_2551_4880.n25 a_2551_4880.t6 60.2505
R13701 a_2551_4880.n80 a_2551_4880.t2 60.2505
R13702 a_2551_4880.n4 a_2551_4880.n88 9.3005
R13703 a_2551_4880.n4 a_2551_4880.n89 9.3005
R13704 a_2551_4880.n4 a_2551_4880.n87 9.3005
R13705 a_2551_4880.n87 a_2551_4880.n86 9.3005
R13706 a_2551_4880.n8 a_2551_4880.n56 9.3005
R13707 a_2551_4880.n10 a_2551_4880.n38 9.3005
R13708 a_2551_4880.n11 a_2551_4880.n34 9.3005
R13709 a_2551_4880.n11 a_2551_4880.n33 9.3005
R13710 a_2551_4880.n11 a_2551_4880.n32 9.3005
R13711 a_2551_4880.n32 a_2551_4880.n31 9.3005
R13712 a_2551_4880.n10 a_2551_4880.n39 9.3005
R13713 a_2551_4880.n10 a_2551_4880.n45 9.3005
R13714 a_2551_4880.n45 a_2551_4880.n44 9.3005
R13715 a_2551_4880.n8 a_2551_4880.n55 9.3005
R13716 a_2551_4880.n8 a_2551_4880.n54 9.3005
R13717 a_2551_4880.n54 a_2551_4880.n53 9.3005
R13718 a_2551_4880.n7 a_2551_4880.n59 9.3005
R13719 a_2551_4880.n7 a_2551_4880.n66 9.3005
R13720 a_2551_4880.n66 a_2551_4880.n65 9.3005
R13721 a_2551_4880.n7 a_2551_4880.n60 9.3005
R13722 a_2551_4880.n5 a_2551_4880.n75 9.3005
R13723 a_2551_4880.n75 a_2551_4880.n74 9.3005
R13724 a_2551_4880.n5 a_2551_4880.n77 9.3005
R13725 a_2551_4880.n5 a_2551_4880.n76 9.3005
R13726 a_2551_4880.n2 a_2551_4880.n94 9.3005
R13727 a_2551_4880.n13 a_2551_4880.n97 9.3005
R13728 a_2551_4880.n12 a_2551_4880.n101 9.3005
R13729 a_2551_4880.n3 a_2551_4880.n105 9.3005
R13730 a_2551_4880.n0 a_2551_4880.n109 9.3005
R13731 a_2551_4880.n0 a_2551_4880.n111 9.3005
R13732 a_2551_4880.n0 a_2551_4880.n108 9.3005
R13733 a_2551_4880.n3 a_2551_4880.n107 9.3005
R13734 a_2551_4880.n3 a_2551_4880.n104 9.3005
R13735 a_2551_4880.n12 a_2551_4880.n103 9.3005
R13736 a_2551_4880.n12 a_2551_4880.n100 9.3005
R13737 a_2551_4880.n13 a_2551_4880.n99 9.3005
R13738 a_2551_4880.n13 a_2551_4880.n96 9.3005
R13739 a_2551_4880.n2 a_2551_4880.n95 9.3005
R13740 a_2551_4880.n2 a_2551_4880.n93 9.3005
R13741 a_2551_4880.n47 a_2551_4880.n46 8.76429
R13742 a_2551_4880.n68 a_2551_4880.n67 8.76429
R13743 a_2551_4880.n30 a_2551_4880.n29 8.21641
R13744 a_2551_4880.n43 a_2551_4880.n42 8.21641
R13745 a_2551_4880.n52 a_2551_4880.n51 8.21641
R13746 a_2551_4880.n85 a_2551_4880.n84 8.21641
R13747 a_2551_4880.n64 a_2551_4880.n63 8.21641
R13748 a_2551_4880.n73 a_2551_4880.n72 8.21641
R13749 a_2551_4880.n19 a_2551_4880.n17 8.0439
R13750 a_2551_4880.n21 a_2551_4880.n20 8.02969
R13751 a_2551_4880.n26 a_2551_4880.n25 6.92242
R13752 a_2551_4880.n81 a_2551_4880.n80 6.92012
R13753 a_2551_4880.n114 a_2551_4880.n1 6.38347
R13754 a_2551_4880.n118 a_2551_4880.n117 6.31608
R13755 a_2551_4880.n28 a_2551_4880.n27 5.64756
R13756 a_2551_4880.n41 a_2551_4880.n40 5.64756
R13757 a_2551_4880.n50 a_2551_4880.n49 5.64756
R13758 a_2551_4880.n83 a_2551_4880.n82 5.64756
R13759 a_2551_4880.n62 a_2551_4880.n61 5.64756
R13760 a_2551_4880.n71 a_2551_4880.n70 5.64756
R13761 a_2551_4880.n119 a_2551_4880.t0 5.5395
R13762 a_2551_4880.t1 a_2551_4880.n119 5.5395
R13763 a_2551_4880.n2 a_2551_4880.n92 5.27461
R13764 a_2551_4880.n36 a_2551_4880.n35 4.76425
R13765 a_2551_4880.n9 a_2551_4880.n37 4.76425
R13766 a_2551_4880.n58 a_2551_4880.n57 4.76425
R13767 a_2551_4880.n90 a_2551_4880.n79 4.76425
R13768 a_2551_4880.n6 a_2551_4880.n24 4.76425
R13769 a_2551_4880.n78 a_2551_4880.n23 4.76425
R13770 a_2551_4880.n48 a_2551_4880.n47 4.6505
R13771 a_2551_4880.n69 a_2551_4880.n68 4.6505
R13772 a_2551_4880.n1 a_2551_4880.n19 4.5005
R13773 a_2551_4880.n1 a_2551_4880.n113 4.5005
R13774 a_2551_4880.n14 a_2551_4880.n116 4.5005
R13775 a_2551_4880.n113 a_2551_4880.n112 3.76521
R13776 a_2551_4880.n116 a_2551_4880.n115 3.76521
R13777 a_2551_4880.n4 a_2551_4880.n81 3.47756
R13778 a_2551_4880.n11 a_2551_4880.n26 3.4767
R13779 a_2551_4880.n19 a_2551_4880.n18 3.38874
R13780 a_2551_4880.n21 a_2551_4880.t5 3.3065
R13781 a_2551_4880.n21 a_2551_4880.t3 3.3065
R13782 a_2551_4880.n16 a_2551_4880.n15 3.01226
R13783 a_2551_4880.n22 a_2551_4880.n21 1.52644
R13784 a_2551_4880.n118 a_2551_4880.n14 1.50792
R13785 a_2551_4880.n14 a_2551_4880.n114 1.13333
R13786 a_2551_4880.n31 a_2551_4880.n30 1.09595
R13787 a_2551_4880.n44 a_2551_4880.n43 1.09595
R13788 a_2551_4880.n53 a_2551_4880.n52 1.09595
R13789 a_2551_4880.n86 a_2551_4880.n85 1.09595
R13790 a_2551_4880.n65 a_2551_4880.n64 1.09595
R13791 a_2551_4880.n74 a_2551_4880.n73 1.09595
R13792 a_2551_4880.n1 a_2551_4880.n22 0.938895
R13793 a_2551_4880.n32 a_2551_4880.n28 0.753441
R13794 a_2551_4880.n45 a_2551_4880.n41 0.753441
R13795 a_2551_4880.n54 a_2551_4880.n50 0.753441
R13796 a_2551_4880.n87 a_2551_4880.n83 0.753441
R13797 a_2551_4880.n66 a_2551_4880.n62 0.753441
R13798 a_2551_4880.n75 a_2551_4880.n71 0.753441
R13799 a_2551_4880.n9 a_2551_4880.n36 0.458354
R13800 a_2551_4880.n6 a_2551_4880.n58 0.458354
R13801 a_2551_4880.n99 a_2551_4880.n98 0.430121
R13802 a_2551_4880.n119 a_2551_4880.n118 0.400734
R13803 a_2551_4880.n103 a_2551_4880.n102 0.398603
R13804 a_2551_4880.n107 a_2551_4880.n106 0.366615
R13805 a_2551_4880.n111 a_2551_4880.n110 0.334147
R13806 a_2551_4880.n14 a_2551_4880.n16 4.77996
R13807 a_2551_4880.n1 a_2551_4880.n0 0.39232
R13808 a_2551_4880.n13 a_2551_4880.n2 0.354994
R13809 a_2551_4880.n91 a_2551_4880.n78 0.229427
R13810 a_2551_4880.n91 a_2551_4880.n90 0.229427
R13811 a_2551_4880.n36 a_2551_4880.n11 0.205546
R13812 a_2551_4880.n10 a_2551_4880.n9 0.205546
R13813 a_2551_4880.n58 a_2551_4880.n8 0.205546
R13814 a_2551_4880.n7 a_2551_4880.n6 0.205546
R13815 a_2551_4880.n78 a_2551_4880.n5 0.205546
R13816 a_2551_4880.n90 a_2551_4880.n4 0.205546
R13817 a_2551_4880.n2 a_2551_4880.n91 0.191391
R13818 a_2551_4880.n3 a_2551_4880.n12 0.190717
R13819 a_2551_4880.n48 a_2551_4880.n10 0.190717
R13820 a_2551_4880.n8 a_2551_4880.n48 0.190717
R13821 a_2551_4880.n69 a_2551_4880.n7 0.190717
R13822 a_2551_4880.n5 a_2551_4880.n69 0.190717
R13823 a_2551_4880.n12 a_2551_4880.n13 0.190717
R13824 a_2551_4880.n0 a_2551_4880.n3 0.190717
R13825 a_8881_1782.n109 a_8881_1782.t2 120.501
R13826 a_8881_1782.n21 a_8881_1782.t0 69.2068
R13827 a_8881_1782.n59 a_8881_1782.t3 60.2505
R13828 a_8881_1782.n46 a_8881_1782.n45 31.4488
R13829 a_8881_1782.n24 a_8881_1782.n23 27.5177
R13830 a_8881_1782.n7 a_8881_1782.n3 26.107
R13831 a_8881_1782.n35 a_8881_1782.n34 23.5867
R13832 a_8881_1782.n13 a_8881_1782.n12 19.6557
R13833 a_8881_1782.n3 a_8881_1782.n2 15.7246
R13834 a_8881_1782.n14 a_8881_1782.n13 13.7591
R13835 a_8881_1782.n36 a_8881_1782.n35 9.82809
R13836 a_8881_1782.n86 a_8881_1782.n85 9.3005
R13837 a_8881_1782.n69 a_8881_1782.n68 9.3005
R13838 a_8881_1782.n123 a_8881_1782.n122 9.3005
R13839 a_8881_1782.n104 a_8881_1782.n103 9.3005
R13840 a_8881_1782.n50 a_8881_1782.n52 9.3005
R13841 a_8881_1782.n15 a_8881_1782.n14 9.3005
R13842 a_8881_1782.n37 a_8881_1782.n36 9.3005
R13843 a_8881_1782.n28 a_8881_1782.n38 9.3005
R13844 a_8881_1782.n26 a_8881_1782.n25 9.3005
R13845 a_8881_1782.n39 a_8881_1782.n41 9.3005
R13846 a_8881_1782.n48 a_8881_1782.n47 9.3005
R13847 a_8881_1782.n1 a_8881_1782.n139 9.3005
R13848 a_8881_1782.n131 a_8881_1782.n146 9.3005
R13849 a_8881_1782.n1 a_8881_1782.n138 9.3005
R13850 a_8881_1782.n0 a_8881_1782.n134 9.3005
R13851 a_8881_1782.n131 a_8881_1782.n145 9.3005
R13852 a_8881_1782.n60 a_8881_1782.n59 8.76429
R13853 a_8881_1782.n110 a_8881_1782.n109 8.76429
R13854 a_8881_1782.n67 a_8881_1782.n66 8.21641
R13855 a_8881_1782.n84 a_8881_1782.n83 8.21641
R13856 a_8881_1782.n102 a_8881_1782.n101 7.45411
R13857 a_8881_1782.n121 a_8881_1782.n120 7.45411
R13858 a_8881_1782.n25 a_8881_1782.n24 5.89705
R13859 a_8881_1782.n150 a_8881_1782.n149 5.38095
R13860 a_8881_1782.n8 a_8881_1782.n7 5.20544
R13861 a_8881_1782.n56 a_8881_1782.n54 4.87224
R13862 a_8881_1782.n89 a_8881_1782.n74 4.86623
R13863 a_8881_1782.n92 a_8881_1782.n90 4.84151
R13864 a_8881_1782.n126 a_8881_1782.n108 4.83995
R13865 a_8881_1782.n111 a_8881_1782.n110 4.6505
R13866 a_8881_1782.n0 a_8881_1782.n133 4.5298
R13867 a_8881_1782.n30 a_8881_1782.n31 4.51815
R13868 a_8881_1782.n33 a_8881_1782.n32 4.51815
R13869 a_8881_1782.n55 a_8881_1782.n70 4.5005
R13870 a_8881_1782.n57 a_8881_1782.n63 4.5005
R13871 a_8881_1782.n77 a_8881_1782.n81 4.5005
R13872 a_8881_1782.n82 a_8881_1782.n88 4.5005
R13873 a_8881_1782.n91 a_8881_1782.n105 4.5005
R13874 a_8881_1782.n93 a_8881_1782.n98 4.5005
R13875 a_8881_1782.n114 a_8881_1782.n118 4.5005
R13876 a_8881_1782.n119 a_8881_1782.n125 4.5005
R13877 a_8881_1782.n8 a_8881_1782.n16 4.5005
R13878 a_8881_1782.n42 a_8881_1782.n49 4.5005
R13879 a_8881_1782.n29 a_8881_1782.n27 4.5005
R13880 a_8881_1782.n94 a_8881_1782.n95 4.5005
R13881 a_8881_1782.n113 a_8881_1782.n112 4.5005
R13882 a_8881_1782.n1 a_8881_1782.n137 4.5005
R13883 a_8881_1782.n130 a_8881_1782.n144 4.5005
R13884 a_8881_1782.n58 a_8881_1782.n60 4.14168
R13885 a_8881_1782.n76 a_8881_1782.n75 4.14168
R13886 a_8881_1782.n49 a_8881_1782.n43 4.14168
R13887 a_8881_1782.n88 a_8881_1782.n86 3.76521
R13888 a_8881_1782.n125 a_8881_1782.n123 3.76521
R13889 a_8881_1782.n16 a_8881_1782.n9 3.76521
R13890 a_8881_1782.n11 a_8881_1782.n10 3.76521
R13891 a_8881_1782.n70 a_8881_1782.n69 3.38874
R13892 a_8881_1782.n105 a_8881_1782.n104 3.38874
R13893 a_8881_1782.n6 a_8881_1782.n5 3.38874
R13894 a_8881_1782.n130 a_8881_1782.n141 3.17178
R13895 a_8881_1782.n70 a_8881_1782.n64 3.01226
R13896 a_8881_1782.n81 a_8881_1782.n80 3.01226
R13897 a_8881_1782.n105 a_8881_1782.n99 3.01226
R13898 a_8881_1782.n98 a_8881_1782.n96 3.01226
R13899 a_8881_1782.n5 a_8881_1782.n4 3.01226
R13900 a_8881_1782.t1 a_8881_1782.n151 2.77
R13901 a_8881_1782.n63 a_8881_1782.n61 2.63579
R13902 a_8881_1782.n88 a_8881_1782.n87 2.63579
R13903 a_8881_1782.n118 a_8881_1782.n117 2.63579
R13904 a_8881_1782.n125 a_8881_1782.n124 2.63579
R13905 a_8881_1782.n16 a_8881_1782.n15 2.63579
R13906 a_8881_1782.n15 a_8881_1782.n11 2.63579
R13907 a_8881_1782.n53 a_8881_1782.n21 2.41452
R13908 a_8881_1782.n107 a_8881_1782.n127 2.28493
R13909 a_8881_1782.n49 a_8881_1782.n48 2.25932
R13910 a_8881_1782.n52 a_8881_1782.n51 2.25932
R13911 a_8881_1782.n47 a_8881_1782.n46 1.96602
R13912 a_8881_1782.n30 a_8881_1782.n37 1.88285
R13913 a_8881_1782.n37 a_8881_1782.n33 1.88285
R13914 a_8881_1782.n151 a_8881_1782.n150 1.84417
R13915 a_8881_1782.n81 a_8881_1782.n78 1.50638
R13916 a_8881_1782.n118 a_8881_1782.n115 1.50638
R13917 a_8881_1782.n117 a_8881_1782.n116 1.50638
R13918 a_8881_1782.n27 a_8881_1782.n26 1.50638
R13919 a_8881_1782.n41 a_8881_1782.n40 1.50638
R13920 a_8881_1782.n151 a_8881_1782.n140 1.32032
R13921 a_8881_1782.n151 a_8881_1782.n148 1.29978
R13922 a_8881_1782.n18 a_8881_1782.n129 1.24675
R13923 a_8881_1782.n107 a_8881_1782.n92 1.21366
R13924 a_8881_1782.n71 a_8881_1782.n89 1.15702
R13925 a_8881_1782.n73 a_8881_1782.n56 1.21147
R13926 a_8881_1782.n106 a_8881_1782.n126 1.15482
R13927 a_8881_1782.n63 a_8881_1782.n62 1.12991
R13928 a_8881_1782.n80 a_8881_1782.n79 1.12991
R13929 a_8881_1782.n98 a_8881_1782.n97 1.12991
R13930 a_8881_1782.n26 a_8881_1782.n22 1.12991
R13931 a_8881_1782.n68 a_8881_1782.n67 1.09595
R13932 a_8881_1782.n85 a_8881_1782.n84 1.09595
R13933 a_8881_1782.n1 a_8881_1782.n132 1.04835
R13934 a_8881_1782.n147 a_8881_1782.n127 0.996877
R13935 a_8881_1782.n103 a_8881_1782.n102 0.994314
R13936 a_8881_1782.n122 a_8881_1782.n121 0.994314
R13937 a_8881_1782.n17 a_8881_1782.n53 0.994096
R13938 a_8881_1782.n72 a_8881_1782.n128 0.963
R13939 a_8881_1782.n69 a_8881_1782.n65 0.753441
R13940 a_8881_1782.n104 a_8881_1782.n100 0.753441
R13941 a_8881_1782.n137 a_8881_1782.n135 0.753441
R13942 a_8881_1782.n140 a_8881_1782.n1 0.418831
R13943 a_8881_1782.n148 a_8881_1782.n147 0.386668
R13944 a_8881_1782.n48 a_8881_1782.n44 0.376971
R13945 a_8881_1782.n144 a_8881_1782.n142 0.376971
R13946 a_8881_1782.n7 a_8881_1782.n6 0.319725
R13947 a_8881_1782.n135 a_8881_1782.n136 0.121922
R13948 a_8881_1782.n142 a_8881_1782.n143 0.110027
R13949 a_8881_1782.n147 a_8881_1782.n131 0.0843535
R13950 a_8881_1782.n53 a_8881_1782.n50 0.0827519
R13951 a_8881_1782.n107 a_8881_1782.n106 0.0590938
R13952 a_8881_1782.n42 a_8881_1782.n39 0.100109
R13953 a_8881_1782.n126 a_8881_1782.n119 0.0371012
R13954 a_8881_1782.n131 a_8881_1782.n130 0.0337031
R13955 a_8881_1782.n20 a_8881_1782.n18 0.0287031
R13956 a_8881_1782.n20 a_8881_1782.n19 0.028
R13957 a_8881_1782.n128 a_8881_1782.n107 0.028
R13958 a_8881_1782.n129 a_8881_1782.n73 0.028
R13959 a_8881_1782.n73 a_8881_1782.n72 0.0276737
R13960 a_8881_1782.n113 a_8881_1782.n111 0.0239375
R13961 a_8881_1782.n77 a_8881_1782.n76 4.5892
R13962 a_8881_1782.n114 a_8881_1782.n113 0.0892218
R13963 a_8881_1782.n93 a_8881_1782.n94 0.0883906
R13964 a_8881_1782.n57 a_8881_1782.n58 4.58839
R13965 a_8881_1782.n20 a_8881_1782.n17 0.119641
R13966 a_8881_1782.n28 a_8881_1782.n30 4.61452
R13967 a_8881_1782.n73 a_8881_1782.n71 0.0590938
R13968 a_8881_1782.n82 a_8881_1782.n77 0.0454219
R13969 a_8881_1782.n119 a_8881_1782.n114 0.0454219
R13970 a_8881_1782.n91 a_8881_1782.n93 0.0454219
R13971 a_8881_1782.n55 a_8881_1782.n57 0.0454219
R13972 a_8881_1782.n92 a_8881_1782.n91 0.0388205
R13973 a_8881_1782.n89 a_8881_1782.n82 0.0385721
R13974 a_8881_1782.n56 a_8881_1782.n55 0.0373496
R13975 a_8881_1782.n50 a_8881_1782.n42 0.0337031
R13976 a_8881_1782.n39 a_8881_1782.n29 0.0337031
R13977 a_8881_1782.n29 a_8881_1782.n28 0.0268395
R13978 a_8881_1782.n20 a_8881_1782.n8 1.5962
R13979 a_8881_1782.n1 a_8881_1782.n0 0.225375
R13980 DVSS.n1176 DVSS.n1174 20457
R13981 DVSS.n2869 DVSS.n2868 13448.3
R13982 DVSS.n1789 DVSS.n1788 11429.2
R13983 DVSS.n2411 DVSS.n2410 10331.4
R13984 DVSS.n538 DVSS.t48 6704.1
R13985 DVSS.n2412 DVSS.n2411 5819.7
R13986 DVSS.n2868 DVSS.n2866 4526.13
R13987 DVSS.n1149 DVSS.n1148 3433.78
R13988 DVSS.n539 DVSS.n538 3379.34
R13989 DVSS.n2870 DVSS.n2869 3274.06
R13990 DVSS.n1762 DVSS.n1761 2954.65
R13991 DVSS.n2973 DVSS.n2972 2607.41
R13992 DVSS.t8 DVSS.t6 2310
R13993 DVSS.n1799 DVSS.n1798 2223.27
R13994 DVSS.n9 DVSS.n8 2223.27
R13995 DVSS.t52 DVSS.t54 2165.3
R13996 DVSS.t48 DVSS.t50 2165.3
R13997 DVSS.n2758 DVSS.n2757 2063.77
R13998 DVSS.n2520 DVSS.n2519 2061.08
R13999 DVSS.n3091 DVSS.n3090 1741.13
R14000 DVSS.n2866 DVSS.n2865 1506.58
R14001 DVSS.n2972 DVSS.n2971 1280.42
R14002 DVSS.n482 DVSS.t8 1265
R14003 DVSS.n2665 DVSS.n2664 1172.41
R14004 DVSS.n1761 DVSS.n1760 1105.62
R14005 DVSS.n2663 DVSS.t52 1068.77
R14006 DVSS.n2140 DVSS.n2003 1013.97
R14007 DVSS.n2138 DVSS.n2004 1013.97
R14008 DVSS.n2130 DVSS.n2129 1013.97
R14009 DVSS.n2132 DVSS.n2124 1013.97
R14010 DVSS.n1522 DVSS.n1385 1013.97
R14011 DVSS.n1520 DVSS.n1386 1013.97
R14012 DVSS.n1512 DVSS.n1511 1013.97
R14013 DVSS.n1514 DVSS.n1506 1013.97
R14014 DVSS.n909 DVSS.n772 1013.97
R14015 DVSS.n907 DVSS.n773 1013.97
R14016 DVSS.n899 DVSS.n898 1013.97
R14017 DVSS.n901 DVSS.n893 1013.97
R14018 DVSS.n320 DVSS.n183 1013.97
R14019 DVSS.n318 DVSS.n184 1013.97
R14020 DVSS.n310 DVSS.n309 1013.97
R14021 DVSS.n312 DVSS.n304 1013.97
R14022 DVSS.n1148 DVSS.n1147 913.518
R14023 DVSS.n530 DVSS.t3 868.74
R14024 DVSS.n2519 DVSS.n1203 794.067
R14025 DVSS.n2757 DVSS.n2756 794.067
R14026 DVSS.n2019 DVSS.n2011 728.663
R14027 DVSS.n2160 DVSS.n1985 728.663
R14028 DVSS.n1401 DVSS.n1393 728.663
R14029 DVSS.n1542 DVSS.n1367 728.663
R14030 DVSS.n788 DVSS.n780 728.663
R14031 DVSS.n929 DVSS.n754 728.663
R14032 DVSS.n199 DVSS.n191 728.663
R14033 DVSS.n340 DVSS.n165 728.663
R14034 DVSS.n2866 DVSS.n481 721.253
R14035 DVSS.n2115 DVSS.n2010 668.5
R14036 DVSS.n2113 DVSS.n2013 668.5
R14037 DVSS.n2162 DVSS.n1982 668.5
R14038 DVSS.n2122 DVSS.n1986 668.5
R14039 DVSS.n2090 DVSS.n2069 668.5
R14040 DVSS.n2094 DVSS.n2071 668.5
R14041 DVSS.n2105 DVSS.n2067 668.5
R14042 DVSS.n2108 DVSS.n2107 668.5
R14043 DVSS.n1935 DVSS.n1907 668.5
R14044 DVSS.n1920 DVSS.n1905 668.5
R14045 DVSS.n2277 DVSS.n2276 668.5
R14046 DVSS.n2292 DVSS.n2291 668.5
R14047 DVSS.n1497 DVSS.n1392 668.5
R14048 DVSS.n1495 DVSS.n1395 668.5
R14049 DVSS.n1544 DVSS.n1364 668.5
R14050 DVSS.n1504 DVSS.n1368 668.5
R14051 DVSS.n1472 DVSS.n1451 668.5
R14052 DVSS.n1476 DVSS.n1453 668.5
R14053 DVSS.n1487 DVSS.n1449 668.5
R14054 DVSS.n1490 DVSS.n1489 668.5
R14055 DVSS.n1317 DVSS.n1289 668.5
R14056 DVSS.n1302 DVSS.n1287 668.5
R14057 DVSS.n1659 DVSS.n1658 668.5
R14058 DVSS.n1674 DVSS.n1673 668.5
R14059 DVSS.n884 DVSS.n779 668.5
R14060 DVSS.n882 DVSS.n782 668.5
R14061 DVSS.n931 DVSS.n751 668.5
R14062 DVSS.n891 DVSS.n755 668.5
R14063 DVSS.n859 DVSS.n838 668.5
R14064 DVSS.n863 DVSS.n840 668.5
R14065 DVSS.n874 DVSS.n836 668.5
R14066 DVSS.n877 DVSS.n876 668.5
R14067 DVSS.n704 DVSS.n676 668.5
R14068 DVSS.n689 DVSS.n674 668.5
R14069 DVSS.n1046 DVSS.n1045 668.5
R14070 DVSS.n1061 DVSS.n1060 668.5
R14071 DVSS.n295 DVSS.n190 668.5
R14072 DVSS.n293 DVSS.n193 668.5
R14073 DVSS.n342 DVSS.n162 668.5
R14074 DVSS.n302 DVSS.n166 668.5
R14075 DVSS.n270 DVSS.n249 668.5
R14076 DVSS.n274 DVSS.n251 668.5
R14077 DVSS.n285 DVSS.n247 668.5
R14078 DVSS.n288 DVSS.n287 668.5
R14079 DVSS.n115 DVSS.n87 668.5
R14080 DVSS.n100 DVSS.n85 668.5
R14081 DVSS.n457 DVSS.n456 668.5
R14082 DVSS.n472 DVSS.n471 668.5
R14083 DVSS.n2868 DVSS.n2867 648.317
R14084 DVSS.t174 DVSS.n482 643.51
R14085 DVSS.n2640 DVSS.n2639 602.423
R14086 DVSS.n2544 DVSS.n2543 579.216
R14087 DVSS.n2204 DVSS.n1869 562.173
R14088 DVSS.n2252 DVSS.n1853 562.173
R14089 DVSS.n1586 DVSS.n1251 562.173
R14090 DVSS.n1634 DVSS.n1235 562.173
R14091 DVSS.n973 DVSS.n638 562.173
R14092 DVSS.n1021 DVSS.n622 562.173
R14093 DVSS.n384 DVSS.n49 562.173
R14094 DVSS.n432 DVSS.n33 562.173
R14095 DVSS.n2865 DVSS.t87 538.777
R14096 DVSS.n2131 DVSS.n2127 535.801
R14097 DVSS.n1513 DVSS.n1509 535.801
R14098 DVSS.n900 DVSS.n896 535.801
R14099 DVSS.n311 DVSS.n307 535.801
R14100 DVSS.n2092 DVSS.n2070 518.471
R14101 DVSS.n2106 DVSS.n2019 518.471
R14102 DVSS.n2114 DVSS.n2011 518.471
R14103 DVSS.n2160 DVSS.n1984 518.471
R14104 DVSS.n1474 DVSS.n1452 518.471
R14105 DVSS.n1488 DVSS.n1401 518.471
R14106 DVSS.n1496 DVSS.n1393 518.471
R14107 DVSS.n1542 DVSS.n1366 518.471
R14108 DVSS.n861 DVSS.n839 518.471
R14109 DVSS.n875 DVSS.n788 518.471
R14110 DVSS.n883 DVSS.n780 518.471
R14111 DVSS.n929 DVSS.n753 518.471
R14112 DVSS.n272 DVSS.n250 518.471
R14113 DVSS.n286 DVSS.n199 518.471
R14114 DVSS.n294 DVSS.n191 518.471
R14115 DVSS.n340 DVSS.n164 518.471
R14116 DVSS.n1934 DVSS.n1906 491.349
R14117 DVSS.n2190 DVSS.n1869 491.349
R14118 DVSS.n1853 DVSS.n1844 491.349
R14119 DVSS.n2274 DVSS.n1838 491.349
R14120 DVSS.n1316 DVSS.n1288 491.349
R14121 DVSS.n1572 DVSS.n1251 491.349
R14122 DVSS.n1235 DVSS.n1226 491.349
R14123 DVSS.n1656 DVSS.n1220 491.349
R14124 DVSS.n703 DVSS.n675 491.349
R14125 DVSS.n959 DVSS.n638 491.349
R14126 DVSS.n622 DVSS.n613 491.349
R14127 DVSS.n1043 DVSS.n607 491.349
R14128 DVSS.n114 DVSS.n86 491.349
R14129 DVSS.n370 DVSS.n49 491.349
R14130 DVSS.n33 DVSS.n24 491.349
R14131 DVSS.n454 DVSS.n18 491.349
R14132 DVSS.n3090 DVSS.n3089 488.889
R14133 DVSS.n2126 DVSS.n1985 448.409
R14134 DVSS.n1508 DVSS.n1367 448.409
R14135 DVSS.n895 DVSS.n754 448.409
R14136 DVSS.n306 DVSS.n165 448.409
R14137 DVSS.n3008 DVSS.t145 403.12
R14138 DVSS.t59 DVSS.t85 394.712
R14139 DVSS.n2124 DVSS.n2004 394
R14140 DVSS.n1506 DVSS.n1386 394
R14141 DVSS.n893 DVSS.n773 394
R14142 DVSS.n304 DVSS.n184 394
R14143 DVSS.t3 DVSS.t90 390.324
R14144 DVSS.n2228 DVSS.n1851 366.841
R14145 DVSS.n2243 DVSS.n1855 366.841
R14146 DVSS.n1882 DVSS.n1868 366.841
R14147 DVSS.n1898 DVSS.n1871 366.841
R14148 DVSS.n1610 DVSS.n1233 366.841
R14149 DVSS.n1625 DVSS.n1237 366.841
R14150 DVSS.n1264 DVSS.n1250 366.841
R14151 DVSS.n1280 DVSS.n1253 366.841
R14152 DVSS.n997 DVSS.n620 366.841
R14153 DVSS.n1012 DVSS.n624 366.841
R14154 DVSS.n651 DVSS.n637 366.841
R14155 DVSS.n667 DVSS.n640 366.841
R14156 DVSS.n408 DVSS.n31 366.841
R14157 DVSS.n423 DVSS.n35 366.841
R14158 DVSS.n62 DVSS.n48 366.841
R14159 DVSS.n78 DVSS.n51 366.841
R14160 DVSS.n3036 DVSS.n3035 359.185
R14161 DVSS.n3036 DVSS.t32 351.022
R14162 DVSS.t85 DVSS.n537 349.909
R14163 DVSS.n1176 DVSS.n1175 343.353
R14164 DVSS.n1158 DVSS.n1157 332.425
R14165 DVSS.n2100 DVSS.n2070 317.623
R14166 DVSS.n2106 DVSS.n2018 317.623
R14167 DVSS.n2114 DVSS.n2012 317.623
R14168 DVSS.n2120 DVSS.n1984 317.623
R14169 DVSS.n1482 DVSS.n1452 317.623
R14170 DVSS.n1488 DVSS.n1400 317.623
R14171 DVSS.n1496 DVSS.n1394 317.623
R14172 DVSS.n1502 DVSS.n1366 317.623
R14173 DVSS.n869 DVSS.n839 317.623
R14174 DVSS.n875 DVSS.n787 317.623
R14175 DVSS.n883 DVSS.n781 317.623
R14176 DVSS.n889 DVSS.n753 317.623
R14177 DVSS.n280 DVSS.n250 317.623
R14178 DVSS.n286 DVSS.n198 317.623
R14179 DVSS.n294 DVSS.n192 317.623
R14180 DVSS.n300 DVSS.n164 317.623
R14181 DVSS.n3017 DVSS.t141 317.349
R14182 DVSS.n2203 DVSS.n1871 306.26
R14183 DVSS.n2251 DVSS.n1855 306.26
R14184 DVSS.n2205 DVSS.n1868 306.26
R14185 DVSS.n2253 DVSS.n1851 306.26
R14186 DVSS.n1585 DVSS.n1253 306.26
R14187 DVSS.n1633 DVSS.n1237 306.26
R14188 DVSS.n1587 DVSS.n1250 306.26
R14189 DVSS.n1635 DVSS.n1233 306.26
R14190 DVSS.n972 DVSS.n640 306.26
R14191 DVSS.n1020 DVSS.n624 306.26
R14192 DVSS.n974 DVSS.n637 306.26
R14193 DVSS.n1022 DVSS.n620 306.26
R14194 DVSS.n383 DVSS.n51 306.26
R14195 DVSS.n431 DVSS.n35 306.26
R14196 DVSS.n385 DVSS.n48 306.26
R14197 DVSS.n433 DVSS.n31 306.26
R14198 DVSS.n2184 DVSS.n1906 301.007
R14199 DVSS.n2190 DVSS.n1902 301.007
R14200 DVSS.n2204 DVSS.n1870 301.007
R14201 DVSS.n2211 DVSS.n1864 301.007
R14202 DVSS.n2252 DVSS.n1852 301.007
R14203 DVSS.n2282 DVSS.n1844 301.007
R14204 DVSS.n1846 DVSS.n1838 301.007
R14205 DVSS.n1566 DVSS.n1288 301.007
R14206 DVSS.n1572 DVSS.n1284 301.007
R14207 DVSS.n1586 DVSS.n1252 301.007
R14208 DVSS.n1593 DVSS.n1246 301.007
R14209 DVSS.n1634 DVSS.n1234 301.007
R14210 DVSS.n1664 DVSS.n1226 301.007
R14211 DVSS.n1228 DVSS.n1220 301.007
R14212 DVSS.n953 DVSS.n675 301.007
R14213 DVSS.n959 DVSS.n671 301.007
R14214 DVSS.n973 DVSS.n639 301.007
R14215 DVSS.n980 DVSS.n633 301.007
R14216 DVSS.n1021 DVSS.n621 301.007
R14217 DVSS.n1051 DVSS.n613 301.007
R14218 DVSS.n615 DVSS.n607 301.007
R14219 DVSS.n364 DVSS.n86 301.007
R14220 DVSS.n370 DVSS.n82 301.007
R14221 DVSS.n384 DVSS.n50 301.007
R14222 DVSS.n391 DVSS.n44 301.007
R14223 DVSS.n432 DVSS.n32 301.007
R14224 DVSS.n462 DVSS.n24 301.007
R14225 DVSS.n26 DVSS.n18 301.007
R14226 DVSS.n2312 DVSS.t73 294.885
R14227 DVSS.n1694 DVSS.t186 294.885
R14228 DVSS.n1081 DVSS.t131 294.885
R14229 DVSS.n2881 DVSS.t25 294.885
R14230 DVSS.n2107 DVSS.n2014 292.5
R14231 DVSS.n2107 DVSS.n2106 292.5
R14232 DVSS.n2123 DVSS.n2122 292.5
R14233 DVSS.n2122 DVSS.n1984 292.5
R14234 DVSS.n2090 DVSS.n2089 292.5
R14235 DVSS.n2088 DVSS.n2077 292.5
R14236 DVSS.n2087 DVSS.n2086 292.5
R14237 DVSS.n2085 DVSS.n2084 292.5
R14238 DVSS.n2083 DVSS.n2082 292.5
R14239 DVSS.n2081 DVSS.n2080 292.5
R14240 DVSS.n2079 DVSS.n2078 292.5
R14241 DVSS.n2073 DVSS.n2072 292.5
R14242 DVSS.n2121 DVSS.n2006 292.5
R14243 DVSS.n2121 DVSS.n2120 292.5
R14244 DVSS.n2111 DVSS.n2007 292.5
R14245 DVSS.n2012 DVSS.n2007 292.5
R14246 DVSS.n2099 DVSS.n2098 292.5
R14247 DVSS.n2100 DVSS.n2099 292.5
R14248 DVSS.n2097 DVSS.n2017 292.5
R14249 DVSS.n2018 DVSS.n2017 292.5
R14250 DVSS.n2113 DVSS.n2112 292.5
R14251 DVSS.n2114 DVSS.n2113 292.5
R14252 DVSS.n2095 DVSS.n2094 292.5
R14253 DVSS.n2096 DVSS.n2071 292.5
R14254 DVSS.n2071 DVSS.n2070 292.5
R14255 DVSS.n2134 DVSS.n2124 292.5
R14256 DVSS.n2127 DVSS.n2124 292.5
R14257 DVSS.n2135 DVSS.n2004 292.5
R14258 DVSS.n2126 DVSS.n2004 292.5
R14259 DVSS.n2133 DVSS.n2132 292.5
R14260 DVSS.n2130 DVSS.n2125 292.5
R14261 DVSS.n2141 DVSS.n2140 292.5
R14262 DVSS.n2143 DVSS.n2142 292.5
R14263 DVSS.n2005 DVSS.n1986 292.5
R14264 DVSS.n2160 DVSS.n1986 292.5
R14265 DVSS.n2138 DVSS.n2137 292.5
R14266 DVSS.n2129 DVSS.n2127 292.5
R14267 DVSS.n2126 DVSS.n2003 292.5
R14268 DVSS.n2001 DVSS.n2000 292.5
R14269 DVSS.n2149 DVSS.n2148 292.5
R14270 DVSS.n2152 DVSS.n2151 292.5
R14271 DVSS.n1995 DVSS.n1994 292.5
R14272 DVSS.n2158 DVSS.n2157 292.5
R14273 DVSS.n1992 DVSS.n1983 292.5
R14274 DVSS.n2163 DVSS.n2162 292.5
R14275 DVSS.n1982 DVSS.n1980 292.5
R14276 DVSS.n1984 DVSS.n1982 292.5
R14277 DVSS.n2119 DVSS.n2118 292.5
R14278 DVSS.n2120 DVSS.n2119 292.5
R14279 DVSS.n2117 DVSS.n2008 292.5
R14280 DVSS.n2012 DVSS.n2008 292.5
R14281 DVSS.n2116 DVSS.n2115 292.5
R14282 DVSS.n2115 DVSS.n2114 292.5
R14283 DVSS.n2069 DVSS.n2068 292.5
R14284 DVSS.n2070 DVSS.n2069 292.5
R14285 DVSS.n2102 DVSS.n2101 292.5
R14286 DVSS.n2101 DVSS.n2100 292.5
R14287 DVSS.n2103 DVSS.n2020 292.5
R14288 DVSS.n2020 DVSS.n2018 292.5
R14289 DVSS.n2105 DVSS.n2104 292.5
R14290 DVSS.n2106 DVSS.n2105 292.5
R14291 DVSS.n2109 DVSS.n2013 292.5
R14292 DVSS.n2067 DVSS.n2066 292.5
R14293 DVSS.n2066 DVSS.n2010 292.5
R14294 DVSS.n2025 DVSS.n2023 292.5
R14295 DVSS.n2030 DVSS.n2023 292.5
R14296 DVSS.n2061 DVSS.n2027 292.5
R14297 DVSS.n2061 DVSS.n2060 292.5
R14298 DVSS.n2035 DVSS.n2032 292.5
R14299 DVSS.n2059 DVSS.n2032 292.5
R14300 DVSS.n2056 DVSS.n2037 292.5
R14301 DVSS.n2057 DVSS.n2056 292.5
R14302 DVSS.n2042 DVSS.n2038 292.5
R14303 DVSS.n2038 DVSS.n2033 292.5
R14304 DVSS.n2051 DVSS.n2044 292.5
R14305 DVSS.n2051 DVSS.n2050 292.5
R14306 DVSS.n2049 DVSS.n2047 292.5
R14307 DVSS.n2047 DVSS.n2046 292.5
R14308 DVSS.n2109 DVSS.n2108 292.5
R14309 DVSS.n1921 DVSS.n1920 292.5
R14310 DVSS.n1912 DVSS.n1911 292.5
R14311 DVSS.n1924 DVSS.n1923 292.5
R14312 DVSS.n1926 DVSS.n1925 292.5
R14313 DVSS.n1928 DVSS.n1927 292.5
R14314 DVSS.n1930 DVSS.n1929 292.5
R14315 DVSS.n1932 DVSS.n1931 292.5
R14316 DVSS.n1922 DVSS.n1919 292.5
R14317 DVSS.n1936 DVSS.n1935 292.5
R14318 DVSS.n1935 DVSS.n1934 292.5
R14319 DVSS.n2228 DVSS.n1848 292.5
R14320 DVSS.n2228 DVSS.n1853 292.5
R14321 DVSS.n2241 DVSS.n2224 292.5
R14322 DVSS.n2240 DVSS.n2239 292.5
R14323 DVSS.n2238 DVSS.n2237 292.5
R14324 DVSS.n2236 DVSS.n2226 292.5
R14325 DVSS.n2234 DVSS.n2233 292.5
R14326 DVSS.n2232 DVSS.n2227 292.5
R14327 DVSS.n2231 DVSS.n2230 292.5
R14328 DVSS.n2244 DVSS.n2243 292.5
R14329 DVSS.n1884 DVSS.n1880 292.5
R14330 DVSS.n1897 DVSS.n1876 292.5
R14331 DVSS.n1895 DVSS.n1894 292.5
R14332 DVSS.n1893 DVSS.n1892 292.5
R14333 DVSS.n1890 DVSS.n1878 292.5
R14334 DVSS.n1888 DVSS.n1887 292.5
R14335 DVSS.n1886 DVSS.n1885 292.5
R14336 DVSS.n1899 DVSS.n1898 292.5
R14337 DVSS.n1898 DVSS.n1869 292.5
R14338 DVSS.n1882 DVSS.n1881 292.5
R14339 DVSS.n2278 DVSS.n2277 292.5
R14340 DVSS.n2277 DVSS.n1838 292.5
R14341 DVSS.n2279 DVSS.n1847 292.5
R14342 DVSS.n1847 DVSS.n1846 292.5
R14343 DVSS.n2281 DVSS.n2280 292.5
R14344 DVSS.n2282 DVSS.n2281 292.5
R14345 DVSS.n2256 DVSS.n1845 292.5
R14346 DVSS.n1845 DVSS.n1844 292.5
R14347 DVSS.n2254 DVSS.n2253 292.5
R14348 DVSS.n2253 DVSS.n2252 292.5
R14349 DVSS.n1850 DVSS.n1849 292.5
R14350 DVSS.n1852 DVSS.n1850 292.5
R14351 DVSS.n2208 DVSS.n1866 292.5
R14352 DVSS.n1866 DVSS.n1864 292.5
R14353 DVSS.n2210 DVSS.n2209 292.5
R14354 DVSS.n2211 DVSS.n2210 292.5
R14355 DVSS.n2207 DVSS.n1865 292.5
R14356 DVSS.n1870 DVSS.n1865 292.5
R14357 DVSS.n2206 DVSS.n2205 292.5
R14358 DVSS.n2205 DVSS.n2204 292.5
R14359 DVSS.n2189 DVSS.n2188 292.5
R14360 DVSS.n2190 DVSS.n2189 292.5
R14361 DVSS.n2187 DVSS.n1903 292.5
R14362 DVSS.n1903 DVSS.n1902 292.5
R14363 DVSS.n2186 DVSS.n2185 292.5
R14364 DVSS.n2185 DVSS.n2184 292.5
R14365 DVSS.n1905 DVSS.n1904 292.5
R14366 DVSS.n1906 DVSS.n1905 292.5
R14367 DVSS.n2276 DVSS.n2257 292.5
R14368 DVSS.n2262 DVSS.n2258 292.5
R14369 DVSS.n2272 DVSS.n2271 292.5
R14370 DVSS.n2270 DVSS.n2261 292.5
R14371 DVSS.n2269 DVSS.n2268 292.5
R14372 DVSS.n2267 DVSS.n2266 292.5
R14373 DVSS.n2265 DVSS.n2264 292.5
R14374 DVSS.n2263 DVSS.n1835 292.5
R14375 DVSS.n2293 DVSS.n2292 292.5
R14376 DVSS.n1489 DVSS.n1396 292.5
R14377 DVSS.n1489 DVSS.n1488 292.5
R14378 DVSS.n1505 DVSS.n1504 292.5
R14379 DVSS.n1504 DVSS.n1366 292.5
R14380 DVSS.n1472 DVSS.n1471 292.5
R14381 DVSS.n1470 DVSS.n1459 292.5
R14382 DVSS.n1469 DVSS.n1468 292.5
R14383 DVSS.n1467 DVSS.n1466 292.5
R14384 DVSS.n1465 DVSS.n1464 292.5
R14385 DVSS.n1463 DVSS.n1462 292.5
R14386 DVSS.n1461 DVSS.n1460 292.5
R14387 DVSS.n1455 DVSS.n1454 292.5
R14388 DVSS.n1503 DVSS.n1388 292.5
R14389 DVSS.n1503 DVSS.n1502 292.5
R14390 DVSS.n1493 DVSS.n1389 292.5
R14391 DVSS.n1394 DVSS.n1389 292.5
R14392 DVSS.n1481 DVSS.n1480 292.5
R14393 DVSS.n1482 DVSS.n1481 292.5
R14394 DVSS.n1479 DVSS.n1399 292.5
R14395 DVSS.n1400 DVSS.n1399 292.5
R14396 DVSS.n1495 DVSS.n1494 292.5
R14397 DVSS.n1496 DVSS.n1495 292.5
R14398 DVSS.n1477 DVSS.n1476 292.5
R14399 DVSS.n1478 DVSS.n1453 292.5
R14400 DVSS.n1453 DVSS.n1452 292.5
R14401 DVSS.n1516 DVSS.n1506 292.5
R14402 DVSS.n1509 DVSS.n1506 292.5
R14403 DVSS.n1517 DVSS.n1386 292.5
R14404 DVSS.n1508 DVSS.n1386 292.5
R14405 DVSS.n1515 DVSS.n1514 292.5
R14406 DVSS.n1512 DVSS.n1507 292.5
R14407 DVSS.n1523 DVSS.n1522 292.5
R14408 DVSS.n1525 DVSS.n1524 292.5
R14409 DVSS.n1387 DVSS.n1368 292.5
R14410 DVSS.n1542 DVSS.n1368 292.5
R14411 DVSS.n1520 DVSS.n1519 292.5
R14412 DVSS.n1511 DVSS.n1509 292.5
R14413 DVSS.n1508 DVSS.n1385 292.5
R14414 DVSS.n1383 DVSS.n1382 292.5
R14415 DVSS.n1531 DVSS.n1530 292.5
R14416 DVSS.n1534 DVSS.n1533 292.5
R14417 DVSS.n1377 DVSS.n1376 292.5
R14418 DVSS.n1540 DVSS.n1539 292.5
R14419 DVSS.n1374 DVSS.n1365 292.5
R14420 DVSS.n1545 DVSS.n1544 292.5
R14421 DVSS.n1364 DVSS.n1362 292.5
R14422 DVSS.n1366 DVSS.n1364 292.5
R14423 DVSS.n1501 DVSS.n1500 292.5
R14424 DVSS.n1502 DVSS.n1501 292.5
R14425 DVSS.n1499 DVSS.n1390 292.5
R14426 DVSS.n1394 DVSS.n1390 292.5
R14427 DVSS.n1498 DVSS.n1497 292.5
R14428 DVSS.n1497 DVSS.n1496 292.5
R14429 DVSS.n1451 DVSS.n1450 292.5
R14430 DVSS.n1452 DVSS.n1451 292.5
R14431 DVSS.n1484 DVSS.n1483 292.5
R14432 DVSS.n1483 DVSS.n1482 292.5
R14433 DVSS.n1485 DVSS.n1402 292.5
R14434 DVSS.n1402 DVSS.n1400 292.5
R14435 DVSS.n1487 DVSS.n1486 292.5
R14436 DVSS.n1488 DVSS.n1487 292.5
R14437 DVSS.n1491 DVSS.n1395 292.5
R14438 DVSS.n1449 DVSS.n1448 292.5
R14439 DVSS.n1448 DVSS.n1392 292.5
R14440 DVSS.n1407 DVSS.n1405 292.5
R14441 DVSS.n1412 DVSS.n1405 292.5
R14442 DVSS.n1443 DVSS.n1409 292.5
R14443 DVSS.n1443 DVSS.n1442 292.5
R14444 DVSS.n1417 DVSS.n1414 292.5
R14445 DVSS.n1441 DVSS.n1414 292.5
R14446 DVSS.n1438 DVSS.n1419 292.5
R14447 DVSS.n1439 DVSS.n1438 292.5
R14448 DVSS.n1424 DVSS.n1420 292.5
R14449 DVSS.n1420 DVSS.n1415 292.5
R14450 DVSS.n1433 DVSS.n1426 292.5
R14451 DVSS.n1433 DVSS.n1432 292.5
R14452 DVSS.n1431 DVSS.n1429 292.5
R14453 DVSS.n1429 DVSS.n1428 292.5
R14454 DVSS.n1491 DVSS.n1490 292.5
R14455 DVSS.n1303 DVSS.n1302 292.5
R14456 DVSS.n1294 DVSS.n1293 292.5
R14457 DVSS.n1306 DVSS.n1305 292.5
R14458 DVSS.n1308 DVSS.n1307 292.5
R14459 DVSS.n1310 DVSS.n1309 292.5
R14460 DVSS.n1312 DVSS.n1311 292.5
R14461 DVSS.n1314 DVSS.n1313 292.5
R14462 DVSS.n1304 DVSS.n1301 292.5
R14463 DVSS.n1318 DVSS.n1317 292.5
R14464 DVSS.n1317 DVSS.n1316 292.5
R14465 DVSS.n1610 DVSS.n1230 292.5
R14466 DVSS.n1610 DVSS.n1235 292.5
R14467 DVSS.n1623 DVSS.n1606 292.5
R14468 DVSS.n1622 DVSS.n1621 292.5
R14469 DVSS.n1620 DVSS.n1619 292.5
R14470 DVSS.n1618 DVSS.n1608 292.5
R14471 DVSS.n1616 DVSS.n1615 292.5
R14472 DVSS.n1614 DVSS.n1609 292.5
R14473 DVSS.n1613 DVSS.n1612 292.5
R14474 DVSS.n1626 DVSS.n1625 292.5
R14475 DVSS.n1266 DVSS.n1262 292.5
R14476 DVSS.n1279 DVSS.n1258 292.5
R14477 DVSS.n1277 DVSS.n1276 292.5
R14478 DVSS.n1275 DVSS.n1274 292.5
R14479 DVSS.n1272 DVSS.n1260 292.5
R14480 DVSS.n1270 DVSS.n1269 292.5
R14481 DVSS.n1268 DVSS.n1267 292.5
R14482 DVSS.n1281 DVSS.n1280 292.5
R14483 DVSS.n1280 DVSS.n1251 292.5
R14484 DVSS.n1264 DVSS.n1263 292.5
R14485 DVSS.n1660 DVSS.n1659 292.5
R14486 DVSS.n1659 DVSS.n1220 292.5
R14487 DVSS.n1661 DVSS.n1229 292.5
R14488 DVSS.n1229 DVSS.n1228 292.5
R14489 DVSS.n1663 DVSS.n1662 292.5
R14490 DVSS.n1664 DVSS.n1663 292.5
R14491 DVSS.n1638 DVSS.n1227 292.5
R14492 DVSS.n1227 DVSS.n1226 292.5
R14493 DVSS.n1636 DVSS.n1635 292.5
R14494 DVSS.n1635 DVSS.n1634 292.5
R14495 DVSS.n1232 DVSS.n1231 292.5
R14496 DVSS.n1234 DVSS.n1232 292.5
R14497 DVSS.n1590 DVSS.n1248 292.5
R14498 DVSS.n1248 DVSS.n1246 292.5
R14499 DVSS.n1592 DVSS.n1591 292.5
R14500 DVSS.n1593 DVSS.n1592 292.5
R14501 DVSS.n1589 DVSS.n1247 292.5
R14502 DVSS.n1252 DVSS.n1247 292.5
R14503 DVSS.n1588 DVSS.n1587 292.5
R14504 DVSS.n1587 DVSS.n1586 292.5
R14505 DVSS.n1571 DVSS.n1570 292.5
R14506 DVSS.n1572 DVSS.n1571 292.5
R14507 DVSS.n1569 DVSS.n1285 292.5
R14508 DVSS.n1285 DVSS.n1284 292.5
R14509 DVSS.n1568 DVSS.n1567 292.5
R14510 DVSS.n1567 DVSS.n1566 292.5
R14511 DVSS.n1287 DVSS.n1286 292.5
R14512 DVSS.n1288 DVSS.n1287 292.5
R14513 DVSS.n1658 DVSS.n1639 292.5
R14514 DVSS.n1644 DVSS.n1640 292.5
R14515 DVSS.n1654 DVSS.n1653 292.5
R14516 DVSS.n1652 DVSS.n1643 292.5
R14517 DVSS.n1651 DVSS.n1650 292.5
R14518 DVSS.n1649 DVSS.n1648 292.5
R14519 DVSS.n1647 DVSS.n1646 292.5
R14520 DVSS.n1645 DVSS.n1217 292.5
R14521 DVSS.n1675 DVSS.n1674 292.5
R14522 DVSS.n876 DVSS.n783 292.5
R14523 DVSS.n876 DVSS.n875 292.5
R14524 DVSS.n892 DVSS.n891 292.5
R14525 DVSS.n891 DVSS.n753 292.5
R14526 DVSS.n859 DVSS.n858 292.5
R14527 DVSS.n857 DVSS.n846 292.5
R14528 DVSS.n856 DVSS.n855 292.5
R14529 DVSS.n854 DVSS.n853 292.5
R14530 DVSS.n852 DVSS.n851 292.5
R14531 DVSS.n850 DVSS.n849 292.5
R14532 DVSS.n848 DVSS.n847 292.5
R14533 DVSS.n842 DVSS.n841 292.5
R14534 DVSS.n890 DVSS.n775 292.5
R14535 DVSS.n890 DVSS.n889 292.5
R14536 DVSS.n880 DVSS.n776 292.5
R14537 DVSS.n781 DVSS.n776 292.5
R14538 DVSS.n868 DVSS.n867 292.5
R14539 DVSS.n869 DVSS.n868 292.5
R14540 DVSS.n866 DVSS.n786 292.5
R14541 DVSS.n787 DVSS.n786 292.5
R14542 DVSS.n882 DVSS.n881 292.5
R14543 DVSS.n883 DVSS.n882 292.5
R14544 DVSS.n864 DVSS.n863 292.5
R14545 DVSS.n865 DVSS.n840 292.5
R14546 DVSS.n840 DVSS.n839 292.5
R14547 DVSS.n903 DVSS.n893 292.5
R14548 DVSS.n896 DVSS.n893 292.5
R14549 DVSS.n904 DVSS.n773 292.5
R14550 DVSS.n895 DVSS.n773 292.5
R14551 DVSS.n902 DVSS.n901 292.5
R14552 DVSS.n899 DVSS.n894 292.5
R14553 DVSS.n910 DVSS.n909 292.5
R14554 DVSS.n912 DVSS.n911 292.5
R14555 DVSS.n774 DVSS.n755 292.5
R14556 DVSS.n929 DVSS.n755 292.5
R14557 DVSS.n907 DVSS.n906 292.5
R14558 DVSS.n898 DVSS.n896 292.5
R14559 DVSS.n895 DVSS.n772 292.5
R14560 DVSS.n770 DVSS.n769 292.5
R14561 DVSS.n918 DVSS.n917 292.5
R14562 DVSS.n921 DVSS.n920 292.5
R14563 DVSS.n764 DVSS.n763 292.5
R14564 DVSS.n927 DVSS.n926 292.5
R14565 DVSS.n761 DVSS.n752 292.5
R14566 DVSS.n932 DVSS.n931 292.5
R14567 DVSS.n751 DVSS.n749 292.5
R14568 DVSS.n753 DVSS.n751 292.5
R14569 DVSS.n888 DVSS.n887 292.5
R14570 DVSS.n889 DVSS.n888 292.5
R14571 DVSS.n886 DVSS.n777 292.5
R14572 DVSS.n781 DVSS.n777 292.5
R14573 DVSS.n885 DVSS.n884 292.5
R14574 DVSS.n884 DVSS.n883 292.5
R14575 DVSS.n838 DVSS.n837 292.5
R14576 DVSS.n839 DVSS.n838 292.5
R14577 DVSS.n871 DVSS.n870 292.5
R14578 DVSS.n870 DVSS.n869 292.5
R14579 DVSS.n872 DVSS.n789 292.5
R14580 DVSS.n789 DVSS.n787 292.5
R14581 DVSS.n874 DVSS.n873 292.5
R14582 DVSS.n875 DVSS.n874 292.5
R14583 DVSS.n878 DVSS.n782 292.5
R14584 DVSS.n836 DVSS.n835 292.5
R14585 DVSS.n835 DVSS.n779 292.5
R14586 DVSS.n794 DVSS.n792 292.5
R14587 DVSS.n799 DVSS.n792 292.5
R14588 DVSS.n830 DVSS.n796 292.5
R14589 DVSS.n830 DVSS.n829 292.5
R14590 DVSS.n804 DVSS.n801 292.5
R14591 DVSS.n828 DVSS.n801 292.5
R14592 DVSS.n825 DVSS.n806 292.5
R14593 DVSS.n826 DVSS.n825 292.5
R14594 DVSS.n811 DVSS.n807 292.5
R14595 DVSS.n807 DVSS.n802 292.5
R14596 DVSS.n820 DVSS.n813 292.5
R14597 DVSS.n820 DVSS.n819 292.5
R14598 DVSS.n818 DVSS.n816 292.5
R14599 DVSS.n816 DVSS.n815 292.5
R14600 DVSS.n878 DVSS.n877 292.5
R14601 DVSS.n690 DVSS.n689 292.5
R14602 DVSS.n681 DVSS.n680 292.5
R14603 DVSS.n693 DVSS.n692 292.5
R14604 DVSS.n695 DVSS.n694 292.5
R14605 DVSS.n697 DVSS.n696 292.5
R14606 DVSS.n699 DVSS.n698 292.5
R14607 DVSS.n701 DVSS.n700 292.5
R14608 DVSS.n691 DVSS.n688 292.5
R14609 DVSS.n705 DVSS.n704 292.5
R14610 DVSS.n704 DVSS.n703 292.5
R14611 DVSS.n997 DVSS.n617 292.5
R14612 DVSS.n997 DVSS.n622 292.5
R14613 DVSS.n1010 DVSS.n993 292.5
R14614 DVSS.n1009 DVSS.n1008 292.5
R14615 DVSS.n1007 DVSS.n1006 292.5
R14616 DVSS.n1005 DVSS.n995 292.5
R14617 DVSS.n1003 DVSS.n1002 292.5
R14618 DVSS.n1001 DVSS.n996 292.5
R14619 DVSS.n1000 DVSS.n999 292.5
R14620 DVSS.n1013 DVSS.n1012 292.5
R14621 DVSS.n653 DVSS.n649 292.5
R14622 DVSS.n666 DVSS.n645 292.5
R14623 DVSS.n664 DVSS.n663 292.5
R14624 DVSS.n662 DVSS.n661 292.5
R14625 DVSS.n659 DVSS.n647 292.5
R14626 DVSS.n657 DVSS.n656 292.5
R14627 DVSS.n655 DVSS.n654 292.5
R14628 DVSS.n668 DVSS.n667 292.5
R14629 DVSS.n667 DVSS.n638 292.5
R14630 DVSS.n651 DVSS.n650 292.5
R14631 DVSS.n1047 DVSS.n1046 292.5
R14632 DVSS.n1046 DVSS.n607 292.5
R14633 DVSS.n1048 DVSS.n616 292.5
R14634 DVSS.n616 DVSS.n615 292.5
R14635 DVSS.n1050 DVSS.n1049 292.5
R14636 DVSS.n1051 DVSS.n1050 292.5
R14637 DVSS.n1025 DVSS.n614 292.5
R14638 DVSS.n614 DVSS.n613 292.5
R14639 DVSS.n1023 DVSS.n1022 292.5
R14640 DVSS.n1022 DVSS.n1021 292.5
R14641 DVSS.n619 DVSS.n618 292.5
R14642 DVSS.n621 DVSS.n619 292.5
R14643 DVSS.n977 DVSS.n635 292.5
R14644 DVSS.n635 DVSS.n633 292.5
R14645 DVSS.n979 DVSS.n978 292.5
R14646 DVSS.n980 DVSS.n979 292.5
R14647 DVSS.n976 DVSS.n634 292.5
R14648 DVSS.n639 DVSS.n634 292.5
R14649 DVSS.n975 DVSS.n974 292.5
R14650 DVSS.n974 DVSS.n973 292.5
R14651 DVSS.n958 DVSS.n957 292.5
R14652 DVSS.n959 DVSS.n958 292.5
R14653 DVSS.n956 DVSS.n672 292.5
R14654 DVSS.n672 DVSS.n671 292.5
R14655 DVSS.n955 DVSS.n954 292.5
R14656 DVSS.n954 DVSS.n953 292.5
R14657 DVSS.n674 DVSS.n673 292.5
R14658 DVSS.n675 DVSS.n674 292.5
R14659 DVSS.n1045 DVSS.n1026 292.5
R14660 DVSS.n1031 DVSS.n1027 292.5
R14661 DVSS.n1041 DVSS.n1040 292.5
R14662 DVSS.n1039 DVSS.n1030 292.5
R14663 DVSS.n1038 DVSS.n1037 292.5
R14664 DVSS.n1036 DVSS.n1035 292.5
R14665 DVSS.n1034 DVSS.n1033 292.5
R14666 DVSS.n1032 DVSS.n604 292.5
R14667 DVSS.n1062 DVSS.n1061 292.5
R14668 DVSS.n287 DVSS.n194 292.5
R14669 DVSS.n287 DVSS.n286 292.5
R14670 DVSS.n303 DVSS.n302 292.5
R14671 DVSS.n302 DVSS.n164 292.5
R14672 DVSS.n270 DVSS.n269 292.5
R14673 DVSS.n268 DVSS.n257 292.5
R14674 DVSS.n267 DVSS.n266 292.5
R14675 DVSS.n265 DVSS.n264 292.5
R14676 DVSS.n263 DVSS.n262 292.5
R14677 DVSS.n261 DVSS.n260 292.5
R14678 DVSS.n259 DVSS.n258 292.5
R14679 DVSS.n253 DVSS.n252 292.5
R14680 DVSS.n301 DVSS.n186 292.5
R14681 DVSS.n301 DVSS.n300 292.5
R14682 DVSS.n291 DVSS.n187 292.5
R14683 DVSS.n192 DVSS.n187 292.5
R14684 DVSS.n279 DVSS.n278 292.5
R14685 DVSS.n280 DVSS.n279 292.5
R14686 DVSS.n277 DVSS.n197 292.5
R14687 DVSS.n198 DVSS.n197 292.5
R14688 DVSS.n293 DVSS.n292 292.5
R14689 DVSS.n294 DVSS.n293 292.5
R14690 DVSS.n275 DVSS.n274 292.5
R14691 DVSS.n276 DVSS.n251 292.5
R14692 DVSS.n251 DVSS.n250 292.5
R14693 DVSS.n314 DVSS.n304 292.5
R14694 DVSS.n307 DVSS.n304 292.5
R14695 DVSS.n315 DVSS.n184 292.5
R14696 DVSS.n306 DVSS.n184 292.5
R14697 DVSS.n313 DVSS.n312 292.5
R14698 DVSS.n310 DVSS.n305 292.5
R14699 DVSS.n321 DVSS.n320 292.5
R14700 DVSS.n323 DVSS.n322 292.5
R14701 DVSS.n185 DVSS.n166 292.5
R14702 DVSS.n340 DVSS.n166 292.5
R14703 DVSS.n318 DVSS.n317 292.5
R14704 DVSS.n309 DVSS.n307 292.5
R14705 DVSS.n306 DVSS.n183 292.5
R14706 DVSS.n181 DVSS.n180 292.5
R14707 DVSS.n329 DVSS.n328 292.5
R14708 DVSS.n332 DVSS.n331 292.5
R14709 DVSS.n175 DVSS.n174 292.5
R14710 DVSS.n338 DVSS.n337 292.5
R14711 DVSS.n172 DVSS.n163 292.5
R14712 DVSS.n343 DVSS.n342 292.5
R14713 DVSS.n162 DVSS.n160 292.5
R14714 DVSS.n164 DVSS.n162 292.5
R14715 DVSS.n299 DVSS.n298 292.5
R14716 DVSS.n300 DVSS.n299 292.5
R14717 DVSS.n297 DVSS.n188 292.5
R14718 DVSS.n192 DVSS.n188 292.5
R14719 DVSS.n296 DVSS.n295 292.5
R14720 DVSS.n295 DVSS.n294 292.5
R14721 DVSS.n249 DVSS.n248 292.5
R14722 DVSS.n250 DVSS.n249 292.5
R14723 DVSS.n282 DVSS.n281 292.5
R14724 DVSS.n281 DVSS.n280 292.5
R14725 DVSS.n283 DVSS.n200 292.5
R14726 DVSS.n200 DVSS.n198 292.5
R14727 DVSS.n285 DVSS.n284 292.5
R14728 DVSS.n286 DVSS.n285 292.5
R14729 DVSS.n289 DVSS.n193 292.5
R14730 DVSS.n247 DVSS.n246 292.5
R14731 DVSS.n246 DVSS.n190 292.5
R14732 DVSS.n205 DVSS.n203 292.5
R14733 DVSS.n210 DVSS.n203 292.5
R14734 DVSS.n241 DVSS.n207 292.5
R14735 DVSS.n241 DVSS.n240 292.5
R14736 DVSS.n215 DVSS.n212 292.5
R14737 DVSS.n239 DVSS.n212 292.5
R14738 DVSS.n236 DVSS.n217 292.5
R14739 DVSS.n237 DVSS.n236 292.5
R14740 DVSS.n222 DVSS.n218 292.5
R14741 DVSS.n218 DVSS.n213 292.5
R14742 DVSS.n231 DVSS.n224 292.5
R14743 DVSS.n231 DVSS.n230 292.5
R14744 DVSS.n229 DVSS.n227 292.5
R14745 DVSS.n227 DVSS.n226 292.5
R14746 DVSS.n289 DVSS.n288 292.5
R14747 DVSS.n101 DVSS.n100 292.5
R14748 DVSS.n92 DVSS.n91 292.5
R14749 DVSS.n104 DVSS.n103 292.5
R14750 DVSS.n106 DVSS.n105 292.5
R14751 DVSS.n108 DVSS.n107 292.5
R14752 DVSS.n110 DVSS.n109 292.5
R14753 DVSS.n112 DVSS.n111 292.5
R14754 DVSS.n102 DVSS.n99 292.5
R14755 DVSS.n116 DVSS.n115 292.5
R14756 DVSS.n115 DVSS.n114 292.5
R14757 DVSS.n408 DVSS.n28 292.5
R14758 DVSS.n408 DVSS.n33 292.5
R14759 DVSS.n421 DVSS.n404 292.5
R14760 DVSS.n420 DVSS.n419 292.5
R14761 DVSS.n418 DVSS.n417 292.5
R14762 DVSS.n416 DVSS.n406 292.5
R14763 DVSS.n414 DVSS.n413 292.5
R14764 DVSS.n412 DVSS.n407 292.5
R14765 DVSS.n411 DVSS.n410 292.5
R14766 DVSS.n424 DVSS.n423 292.5
R14767 DVSS.n64 DVSS.n60 292.5
R14768 DVSS.n77 DVSS.n56 292.5
R14769 DVSS.n75 DVSS.n74 292.5
R14770 DVSS.n73 DVSS.n72 292.5
R14771 DVSS.n70 DVSS.n58 292.5
R14772 DVSS.n68 DVSS.n67 292.5
R14773 DVSS.n66 DVSS.n65 292.5
R14774 DVSS.n79 DVSS.n78 292.5
R14775 DVSS.n78 DVSS.n49 292.5
R14776 DVSS.n62 DVSS.n61 292.5
R14777 DVSS.n458 DVSS.n457 292.5
R14778 DVSS.n457 DVSS.n18 292.5
R14779 DVSS.n459 DVSS.n27 292.5
R14780 DVSS.n27 DVSS.n26 292.5
R14781 DVSS.n461 DVSS.n460 292.5
R14782 DVSS.n462 DVSS.n461 292.5
R14783 DVSS.n436 DVSS.n25 292.5
R14784 DVSS.n25 DVSS.n24 292.5
R14785 DVSS.n434 DVSS.n433 292.5
R14786 DVSS.n433 DVSS.n432 292.5
R14787 DVSS.n30 DVSS.n29 292.5
R14788 DVSS.n32 DVSS.n30 292.5
R14789 DVSS.n388 DVSS.n46 292.5
R14790 DVSS.n46 DVSS.n44 292.5
R14791 DVSS.n390 DVSS.n389 292.5
R14792 DVSS.n391 DVSS.n390 292.5
R14793 DVSS.n387 DVSS.n45 292.5
R14794 DVSS.n50 DVSS.n45 292.5
R14795 DVSS.n386 DVSS.n385 292.5
R14796 DVSS.n385 DVSS.n384 292.5
R14797 DVSS.n369 DVSS.n368 292.5
R14798 DVSS.n370 DVSS.n369 292.5
R14799 DVSS.n367 DVSS.n83 292.5
R14800 DVSS.n83 DVSS.n82 292.5
R14801 DVSS.n366 DVSS.n365 292.5
R14802 DVSS.n365 DVSS.n364 292.5
R14803 DVSS.n85 DVSS.n84 292.5
R14804 DVSS.n86 DVSS.n85 292.5
R14805 DVSS.n456 DVSS.n437 292.5
R14806 DVSS.n442 DVSS.n438 292.5
R14807 DVSS.n452 DVSS.n451 292.5
R14808 DVSS.n450 DVSS.n441 292.5
R14809 DVSS.n449 DVSS.n448 292.5
R14810 DVSS.n447 DVSS.n446 292.5
R14811 DVSS.n445 DVSS.n444 292.5
R14812 DVSS.n443 DVSS.n15 292.5
R14813 DVSS.n473 DVSS.n472 292.5
R14814 DVSS.n2191 DVSS.n1871 270.034
R14815 DVSS.n1851 DVSS.n1845 270.034
R14816 DVSS.n1855 DVSS.n1843 270.034
R14817 DVSS.n2189 DVSS.n1868 270.034
R14818 DVSS.n1573 DVSS.n1253 270.034
R14819 DVSS.n1233 DVSS.n1227 270.034
R14820 DVSS.n1237 DVSS.n1225 270.034
R14821 DVSS.n1571 DVSS.n1250 270.034
R14822 DVSS.n960 DVSS.n640 270.034
R14823 DVSS.n620 DVSS.n614 270.034
R14824 DVSS.n624 DVSS.n612 270.034
R14825 DVSS.n958 DVSS.n637 270.034
R14826 DVSS.n371 DVSS.n51 270.034
R14827 DVSS.n31 DVSS.n25 270.034
R14828 DVSS.n35 DVSS.n23 270.034
R14829 DVSS.n369 DVSS.n48 270.034
R14830 DVSS.n2757 DVSS.n559 267.663
R14831 DVSS.n2519 DVSS.n2518 267.094
R14832 DVSS.n3063 DVSS.t36 265.887
R14833 DVSS.n1814 DVSS.n1813 261.063
R14834 DVSS.n572 DVSS.n571 261.063
R14835 DVSS.n3059 DVSS.t34 248.733
R14836 DVSS.n1877 DVSS.n1869 248.683
R14837 DVSS.n1891 DVSS.n1869 248.683
R14838 DVSS.n1889 DVSS.n1869 248.683
R14839 DVSS.n1259 DVSS.n1251 248.683
R14840 DVSS.n1273 DVSS.n1251 248.683
R14841 DVSS.n1271 DVSS.n1251 248.683
R14842 DVSS.n646 DVSS.n638 248.683
R14843 DVSS.n660 DVSS.n638 248.683
R14844 DVSS.n658 DVSS.n638 248.683
R14845 DVSS.n57 DVSS.n49 248.683
R14846 DVSS.n71 DVSS.n49 248.683
R14847 DVSS.n69 DVSS.n49 248.683
R14848 DVSS.n2160 DVSS.n1988 245.512
R14849 DVSS.n2160 DVSS.n1989 245.512
R14850 DVSS.n2160 DVSS.n1990 245.512
R14851 DVSS.n2160 DVSS.n1991 245.512
R14852 DVSS.n2160 DVSS.n2159 245.512
R14853 DVSS.n1934 DVSS.n1915 245.512
R14854 DVSS.n1934 DVSS.n1916 245.512
R14855 DVSS.n1934 DVSS.n1917 245.512
R14856 DVSS.n1934 DVSS.n1918 245.512
R14857 DVSS.n1934 DVSS.n1933 245.512
R14858 DVSS.n1542 DVSS.n1370 245.512
R14859 DVSS.n1542 DVSS.n1371 245.512
R14860 DVSS.n1542 DVSS.n1372 245.512
R14861 DVSS.n1542 DVSS.n1373 245.512
R14862 DVSS.n1542 DVSS.n1541 245.512
R14863 DVSS.n1316 DVSS.n1297 245.512
R14864 DVSS.n1316 DVSS.n1298 245.512
R14865 DVSS.n1316 DVSS.n1299 245.512
R14866 DVSS.n1316 DVSS.n1300 245.512
R14867 DVSS.n1316 DVSS.n1315 245.512
R14868 DVSS.n929 DVSS.n757 245.512
R14869 DVSS.n929 DVSS.n758 245.512
R14870 DVSS.n929 DVSS.n759 245.512
R14871 DVSS.n929 DVSS.n760 245.512
R14872 DVSS.n929 DVSS.n928 245.512
R14873 DVSS.n703 DVSS.n684 245.512
R14874 DVSS.n703 DVSS.n685 245.512
R14875 DVSS.n703 DVSS.n686 245.512
R14876 DVSS.n703 DVSS.n687 245.512
R14877 DVSS.n703 DVSS.n702 245.512
R14878 DVSS.n340 DVSS.n168 245.512
R14879 DVSS.n340 DVSS.n169 245.512
R14880 DVSS.n340 DVSS.n170 245.512
R14881 DVSS.n340 DVSS.n171 245.512
R14882 DVSS.n340 DVSS.n339 245.512
R14883 DVSS.n114 DVSS.n95 245.512
R14884 DVSS.n114 DVSS.n96 245.512
R14885 DVSS.n114 DVSS.n97 245.512
R14886 DVSS.n114 DVSS.n98 245.512
R14887 DVSS.n114 DVSS.n113 245.512
R14888 DVSS.n1818 DVSS.t123 233.869
R14889 DVSS.n576 DVSS.t23 233.869
R14890 DVSS.n2060 DVSS.n2059 223.931
R14891 DVSS.n2057 DVSS.n2033 223.931
R14892 DVSS.n2050 DVSS.n2049 223.931
R14893 DVSS.n2115 DVSS.n2008 223.931
R14894 DVSS.n2119 DVSS.n2008 223.931
R14895 DVSS.n2119 DVSS.n1982 223.931
R14896 DVSS.n2142 DVSS.n1986 223.931
R14897 DVSS.n2113 DVSS.n2007 223.931
R14898 DVSS.n2121 DVSS.n2007 223.931
R14899 DVSS.n2122 DVSS.n2121 223.931
R14900 DVSS.n2086 DVSS.n2085 223.931
R14901 DVSS.n2082 DVSS.n2081 223.931
R14902 DVSS.n2078 DVSS.n2073 223.931
R14903 DVSS.n2101 DVSS.n2069 223.931
R14904 DVSS.n2101 DVSS.n2020 223.931
R14905 DVSS.n2105 DVSS.n2020 223.931
R14906 DVSS.n2035 DVSS.n2027 223.931
R14907 DVSS.n2042 DVSS.n2037 223.931
R14908 DVSS.n2046 DVSS.n2044 223.931
R14909 DVSS.n2099 DVSS.n2071 223.931
R14910 DVSS.n2099 DVSS.n2017 223.931
R14911 DVSS.n2107 DVSS.n2017 223.931
R14912 DVSS.n2183 DVSS.n1907 223.931
R14913 DVSS.n2183 DVSS.n1901 223.931
R14914 DVSS.n2191 DVSS.n1901 223.931
R14915 DVSS.n1935 DVSS.n1912 223.931
R14916 DVSS.n2281 DVSS.n1845 223.931
R14917 DVSS.n2281 DVSS.n1847 223.931
R14918 DVSS.n2277 DVSS.n1847 223.931
R14919 DVSS.n2272 DVSS.n2261 223.931
R14920 DVSS.n2268 DVSS.n2267 223.931
R14921 DVSS.n2264 DVSS.n2263 223.931
R14922 DVSS.n2283 DVSS.n1843 223.931
R14923 DVSS.n2283 DVSS.n1837 223.931
R14924 DVSS.n2291 DVSS.n1837 223.931
R14925 DVSS.n2203 DVSS.n1862 223.931
R14926 DVSS.n2212 DVSS.n1862 223.931
R14927 DVSS.n2212 DVSS.n1863 223.931
R14928 DVSS.n1863 DVSS.n1854 223.931
R14929 DVSS.n2251 DVSS.n1854 223.931
R14930 DVSS.n2205 DVSS.n1865 223.931
R14931 DVSS.n2210 DVSS.n1865 223.931
R14932 DVSS.n2210 DVSS.n1866 223.931
R14933 DVSS.n1866 DVSS.n1850 223.931
R14934 DVSS.n2253 DVSS.n1850 223.931
R14935 DVSS.n2185 DVSS.n1905 223.931
R14936 DVSS.n2185 DVSS.n1903 223.931
R14937 DVSS.n2189 DVSS.n1903 223.931
R14938 DVSS.n1442 DVSS.n1441 223.931
R14939 DVSS.n1439 DVSS.n1415 223.931
R14940 DVSS.n1432 DVSS.n1431 223.931
R14941 DVSS.n1497 DVSS.n1390 223.931
R14942 DVSS.n1501 DVSS.n1390 223.931
R14943 DVSS.n1501 DVSS.n1364 223.931
R14944 DVSS.n1524 DVSS.n1368 223.931
R14945 DVSS.n1495 DVSS.n1389 223.931
R14946 DVSS.n1503 DVSS.n1389 223.931
R14947 DVSS.n1504 DVSS.n1503 223.931
R14948 DVSS.n1468 DVSS.n1467 223.931
R14949 DVSS.n1464 DVSS.n1463 223.931
R14950 DVSS.n1460 DVSS.n1455 223.931
R14951 DVSS.n1483 DVSS.n1451 223.931
R14952 DVSS.n1483 DVSS.n1402 223.931
R14953 DVSS.n1487 DVSS.n1402 223.931
R14954 DVSS.n1417 DVSS.n1409 223.931
R14955 DVSS.n1424 DVSS.n1419 223.931
R14956 DVSS.n1428 DVSS.n1426 223.931
R14957 DVSS.n1481 DVSS.n1453 223.931
R14958 DVSS.n1481 DVSS.n1399 223.931
R14959 DVSS.n1489 DVSS.n1399 223.931
R14960 DVSS.n1565 DVSS.n1289 223.931
R14961 DVSS.n1565 DVSS.n1283 223.931
R14962 DVSS.n1573 DVSS.n1283 223.931
R14963 DVSS.n1317 DVSS.n1294 223.931
R14964 DVSS.n1663 DVSS.n1227 223.931
R14965 DVSS.n1663 DVSS.n1229 223.931
R14966 DVSS.n1659 DVSS.n1229 223.931
R14967 DVSS.n1654 DVSS.n1643 223.931
R14968 DVSS.n1650 DVSS.n1649 223.931
R14969 DVSS.n1646 DVSS.n1645 223.931
R14970 DVSS.n1665 DVSS.n1225 223.931
R14971 DVSS.n1665 DVSS.n1219 223.931
R14972 DVSS.n1673 DVSS.n1219 223.931
R14973 DVSS.n1585 DVSS.n1244 223.931
R14974 DVSS.n1594 DVSS.n1244 223.931
R14975 DVSS.n1594 DVSS.n1245 223.931
R14976 DVSS.n1245 DVSS.n1236 223.931
R14977 DVSS.n1633 DVSS.n1236 223.931
R14978 DVSS.n1587 DVSS.n1247 223.931
R14979 DVSS.n1592 DVSS.n1247 223.931
R14980 DVSS.n1592 DVSS.n1248 223.931
R14981 DVSS.n1248 DVSS.n1232 223.931
R14982 DVSS.n1635 DVSS.n1232 223.931
R14983 DVSS.n1567 DVSS.n1287 223.931
R14984 DVSS.n1567 DVSS.n1285 223.931
R14985 DVSS.n1571 DVSS.n1285 223.931
R14986 DVSS.n829 DVSS.n828 223.931
R14987 DVSS.n826 DVSS.n802 223.931
R14988 DVSS.n819 DVSS.n818 223.931
R14989 DVSS.n884 DVSS.n777 223.931
R14990 DVSS.n888 DVSS.n777 223.931
R14991 DVSS.n888 DVSS.n751 223.931
R14992 DVSS.n911 DVSS.n755 223.931
R14993 DVSS.n882 DVSS.n776 223.931
R14994 DVSS.n890 DVSS.n776 223.931
R14995 DVSS.n891 DVSS.n890 223.931
R14996 DVSS.n855 DVSS.n854 223.931
R14997 DVSS.n851 DVSS.n850 223.931
R14998 DVSS.n847 DVSS.n842 223.931
R14999 DVSS.n870 DVSS.n838 223.931
R15000 DVSS.n870 DVSS.n789 223.931
R15001 DVSS.n874 DVSS.n789 223.931
R15002 DVSS.n804 DVSS.n796 223.931
R15003 DVSS.n811 DVSS.n806 223.931
R15004 DVSS.n815 DVSS.n813 223.931
R15005 DVSS.n868 DVSS.n840 223.931
R15006 DVSS.n868 DVSS.n786 223.931
R15007 DVSS.n876 DVSS.n786 223.931
R15008 DVSS.n952 DVSS.n676 223.931
R15009 DVSS.n952 DVSS.n670 223.931
R15010 DVSS.n960 DVSS.n670 223.931
R15011 DVSS.n704 DVSS.n681 223.931
R15012 DVSS.n1050 DVSS.n614 223.931
R15013 DVSS.n1050 DVSS.n616 223.931
R15014 DVSS.n1046 DVSS.n616 223.931
R15015 DVSS.n1041 DVSS.n1030 223.931
R15016 DVSS.n1037 DVSS.n1036 223.931
R15017 DVSS.n1033 DVSS.n1032 223.931
R15018 DVSS.n1052 DVSS.n612 223.931
R15019 DVSS.n1052 DVSS.n606 223.931
R15020 DVSS.n1060 DVSS.n606 223.931
R15021 DVSS.n972 DVSS.n631 223.931
R15022 DVSS.n981 DVSS.n631 223.931
R15023 DVSS.n981 DVSS.n632 223.931
R15024 DVSS.n632 DVSS.n623 223.931
R15025 DVSS.n1020 DVSS.n623 223.931
R15026 DVSS.n974 DVSS.n634 223.931
R15027 DVSS.n979 DVSS.n634 223.931
R15028 DVSS.n979 DVSS.n635 223.931
R15029 DVSS.n635 DVSS.n619 223.931
R15030 DVSS.n1022 DVSS.n619 223.931
R15031 DVSS.n954 DVSS.n674 223.931
R15032 DVSS.n954 DVSS.n672 223.931
R15033 DVSS.n958 DVSS.n672 223.931
R15034 DVSS.n240 DVSS.n239 223.931
R15035 DVSS.n237 DVSS.n213 223.931
R15036 DVSS.n230 DVSS.n229 223.931
R15037 DVSS.n295 DVSS.n188 223.931
R15038 DVSS.n299 DVSS.n188 223.931
R15039 DVSS.n299 DVSS.n162 223.931
R15040 DVSS.n322 DVSS.n166 223.931
R15041 DVSS.n293 DVSS.n187 223.931
R15042 DVSS.n301 DVSS.n187 223.931
R15043 DVSS.n302 DVSS.n301 223.931
R15044 DVSS.n266 DVSS.n265 223.931
R15045 DVSS.n262 DVSS.n261 223.931
R15046 DVSS.n258 DVSS.n253 223.931
R15047 DVSS.n281 DVSS.n249 223.931
R15048 DVSS.n281 DVSS.n200 223.931
R15049 DVSS.n285 DVSS.n200 223.931
R15050 DVSS.n215 DVSS.n207 223.931
R15051 DVSS.n222 DVSS.n217 223.931
R15052 DVSS.n226 DVSS.n224 223.931
R15053 DVSS.n279 DVSS.n251 223.931
R15054 DVSS.n279 DVSS.n197 223.931
R15055 DVSS.n287 DVSS.n197 223.931
R15056 DVSS.n363 DVSS.n87 223.931
R15057 DVSS.n363 DVSS.n81 223.931
R15058 DVSS.n371 DVSS.n81 223.931
R15059 DVSS.n115 DVSS.n92 223.931
R15060 DVSS.n461 DVSS.n25 223.931
R15061 DVSS.n461 DVSS.n27 223.931
R15062 DVSS.n457 DVSS.n27 223.931
R15063 DVSS.n452 DVSS.n441 223.931
R15064 DVSS.n448 DVSS.n447 223.931
R15065 DVSS.n444 DVSS.n443 223.931
R15066 DVSS.n463 DVSS.n23 223.931
R15067 DVSS.n463 DVSS.n17 223.931
R15068 DVSS.n471 DVSS.n17 223.931
R15069 DVSS.n383 DVSS.n42 223.931
R15070 DVSS.n392 DVSS.n42 223.931
R15071 DVSS.n392 DVSS.n43 223.931
R15072 DVSS.n43 DVSS.n34 223.931
R15073 DVSS.n431 DVSS.n34 223.931
R15074 DVSS.n385 DVSS.n45 223.931
R15075 DVSS.n390 DVSS.n45 223.931
R15076 DVSS.n390 DVSS.n46 223.931
R15077 DVSS.n46 DVSS.n30 223.931
R15078 DVSS.n433 DVSS.n30 223.931
R15079 DVSS.n365 DVSS.n85 223.931
R15080 DVSS.n365 DVSS.n83 223.931
R15081 DVSS.n369 DVSS.n83 223.931
R15082 DVSS.n2763 DVSS.t148 219.49
R15083 DVSS.n2526 DVSS.t75 218.476
R15084 DVSS.n2362 DVSS.t112 212.382
R15085 DVSS.n2931 DVSS.t135 212.382
R15086 DVSS.n1131 DVSS.t93 212.382
R15087 DVSS.n1744 DVSS.t166 212.382
R15088 DVSS.n2230 DVSS.n2228 206.16
R15089 DVSS.n2234 DVSS.n2227 206.16
R15090 DVSS.n2237 DVSS.n2236 206.16
R15091 DVSS.n2241 DVSS.n2240 206.16
R15092 DVSS.n1885 DVSS.n1884 206.16
R15093 DVSS.n1898 DVSS.n1897 206.16
R15094 DVSS.n1612 DVSS.n1610 206.16
R15095 DVSS.n1616 DVSS.n1609 206.16
R15096 DVSS.n1619 DVSS.n1618 206.16
R15097 DVSS.n1623 DVSS.n1622 206.16
R15098 DVSS.n1267 DVSS.n1266 206.16
R15099 DVSS.n1280 DVSS.n1279 206.16
R15100 DVSS.n999 DVSS.n997 206.16
R15101 DVSS.n1003 DVSS.n996 206.16
R15102 DVSS.n1006 DVSS.n1005 206.16
R15103 DVSS.n1010 DVSS.n1009 206.16
R15104 DVSS.n654 DVSS.n653 206.16
R15105 DVSS.n667 DVSS.n666 206.16
R15106 DVSS.n410 DVSS.n408 206.16
R15107 DVSS.n414 DVSS.n407 206.16
R15108 DVSS.n417 DVSS.n416 206.16
R15109 DVSS.n421 DVSS.n420 206.16
R15110 DVSS.n65 DVSS.n64 206.16
R15111 DVSS.n78 DVSS.n77 206.16
R15112 DVSS.n1763 DVSS.n1762 203.149
R15113 DVSS.n2341 DVSS.t116 201.764
R15114 DVSS.n2910 DVSS.t139 201.764
R15115 DVSS.n2211 DVSS.t58 199.196
R15116 DVSS.n1864 DVSS.t57 199.196
R15117 DVSS.n1593 DVSS.t147 199.196
R15118 DVSS.n1246 DVSS.t121 199.196
R15119 DVSS.n980 DVSS.t122 199.196
R15120 DVSS.n633 DVSS.t27 199.196
R15121 DVSS.n391 DVSS.t44 199.196
R15122 DVSS.n44 DVSS.t118 199.196
R15123 DVSS.n1974 DVSS.n1961 185
R15124 DVSS.n1976 DVSS.n1975 185
R15125 DVSS.n1953 DVSS.n1940 185
R15126 DVSS.n1955 DVSS.n1954 185
R15127 DVSS.n1356 DVSS.n1343 185
R15128 DVSS.n1358 DVSS.n1357 185
R15129 DVSS.n1335 DVSS.n1322 185
R15130 DVSS.n1337 DVSS.n1336 185
R15131 DVSS.n743 DVSS.n730 185
R15132 DVSS.n745 DVSS.n744 185
R15133 DVSS.n722 DVSS.n709 185
R15134 DVSS.n724 DVSS.n723 185
R15135 DVSS.n154 DVSS.n141 185
R15136 DVSS.n156 DVSS.n155 185
R15137 DVSS.n133 DVSS.n120 185
R15138 DVSS.n135 DVSS.n134 185
R15139 DVSS.n2846 DVSS.n2844 184.572
R15140 DVSS.n533 DVSS.n531 184.572
R15141 DVSS.n2849 DVSS.n2847 184.572
R15142 DVSS.n2378 DVSS.t110 170.724
R15143 DVSS.n2947 DVSS.t143 170.724
R15144 DVSS.n2666 DVSS.n2665 169.05
R15145 DVSS.n2100 DVSS.t79 158.811
R15146 DVSS.t79 DVSS.n2018 158.811
R15147 DVSS.n2012 DVSS.t83 158.811
R15148 DVSS.n2120 DVSS.t83 158.811
R15149 DVSS.t81 DVSS.n2126 158.811
R15150 DVSS.n2127 DVSS.t81 158.811
R15151 DVSS.n1482 DVSS.t15 158.811
R15152 DVSS.t15 DVSS.n1400 158.811
R15153 DVSS.n1394 DVSS.t188 158.811
R15154 DVSS.n1502 DVSS.t188 158.811
R15155 DVSS.t17 DVSS.n1508 158.811
R15156 DVSS.n1509 DVSS.t17 158.811
R15157 DVSS.n869 DVSS.t10 158.811
R15158 DVSS.t10 DVSS.n787 158.811
R15159 DVSS.n781 DVSS.t28 158.811
R15160 DVSS.n889 DVSS.t28 158.811
R15161 DVSS.t12 DVSS.n895 158.811
R15162 DVSS.n896 DVSS.t12 158.811
R15163 DVSS.n280 DVSS.t45 158.811
R15164 DVSS.t45 DVSS.n198 158.811
R15165 DVSS.n192 DVSS.t13 158.811
R15166 DVSS.n300 DVSS.t13 158.811
R15167 DVSS.t47 DVSS.n306 158.811
R15168 DVSS.n307 DVSS.t47 158.811
R15169 DVSS.n1879 DVSS.n1869 157.904
R15170 DVSS.n1261 DVSS.n1251 157.904
R15171 DVSS.n648 DVSS.n638 157.904
R15172 DVSS.n59 DVSS.n49 157.904
R15173 DVSS.n1896 DVSS.n1869 157.904
R15174 DVSS.n1278 DVSS.n1251 157.904
R15175 DVSS.n665 DVSS.n638 157.904
R15176 DVSS.n76 DVSS.n49 157.904
R15177 DVSS.n2161 DVSS.n2160 155.356
R15178 DVSS.n1543 DVSS.n1542 155.356
R15179 DVSS.n930 DVSS.n929 155.356
R15180 DVSS.n341 DVSS.n340 155.356
R15181 DVSS.n2092 DVSS.n2091 155.356
R15182 DVSS.n2092 DVSS.n2076 155.356
R15183 DVSS.n2160 DVSS.n1987 155.356
R15184 DVSS.n2021 DVSS.n2019 155.356
R15185 DVSS.n2029 DVSS.n2011 155.356
R15186 DVSS.n2026 DVSS.n2019 155.356
R15187 DVSS.n2031 DVSS.n2011 155.356
R15188 DVSS.n1934 DVSS.n1913 155.356
R15189 DVSS.n1934 DVSS.n1914 155.356
R15190 DVSS.n2275 DVSS.n2274 155.356
R15191 DVSS.n2274 DVSS.n2273 155.356
R15192 DVSS.n1474 DVSS.n1473 155.356
R15193 DVSS.n1474 DVSS.n1458 155.356
R15194 DVSS.n1542 DVSS.n1369 155.356
R15195 DVSS.n1403 DVSS.n1401 155.356
R15196 DVSS.n1411 DVSS.n1393 155.356
R15197 DVSS.n1408 DVSS.n1401 155.356
R15198 DVSS.n1413 DVSS.n1393 155.356
R15199 DVSS.n1316 DVSS.n1295 155.356
R15200 DVSS.n1316 DVSS.n1296 155.356
R15201 DVSS.n1657 DVSS.n1656 155.356
R15202 DVSS.n1656 DVSS.n1655 155.356
R15203 DVSS.n861 DVSS.n860 155.356
R15204 DVSS.n861 DVSS.n845 155.356
R15205 DVSS.n929 DVSS.n756 155.356
R15206 DVSS.n790 DVSS.n788 155.356
R15207 DVSS.n798 DVSS.n780 155.356
R15208 DVSS.n795 DVSS.n788 155.356
R15209 DVSS.n800 DVSS.n780 155.356
R15210 DVSS.n703 DVSS.n682 155.356
R15211 DVSS.n703 DVSS.n683 155.356
R15212 DVSS.n1044 DVSS.n1043 155.356
R15213 DVSS.n1043 DVSS.n1042 155.356
R15214 DVSS.n272 DVSS.n271 155.356
R15215 DVSS.n272 DVSS.n256 155.356
R15216 DVSS.n340 DVSS.n167 155.356
R15217 DVSS.n201 DVSS.n199 155.356
R15218 DVSS.n209 DVSS.n191 155.356
R15219 DVSS.n206 DVSS.n199 155.356
R15220 DVSS.n211 DVSS.n191 155.356
R15221 DVSS.n114 DVSS.n93 155.356
R15222 DVSS.n114 DVSS.n94 155.356
R15223 DVSS.n455 DVSS.n454 155.356
R15224 DVSS.n454 DVSS.n453 155.356
R15225 DVSS.n2184 DVSS.t0 150.504
R15226 DVSS.t0 DVSS.n1902 150.504
R15227 DVSS.n2282 DVSS.t56 150.504
R15228 DVSS.n1846 DVSS.t56 150.504
R15229 DVSS.n1566 DVSS.t105 150.504
R15230 DVSS.t105 DVSS.n1284 150.504
R15231 DVSS.n1664 DVSS.t82 150.504
R15232 DVSS.n1228 DVSS.t82 150.504
R15233 DVSS.n953 DVSS.t190 150.504
R15234 DVSS.t190 DVSS.n671 150.504
R15235 DVSS.n1051 DVSS.t18 150.504
R15236 DVSS.n615 DVSS.t18 150.504
R15237 DVSS.n364 DVSS.t130 150.504
R15238 DVSS.t130 DVSS.n82 150.504
R15239 DVSS.n462 DVSS.t129 150.504
R15240 DVSS.n26 DVSS.t129 150.504
R15241 DVSS.n2375 DVSS.n2374 131.416
R15242 DVSS.n2944 DVSS.n2943 131.416
R15243 DVSS.t116 DVSS.n2340 125.389
R15244 DVSS.t139 DVSS.n2909 125.389
R15245 DVSS.n1110 DVSS.t101 120.043
R15246 DVSS.n1723 DVSS.t172 120.043
R15247 DVSS.n1969 DVSS.t84 119.998
R15248 DVSS.n1948 DVSS.t80 119.998
R15249 DVSS.n1351 DVSS.t189 119.998
R15250 DVSS.n1330 DVSS.t16 119.998
R15251 DVSS.n738 DVSS.t29 119.998
R15252 DVSS.n717 DVSS.t11 119.998
R15253 DVSS.n149 DVSS.t14 119.998
R15254 DVSS.n128 DVSS.t46 119.998
R15255 DVSS.n2161 DVSS.n1983 118.938
R15256 DVSS.n1543 DVSS.n1365 118.938
R15257 DVSS.n930 DVSS.n752 118.938
R15258 DVSS.n341 DVSS.n163 118.938
R15259 DVSS.n2091 DVSS.n2077 118.936
R15260 DVSS.n2077 DVSS.n2076 118.936
R15261 DVSS.n2000 DVSS.n1987 118.936
R15262 DVSS.n2025 DVSS.n2021 118.936
R15263 DVSS.n2030 DVSS.n2029 118.936
R15264 DVSS.n2026 DVSS.n2025 118.936
R15265 DVSS.n2031 DVSS.n2030 118.936
R15266 DVSS.n1919 DVSS.n1913 118.936
R15267 DVSS.n1923 DVSS.n1914 118.936
R15268 DVSS.n2275 DVSS.n2258 118.936
R15269 DVSS.n2273 DVSS.n2258 118.936
R15270 DVSS.n1473 DVSS.n1459 118.936
R15271 DVSS.n1459 DVSS.n1458 118.936
R15272 DVSS.n1382 DVSS.n1369 118.936
R15273 DVSS.n1407 DVSS.n1403 118.936
R15274 DVSS.n1412 DVSS.n1411 118.936
R15275 DVSS.n1408 DVSS.n1407 118.936
R15276 DVSS.n1413 DVSS.n1412 118.936
R15277 DVSS.n1301 DVSS.n1295 118.936
R15278 DVSS.n1305 DVSS.n1296 118.936
R15279 DVSS.n1657 DVSS.n1640 118.936
R15280 DVSS.n1655 DVSS.n1640 118.936
R15281 DVSS.n860 DVSS.n846 118.936
R15282 DVSS.n846 DVSS.n845 118.936
R15283 DVSS.n769 DVSS.n756 118.936
R15284 DVSS.n794 DVSS.n790 118.936
R15285 DVSS.n799 DVSS.n798 118.936
R15286 DVSS.n795 DVSS.n794 118.936
R15287 DVSS.n800 DVSS.n799 118.936
R15288 DVSS.n688 DVSS.n682 118.936
R15289 DVSS.n692 DVSS.n683 118.936
R15290 DVSS.n1044 DVSS.n1027 118.936
R15291 DVSS.n1042 DVSS.n1027 118.936
R15292 DVSS.n271 DVSS.n257 118.936
R15293 DVSS.n257 DVSS.n256 118.936
R15294 DVSS.n180 DVSS.n167 118.936
R15295 DVSS.n205 DVSS.n201 118.936
R15296 DVSS.n210 DVSS.n209 118.936
R15297 DVSS.n206 DVSS.n205 118.936
R15298 DVSS.n211 DVSS.n210 118.936
R15299 DVSS.n99 DVSS.n93 118.936
R15300 DVSS.n103 DVSS.n94 118.936
R15301 DVSS.n455 DVSS.n438 118.936
R15302 DVSS.n453 DVSS.n438 118.936
R15303 DVSS.n2132 DVSS.n2131 117.719
R15304 DVSS.n2140 DVSS.n2139 117.719
R15305 DVSS.n2129 DVSS.n2128 117.719
R15306 DVSS.n1514 DVSS.n1513 117.719
R15307 DVSS.n1522 DVSS.n1521 117.719
R15308 DVSS.n1511 DVSS.n1510 117.719
R15309 DVSS.n901 DVSS.n900 117.719
R15310 DVSS.n909 DVSS.n908 117.719
R15311 DVSS.n898 DVSS.n897 117.719
R15312 DVSS.n312 DVSS.n311 117.719
R15313 DVSS.n320 DVSS.n319 117.719
R15314 DVSS.n309 DVSS.n308 117.719
R15315 DVSS.n2139 DVSS.n2138 117.719
R15316 DVSS.n2128 DVSS.n2003 117.719
R15317 DVSS.n1521 DVSS.n1520 117.719
R15318 DVSS.n1510 DVSS.n1385 117.719
R15319 DVSS.n908 DVSS.n907 117.719
R15320 DVSS.n897 DVSS.n772 117.719
R15321 DVSS.n319 DVSS.n318 117.719
R15322 DVSS.n308 DVSS.n183 117.719
R15323 DVSS.n2131 DVSS.n2130 117.719
R15324 DVSS.n1513 DVSS.n1512 117.719
R15325 DVSS.n900 DVSS.n899 117.719
R15326 DVSS.n311 DVSS.n310 117.719
R15327 DVSS.n2826 DVSS.t86 115.689
R15328 DVSS.n543 DVSS.t49 114.245
R15329 DVSS.n2776 DVSS.t31 114.245
R15330 DVSS.n566 DVSS.t22 114.245
R15331 DVSS.n1808 DVSS.t126 114.245
R15332 DVSS.n2659 DVSS.t53 114.245
R15333 DVSS.n2539 DVSS.t2 114.245
R15334 DVSS.n483 DVSS.t7 113.74
R15335 DVSS.n1977 DVSS.n1976 112.831
R15336 DVSS.n1956 DVSS.n1955 112.831
R15337 DVSS.n1359 DVSS.n1358 112.831
R15338 DVSS.n1338 DVSS.n1337 112.831
R15339 DVSS.n746 DVSS.n745 112.831
R15340 DVSS.n725 DVSS.n724 112.831
R15341 DVSS.n157 DVSS.n156 112.831
R15342 DVSS.n136 DVSS.n135 112.831
R15343 DVSS.n1888 DVSS.n1879 111.293
R15344 DVSS.n1270 DVSS.n1261 111.293
R15345 DVSS.n657 DVSS.n648 111.293
R15346 DVSS.n68 DVSS.n59 111.293
R15347 DVSS.n1896 DVSS.n1895 111.293
R15348 DVSS.n1278 DVSS.n1277 111.293
R15349 DVSS.n665 DVSS.n664 111.293
R15350 DVSS.n76 DVSS.n75 111.293
R15351 DVSS.n1775 DVSS.n1774 110.808
R15352 DVSS.n2675 DVSS.t42 110.353
R15353 DVSS.n2442 DVSS.t127 110.118
R15354 DVSS.n2561 DVSS.t119 108.9
R15355 DVSS.n1883 DVSS.n1869 108.141
R15356 DVSS.n1265 DVSS.n1251 108.141
R15357 DVSS.n652 DVSS.n638 108.141
R15358 DVSS.n63 DVSS.n49 108.141
R15359 DVSS.n2229 DVSS.n1853 108.141
R15360 DVSS.n2235 DVSS.n1853 108.141
R15361 DVSS.n2225 DVSS.n1853 108.141
R15362 DVSS.n2242 DVSS.n1853 108.141
R15363 DVSS.n1611 DVSS.n1235 108.141
R15364 DVSS.n1617 DVSS.n1235 108.141
R15365 DVSS.n1607 DVSS.n1235 108.141
R15366 DVSS.n1624 DVSS.n1235 108.141
R15367 DVSS.n998 DVSS.n622 108.141
R15368 DVSS.n1004 DVSS.n622 108.141
R15369 DVSS.n994 DVSS.n622 108.141
R15370 DVSS.n1011 DVSS.n622 108.141
R15371 DVSS.n409 DVSS.n33 108.141
R15372 DVSS.n415 DVSS.n33 108.141
R15373 DVSS.n405 DVSS.n33 108.141
R15374 DVSS.n422 DVSS.n33 108.141
R15375 DVSS.n501 DVSS.t175 108.037
R15376 DVSS.n2048 DVSS.n2011 105.766
R15377 DVSS.n1430 DVSS.n1393 105.766
R15378 DVSS.n817 DVSS.n780 105.766
R15379 DVSS.n228 DVSS.n191 105.766
R15380 DVSS.n2092 DVSS.n2075 105.766
R15381 DVSS.n2092 DVSS.n2074 105.766
R15382 DVSS.n2093 DVSS.n2092 105.766
R15383 DVSS.n2036 DVSS.n2019 105.766
R15384 DVSS.n2058 DVSS.n2011 105.766
R15385 DVSS.n2043 DVSS.n2019 105.766
R15386 DVSS.n2045 DVSS.n2011 105.766
R15387 DVSS.n2019 DVSS.n2016 105.766
R15388 DVSS.n2274 DVSS.n2260 105.766
R15389 DVSS.n2274 DVSS.n2259 105.766
R15390 DVSS.n2274 DVSS.n1836 105.766
R15391 DVSS.n1474 DVSS.n1457 105.766
R15392 DVSS.n1474 DVSS.n1456 105.766
R15393 DVSS.n1475 DVSS.n1474 105.766
R15394 DVSS.n1418 DVSS.n1401 105.766
R15395 DVSS.n1440 DVSS.n1393 105.766
R15396 DVSS.n1425 DVSS.n1401 105.766
R15397 DVSS.n1427 DVSS.n1393 105.766
R15398 DVSS.n1401 DVSS.n1398 105.766
R15399 DVSS.n1656 DVSS.n1642 105.766
R15400 DVSS.n1656 DVSS.n1641 105.766
R15401 DVSS.n1656 DVSS.n1218 105.766
R15402 DVSS.n861 DVSS.n844 105.766
R15403 DVSS.n861 DVSS.n843 105.766
R15404 DVSS.n862 DVSS.n861 105.766
R15405 DVSS.n805 DVSS.n788 105.766
R15406 DVSS.n827 DVSS.n780 105.766
R15407 DVSS.n812 DVSS.n788 105.766
R15408 DVSS.n814 DVSS.n780 105.766
R15409 DVSS.n788 DVSS.n785 105.766
R15410 DVSS.n1043 DVSS.n1029 105.766
R15411 DVSS.n1043 DVSS.n1028 105.766
R15412 DVSS.n1043 DVSS.n605 105.766
R15413 DVSS.n272 DVSS.n255 105.766
R15414 DVSS.n272 DVSS.n254 105.766
R15415 DVSS.n273 DVSS.n272 105.766
R15416 DVSS.n216 DVSS.n199 105.766
R15417 DVSS.n238 DVSS.n191 105.766
R15418 DVSS.n223 DVSS.n199 105.766
R15419 DVSS.n225 DVSS.n191 105.766
R15420 DVSS.n199 DVSS.n196 105.766
R15421 DVSS.n454 DVSS.n440 105.766
R15422 DVSS.n454 DVSS.n439 105.766
R15423 DVSS.n454 DVSS.n16 105.766
R15424 DVSS.n1972 DVSS.n1971 104.172
R15425 DVSS.n1951 DVSS.n1950 104.172
R15426 DVSS.n1354 DVSS.n1353 104.172
R15427 DVSS.n1333 DVSS.n1332 104.172
R15428 DVSS.n741 DVSS.n740 104.172
R15429 DVSS.n720 DVSS.n719 104.172
R15430 DVSS.n152 DVSS.n151 104.172
R15431 DVSS.n131 DVSS.n130 104.172
R15432 DVSS.n1870 DVSS.t58 101.811
R15433 DVSS.t57 DVSS.n1852 101.811
R15434 DVSS.n1252 DVSS.t147 101.811
R15435 DVSS.t121 DVSS.n1234 101.811
R15436 DVSS.n639 DVSS.t122 101.811
R15437 DVSS.t27 DVSS.n621 101.811
R15438 DVSS.n50 DVSS.t44 101.811
R15439 DVSS.t118 DVSS.n32 101.811
R15440 DVSS.n2467 DVSS.n2466 101.681
R15441 DVSS.n1150 DVSS.t95 101.575
R15442 DVSS.n1763 DVSS.t164 101.575
R15443 DVSS.n4 DVSS.t51 101.038
R15444 DVSS.n557 DVSS.t149 101.038
R15445 DVSS.n581 DVSS.t24 101.038
R15446 DVSS.n1823 DVSS.t124 101.038
R15447 DVSS.n1192 DVSS.t55 101.038
R15448 DVSS.n1202 DVSS.t76 101.038
R15449 DVSS.n2467 DVSS.t154 99.3708
R15450 DVSS.n2586 DVSS.t71 98.2867
R15451 DVSS.n2159 DVSS.n2158 93.9796
R15452 DVSS.n1994 DVSS.n1991 93.9796
R15453 DVSS.n2151 DVSS.n1990 93.9796
R15454 DVSS.n2148 DVSS.n1989 93.9796
R15455 DVSS.n2000 DVSS.n1988 93.9796
R15456 DVSS.n2148 DVSS.n1988 93.9796
R15457 DVSS.n2151 DVSS.n1989 93.9796
R15458 DVSS.n1994 DVSS.n1990 93.9796
R15459 DVSS.n2158 DVSS.n1991 93.9796
R15460 DVSS.n2159 DVSS.n1983 93.9796
R15461 DVSS.n1933 DVSS.n1932 93.9796
R15462 DVSS.n1929 DVSS.n1918 93.9796
R15463 DVSS.n1927 DVSS.n1917 93.9796
R15464 DVSS.n1925 DVSS.n1916 93.9796
R15465 DVSS.n1923 DVSS.n1915 93.9796
R15466 DVSS.n1932 DVSS.n1918 93.9796
R15467 DVSS.n1929 DVSS.n1917 93.9796
R15468 DVSS.n1927 DVSS.n1916 93.9796
R15469 DVSS.n1925 DVSS.n1915 93.9796
R15470 DVSS.n1933 DVSS.n1919 93.9796
R15471 DVSS.n1541 DVSS.n1540 93.9796
R15472 DVSS.n1376 DVSS.n1373 93.9796
R15473 DVSS.n1533 DVSS.n1372 93.9796
R15474 DVSS.n1530 DVSS.n1371 93.9796
R15475 DVSS.n1382 DVSS.n1370 93.9796
R15476 DVSS.n1530 DVSS.n1370 93.9796
R15477 DVSS.n1533 DVSS.n1371 93.9796
R15478 DVSS.n1376 DVSS.n1372 93.9796
R15479 DVSS.n1540 DVSS.n1373 93.9796
R15480 DVSS.n1541 DVSS.n1365 93.9796
R15481 DVSS.n1315 DVSS.n1314 93.9796
R15482 DVSS.n1311 DVSS.n1300 93.9796
R15483 DVSS.n1309 DVSS.n1299 93.9796
R15484 DVSS.n1307 DVSS.n1298 93.9796
R15485 DVSS.n1305 DVSS.n1297 93.9796
R15486 DVSS.n1314 DVSS.n1300 93.9796
R15487 DVSS.n1311 DVSS.n1299 93.9796
R15488 DVSS.n1309 DVSS.n1298 93.9796
R15489 DVSS.n1307 DVSS.n1297 93.9796
R15490 DVSS.n1315 DVSS.n1301 93.9796
R15491 DVSS.n928 DVSS.n927 93.9796
R15492 DVSS.n763 DVSS.n760 93.9796
R15493 DVSS.n920 DVSS.n759 93.9796
R15494 DVSS.n917 DVSS.n758 93.9796
R15495 DVSS.n769 DVSS.n757 93.9796
R15496 DVSS.n917 DVSS.n757 93.9796
R15497 DVSS.n920 DVSS.n758 93.9796
R15498 DVSS.n763 DVSS.n759 93.9796
R15499 DVSS.n927 DVSS.n760 93.9796
R15500 DVSS.n928 DVSS.n752 93.9796
R15501 DVSS.n702 DVSS.n701 93.9796
R15502 DVSS.n698 DVSS.n687 93.9796
R15503 DVSS.n696 DVSS.n686 93.9796
R15504 DVSS.n694 DVSS.n685 93.9796
R15505 DVSS.n692 DVSS.n684 93.9796
R15506 DVSS.n701 DVSS.n687 93.9796
R15507 DVSS.n698 DVSS.n686 93.9796
R15508 DVSS.n696 DVSS.n685 93.9796
R15509 DVSS.n694 DVSS.n684 93.9796
R15510 DVSS.n702 DVSS.n688 93.9796
R15511 DVSS.n339 DVSS.n338 93.9796
R15512 DVSS.n174 DVSS.n171 93.9796
R15513 DVSS.n331 DVSS.n170 93.9796
R15514 DVSS.n328 DVSS.n169 93.9796
R15515 DVSS.n180 DVSS.n168 93.9796
R15516 DVSS.n328 DVSS.n168 93.9796
R15517 DVSS.n331 DVSS.n169 93.9796
R15518 DVSS.n174 DVSS.n170 93.9796
R15519 DVSS.n338 DVSS.n171 93.9796
R15520 DVSS.n339 DVSS.n163 93.9796
R15521 DVSS.n113 DVSS.n112 93.9796
R15522 DVSS.n109 DVSS.n98 93.9796
R15523 DVSS.n107 DVSS.n97 93.9796
R15524 DVSS.n105 DVSS.n96 93.9796
R15525 DVSS.n103 DVSS.n95 93.9796
R15526 DVSS.n112 DVSS.n98 93.9796
R15527 DVSS.n109 DVSS.n97 93.9796
R15528 DVSS.n107 DVSS.n96 93.9796
R15529 DVSS.n105 DVSS.n95 93.9796
R15530 DVSS.n113 DVSS.n99 93.9796
R15531 DVSS.n1971 DVSS.n1970 92.5005
R15532 DVSS.n1950 DVSS.n1949 92.5005
R15533 DVSS.n1353 DVSS.n1352 92.5005
R15534 DVSS.n1332 DVSS.n1331 92.5005
R15535 DVSS.n740 DVSS.n739 92.5005
R15536 DVSS.n719 DVSS.n718 92.5005
R15537 DVSS.n151 DVSS.n150 92.5005
R15538 DVSS.n130 DVSS.n129 92.5005
R15539 DVSS.n1150 DVSS.n1149 92.3405
R15540 DVSS.n484 DVSS.t4 91.1965
R15541 DVSS.n483 DVSS.t9 91.1965
R15542 DVSS.n2704 DVSS.t177 90.704
R15543 DVSS.n3040 DVSS.t33 90.704
R15544 DVSS.n2590 DVSS.t72 90.704
R15545 DVSS.n1828 DVSS.t155 90.704
R15546 DVSS.n1767 DVSS.t165 90.703
R15547 DVSS.n2382 DVSS.t111 90.703
R15548 DVSS.n1154 DVSS.t96 90.703
R15549 DVSS.n2951 DVSS.t144 90.703
R15550 DVSS.n1890 DVSS.n1889 87.6383
R15551 DVSS.n1892 DVSS.n1891 87.6383
R15552 DVSS.n1895 DVSS.n1877 87.6383
R15553 DVSS.n1889 DVSS.n1888 87.6383
R15554 DVSS.n1891 DVSS.n1890 87.6383
R15555 DVSS.n1892 DVSS.n1877 87.6383
R15556 DVSS.n1272 DVSS.n1271 87.6383
R15557 DVSS.n1274 DVSS.n1273 87.6383
R15558 DVSS.n1277 DVSS.n1259 87.6383
R15559 DVSS.n1271 DVSS.n1270 87.6383
R15560 DVSS.n1273 DVSS.n1272 87.6383
R15561 DVSS.n1274 DVSS.n1259 87.6383
R15562 DVSS.n659 DVSS.n658 87.6383
R15563 DVSS.n661 DVSS.n660 87.6383
R15564 DVSS.n664 DVSS.n646 87.6383
R15565 DVSS.n658 DVSS.n657 87.6383
R15566 DVSS.n660 DVSS.n659 87.6383
R15567 DVSS.n661 DVSS.n646 87.6383
R15568 DVSS.n70 DVSS.n69 87.6383
R15569 DVSS.n72 DVSS.n71 87.6383
R15570 DVSS.n75 DVSS.n57 87.6383
R15571 DVSS.n69 DVSS.n68 87.6383
R15572 DVSS.n71 DVSS.n70 87.6383
R15573 DVSS.n72 DVSS.n57 87.6383
R15574 DVSS.n2139 DVSS.n1985 87.3927
R15575 DVSS.n2128 DVSS.n1998 87.3927
R15576 DVSS.n1521 DVSS.n1367 87.3927
R15577 DVSS.n1510 DVSS.n1380 87.3927
R15578 DVSS.n908 DVSS.n754 87.3927
R15579 DVSS.n897 DVSS.n767 87.3927
R15580 DVSS.n319 DVSS.n165 87.3927
R15581 DVSS.n308 DVSS.n178 87.3927
R15582 DVSS.n2681 DVSS.t103 86.8735
R15583 DVSS.n2448 DVSS.t114 86.6885
R15584 DVSS.n2567 DVSS.t162 85.7298
R15585 DVSS.n2300 DVSS.t150 85.3621
R15586 DVSS.n1680 DVSS.t61 85.3621
R15587 DVSS.n1067 DVSS.t19 85.3621
R15588 DVSS.n478 DVSS.t77 85.3621
R15589 DVSS.t87 DVSS.t59 82.3134
R15590 DVSS.n2699 DVSS.t176 81.0531
R15591 DVSS.n2048 DVSS.n2013 80.9725
R15592 DVSS.n1430 DVSS.n1395 80.9725
R15593 DVSS.n817 DVSS.n782 80.9725
R15594 DVSS.n228 DVSS.n193 80.9725
R15595 DVSS.n2049 DVSS.n2048 80.9721
R15596 DVSS.n1431 DVSS.n1430 80.9721
R15597 DVSS.n818 DVSS.n817 80.9721
R15598 DVSS.n229 DVSS.n228 80.9721
R15599 DVSS.n2058 DVSS.n2057 80.9719
R15600 DVSS.n2050 DVSS.n2045 80.9719
R15601 DVSS.n2082 DVSS.n2075 80.9719
R15602 DVSS.n2078 DVSS.n2074 80.9719
R15603 DVSS.n2094 DVSS.n2093 80.9719
R15604 DVSS.n2037 DVSS.n2036 80.9719
R15605 DVSS.n2044 DVSS.n2043 80.9719
R15606 DVSS.n2108 DVSS.n2016 80.9719
R15607 DVSS.n2085 DVSS.n2075 80.9719
R15608 DVSS.n2081 DVSS.n2074 80.9719
R15609 DVSS.n2093 DVSS.n2073 80.9719
R15610 DVSS.n2036 DVSS.n2035 80.9719
R15611 DVSS.n2059 DVSS.n2058 80.9719
R15612 DVSS.n2043 DVSS.n2042 80.9719
R15613 DVSS.n2045 DVSS.n2033 80.9719
R15614 DVSS.n2046 DVSS.n2016 80.9719
R15615 DVSS.n2268 DVSS.n2260 80.9719
R15616 DVSS.n2264 DVSS.n2259 80.9719
R15617 DVSS.n2292 DVSS.n1836 80.9719
R15618 DVSS.n2261 DVSS.n2260 80.9719
R15619 DVSS.n2267 DVSS.n2259 80.9719
R15620 DVSS.n2263 DVSS.n1836 80.9719
R15621 DVSS.n1440 DVSS.n1439 80.9719
R15622 DVSS.n1432 DVSS.n1427 80.9719
R15623 DVSS.n1464 DVSS.n1457 80.9719
R15624 DVSS.n1460 DVSS.n1456 80.9719
R15625 DVSS.n1476 DVSS.n1475 80.9719
R15626 DVSS.n1419 DVSS.n1418 80.9719
R15627 DVSS.n1426 DVSS.n1425 80.9719
R15628 DVSS.n1490 DVSS.n1398 80.9719
R15629 DVSS.n1467 DVSS.n1457 80.9719
R15630 DVSS.n1463 DVSS.n1456 80.9719
R15631 DVSS.n1475 DVSS.n1455 80.9719
R15632 DVSS.n1418 DVSS.n1417 80.9719
R15633 DVSS.n1441 DVSS.n1440 80.9719
R15634 DVSS.n1425 DVSS.n1424 80.9719
R15635 DVSS.n1427 DVSS.n1415 80.9719
R15636 DVSS.n1428 DVSS.n1398 80.9719
R15637 DVSS.n1650 DVSS.n1642 80.9719
R15638 DVSS.n1646 DVSS.n1641 80.9719
R15639 DVSS.n1674 DVSS.n1218 80.9719
R15640 DVSS.n1643 DVSS.n1642 80.9719
R15641 DVSS.n1649 DVSS.n1641 80.9719
R15642 DVSS.n1645 DVSS.n1218 80.9719
R15643 DVSS.n827 DVSS.n826 80.9719
R15644 DVSS.n819 DVSS.n814 80.9719
R15645 DVSS.n851 DVSS.n844 80.9719
R15646 DVSS.n847 DVSS.n843 80.9719
R15647 DVSS.n863 DVSS.n862 80.9719
R15648 DVSS.n806 DVSS.n805 80.9719
R15649 DVSS.n813 DVSS.n812 80.9719
R15650 DVSS.n877 DVSS.n785 80.9719
R15651 DVSS.n854 DVSS.n844 80.9719
R15652 DVSS.n850 DVSS.n843 80.9719
R15653 DVSS.n862 DVSS.n842 80.9719
R15654 DVSS.n805 DVSS.n804 80.9719
R15655 DVSS.n828 DVSS.n827 80.9719
R15656 DVSS.n812 DVSS.n811 80.9719
R15657 DVSS.n814 DVSS.n802 80.9719
R15658 DVSS.n815 DVSS.n785 80.9719
R15659 DVSS.n1037 DVSS.n1029 80.9719
R15660 DVSS.n1033 DVSS.n1028 80.9719
R15661 DVSS.n1061 DVSS.n605 80.9719
R15662 DVSS.n1030 DVSS.n1029 80.9719
R15663 DVSS.n1036 DVSS.n1028 80.9719
R15664 DVSS.n1032 DVSS.n605 80.9719
R15665 DVSS.n238 DVSS.n237 80.9719
R15666 DVSS.n230 DVSS.n225 80.9719
R15667 DVSS.n262 DVSS.n255 80.9719
R15668 DVSS.n258 DVSS.n254 80.9719
R15669 DVSS.n274 DVSS.n273 80.9719
R15670 DVSS.n217 DVSS.n216 80.9719
R15671 DVSS.n224 DVSS.n223 80.9719
R15672 DVSS.n288 DVSS.n196 80.9719
R15673 DVSS.n265 DVSS.n255 80.9719
R15674 DVSS.n261 DVSS.n254 80.9719
R15675 DVSS.n273 DVSS.n253 80.9719
R15676 DVSS.n216 DVSS.n215 80.9719
R15677 DVSS.n239 DVSS.n238 80.9719
R15678 DVSS.n223 DVSS.n222 80.9719
R15679 DVSS.n225 DVSS.n213 80.9719
R15680 DVSS.n226 DVSS.n196 80.9719
R15681 DVSS.n448 DVSS.n440 80.9719
R15682 DVSS.n444 DVSS.n439 80.9719
R15683 DVSS.n472 DVSS.n16 80.9719
R15684 DVSS.n441 DVSS.n440 80.9719
R15685 DVSS.n447 DVSS.n439 80.9719
R15686 DVSS.n443 DVSS.n16 80.9719
R15687 DVSS.n2353 DVSS.t108 77.6019
R15688 DVSS.n2922 DVSS.t137 77.6019
R15689 DVSS.n2866 DVSS.n530 76.4173
R15690 DVSS.n1884 DVSS.n1883 76.2208
R15691 DVSS.n1266 DVSS.n1265 76.2208
R15692 DVSS.n653 DVSS.n652 76.2208
R15693 DVSS.n64 DVSS.n63 76.2208
R15694 DVSS.n1883 DVSS.n1882 76.2204
R15695 DVSS.n1265 DVSS.n1264 76.2204
R15696 DVSS.n652 DVSS.n651 76.2204
R15697 DVSS.n63 DVSS.n62 76.2204
R15698 DVSS.n2229 DVSS.n2227 76.2201
R15699 DVSS.n2236 DVSS.n2235 76.2201
R15700 DVSS.n2240 DVSS.n2225 76.2201
R15701 DVSS.n2243 DVSS.n2242 76.2201
R15702 DVSS.n2230 DVSS.n2229 76.2201
R15703 DVSS.n2235 DVSS.n2234 76.2201
R15704 DVSS.n2237 DVSS.n2225 76.2201
R15705 DVSS.n2242 DVSS.n2241 76.2201
R15706 DVSS.n1611 DVSS.n1609 76.2201
R15707 DVSS.n1618 DVSS.n1617 76.2201
R15708 DVSS.n1622 DVSS.n1607 76.2201
R15709 DVSS.n1625 DVSS.n1624 76.2201
R15710 DVSS.n1612 DVSS.n1611 76.2201
R15711 DVSS.n1617 DVSS.n1616 76.2201
R15712 DVSS.n1619 DVSS.n1607 76.2201
R15713 DVSS.n1624 DVSS.n1623 76.2201
R15714 DVSS.n998 DVSS.n996 76.2201
R15715 DVSS.n1005 DVSS.n1004 76.2201
R15716 DVSS.n1009 DVSS.n994 76.2201
R15717 DVSS.n1012 DVSS.n1011 76.2201
R15718 DVSS.n999 DVSS.n998 76.2201
R15719 DVSS.n1004 DVSS.n1003 76.2201
R15720 DVSS.n1006 DVSS.n994 76.2201
R15721 DVSS.n1011 DVSS.n1010 76.2201
R15722 DVSS.n409 DVSS.n407 76.2201
R15723 DVSS.n416 DVSS.n415 76.2201
R15724 DVSS.n420 DVSS.n405 76.2201
R15725 DVSS.n423 DVSS.n422 76.2201
R15726 DVSS.n410 DVSS.n409 76.2201
R15727 DVSS.n415 DVSS.n414 76.2201
R15728 DVSS.n417 DVSS.n405 76.2201
R15729 DVSS.n422 DVSS.n421 76.2201
R15730 DVSS.n2727 DVSS.t182 72.786
R15731 DVSS.n2493 DVSS.t158 72.631
R15732 DVSS.n2613 DVSS.t67 71.8278
R15733 DVSS.n3052 DVSS.n3051 69.6175
R15734 DVSS.n586 DVSS.n584 69.3226
R15735 DVSS.n3015 DVSS.n3013 69.3226
R15736 DVSS.n1198 DVSS.n1196 69.3226
R15737 DVSS.n1831 DVSS.n1829 69.3226
R15738 DVSS.n3069 DVSS.n3068 69.1308
R15739 DVSS.n2723 DVSS.t180 68.0901
R15740 DVSS.n2489 DVSS.t156 67.9451
R15741 DVSS.n2609 DVSS.t65 67.1938
R15742 DVSS.n1971 DVSS.t84 66.8281
R15743 DVSS.n1950 DVSS.t80 66.8281
R15744 DVSS.n1353 DVSS.t189 66.8281
R15745 DVSS.n1332 DVSS.t16 66.8281
R15746 DVSS.n740 DVSS.t29 66.8281
R15747 DVSS.n719 DVSS.t11 66.8281
R15748 DVSS.n151 DVSS.t14 66.8281
R15749 DVSS.n130 DVSS.t46 66.8281
R15750 DVSS.n2370 DVSS.t106 64.639
R15751 DVSS.n2939 DVSS.t133 64.639
R15752 DVSS.n1139 DVSS.t97 64.6385
R15753 DVSS.n1752 DVSS.t168 64.6385
R15754 DVSS.n3046 DVSS.t40 60.0395
R15755 DVSS.n2162 DVSS.n2161 59.4692
R15756 DVSS.n1544 DVSS.n1543 59.4692
R15757 DVSS.n931 DVSS.n930 59.4692
R15758 DVSS.n342 DVSS.n341 59.4692
R15759 DVSS.n2029 DVSS.n2010 59.4689
R15760 DVSS.n2060 DVSS.n2031 59.4689
R15761 DVSS.n2142 DVSS.n1987 59.4689
R15762 DVSS.n2091 DVSS.n2090 59.4689
R15763 DVSS.n2086 DVSS.n2076 59.4689
R15764 DVSS.n2067 DVSS.n2021 59.4689
R15765 DVSS.n2027 DVSS.n2026 59.4689
R15766 DVSS.n1920 DVSS.n1913 59.4689
R15767 DVSS.n1914 DVSS.n1912 59.4689
R15768 DVSS.n2276 DVSS.n2275 59.4689
R15769 DVSS.n2273 DVSS.n2272 59.4689
R15770 DVSS.n1411 DVSS.n1392 59.4689
R15771 DVSS.n1442 DVSS.n1413 59.4689
R15772 DVSS.n1524 DVSS.n1369 59.4689
R15773 DVSS.n1473 DVSS.n1472 59.4689
R15774 DVSS.n1468 DVSS.n1458 59.4689
R15775 DVSS.n1449 DVSS.n1403 59.4689
R15776 DVSS.n1409 DVSS.n1408 59.4689
R15777 DVSS.n1302 DVSS.n1295 59.4689
R15778 DVSS.n1296 DVSS.n1294 59.4689
R15779 DVSS.n1658 DVSS.n1657 59.4689
R15780 DVSS.n1655 DVSS.n1654 59.4689
R15781 DVSS.n798 DVSS.n779 59.4689
R15782 DVSS.n829 DVSS.n800 59.4689
R15783 DVSS.n911 DVSS.n756 59.4689
R15784 DVSS.n860 DVSS.n859 59.4689
R15785 DVSS.n855 DVSS.n845 59.4689
R15786 DVSS.n836 DVSS.n790 59.4689
R15787 DVSS.n796 DVSS.n795 59.4689
R15788 DVSS.n689 DVSS.n682 59.4689
R15789 DVSS.n683 DVSS.n681 59.4689
R15790 DVSS.n1045 DVSS.n1044 59.4689
R15791 DVSS.n1042 DVSS.n1041 59.4689
R15792 DVSS.n209 DVSS.n190 59.4689
R15793 DVSS.n240 DVSS.n211 59.4689
R15794 DVSS.n322 DVSS.n167 59.4689
R15795 DVSS.n271 DVSS.n270 59.4689
R15796 DVSS.n266 DVSS.n256 59.4689
R15797 DVSS.n247 DVSS.n201 59.4689
R15798 DVSS.n207 DVSS.n206 59.4689
R15799 DVSS.n100 DVSS.n93 59.4689
R15800 DVSS.n94 DVSS.n92 59.4689
R15801 DVSS.n456 DVSS.n455 59.4689
R15802 DVSS.n453 DVSS.n452 59.4689
R15803 DVSS.n2790 DVSS.n2789 59.3519
R15804 DVSS.n2812 DVSS.n2811 59.3519
R15805 DVSS.n1885 DVSS.n1879 55.6474
R15806 DVSS.n1267 DVSS.n1261 55.6474
R15807 DVSS.n654 DVSS.n648 55.6474
R15808 DVSS.n65 DVSS.n59 55.6474
R15809 DVSS.n1897 DVSS.n1896 55.6471
R15810 DVSS.n1279 DVSS.n1278 55.6471
R15811 DVSS.n666 DVSS.n665 55.6471
R15812 DVSS.n77 DVSS.n76 55.6471
R15813 DVSS.n2545 DVSS.n2544 55.6087
R15814 DVSS.n1692 DVSS.n1691 52.3069
R15815 DVSS.n2310 DVSS.n2309 52.3069
R15816 DVSS.n1079 DVSS.n1078 52.3069
R15817 DVSS.n2879 DVSS.n2878 52.3069
R15818 DVSS.t101 DVSS.n1109 50.7875
R15819 DVSS.t172 DVSS.n1722 50.7875
R15820 DVSS.n2371 DVSS.n2370 47.1783
R15821 DVSS.n2940 DVSS.n2939 47.1783
R15822 DVSS.n1122 DVSS.t99 46.1705
R15823 DVSS.n1735 DVSS.t170 46.1705
R15824 DVSS.n2089 DVSS.n2068 45.5782
R15825 DVSS.n2096 DVSS.n2095 45.5782
R15826 DVSS.n1471 DVSS.n1450 45.5782
R15827 DVSS.n1478 DVSS.n1477 45.5782
R15828 DVSS.n858 DVSS.n837 45.5782
R15829 DVSS.n865 DVSS.n864 45.5782
R15830 DVSS.n269 DVSS.n248 45.5782
R15831 DVSS.n276 DVSS.n275 45.5782
R15832 DVSS.n2826 DVSS.n2825 43.8838
R15833 DVSS.n3073 DVSS.t38 42.8855
R15834 DVSS.n2134 DVSS.n2133 42.4097
R15835 DVSS.n1516 DVSS.n1515 42.4097
R15836 DVSS.n903 DVSS.n902 42.4097
R15837 DVSS.n314 DVSS.n313 42.4097
R15838 DVSS.n1774 DVSS.n1773 38.7626
R15839 DVSS.n1809 DVSS.t125 38.0722
R15840 DVSS.n567 DVSS.t21 38.0722
R15841 DVSS.n2164 DVSS.n1980 36.7611
R15842 DVSS.n1546 DVSS.n1362 36.7611
R15843 DVSS.n933 DVSS.n749 36.7611
R15844 DVSS.n344 DVSS.n160 36.7611
R15845 DVSS.n2586 DVSS.n2585 36.5724
R15846 DVSS.t3 DVSS.t174 36.1979
R15847 DVSS.n2436 DVSS.n2433 36.1417
R15848 DVSS.n2669 DVSS.n2668 36.1417
R15849 DVSS.n3002 DVSS.n2999 36.1417
R15850 DVSS.n2772 DVSS.t30 35.7314
R15851 DVSS.n2535 DVSS.t1 35.5663
R15852 DVSS.n2112 DVSS.n2110 35.3887
R15853 DVSS.n2136 DVSS.n2123 35.3887
R15854 DVSS.n2110 DVSS.n2014 35.3887
R15855 DVSS.n2116 DVSS.n2009 35.3887
R15856 DVSS.n2104 DVSS.n2009 35.3887
R15857 DVSS.n1494 DVSS.n1492 35.3887
R15858 DVSS.n1518 DVSS.n1505 35.3887
R15859 DVSS.n1492 DVSS.n1396 35.3887
R15860 DVSS.n1498 DVSS.n1391 35.3887
R15861 DVSS.n1486 DVSS.n1391 35.3887
R15862 DVSS.n881 DVSS.n879 35.3887
R15863 DVSS.n905 DVSS.n892 35.3887
R15864 DVSS.n879 DVSS.n783 35.3887
R15865 DVSS.n885 DVSS.n778 35.3887
R15866 DVSS.n873 DVSS.n778 35.3887
R15867 DVSS.n292 DVSS.n290 35.3887
R15868 DVSS.n316 DVSS.n303 35.3887
R15869 DVSS.n290 DVSS.n194 35.3887
R15870 DVSS.n296 DVSS.n189 35.3887
R15871 DVSS.n284 DVSS.n189 35.3887
R15872 DVSS.n2789 DVSS.t91 35.0689
R15873 DVSS.n2811 DVSS.t60 35.0689
R15874 DVSS.n2255 DVSS.n1848 34.1338
R15875 DVSS.n1881 DVSS.n1867 34.1338
R15876 DVSS.n1637 DVSS.n1230 34.1338
R15877 DVSS.n1263 DVSS.n1249 34.1338
R15878 DVSS.n1024 DVSS.n617 34.1338
R15879 DVSS.n650 DVSS.n636 34.1338
R15880 DVSS.n435 DVSS.n28 34.1338
R15881 DVSS.n61 DVSS.n47 34.1338
R15882 DVSS.n2721 DVSS.n2719 33.5205
R15883 DVSS.n583 DVSS.n582 33.5205
R15884 DVSS.n3057 DVSS.n3055 33.5205
R15885 DVSS.n7 DVSS.n6 33.5205
R15886 DVSS.n1733 DVSS.n1732 33.5205
R15887 DVSS.n1750 DVSS.n1749 33.5205
R15888 DVSS.n2607 DVSS.n2605 33.5205
R15889 DVSS.n1195 DVSS.n1194 33.5205
R15890 DVSS.n2503 DVSS.n2502 33.5205
R15891 DVSS.n2487 DVSS.n2485 33.5205
R15892 DVSS.n2351 DVSS.n2350 33.5205
R15893 DVSS.n2368 DVSS.n2367 33.5205
R15894 DVSS.n1120 DVSS.n1119 33.5205
R15895 DVSS.n1137 DVSS.n1136 33.5205
R15896 DVSS.n2920 DVSS.n2919 33.5205
R15897 DVSS.n2937 DVSS.n2936 33.5205
R15898 DVSS.n484 DVSS.n483 30.5709
R15899 DVSS.n2136 DVSS.n2135 29.7417
R15900 DVSS.n1518 DVSS.n1517 29.7417
R15901 DVSS.n905 DVSS.n904 29.7417
R15902 DVSS.n316 DVSS.n315 29.7417
R15903 DVSS.n1972 DVSS.n1961 29.4833
R15904 DVSS.n1951 DVSS.n1940 29.4833
R15905 DVSS.n1354 DVSS.n1343 29.4833
R15906 DVSS.n1333 DVSS.n1322 29.4833
R15907 DVSS.n741 DVSS.n730 29.4833
R15908 DVSS.n720 DVSS.n709 29.4833
R15909 DVSS.n152 DVSS.n141 29.4833
R15910 DVSS.n131 DVSS.n120 29.4833
R15911 DVSS.n1921 DVSS.n1904 29.1989
R15912 DVSS.n2278 DVSS.n2257 29.1989
R15913 DVSS.n1303 DVSS.n1286 29.1989
R15914 DVSS.n1660 DVSS.n1639 29.1989
R15915 DVSS.n690 DVSS.n673 29.1989
R15916 DVSS.n1047 DVSS.n1026 29.1989
R15917 DVSS.n101 DVSS.n84 29.1989
R15918 DVSS.n458 DVSS.n437 29.1989
R15919 DVSS.n2779 DVSS.n2778 28.2915
R15920 DVSS.n2363 DVSS.n2362 28.2515
R15921 DVSS.n2932 DVSS.n2931 28.2515
R15922 DVSS.n1691 DVSS.t187 28.1205
R15923 DVSS.n2309 DVSS.t74 28.1205
R15924 DVSS.n1078 DVSS.t132 28.1205
R15925 DVSS.n2878 DVSS.t26 28.1205
R15926 DVSS.n2664 DVSS.n2663 27.8046
R15927 DVSS.n2112 DVSS.n2111 25.6005
R15928 DVSS.n2111 DVSS.n2006 25.6005
R15929 DVSS.n2123 DVSS.n2006 25.6005
R15930 DVSS.n2098 DVSS.n2096 25.6005
R15931 DVSS.n2098 DVSS.n2097 25.6005
R15932 DVSS.n2097 DVSS.n2014 25.6005
R15933 DVSS.n2135 DVSS.n2134 25.6005
R15934 DVSS.n2117 DVSS.n2116 25.6005
R15935 DVSS.n2118 DVSS.n2117 25.6005
R15936 DVSS.n2118 DVSS.n1980 25.6005
R15937 DVSS.n2102 DVSS.n2068 25.6005
R15938 DVSS.n2103 DVSS.n2102 25.6005
R15939 DVSS.n2104 DVSS.n2103 25.6005
R15940 DVSS.n1494 DVSS.n1493 25.6005
R15941 DVSS.n1493 DVSS.n1388 25.6005
R15942 DVSS.n1505 DVSS.n1388 25.6005
R15943 DVSS.n1480 DVSS.n1478 25.6005
R15944 DVSS.n1480 DVSS.n1479 25.6005
R15945 DVSS.n1479 DVSS.n1396 25.6005
R15946 DVSS.n1517 DVSS.n1516 25.6005
R15947 DVSS.n1499 DVSS.n1498 25.6005
R15948 DVSS.n1500 DVSS.n1499 25.6005
R15949 DVSS.n1500 DVSS.n1362 25.6005
R15950 DVSS.n1484 DVSS.n1450 25.6005
R15951 DVSS.n1485 DVSS.n1484 25.6005
R15952 DVSS.n1486 DVSS.n1485 25.6005
R15953 DVSS.n881 DVSS.n880 25.6005
R15954 DVSS.n880 DVSS.n775 25.6005
R15955 DVSS.n892 DVSS.n775 25.6005
R15956 DVSS.n867 DVSS.n865 25.6005
R15957 DVSS.n867 DVSS.n866 25.6005
R15958 DVSS.n866 DVSS.n783 25.6005
R15959 DVSS.n904 DVSS.n903 25.6005
R15960 DVSS.n886 DVSS.n885 25.6005
R15961 DVSS.n887 DVSS.n886 25.6005
R15962 DVSS.n887 DVSS.n749 25.6005
R15963 DVSS.n871 DVSS.n837 25.6005
R15964 DVSS.n872 DVSS.n871 25.6005
R15965 DVSS.n873 DVSS.n872 25.6005
R15966 DVSS.n292 DVSS.n291 25.6005
R15967 DVSS.n291 DVSS.n186 25.6005
R15968 DVSS.n303 DVSS.n186 25.6005
R15969 DVSS.n278 DVSS.n276 25.6005
R15970 DVSS.n278 DVSS.n277 25.6005
R15971 DVSS.n277 DVSS.n194 25.6005
R15972 DVSS.n315 DVSS.n314 25.6005
R15973 DVSS.n297 DVSS.n296 25.6005
R15974 DVSS.n298 DVSS.n297 25.6005
R15975 DVSS.n298 DVSS.n160 25.6005
R15976 DVSS.n282 DVSS.n248 25.6005
R15977 DVSS.n283 DVSS.n282 25.6005
R15978 DVSS.n284 DVSS.n283 25.6005
R15979 DVSS.n2231 DVSS.n1848 22.3184
R15980 DVSS.n2232 DVSS.n2231 22.3184
R15981 DVSS.n2233 DVSS.n2232 22.3184
R15982 DVSS.n2233 DVSS.n2226 22.3184
R15983 DVSS.n2238 DVSS.n2226 22.3184
R15984 DVSS.n2239 DVSS.n2238 22.3184
R15985 DVSS.n2239 DVSS.n2224 22.3184
R15986 DVSS.n2244 DVSS.n2224 22.3184
R15987 DVSS.n1881 DVSS.n1880 22.3184
R15988 DVSS.n1886 DVSS.n1880 22.3184
R15989 DVSS.n1887 DVSS.n1886 22.3184
R15990 DVSS.n1887 DVSS.n1878 22.3184
R15991 DVSS.n1893 DVSS.n1878 22.3184
R15992 DVSS.n1894 DVSS.n1893 22.3184
R15993 DVSS.n1894 DVSS.n1876 22.3184
R15994 DVSS.n1899 DVSS.n1876 22.3184
R15995 DVSS.n1613 DVSS.n1230 22.3184
R15996 DVSS.n1614 DVSS.n1613 22.3184
R15997 DVSS.n1615 DVSS.n1614 22.3184
R15998 DVSS.n1615 DVSS.n1608 22.3184
R15999 DVSS.n1620 DVSS.n1608 22.3184
R16000 DVSS.n1621 DVSS.n1620 22.3184
R16001 DVSS.n1621 DVSS.n1606 22.3184
R16002 DVSS.n1626 DVSS.n1606 22.3184
R16003 DVSS.n1263 DVSS.n1262 22.3184
R16004 DVSS.n1268 DVSS.n1262 22.3184
R16005 DVSS.n1269 DVSS.n1268 22.3184
R16006 DVSS.n1269 DVSS.n1260 22.3184
R16007 DVSS.n1275 DVSS.n1260 22.3184
R16008 DVSS.n1276 DVSS.n1275 22.3184
R16009 DVSS.n1276 DVSS.n1258 22.3184
R16010 DVSS.n1281 DVSS.n1258 22.3184
R16011 DVSS.n1000 DVSS.n617 22.3184
R16012 DVSS.n1001 DVSS.n1000 22.3184
R16013 DVSS.n1002 DVSS.n1001 22.3184
R16014 DVSS.n1002 DVSS.n995 22.3184
R16015 DVSS.n1007 DVSS.n995 22.3184
R16016 DVSS.n1008 DVSS.n1007 22.3184
R16017 DVSS.n1008 DVSS.n993 22.3184
R16018 DVSS.n1013 DVSS.n993 22.3184
R16019 DVSS.n650 DVSS.n649 22.3184
R16020 DVSS.n655 DVSS.n649 22.3184
R16021 DVSS.n656 DVSS.n655 22.3184
R16022 DVSS.n656 DVSS.n647 22.3184
R16023 DVSS.n662 DVSS.n647 22.3184
R16024 DVSS.n663 DVSS.n662 22.3184
R16025 DVSS.n663 DVSS.n645 22.3184
R16026 DVSS.n668 DVSS.n645 22.3184
R16027 DVSS.n411 DVSS.n28 22.3184
R16028 DVSS.n412 DVSS.n411 22.3184
R16029 DVSS.n413 DVSS.n412 22.3184
R16030 DVSS.n413 DVSS.n406 22.3184
R16031 DVSS.n418 DVSS.n406 22.3184
R16032 DVSS.n419 DVSS.n418 22.3184
R16033 DVSS.n419 DVSS.n404 22.3184
R16034 DVSS.n424 DVSS.n404 22.3184
R16035 DVSS.n61 DVSS.n60 22.3184
R16036 DVSS.n66 DVSS.n60 22.3184
R16037 DVSS.n67 DVSS.n66 22.3184
R16038 DVSS.n67 DVSS.n58 22.3184
R16039 DVSS.n73 DVSS.n58 22.3184
R16040 DVSS.n74 DVSS.n73 22.3184
R16041 DVSS.n74 DVSS.n56 22.3184
R16042 DVSS.n79 DVSS.n56 22.3184
R16043 DVSS.n2789 DVSS.t5 22.2377
R16044 DVSS.n2811 DVSS.t92 22.2377
R16045 DVSS.n1691 DVSS.t62 21.2805
R16046 DVSS.n2309 DVSS.t151 21.2805
R16047 DVSS.n1078 DVSS.t20 21.2805
R16048 DVSS.n2825 DVSS.t88 21.2805
R16049 DVSS.n2825 DVSS.t89 21.2805
R16050 DVSS.n2878 DVSS.t78 21.2805
R16051 DVSS.n2245 DVSS.n2244 20.3492
R16052 DVSS.n1900 DVSS.n1899 20.3492
R16053 DVSS.n1627 DVSS.n1626 20.3492
R16054 DVSS.n1282 DVSS.n1281 20.3492
R16055 DVSS.n1014 DVSS.n1013 20.3492
R16056 DVSS.n669 DVSS.n668 20.3492
R16057 DVSS.n425 DVSS.n424 20.3492
R16058 DVSS.n80 DVSS.n79 20.3492
R16059 DVSS.n584 DVSS.t104 20.0005
R16060 DVSS.n584 DVSS.t43 20.0005
R16061 DVSS.n3013 DVSS.t142 20.0005
R16062 DVSS.n3013 DVSS.t146 20.0005
R16063 DVSS.n1196 DVSS.t163 20.0005
R16064 DVSS.n1196 DVSS.t120 20.0005
R16065 DVSS.n1829 DVSS.t115 20.0005
R16066 DVSS.n1829 DVSS.t128 20.0005
R16067 DVSS.n2700 DVSS.n2699 18.7839
R16068 DVSS.n3037 DVSS.n3036 18.153
R16069 DVSS.n1178 DVSS.n1177 18.0103
R16070 DVSS.n1791 DVSS.n1790 18.0103
R16071 DVSS.n2810 DVSS.n2806 18.0093
R16072 DVSS.n2864 DVSS.n2863 17.2422
R16073 DVSS.n2255 DVSS.n2254 17.0218
R16074 DVSS.n1637 DVSS.n1636 17.0218
R16075 DVSS.n1024 DVSS.n1023 17.0218
R16076 DVSS.n435 DVSS.n434 17.0218
R16077 DVSS.n2206 DVSS.n1867 16.8856
R16078 DVSS.n1588 DVSS.n1249 16.8856
R16079 DVSS.n975 DVSS.n636 16.8856
R16080 DVSS.n386 DVSS.n47 16.8856
R16081 DVSS.n2710 DVSS.t178 16.4359
R16082 DVSS.n2476 DVSS.t152 16.4009
R16083 DVSS.n2596 DVSS.t63 16.2196
R16084 DVSS.n2188 DVSS.n1867 15.5239
R16085 DVSS.n1570 DVSS.n1249 15.5239
R16086 DVSS.n957 DVSS.n636 15.5239
R16087 DVSS.n368 DVSS.n47 15.5239
R16088 DVSS.n1970 DVSS.n1969 15.463
R16089 DVSS.n1949 DVSS.n1948 15.463
R16090 DVSS.n1352 DVSS.n1351 15.463
R16091 DVSS.n1331 DVSS.n1330 15.463
R16092 DVSS.n739 DVSS.n738 15.463
R16093 DVSS.n718 DVSS.n717 15.463
R16094 DVSS.n150 DVSS.n149 15.463
R16095 DVSS.n129 DVSS.n128 15.463
R16096 DVSS.n2256 DVSS.n2255 15.3877
R16097 DVSS.n1638 DVSS.n1637 15.3877
R16098 DVSS.n1025 DVSS.n1024 15.3877
R16099 DVSS.n436 DVSS.n435 15.3877
R16100 DVSS.n2534 DVSS 15.0005
R16101 DVSS.n485 DVSS.n484 14.4554
R16102 DVSS.n2827 DVSS.n2826 14.4288
R16103 DVSS.n2716 DVSS.n2715 14.387
R16104 DVSS.n2482 DVSS.n2481 14.3654
R16105 DVSS.n2733 DVSS.n2732 14.3449
R16106 DVSS.n2499 DVSS.n2498 14.3234
R16107 DVSS.n2602 DVSS.n2601 14.2541
R16108 DVSS.n2619 DVSS.n2618 14.213
R16109 DVSS.n1975 DVSS.n1962 13.5534
R16110 DVSS.n1970 DVSS.n1966 13.5534
R16111 DVSS.n1954 DVSS.n1941 13.5534
R16112 DVSS.n1949 DVSS.n1945 13.5534
R16113 DVSS.n1357 DVSS.n1344 13.5534
R16114 DVSS.n1352 DVSS.n1348 13.5534
R16115 DVSS.n1336 DVSS.n1323 13.5534
R16116 DVSS.n1331 DVSS.n1327 13.5534
R16117 DVSS.n744 DVSS.n731 13.5534
R16118 DVSS.n739 DVSS.n735 13.5534
R16119 DVSS.n723 DVSS.n710 13.5534
R16120 DVSS.n718 DVSS.n714 13.5534
R16121 DVSS.n155 DVSS.n142 13.5534
R16122 DVSS.n150 DVSS.n146 13.5534
R16123 DVSS.n134 DVSS.n121 13.5534
R16124 DVSS.n129 DVSS.n125 13.5534
R16125 DVSS.n2802 DVSS.n2801 13.5112
R16126 DVSS.n2303 DVSS.n2299 12.8977
R16127 DVSS.n1685 DVSS.n1684 12.8977
R16128 DVSS.n1072 DVSS.n1071 12.8977
R16129 DVSS.n2872 DVSS.n2871 12.8977
R16130 DVSS.n525 DVSS.n521 12.8862
R16131 DVSS.n2737 DVSS.t184 11.7401
R16132 DVSS.n2505 DVSS.t160 11.7151
R16133 DVSS.n2623 DVSS.t69 11.5855
R16134 DVSS.n582 DVSS.t185 10.6405
R16135 DVSS.n582 DVSS.t183 10.6405
R16136 DVSS.n2719 DVSS.t181 10.6405
R16137 DVSS.n2719 DVSS.t179 10.6405
R16138 DVSS.n6 DVSS.t39 10.6405
R16139 DVSS.n6 DVSS.t37 10.6405
R16140 DVSS.n3055 DVSS.t35 10.6405
R16141 DVSS.n3055 DVSS.t41 10.6405
R16142 DVSS.n1732 DVSS.t173 10.6405
R16143 DVSS.n1732 DVSS.t171 10.6405
R16144 DVSS.n1749 DVSS.t167 10.6405
R16145 DVSS.n1749 DVSS.t169 10.6405
R16146 DVSS.n1194 DVSS.t70 10.6405
R16147 DVSS.n1194 DVSS.t68 10.6405
R16148 DVSS.n2605 DVSS.t66 10.6405
R16149 DVSS.n2605 DVSS.t64 10.6405
R16150 DVSS.n2502 DVSS.t161 10.6405
R16151 DVSS.n2502 DVSS.t159 10.6405
R16152 DVSS.n2485 DVSS.t157 10.6405
R16153 DVSS.n2485 DVSS.t153 10.6405
R16154 DVSS.n2350 DVSS.t117 10.6405
R16155 DVSS.n2350 DVSS.t109 10.6405
R16156 DVSS.n2367 DVSS.t113 10.6405
R16157 DVSS.n2367 DVSS.t107 10.6405
R16158 DVSS.n1119 DVSS.t102 10.6405
R16159 DVSS.n1119 DVSS.t100 10.6405
R16160 DVSS.n1136 DVSS.t94 10.6405
R16161 DVSS.n1136 DVSS.t98 10.6405
R16162 DVSS.n2919 DVSS.t140 10.6405
R16163 DVSS.n2919 DVSS.t138 10.6405
R16164 DVSS.n2936 DVSS.t136 10.6405
R16165 DVSS.n2936 DVSS.t134 10.6405
R16166 DVSS.n2125 DVSS.n2002 10.4252
R16167 DVSS.n1507 DVSS.n1384 10.4252
R16168 DVSS.n894 DVSS.n771 10.4252
R16169 DVSS.n305 DVSS.n182 10.4252
R16170 DVSS.n2468 DVSS.n2467 9.85124
R16171 DVSS.n2587 DVSS.n2586 9.5204
R16172 DVSS.n2295 DVSS.n2294 9.31763
R16173 DVSS.n1677 DVSS.n1676 9.31763
R16174 DVSS.n1064 DVSS.n1063 9.31763
R16175 DVSS.n475 DVSS.n474 9.31763
R16176 DVSS.n2393 DVSS.n2392 9.3005
R16177 DVSS.n1960 DVSS.n1959 9.3005
R16178 DVSS.n1967 DVSS.n1963 9.3005
R16179 DVSS.n1968 DVSS.n1966 9.3005
R16180 DVSS.n1973 DVSS.n1965 9.3005
R16181 DVSS.n1973 DVSS.n1972 9.3005
R16182 DVSS.n1964 DVSS.n1962 9.3005
R16183 DVSS.n1978 DVSS.n1977 9.3005
R16184 DVSS.n1939 DVSS.n1938 9.3005
R16185 DVSS.n1946 DVSS.n1942 9.3005
R16186 DVSS.n1947 DVSS.n1945 9.3005
R16187 DVSS.n1952 DVSS.n1944 9.3005
R16188 DVSS.n1952 DVSS.n1951 9.3005
R16189 DVSS.n1943 DVSS.n1941 9.3005
R16190 DVSS.n1957 DVSS.n1956 9.3005
R16191 DVSS.n2173 DVSS.n2172 9.3005
R16192 DVSS.n2176 DVSS.n2175 9.3005
R16193 DVSS.n2177 DVSS.n1908 9.3005
R16194 DVSS.n2182 DVSS.n2181 9.3005
R16195 DVSS.n2180 DVSS.n1909 9.3005
R16196 DVSS.n2179 DVSS.n2178 9.3005
R16197 DVSS.n1875 DVSS.n1874 9.3005
R16198 DVSS.n2193 DVSS.n2192 9.3005
R16199 DVSS.n2194 DVSS.n1872 9.3005
R16200 DVSS.n2202 DVSS.n2201 9.3005
R16201 DVSS.n2200 DVSS.n1873 9.3005
R16202 DVSS.n2197 DVSS.n2196 9.3005
R16203 DVSS.n2195 DVSS.n1861 9.3005
R16204 DVSS.n2213 DVSS.n1860 9.3005
R16205 DVSS.n2215 DVSS.n2214 9.3005
R16206 DVSS.n2216 DVSS.n1859 9.3005
R16207 DVSS.n2219 DVSS.n1858 9.3005
R16208 DVSS.n2221 DVSS.n2220 9.3005
R16209 DVSS.n2222 DVSS.n1856 9.3005
R16210 DVSS.n2250 DVSS.n2249 9.3005
R16211 DVSS.n2248 DVSS.n1857 9.3005
R16212 DVSS.n2247 DVSS.n2246 9.3005
R16213 DVSS.n2223 DVSS.n1841 9.3005
R16214 DVSS.n2284 DVSS.n1842 9.3005
R16215 DVSS.n2285 DVSS.n1840 9.3005
R16216 DVSS.n2287 DVSS.n2286 9.3005
R16217 DVSS.n2288 DVSS.n1839 9.3005
R16218 DVSS.n2290 DVSS.n2289 9.3005
R16219 DVSS.n2425 DVSS.n2424 9.3005
R16220 DVSS.n1200 DVSS.n1199 9.3005
R16221 DVSS.n1211 DVSS.n1210 9.3005
R16222 DVSS.n1342 DVSS.n1341 9.3005
R16223 DVSS.n1349 DVSS.n1345 9.3005
R16224 DVSS.n1350 DVSS.n1348 9.3005
R16225 DVSS.n1355 DVSS.n1347 9.3005
R16226 DVSS.n1355 DVSS.n1354 9.3005
R16227 DVSS.n1346 DVSS.n1344 9.3005
R16228 DVSS.n1360 DVSS.n1359 9.3005
R16229 DVSS.n1321 DVSS.n1320 9.3005
R16230 DVSS.n1328 DVSS.n1324 9.3005
R16231 DVSS.n1329 DVSS.n1327 9.3005
R16232 DVSS.n1334 DVSS.n1326 9.3005
R16233 DVSS.n1334 DVSS.n1333 9.3005
R16234 DVSS.n1325 DVSS.n1323 9.3005
R16235 DVSS.n1339 DVSS.n1338 9.3005
R16236 DVSS.n1555 DVSS.n1554 9.3005
R16237 DVSS.n1558 DVSS.n1557 9.3005
R16238 DVSS.n1559 DVSS.n1290 9.3005
R16239 DVSS.n1564 DVSS.n1563 9.3005
R16240 DVSS.n1562 DVSS.n1291 9.3005
R16241 DVSS.n1561 DVSS.n1560 9.3005
R16242 DVSS.n1257 DVSS.n1256 9.3005
R16243 DVSS.n1575 DVSS.n1574 9.3005
R16244 DVSS.n1576 DVSS.n1254 9.3005
R16245 DVSS.n1584 DVSS.n1583 9.3005
R16246 DVSS.n1582 DVSS.n1255 9.3005
R16247 DVSS.n1579 DVSS.n1578 9.3005
R16248 DVSS.n1577 DVSS.n1243 9.3005
R16249 DVSS.n1595 DVSS.n1242 9.3005
R16250 DVSS.n1597 DVSS.n1596 9.3005
R16251 DVSS.n1598 DVSS.n1241 9.3005
R16252 DVSS.n1601 DVSS.n1240 9.3005
R16253 DVSS.n1603 DVSS.n1602 9.3005
R16254 DVSS.n1604 DVSS.n1238 9.3005
R16255 DVSS.n1632 DVSS.n1631 9.3005
R16256 DVSS.n1630 DVSS.n1239 9.3005
R16257 DVSS.n1629 DVSS.n1628 9.3005
R16258 DVSS.n1605 DVSS.n1223 9.3005
R16259 DVSS.n1666 DVSS.n1224 9.3005
R16260 DVSS.n1667 DVSS.n1222 9.3005
R16261 DVSS.n1669 DVSS.n1668 9.3005
R16262 DVSS.n1670 DVSS.n1221 9.3005
R16263 DVSS.n1672 DVSS.n1671 9.3005
R16264 DVSS.n1780 DVSS.n1779 9.3005
R16265 DVSS.n729 DVSS.n728 9.3005
R16266 DVSS.n736 DVSS.n732 9.3005
R16267 DVSS.n737 DVSS.n735 9.3005
R16268 DVSS.n742 DVSS.n734 9.3005
R16269 DVSS.n742 DVSS.n741 9.3005
R16270 DVSS.n733 DVSS.n731 9.3005
R16271 DVSS.n747 DVSS.n746 9.3005
R16272 DVSS.n708 DVSS.n707 9.3005
R16273 DVSS.n715 DVSS.n711 9.3005
R16274 DVSS.n716 DVSS.n714 9.3005
R16275 DVSS.n721 DVSS.n713 9.3005
R16276 DVSS.n721 DVSS.n720 9.3005
R16277 DVSS.n712 DVSS.n710 9.3005
R16278 DVSS.n726 DVSS.n725 9.3005
R16279 DVSS.n942 DVSS.n941 9.3005
R16280 DVSS.n945 DVSS.n944 9.3005
R16281 DVSS.n946 DVSS.n677 9.3005
R16282 DVSS.n951 DVSS.n950 9.3005
R16283 DVSS.n949 DVSS.n678 9.3005
R16284 DVSS.n948 DVSS.n947 9.3005
R16285 DVSS.n644 DVSS.n643 9.3005
R16286 DVSS.n962 DVSS.n961 9.3005
R16287 DVSS.n963 DVSS.n641 9.3005
R16288 DVSS.n971 DVSS.n970 9.3005
R16289 DVSS.n969 DVSS.n642 9.3005
R16290 DVSS.n966 DVSS.n965 9.3005
R16291 DVSS.n964 DVSS.n630 9.3005
R16292 DVSS.n982 DVSS.n629 9.3005
R16293 DVSS.n984 DVSS.n983 9.3005
R16294 DVSS.n985 DVSS.n628 9.3005
R16295 DVSS.n988 DVSS.n627 9.3005
R16296 DVSS.n990 DVSS.n989 9.3005
R16297 DVSS.n991 DVSS.n625 9.3005
R16298 DVSS.n1019 DVSS.n1018 9.3005
R16299 DVSS.n1017 DVSS.n626 9.3005
R16300 DVSS.n1016 DVSS.n1015 9.3005
R16301 DVSS.n992 DVSS.n610 9.3005
R16302 DVSS.n1053 DVSS.n611 9.3005
R16303 DVSS.n1054 DVSS.n609 9.3005
R16304 DVSS.n1056 DVSS.n1055 9.3005
R16305 DVSS.n1057 DVSS.n608 9.3005
R16306 DVSS.n1059 DVSS.n1058 9.3005
R16307 DVSS.n1166 DVSS.n1165 9.3005
R16308 DVSS.n1169 DVSS.n1168 9.3005
R16309 DVSS.n1783 DVSS.n1782 9.3005
R16310 DVSS.n2423 DVSS.n2422 9.3005
R16311 DVSS.n2397 DVSS.n2396 9.3005
R16312 DVSS.n140 DVSS.n139 9.3005
R16313 DVSS.n147 DVSS.n143 9.3005
R16314 DVSS.n148 DVSS.n146 9.3005
R16315 DVSS.n153 DVSS.n145 9.3005
R16316 DVSS.n153 DVSS.n152 9.3005
R16317 DVSS.n144 DVSS.n142 9.3005
R16318 DVSS.n158 DVSS.n157 9.3005
R16319 DVSS.n119 DVSS.n118 9.3005
R16320 DVSS.n126 DVSS.n122 9.3005
R16321 DVSS.n127 DVSS.n125 9.3005
R16322 DVSS.n132 DVSS.n124 9.3005
R16323 DVSS.n132 DVSS.n131 9.3005
R16324 DVSS.n123 DVSS.n121 9.3005
R16325 DVSS.n137 DVSS.n136 9.3005
R16326 DVSS.n353 DVSS.n352 9.3005
R16327 DVSS.n356 DVSS.n355 9.3005
R16328 DVSS.n357 DVSS.n88 9.3005
R16329 DVSS.n362 DVSS.n361 9.3005
R16330 DVSS.n360 DVSS.n89 9.3005
R16331 DVSS.n359 DVSS.n358 9.3005
R16332 DVSS.n55 DVSS.n54 9.3005
R16333 DVSS.n373 DVSS.n372 9.3005
R16334 DVSS.n374 DVSS.n52 9.3005
R16335 DVSS.n382 DVSS.n381 9.3005
R16336 DVSS.n380 DVSS.n53 9.3005
R16337 DVSS.n377 DVSS.n376 9.3005
R16338 DVSS.n375 DVSS.n41 9.3005
R16339 DVSS.n393 DVSS.n40 9.3005
R16340 DVSS.n395 DVSS.n394 9.3005
R16341 DVSS.n396 DVSS.n39 9.3005
R16342 DVSS.n399 DVSS.n38 9.3005
R16343 DVSS.n401 DVSS.n400 9.3005
R16344 DVSS.n402 DVSS.n36 9.3005
R16345 DVSS.n430 DVSS.n429 9.3005
R16346 DVSS.n428 DVSS.n37 9.3005
R16347 DVSS.n427 DVSS.n426 9.3005
R16348 DVSS.n403 DVSS.n21 9.3005
R16349 DVSS.n464 DVSS.n22 9.3005
R16350 DVSS.n465 DVSS.n20 9.3005
R16351 DVSS.n467 DVSS.n466 9.3005
R16352 DVSS.n468 DVSS.n19 9.3005
R16353 DVSS.n470 DVSS.n469 9.3005
R16354 DVSS.n2962 DVSS.n2961 9.3005
R16355 DVSS.n2966 DVSS.n2965 9.3005
R16356 DVSS.n2990 DVSS.n2989 9.3005
R16357 DVSS.n2988 DVSS.n2987 9.3005
R16358 DVSS.n594 DVSS.n593 9.3005
R16359 DVSS.n597 DVSS.n596 9.3005
R16360 DVSS.n2186 DVSS.n1904 9.26007
R16361 DVSS.n2187 DVSS.n2186 9.26007
R16362 DVSS.n2188 DVSS.n2187 9.26007
R16363 DVSS.n2207 DVSS.n2206 9.26007
R16364 DVSS.n2209 DVSS.n2207 9.26007
R16365 DVSS.n2209 DVSS.n2208 9.26007
R16366 DVSS.n2208 DVSS.n1849 9.26007
R16367 DVSS.n2254 DVSS.n1849 9.26007
R16368 DVSS.n2280 DVSS.n2256 9.26007
R16369 DVSS.n2280 DVSS.n2279 9.26007
R16370 DVSS.n2279 DVSS.n2278 9.26007
R16371 DVSS.n1568 DVSS.n1286 9.26007
R16372 DVSS.n1569 DVSS.n1568 9.26007
R16373 DVSS.n1570 DVSS.n1569 9.26007
R16374 DVSS.n1589 DVSS.n1588 9.26007
R16375 DVSS.n1591 DVSS.n1589 9.26007
R16376 DVSS.n1591 DVSS.n1590 9.26007
R16377 DVSS.n1590 DVSS.n1231 9.26007
R16378 DVSS.n1636 DVSS.n1231 9.26007
R16379 DVSS.n1662 DVSS.n1638 9.26007
R16380 DVSS.n1662 DVSS.n1661 9.26007
R16381 DVSS.n1661 DVSS.n1660 9.26007
R16382 DVSS.n955 DVSS.n673 9.26007
R16383 DVSS.n956 DVSS.n955 9.26007
R16384 DVSS.n957 DVSS.n956 9.26007
R16385 DVSS.n976 DVSS.n975 9.26007
R16386 DVSS.n978 DVSS.n976 9.26007
R16387 DVSS.n978 DVSS.n977 9.26007
R16388 DVSS.n977 DVSS.n618 9.26007
R16389 DVSS.n1023 DVSS.n618 9.26007
R16390 DVSS.n1049 DVSS.n1025 9.26007
R16391 DVSS.n1049 DVSS.n1048 9.26007
R16392 DVSS.n1048 DVSS.n1047 9.26007
R16393 DVSS.n366 DVSS.n84 9.26007
R16394 DVSS.n367 DVSS.n366 9.26007
R16395 DVSS.n368 DVSS.n367 9.26007
R16396 DVSS.n387 DVSS.n386 9.26007
R16397 DVSS.n389 DVSS.n387 9.26007
R16398 DVSS.n389 DVSS.n388 9.26007
R16399 DVSS.n388 DVSS.n29 9.26007
R16400 DVSS.n434 DVSS.n29 9.26007
R16401 DVSS.n460 DVSS.n436 9.26007
R16402 DVSS.n460 DVSS.n459 9.26007
R16403 DVSS.n459 DVSS.n458 9.26007
R16404 DVSS.n2299 DVSS.n2298 9.15497
R16405 DVSS.n2302 DVSS.n2301 9.15497
R16406 DVSS.n2301 DVSS.n2300 9.15497
R16407 DVSS.n2307 DVSS.n2306 9.15497
R16408 DVSS.n2306 DVSS.n2305 9.15497
R16409 DVSS.n2314 DVSS.n2313 9.15497
R16410 DVSS.n2313 DVSS.n2312 9.15497
R16411 DVSS.n2318 DVSS.n2317 9.15497
R16412 DVSS.n2317 DVSS.n2316 9.15497
R16413 DVSS.n2322 DVSS.n2321 9.15497
R16414 DVSS.n2321 DVSS.n2320 9.15497
R16415 DVSS.n2326 DVSS.n2325 9.15497
R16416 DVSS.n2325 DVSS.n2324 9.15497
R16417 DVSS.n2330 DVSS.n2329 9.15497
R16418 DVSS.n2329 DVSS.n2328 9.15497
R16419 DVSS.n2334 DVSS.n2333 9.15497
R16420 DVSS.n2333 DVSS.n2332 9.15497
R16421 DVSS.n1801 DVSS.n1800 9.15497
R16422 DVSS.n1800 DVSS.n1799 9.15497
R16423 DVSS.n2522 DVSS.n2521 9.15497
R16424 DVSS.n2521 DVSS.n2520 9.15497
R16425 DVSS.n2528 DVSS.n2527 9.15497
R16426 DVSS.n2527 DVSS.n2526 9.15497
R16427 DVSS.n2533 DVSS.n2532 9.15497
R16428 DVSS.n2532 DVSS.n2531 9.15497
R16429 DVSS.n2537 DVSS.n2536 9.15497
R16430 DVSS.n2536 DVSS.n2535 9.15497
R16431 DVSS.n2542 DVSS.n2541 9.15497
R16432 DVSS.n2543 DVSS.n2542 9.15497
R16433 DVSS.n1210 DVSS.n1209 9.15497
R16434 DVSS.n1209 DVSS.n1208 9.15497
R16435 DVSS.n1684 DVSS.n1683 9.15497
R16436 DVSS.n1682 DVSS.n1681 9.15497
R16437 DVSS.n1681 DVSS.n1680 9.15497
R16438 DVSS.n1689 DVSS.n1688 9.15497
R16439 DVSS.n1688 DVSS.n1687 9.15497
R16440 DVSS.n1696 DVSS.n1695 9.15497
R16441 DVSS.n1695 DVSS.n1694 9.15497
R16442 DVSS.n1700 DVSS.n1699 9.15497
R16443 DVSS.n1699 DVSS.n1698 9.15497
R16444 DVSS.n1704 DVSS.n1703 9.15497
R16445 DVSS.n1703 DVSS.n1702 9.15497
R16446 DVSS.n1708 DVSS.n1707 9.15497
R16447 DVSS.n1707 DVSS.n1706 9.15497
R16448 DVSS.n1712 DVSS.n1711 9.15497
R16449 DVSS.n1711 DVSS.n1710 9.15497
R16450 DVSS.n1716 DVSS.n1715 9.15497
R16451 DVSS.n1715 DVSS.n1714 9.15497
R16452 DVSS.n1071 DVSS.n1070 9.15497
R16453 DVSS.n1069 DVSS.n1068 9.15497
R16454 DVSS.n1068 DVSS.n1067 9.15497
R16455 DVSS.n1076 DVSS.n1075 9.15497
R16456 DVSS.n1075 DVSS.n1074 9.15497
R16457 DVSS.n1083 DVSS.n1082 9.15497
R16458 DVSS.n1082 DVSS.n1081 9.15497
R16459 DVSS.n1087 DVSS.n1086 9.15497
R16460 DVSS.n1086 DVSS.n1085 9.15497
R16461 DVSS.n1091 DVSS.n1090 9.15497
R16462 DVSS.n1090 DVSS.n1089 9.15497
R16463 DVSS.n1095 DVSS.n1094 9.15497
R16464 DVSS.n1094 DVSS.n1093 9.15497
R16465 DVSS.n1099 DVSS.n1098 9.15497
R16466 DVSS.n1098 DVSS.n1097 9.15497
R16467 DVSS.n1103 DVSS.n1102 9.15497
R16468 DVSS.n1102 DVSS.n1101 9.15497
R16469 DVSS.n591 DVSS.n590 9.15497
R16470 DVSS.n1107 DVSS.n1106 9.15497
R16471 DVSS.n1106 DVSS.n1105 9.15497
R16472 DVSS.n1112 DVSS.n1111 9.15497
R16473 DVSS.n1111 DVSS.n1110 9.15497
R16474 DVSS.n1117 DVSS.n1116 9.15497
R16475 DVSS.n1116 DVSS.n1115 9.15497
R16476 DVSS.n1124 DVSS.n1123 9.15497
R16477 DVSS.n1123 DVSS.n1122 9.15497
R16478 DVSS.n1128 DVSS.n1127 9.15497
R16479 DVSS.n1127 DVSS.n1126 9.15497
R16480 DVSS.n1133 DVSS.n1132 9.15497
R16481 DVSS.n1132 DVSS.n1131 9.15497
R16482 DVSS.n1141 DVSS.n1140 9.15497
R16483 DVSS.n1140 DVSS.n1139 9.15497
R16484 DVSS.n1145 DVSS.n1144 9.15497
R16485 DVSS.n1144 DVSS.n1143 9.15497
R16486 DVSS.n1152 DVSS.n1151 9.15497
R16487 DVSS.n1151 DVSS.n1150 9.15497
R16488 DVSS.n1160 DVSS.n1159 9.15497
R16489 DVSS.n1159 DVSS.n1158 9.15497
R16490 DVSS.n1163 DVSS.n1162 9.15497
R16491 DVSS.n1168 DVSS.n1167 9.15497
R16492 DVSS.n2662 DVSS.n2661 9.15497
R16493 DVSS.n2664 DVSS.n2662 9.15497
R16494 DVSS.n2656 DVSS.n2655 9.15497
R16495 DVSS.n2655 DVSS.n2654 9.15497
R16496 DVSS.n2652 DVSS.n2651 9.15497
R16497 DVSS.n2651 DVSS.n2650 9.15497
R16498 DVSS.n2647 DVSS.n2646 9.15497
R16499 DVSS.n2646 DVSS.n2645 9.15497
R16500 DVSS.n2642 DVSS.n2641 9.15497
R16501 DVSS.n2641 DVSS.n2640 9.15497
R16502 DVSS.n2547 DVSS.n2546 9.15497
R16503 DVSS.n2546 DVSS.n2545 9.15497
R16504 DVSS.n2551 DVSS.n2550 9.15497
R16505 DVSS.n2550 DVSS.n2549 9.15497
R16506 DVSS.n2555 DVSS.n2554 9.15497
R16507 DVSS.n2554 DVSS.n2553 9.15497
R16508 DVSS.n2559 DVSS.n2558 9.15497
R16509 DVSS.n2558 DVSS.n2557 9.15497
R16510 DVSS.n2563 DVSS.n2562 9.15497
R16511 DVSS.n2562 DVSS.n2561 9.15497
R16512 DVSS.n2569 DVSS.n2568 9.15497
R16513 DVSS.n2568 DVSS.n2567 9.15497
R16514 DVSS.n2574 DVSS.n2573 9.15497
R16515 DVSS.n2573 DVSS.n2572 9.15497
R16516 DVSS.n2578 DVSS.n2577 9.15497
R16517 DVSS.n2577 DVSS.n2576 9.15497
R16518 DVSS.n2582 DVSS.n2581 9.15497
R16519 DVSS.n2581 DVSS.n2580 9.15497
R16520 DVSS.n2588 DVSS.n2587 9.15497
R16521 DVSS.n2594 DVSS.n2593 9.15497
R16522 DVSS.n2593 DVSS.n2592 9.15497
R16523 DVSS.n2598 DVSS.n2597 9.15497
R16524 DVSS.n2597 DVSS.n2596 9.15497
R16525 DVSS.n2603 DVSS.n2602 9.15497
R16526 DVSS.n2611 DVSS.n2610 9.15497
R16527 DVSS.n2610 DVSS.n2609 9.15497
R16528 DVSS.n2615 DVSS.n2614 9.15497
R16529 DVSS.n2614 DVSS.n2613 9.15497
R16530 DVSS.n2620 DVSS.n2619 9.15497
R16531 DVSS.n2625 DVSS.n2624 9.15497
R16532 DVSS.n2624 DVSS.n2623 9.15497
R16533 DVSS.n2629 DVSS.n2628 9.15497
R16534 DVSS.n2628 DVSS.n2627 9.15497
R16535 DVSS.n2633 DVSS.n2632 9.15497
R16536 DVSS.n2632 DVSS.n2631 9.15497
R16537 DVSS.n2638 DVSS.n2637 9.15497
R16538 DVSS.n2639 DVSS.n2638 9.15497
R16539 DVSS.n1720 DVSS.n1719 9.15497
R16540 DVSS.n1719 DVSS.n1718 9.15497
R16541 DVSS.n1725 DVSS.n1724 9.15497
R16542 DVSS.n1724 DVSS.n1723 9.15497
R16543 DVSS.n1730 DVSS.n1729 9.15497
R16544 DVSS.n1729 DVSS.n1728 9.15497
R16545 DVSS.n1737 DVSS.n1736 9.15497
R16546 DVSS.n1736 DVSS.n1735 9.15497
R16547 DVSS.n1741 DVSS.n1740 9.15497
R16548 DVSS.n1740 DVSS.n1739 9.15497
R16549 DVSS.n1746 DVSS.n1745 9.15497
R16550 DVSS.n1745 DVSS.n1744 9.15497
R16551 DVSS.n1754 DVSS.n1753 9.15497
R16552 DVSS.n1753 DVSS.n1752 9.15497
R16553 DVSS.n1758 DVSS.n1757 9.15497
R16554 DVSS.n1757 DVSS.n1756 9.15497
R16555 DVSS.n1765 DVSS.n1764 9.15497
R16556 DVSS.n1764 DVSS.n1763 9.15497
R16557 DVSS.n1771 DVSS.n1770 9.15497
R16558 DVSS.n1770 DVSS.n1769 9.15497
R16559 DVSS.n1776 DVSS.n1775 9.15497
R16560 DVSS.n1777 DVSS.n1776 9.15497
R16561 DVSS.n1782 DVSS.n1781 9.15497
R16562 DVSS.n1806 DVSS.n1805 9.15497
R16563 DVSS.n1805 DVSS.n1804 9.15497
R16564 DVSS.n1811 DVSS.n1810 9.15497
R16565 DVSS.n1810 DVSS.n1809 9.15497
R16566 DVSS.n1816 DVSS.n1815 9.15497
R16567 DVSS.n1815 DVSS.n1814 9.15497
R16568 DVSS.n1820 DVSS.n1819 9.15497
R16569 DVSS.n1819 DVSS.n1818 9.15497
R16570 DVSS.n1205 DVSS.n1204 9.15497
R16571 DVSS.n1204 DVSS.n1203 9.15497
R16572 DVSS.n2517 DVSS.n2516 9.15497
R16573 DVSS.n2518 DVSS.n2517 9.15497
R16574 DVSS.n1827 DVSS.n1826 9.15497
R16575 DVSS.n1826 DVSS.n1825 9.15497
R16576 DVSS.n2511 DVSS.n2510 9.15497
R16577 DVSS.n2510 DVSS.n2509 9.15497
R16578 DVSS.n2507 DVSS.n2506 9.15497
R16579 DVSS.n2506 DVSS.n2505 9.15497
R16580 DVSS.n2500 DVSS.n2499 9.15497
R16581 DVSS.n2495 DVSS.n2494 9.15497
R16582 DVSS.n2494 DVSS.n2493 9.15497
R16583 DVSS.n2491 DVSS.n2490 9.15497
R16584 DVSS.n2490 DVSS.n2489 9.15497
R16585 DVSS.n2483 DVSS.n2482 9.15497
R16586 DVSS.n2478 DVSS.n2477 9.15497
R16587 DVSS.n2477 DVSS.n2476 9.15497
R16588 DVSS.n2474 DVSS.n2473 9.15497
R16589 DVSS.n2473 DVSS.n2472 9.15497
R16590 DVSS.n2469 DVSS.n2468 9.15497
R16591 DVSS.n2463 DVSS.n2462 9.15497
R16592 DVSS.n2462 DVSS.n2461 9.15497
R16593 DVSS.n2459 DVSS.n2458 9.15497
R16594 DVSS.n2458 DVSS.n2457 9.15497
R16595 DVSS.n2455 DVSS.n2454 9.15497
R16596 DVSS.n2454 DVSS.n2453 9.15497
R16597 DVSS.n2450 DVSS.n2449 9.15497
R16598 DVSS.n2449 DVSS.n2448 9.15497
R16599 DVSS.n2444 DVSS.n2443 9.15497
R16600 DVSS.n2443 DVSS.n2442 9.15497
R16601 DVSS.n2440 DVSS.n2439 9.15497
R16602 DVSS.n2439 DVSS.n2438 9.15497
R16603 DVSS.n2436 DVSS.n2435 9.15497
R16604 DVSS.n2435 DVSS.n2434 9.15497
R16605 DVSS.n2433 DVSS.n2432 9.15497
R16606 DVSS.n2432 DVSS.n2431 9.15497
R16607 DVSS.n2428 DVSS.n2427 9.15497
R16608 DVSS.n2427 DVSS.n2426 9.15497
R16609 DVSS.n2422 DVSS.n2421 9.15497
R16610 DVSS.n2421 DVSS.n2420 9.15497
R16611 DVSS.n2414 DVSS.n2413 9.15497
R16612 DVSS.n2413 DVSS.n2412 9.15497
R16613 DVSS.n2404 DVSS.n2403 9.15497
R16614 DVSS.n2403 DVSS.n2402 9.15497
R16615 DVSS.n2338 DVSS.n2337 9.15497
R16616 DVSS.n2337 DVSS.n2336 9.15497
R16617 DVSS.n2343 DVSS.n2342 9.15497
R16618 DVSS.n2342 DVSS.n2341 9.15497
R16619 DVSS.n2348 DVSS.n2347 9.15497
R16620 DVSS.n2347 DVSS.n2346 9.15497
R16621 DVSS.n2355 DVSS.n2354 9.15497
R16622 DVSS.n2354 DVSS.n2353 9.15497
R16623 DVSS.n2359 DVSS.n2358 9.15497
R16624 DVSS.n2358 DVSS.n2357 9.15497
R16625 DVSS.n2364 DVSS.n2363 9.15497
R16626 DVSS.n2372 DVSS.n2371 9.15497
R16627 DVSS.n2376 DVSS.n2375 9.15497
R16628 DVSS.n2380 DVSS.n2379 9.15497
R16629 DVSS.n2379 DVSS.n2378 9.15497
R16630 DVSS.n2386 DVSS.n2385 9.15497
R16631 DVSS.n2385 DVSS.n2384 9.15497
R16632 DVSS.n2390 DVSS.n2389 9.15497
R16633 DVSS.n2389 DVSS.n2388 9.15497
R16634 DVSS.n2396 DVSS.n2395 9.15497
R16635 DVSS.n2395 DVSS.n2394 9.15497
R16636 DVSS.n524 DVSS.n523 9.15497
R16637 DVSS.n523 DVSS.n522 9.15497
R16638 DVSS.n521 DVSS.n520 9.15497
R16639 DVSS.n528 DVSS.n527 9.15497
R16640 DVSS.n519 DVSS.n518 9.15497
R16641 DVSS.n515 DVSS.n514 9.15497
R16642 DVSS.n512 DVSS.n511 9.15497
R16643 DVSS.n508 DVSS.n507 9.15497
R16644 DVSS.n505 DVSS.n504 9.15497
R16645 DVSS.n499 DVSS.n498 9.15497
R16646 DVSS.n495 DVSS.n494 9.15497
R16647 DVSS.n491 DVSS.n490 9.15497
R16648 DVSS.n488 DVSS.n487 9.15497
R16649 DVSS.n2784 DVSS.n2783 9.15497
R16650 DVSS.n2787 DVSS.n2786 9.15497
R16651 DVSS.n535 DVSS.n534 9.15497
R16652 DVSS.n533 DVSS.n532 9.15497
R16653 DVSS.n2842 DVSS.n2841 9.15497
R16654 DVSS.n2840 DVSS.n2839 9.15497
R16655 DVSS.n2849 DVSS.n2848 9.15497
R16656 DVSS.n2846 DVSS.n2845 9.15497
R16657 DVSS.n2854 DVSS.n2853 9.15497
R16658 DVSS.n2852 DVSS.n2851 9.15497
R16659 DVSS.n2837 DVSS.n2836 9.15497
R16660 DVSS.n2809 DVSS.n2808 9.15497
R16661 DVSS.n2817 DVSS.n2816 9.15497
R16662 DVSS.n2820 DVSS.n2819 9.15497
R16663 DVSS.n2824 DVSS.n2823 9.15497
R16664 DVSS.n2830 DVSS.n2829 9.15497
R16665 DVSS.n2834 DVSS.n2833 9.15497
R16666 DVSS.n2795 DVSS.n2794 9.15497
R16667 DVSS.n2799 DVSS.n2798 9.15497
R16668 DVSS.n2871 DVSS.n2870 9.15497
R16669 DVSS.n480 DVSS.n479 9.15497
R16670 DVSS.n479 DVSS.n478 9.15497
R16671 DVSS.n2876 DVSS.n2875 9.15497
R16672 DVSS.n2875 DVSS.n2874 9.15497
R16673 DVSS.n2883 DVSS.n2882 9.15497
R16674 DVSS.n2882 DVSS.n2881 9.15497
R16675 DVSS.n2887 DVSS.n2886 9.15497
R16676 DVSS.n2886 DVSS.n2885 9.15497
R16677 DVSS.n2891 DVSS.n2890 9.15497
R16678 DVSS.n2890 DVSS.n2889 9.15497
R16679 DVSS.n2895 DVSS.n2894 9.15497
R16680 DVSS.n2894 DVSS.n2893 9.15497
R16681 DVSS.n2899 DVSS.n2898 9.15497
R16682 DVSS.n2898 DVSS.n2897 9.15497
R16683 DVSS.n2903 DVSS.n2902 9.15497
R16684 DVSS.n2902 DVSS.n2901 9.15497
R16685 DVSS.n2975 DVSS.n2974 9.15497
R16686 DVSS.n2974 DVSS.n2973 9.15497
R16687 DVSS.n2907 DVSS.n2906 9.15497
R16688 DVSS.n2906 DVSS.n2905 9.15497
R16689 DVSS.n2912 DVSS.n2911 9.15497
R16690 DVSS.n2911 DVSS.n2910 9.15497
R16691 DVSS.n2917 DVSS.n2916 9.15497
R16692 DVSS.n2916 DVSS.n2915 9.15497
R16693 DVSS.n2924 DVSS.n2923 9.15497
R16694 DVSS.n2923 DVSS.n2922 9.15497
R16695 DVSS.n2928 DVSS.n2927 9.15497
R16696 DVSS.n2927 DVSS.n2926 9.15497
R16697 DVSS.n2933 DVSS.n2932 9.15497
R16698 DVSS.n2941 DVSS.n2940 9.15497
R16699 DVSS.n2945 DVSS.n2944 9.15497
R16700 DVSS.n2949 DVSS.n2948 9.15497
R16701 DVSS.n2948 DVSS.n2947 9.15497
R16702 DVSS.n2955 DVSS.n2954 9.15497
R16703 DVSS.n2954 DVSS.n2953 9.15497
R16704 DVSS.n2959 DVSS.n2958 9.15497
R16705 DVSS.n2958 DVSS.n2957 9.15497
R16706 DVSS.n2965 DVSS.n2964 9.15497
R16707 DVSS.n2964 DVSS.n2963 9.15497
R16708 DVSS.n564 DVSS.n563 9.15497
R16709 DVSS.n563 DVSS.n562 9.15497
R16710 DVSS.n556 DVSS.n555 9.15497
R16711 DVSS.n555 DVSS.n554 9.15497
R16712 DVSS.n541 DVSS.n540 9.15497
R16713 DVSS.n540 DVSS.n539 9.15497
R16714 DVSS.n11 DVSS.n10 9.15497
R16715 DVSS.n10 DVSS.n9 9.15497
R16716 DVSS.n3088 DVSS.n3087 9.15497
R16717 DVSS.n3089 DVSS.n3088 9.15497
R16718 DVSS.n2999 DVSS.n2998 9.15497
R16719 DVSS.n2998 DVSS.n2997 9.15497
R16720 DVSS.n3002 DVSS.n3001 9.15497
R16721 DVSS.n3001 DVSS.n3000 9.15497
R16722 DVSS.n3006 DVSS.n3005 9.15497
R16723 DVSS.n3005 DVSS.n3004 9.15497
R16724 DVSS.n3010 DVSS.n3009 9.15497
R16725 DVSS.n3009 DVSS.n3008 9.15497
R16726 DVSS.n3019 DVSS.n3018 9.15497
R16727 DVSS.n3018 DVSS.n3017 9.15497
R16728 DVSS.n3024 DVSS.n3023 9.15497
R16729 DVSS.n3023 DVSS.n3022 9.15497
R16730 DVSS.n3028 DVSS.n3027 9.15497
R16731 DVSS.n3027 DVSS.n3026 9.15497
R16732 DVSS.n3032 DVSS.n3031 9.15497
R16733 DVSS.n3031 DVSS.n3030 9.15497
R16734 DVSS.n3038 DVSS.n3037 9.15497
R16735 DVSS.n3044 DVSS.n3043 9.15497
R16736 DVSS.n3043 DVSS.n3042 9.15497
R16737 DVSS.n3048 DVSS.n3047 9.15497
R16738 DVSS.n3047 DVSS.n3046 9.15497
R16739 DVSS.n3053 DVSS.n3052 9.15497
R16740 DVSS.n3061 DVSS.n3060 9.15497
R16741 DVSS.n3060 DVSS.n3059 9.15497
R16742 DVSS.n3065 DVSS.n3064 9.15497
R16743 DVSS.n3064 DVSS.n3063 9.15497
R16744 DVSS.n3070 DVSS.n3069 9.15497
R16745 DVSS.n3075 DVSS.n3074 9.15497
R16746 DVSS.n3074 DVSS.n3073 9.15497
R16747 DVSS.n3079 DVSS.n3078 9.15497
R16748 DVSS.n3078 DVSS.n3077 9.15497
R16749 DVSS.n3083 DVSS.n3082 9.15497
R16750 DVSS.n3082 DVSS.n3081 9.15497
R16751 DVSS.n2987 DVSS.n2986 9.15497
R16752 DVSS.n2986 DVSS.n2985 9.15497
R16753 DVSS.n2993 DVSS.n2992 9.15497
R16754 DVSS.n2992 DVSS.n2991 9.15497
R16755 DVSS.n569 DVSS.n568 9.15497
R16756 DVSS.n568 DVSS.n567 9.15497
R16757 DVSS.n574 DVSS.n573 9.15497
R16758 DVSS.n573 DVSS.n572 9.15497
R16759 DVSS.n578 DVSS.n577 9.15497
R16760 DVSS.n577 DVSS.n576 9.15497
R16761 DVSS.n2755 DVSS.n2754 9.15497
R16762 DVSS.n2756 DVSS.n2755 9.15497
R16763 DVSS.n2750 DVSS.n2749 9.15497
R16764 DVSS.n2749 DVSS.n559 9.15497
R16765 DVSS.n2747 DVSS.n2746 9.15497
R16766 DVSS.n2746 DVSS.n2745 9.15497
R16767 DVSS.n2743 DVSS.n2742 9.15497
R16768 DVSS.n2742 DVSS.n2741 9.15497
R16769 DVSS.n2739 DVSS.n2738 9.15497
R16770 DVSS.n2738 DVSS.n2737 9.15497
R16771 DVSS.n2734 DVSS.n2733 9.15497
R16772 DVSS.n2729 DVSS.n2728 9.15497
R16773 DVSS.n2728 DVSS.n2727 9.15497
R16774 DVSS.n2725 DVSS.n2724 9.15497
R16775 DVSS.n2724 DVSS.n2723 9.15497
R16776 DVSS.n2717 DVSS.n2716 9.15497
R16777 DVSS.n2712 DVSS.n2711 9.15497
R16778 DVSS.n2711 DVSS.n2710 9.15497
R16779 DVSS.n2708 DVSS.n2707 9.15497
R16780 DVSS.n2707 DVSS.n2706 9.15497
R16781 DVSS.n2702 DVSS.n2701 9.15497
R16782 DVSS.n2701 DVSS.n2700 9.15497
R16783 DVSS.n2696 DVSS.n2695 9.15497
R16784 DVSS.n2695 DVSS.n2694 9.15497
R16785 DVSS.n2692 DVSS.n2691 9.15497
R16786 DVSS.n2691 DVSS.n2690 9.15497
R16787 DVSS.n2688 DVSS.n2687 9.15497
R16788 DVSS.n2687 DVSS.n2686 9.15497
R16789 DVSS.n2683 DVSS.n2682 9.15497
R16790 DVSS.n2682 DVSS.n2681 9.15497
R16791 DVSS.n2677 DVSS.n2676 9.15497
R16792 DVSS.n2676 DVSS.n2675 9.15497
R16793 DVSS.n2673 DVSS.n2672 9.15497
R16794 DVSS.n2672 DVSS.n2671 9.15497
R16795 DVSS.n2669 DVSS.n588 9.15497
R16796 DVSS.n588 DVSS.n587 9.15497
R16797 DVSS.n2668 DVSS.n2667 9.15497
R16798 DVSS.n2667 DVSS.n2666 9.15497
R16799 DVSS.n596 DVSS.n595 9.15497
R16800 DVSS.n1187 DVSS.n1186 9.15497
R16801 DVSS.n1186 DVSS.n1185 9.15497
R16802 DVSS.n2774 DVSS.n2773 9.15497
R16803 DVSS.n2773 DVSS.n2772 9.15497
R16804 DVSS.n2770 DVSS.n2769 9.15497
R16805 DVSS.n2769 DVSS.n2768 9.15497
R16806 DVSS.n2765 DVSS.n2764 9.15497
R16807 DVSS.n2764 DVSS.n2763 9.15497
R16808 DVSS.n2760 DVSS.n2759 9.15497
R16809 DVSS.n2759 DVSS.n2758 9.15497
R16810 DVSS.n551 DVSS.n550 9.15497
R16811 DVSS.n550 DVSS.n549 9.15497
R16812 DVSS.n547 DVSS.n546 9.15497
R16813 DVSS.n546 DVSS.n545 9.15497
R16814 DVSS.n2 DVSS.n1 9.15497
R16815 DVSS.n1 DVSS.n0 9.15497
R16816 DVSS.n3093 DVSS.n3092 9.15497
R16817 DVSS.n3092 DVSS.n3091 9.15497
R16818 DVSS.n2291 DVSS.n1838 9.01392
R16819 DVSS.n1846 DVSS.n1837 9.01392
R16820 DVSS.n2283 DVSS.n2282 9.01392
R16821 DVSS.n1844 DVSS.n1843 9.01392
R16822 DVSS.n2252 DVSS.n2251 9.01392
R16823 DVSS.n1854 DVSS.n1852 9.01392
R16824 DVSS.n1864 DVSS.n1863 9.01392
R16825 DVSS.n2212 DVSS.n2211 9.01392
R16826 DVSS.n1870 DVSS.n1862 9.01392
R16827 DVSS.n2204 DVSS.n2203 9.01392
R16828 DVSS.n2191 DVSS.n2190 9.01392
R16829 DVSS.n1902 DVSS.n1901 9.01392
R16830 DVSS.n2184 DVSS.n2183 9.01392
R16831 DVSS.n1907 DVSS.n1906 9.01392
R16832 DVSS.n1673 DVSS.n1220 9.01392
R16833 DVSS.n1228 DVSS.n1219 9.01392
R16834 DVSS.n1665 DVSS.n1664 9.01392
R16835 DVSS.n1226 DVSS.n1225 9.01392
R16836 DVSS.n1634 DVSS.n1633 9.01392
R16837 DVSS.n1236 DVSS.n1234 9.01392
R16838 DVSS.n1246 DVSS.n1245 9.01392
R16839 DVSS.n1594 DVSS.n1593 9.01392
R16840 DVSS.n1252 DVSS.n1244 9.01392
R16841 DVSS.n1586 DVSS.n1585 9.01392
R16842 DVSS.n1573 DVSS.n1572 9.01392
R16843 DVSS.n1284 DVSS.n1283 9.01392
R16844 DVSS.n1566 DVSS.n1565 9.01392
R16845 DVSS.n1289 DVSS.n1288 9.01392
R16846 DVSS.n1060 DVSS.n607 9.01392
R16847 DVSS.n615 DVSS.n606 9.01392
R16848 DVSS.n1052 DVSS.n1051 9.01392
R16849 DVSS.n613 DVSS.n612 9.01392
R16850 DVSS.n1021 DVSS.n1020 9.01392
R16851 DVSS.n623 DVSS.n621 9.01392
R16852 DVSS.n633 DVSS.n632 9.01392
R16853 DVSS.n981 DVSS.n980 9.01392
R16854 DVSS.n639 DVSS.n631 9.01392
R16855 DVSS.n973 DVSS.n972 9.01392
R16856 DVSS.n960 DVSS.n959 9.01392
R16857 DVSS.n671 DVSS.n670 9.01392
R16858 DVSS.n953 DVSS.n952 9.01392
R16859 DVSS.n676 DVSS.n675 9.01392
R16860 DVSS.n471 DVSS.n18 9.01392
R16861 DVSS.n26 DVSS.n17 9.01392
R16862 DVSS.n463 DVSS.n462 9.01392
R16863 DVSS.n24 DVSS.n23 9.01392
R16864 DVSS.n432 DVSS.n431 9.01392
R16865 DVSS.n34 DVSS.n32 9.01392
R16866 DVSS.n44 DVSS.n43 9.01392
R16867 DVSS.n392 DVSS.n391 9.01392
R16868 DVSS.n50 DVSS.n42 9.01392
R16869 DVSS.n384 DVSS.n383 9.01392
R16870 DVSS.n371 DVSS.n370 9.01392
R16871 DVSS.n82 DVSS.n81 9.01392
R16872 DVSS.n364 DVSS.n363 9.01392
R16873 DVSS.n87 DVSS.n86 9.01392
R16874 DVSS.n2175 DVSS.n1907 9.01392
R16875 DVSS.n2183 DVSS.n2182 9.01392
R16876 DVSS.n2178 DVSS.n1901 9.01392
R16877 DVSS.n2192 DVSS.n2191 9.01392
R16878 DVSS.n2203 DVSS.n2202 9.01392
R16879 DVSS.n2197 DVSS.n1862 9.01392
R16880 DVSS.n2213 DVSS.n2212 9.01392
R16881 DVSS.n1863 DVSS.n1859 9.01392
R16882 DVSS.n2220 DVSS.n1854 9.01392
R16883 DVSS.n2251 DVSS.n2250 9.01392
R16884 DVSS.n2246 DVSS.n1843 9.01392
R16885 DVSS.n2284 DVSS.n2283 9.01392
R16886 DVSS.n2286 DVSS.n1837 9.01392
R16887 DVSS.n2291 DVSS.n2290 9.01392
R16888 DVSS.n1557 DVSS.n1289 9.01392
R16889 DVSS.n1565 DVSS.n1564 9.01392
R16890 DVSS.n1560 DVSS.n1283 9.01392
R16891 DVSS.n1574 DVSS.n1573 9.01392
R16892 DVSS.n1585 DVSS.n1584 9.01392
R16893 DVSS.n1579 DVSS.n1244 9.01392
R16894 DVSS.n1595 DVSS.n1594 9.01392
R16895 DVSS.n1245 DVSS.n1241 9.01392
R16896 DVSS.n1602 DVSS.n1236 9.01392
R16897 DVSS.n1633 DVSS.n1632 9.01392
R16898 DVSS.n1628 DVSS.n1225 9.01392
R16899 DVSS.n1666 DVSS.n1665 9.01392
R16900 DVSS.n1668 DVSS.n1219 9.01392
R16901 DVSS.n1673 DVSS.n1672 9.01392
R16902 DVSS.n944 DVSS.n676 9.01392
R16903 DVSS.n952 DVSS.n951 9.01392
R16904 DVSS.n947 DVSS.n670 9.01392
R16905 DVSS.n961 DVSS.n960 9.01392
R16906 DVSS.n972 DVSS.n971 9.01392
R16907 DVSS.n966 DVSS.n631 9.01392
R16908 DVSS.n982 DVSS.n981 9.01392
R16909 DVSS.n632 DVSS.n628 9.01392
R16910 DVSS.n989 DVSS.n623 9.01392
R16911 DVSS.n1020 DVSS.n1019 9.01392
R16912 DVSS.n1015 DVSS.n612 9.01392
R16913 DVSS.n1053 DVSS.n1052 9.01392
R16914 DVSS.n1055 DVSS.n606 9.01392
R16915 DVSS.n1060 DVSS.n1059 9.01392
R16916 DVSS.n355 DVSS.n87 9.01392
R16917 DVSS.n363 DVSS.n362 9.01392
R16918 DVSS.n358 DVSS.n81 9.01392
R16919 DVSS.n372 DVSS.n371 9.01392
R16920 DVSS.n383 DVSS.n382 9.01392
R16921 DVSS.n377 DVSS.n42 9.01392
R16922 DVSS.n393 DVSS.n392 9.01392
R16923 DVSS.n43 DVSS.n39 9.01392
R16924 DVSS.n400 DVSS.n34 9.01392
R16925 DVSS.n431 DVSS.n430 9.01392
R16926 DVSS.n426 DVSS.n23 9.01392
R16927 DVSS.n464 DVSS.n463 9.01392
R16928 DVSS.n466 DVSS.n17 9.01392
R16929 DVSS.n471 DVSS.n470 9.01392
R16930 DVSS.n536 DVSS.n533 8.99329
R16931 DVSS.n2855 DVSS.n2854 8.99094
R16932 DVSS.n2850 DVSS.n2849 8.99094
R16933 DVSS.n2843 DVSS.n2842 8.99094
R16934 DVSS.n2843 DVSS.n2840 8.99094
R16935 DVSS.n2850 DVSS.n2846 8.99094
R16936 DVSS.n2855 DVSS.n2852 8.99094
R16937 DVSS.n2133 DVSS.n2125 8.9737
R16938 DVSS.n1515 DVSS.n1507 8.9737
R16939 DVSS.n902 DVSS.n894 8.9737
R16940 DVSS.n313 DVSS.n305 8.9737
R16941 DVSS.n2173 DVSS.n1936 8.8706
R16942 DVSS.n1555 DVSS.n1318 8.8706
R16943 DVSS.n942 DVSS.n705 8.8706
R16944 DVSS.n353 DVSS.n116 8.8706
R16945 DVSS.n529 DVSS.n528 8.85539
R16946 DVSS.n529 DVSS.n519 8.85536
R16947 DVSS.n2838 DVSS.n2834 8.85488
R16948 DVSS.n2831 DVSS.n2824 8.85488
R16949 DVSS.n2821 DVSS.n2817 8.85488
R16950 DVSS.n516 DVSS.n512 8.85488
R16951 DVSS.n509 DVSS.n505 8.85488
R16952 DVSS.n500 DVSS.n495 8.85488
R16953 DVSS.n492 DVSS.n488 8.85488
R16954 DVSS.n2786 DVSS.n2785 8.85488
R16955 DVSS.n516 DVSS.n515 8.85488
R16956 DVSS.n509 DVSS.n508 8.85488
R16957 DVSS.n500 DVSS.n499 8.85488
R16958 DVSS.n492 DVSS.n491 8.85488
R16959 DVSS.n2785 DVSS.n2784 8.85488
R16960 DVSS.n2838 DVSS.n2837 8.85488
R16961 DVSS.n2810 DVSS.n2809 8.85488
R16962 DVSS.n2821 DVSS.n2820 8.85488
R16963 DVSS.n2831 DVSS.n2830 8.85488
R16964 DVSS.n536 DVSS.n535 8.85257
R16965 DVSS.n2794 DVSS.n2793 8.85257
R16966 DVSS.n2110 DVSS.n2109 8.15208
R16967 DVSS.n1492 DVSS.n1491 8.15208
R16968 DVSS.n879 DVSS.n878 8.15208
R16969 DVSS.n290 DVSS.n289 8.15208
R16970 DVSS.n1922 DVSS.n1921 7.5692
R16971 DVSS.n1931 DVSS.n1922 7.5692
R16972 DVSS.n1931 DVSS.n1930 7.5692
R16973 DVSS.n1930 DVSS.n1928 7.5692
R16974 DVSS.n1928 DVSS.n1926 7.5692
R16975 DVSS.n1926 DVSS.n1924 7.5692
R16976 DVSS.n1924 DVSS.n1911 7.5692
R16977 DVSS.n1936 DVSS.n1911 7.5692
R16978 DVSS.n2262 DVSS.n2257 7.5692
R16979 DVSS.n2271 DVSS.n2262 7.5692
R16980 DVSS.n2271 DVSS.n2270 7.5692
R16981 DVSS.n2270 DVSS.n2269 7.5692
R16982 DVSS.n2269 DVSS.n2266 7.5692
R16983 DVSS.n2266 DVSS.n2265 7.5692
R16984 DVSS.n2265 DVSS.n1835 7.5692
R16985 DVSS.n2293 DVSS.n1835 7.5692
R16986 DVSS.n1304 DVSS.n1303 7.5692
R16987 DVSS.n1313 DVSS.n1304 7.5692
R16988 DVSS.n1313 DVSS.n1312 7.5692
R16989 DVSS.n1312 DVSS.n1310 7.5692
R16990 DVSS.n1310 DVSS.n1308 7.5692
R16991 DVSS.n1308 DVSS.n1306 7.5692
R16992 DVSS.n1306 DVSS.n1293 7.5692
R16993 DVSS.n1318 DVSS.n1293 7.5692
R16994 DVSS.n1644 DVSS.n1639 7.5692
R16995 DVSS.n1653 DVSS.n1644 7.5692
R16996 DVSS.n1653 DVSS.n1652 7.5692
R16997 DVSS.n1652 DVSS.n1651 7.5692
R16998 DVSS.n1651 DVSS.n1648 7.5692
R16999 DVSS.n1648 DVSS.n1647 7.5692
R17000 DVSS.n1647 DVSS.n1217 7.5692
R17001 DVSS.n1675 DVSS.n1217 7.5692
R17002 DVSS.n691 DVSS.n690 7.5692
R17003 DVSS.n700 DVSS.n691 7.5692
R17004 DVSS.n700 DVSS.n699 7.5692
R17005 DVSS.n699 DVSS.n697 7.5692
R17006 DVSS.n697 DVSS.n695 7.5692
R17007 DVSS.n695 DVSS.n693 7.5692
R17008 DVSS.n693 DVSS.n680 7.5692
R17009 DVSS.n705 DVSS.n680 7.5692
R17010 DVSS.n1031 DVSS.n1026 7.5692
R17011 DVSS.n1040 DVSS.n1031 7.5692
R17012 DVSS.n1040 DVSS.n1039 7.5692
R17013 DVSS.n1039 DVSS.n1038 7.5692
R17014 DVSS.n1038 DVSS.n1035 7.5692
R17015 DVSS.n1035 DVSS.n1034 7.5692
R17016 DVSS.n1034 DVSS.n604 7.5692
R17017 DVSS.n1062 DVSS.n604 7.5692
R17018 DVSS.n102 DVSS.n101 7.5692
R17019 DVSS.n111 DVSS.n102 7.5692
R17020 DVSS.n111 DVSS.n110 7.5692
R17021 DVSS.n110 DVSS.n108 7.5692
R17022 DVSS.n108 DVSS.n106 7.5692
R17023 DVSS.n106 DVSS.n104 7.5692
R17024 DVSS.n104 DVSS.n91 7.5692
R17025 DVSS.n116 DVSS.n91 7.5692
R17026 DVSS.n442 DVSS.n437 7.5692
R17027 DVSS.n451 DVSS.n442 7.5692
R17028 DVSS.n451 DVSS.n450 7.5692
R17029 DVSS.n450 DVSS.n449 7.5692
R17030 DVSS.n449 DVSS.n446 7.5692
R17031 DVSS.n446 DVSS.n445 7.5692
R17032 DVSS.n445 DVSS.n15 7.5692
R17033 DVSS.n473 DVSS.n15 7.5692
R17034 DVSS.n2294 DVSS.n2293 7.1358
R17035 DVSS.n1676 DVSS.n1675 7.1358
R17036 DVSS.n1063 DVSS.n1062 7.1358
R17037 DVSS.n474 DVSS.n473 7.1358
R17038 DVSS.n2294 DVSS.n1834 6.65838
R17039 DVSS.n1676 DVSS.n1216 6.65838
R17040 DVSS.n1063 DVSS.n603 6.65838
R17041 DVSS.n474 DVSS.n14 6.65838
R17042 DVSS.n2137 DVSS.n2136 6.46787
R17043 DVSS.n1519 DVSS.n1518 6.46787
R17044 DVSS.n906 DVSS.n905 6.46787
R17045 DVSS.n317 DVSS.n316 6.46787
R17046 DVSS.n2089 DVSS.n2088 5.72682
R17047 DVSS.n2088 DVSS.n2087 5.72682
R17048 DVSS.n2087 DVSS.n2084 5.72682
R17049 DVSS.n2084 DVSS.n2083 5.72682
R17050 DVSS.n2083 DVSS.n2080 5.72682
R17051 DVSS.n2080 DVSS.n2079 5.72682
R17052 DVSS.n2079 DVSS.n2072 5.72682
R17053 DVSS.n2095 DVSS.n2072 5.72682
R17054 DVSS.n1471 DVSS.n1470 5.72682
R17055 DVSS.n1470 DVSS.n1469 5.72682
R17056 DVSS.n1469 DVSS.n1466 5.72682
R17057 DVSS.n1466 DVSS.n1465 5.72682
R17058 DVSS.n1465 DVSS.n1462 5.72682
R17059 DVSS.n1462 DVSS.n1461 5.72682
R17060 DVSS.n1461 DVSS.n1454 5.72682
R17061 DVSS.n1477 DVSS.n1454 5.72682
R17062 DVSS.n858 DVSS.n857 5.72682
R17063 DVSS.n857 DVSS.n856 5.72682
R17064 DVSS.n856 DVSS.n853 5.72682
R17065 DVSS.n853 DVSS.n852 5.72682
R17066 DVSS.n852 DVSS.n849 5.72682
R17067 DVSS.n849 DVSS.n848 5.72682
R17068 DVSS.n848 DVSS.n841 5.72682
R17069 DVSS.n864 DVSS.n841 5.72682
R17070 DVSS.n269 DVSS.n268 5.72682
R17071 DVSS.n268 DVSS.n267 5.72682
R17072 DVSS.n267 DVSS.n264 5.72682
R17073 DVSS.n264 DVSS.n263 5.72682
R17074 DVSS.n263 DVSS.n260 5.72682
R17075 DVSS.n260 DVSS.n259 5.72682
R17076 DVSS.n259 DVSS.n252 5.72682
R17077 DVSS.n275 DVSS.n252 5.72682
R17078 DVSS.n1974 DVSS.n1973 5.64756
R17079 DVSS.n1973 DVSS.n1963 5.64756
R17080 DVSS.n1953 DVSS.n1952 5.64756
R17081 DVSS.n1952 DVSS.n1942 5.64756
R17082 DVSS.n1356 DVSS.n1355 5.64756
R17083 DVSS.n1355 DVSS.n1345 5.64756
R17084 DVSS.n1335 DVSS.n1334 5.64756
R17085 DVSS.n1334 DVSS.n1324 5.64756
R17086 DVSS.n743 DVSS.n742 5.64756
R17087 DVSS.n742 DVSS.n732 5.64756
R17088 DVSS.n722 DVSS.n721 5.64756
R17089 DVSS.n721 DVSS.n711 5.64756
R17090 DVSS.n154 DVSS.n153 5.64756
R17091 DVSS.n153 DVSS.n143 5.64756
R17092 DVSS.n133 DVSS.n132 5.64756
R17093 DVSS.n132 DVSS.n122 5.64756
R17094 DVSS.n2202 DVSS.n1872 5.57999
R17095 DVSS.n2250 DVSS.n1857 5.57999
R17096 DVSS.n1584 DVSS.n1254 5.57999
R17097 DVSS.n1632 DVSS.n1239 5.57999
R17098 DVSS.n971 DVSS.n641 5.57999
R17099 DVSS.n1019 DVSS.n626 5.57999
R17100 DVSS.n382 DVSS.n52 5.57999
R17101 DVSS.n430 DVSS.n37 5.57999
R17102 DVSS.n2192 DVSS.n1900 5.34556
R17103 DVSS.n1574 DVSS.n1282 5.34556
R17104 DVSS.n961 DVSS.n669 5.34556
R17105 DVSS.n372 DVSS.n80 5.34556
R17106 DVSS.n2246 DVSS.n2245 5.29867
R17107 DVSS.n1628 DVSS.n1627 5.29867
R17108 DVSS.n1015 DVSS.n1014 5.29867
R17109 DVSS.n426 DVSS.n425 5.29867
R17110 DVSS.n1977 DVSS.n1960 4.89462
R17111 DVSS.n1956 DVSS.n1939 4.89462
R17112 DVSS.n1359 DVSS.n1342 4.89462
R17113 DVSS.n1338 DVSS.n1321 4.89462
R17114 DVSS.n746 DVSS.n729 4.89462
R17115 DVSS.n725 DVSS.n708 4.89462
R17116 DVSS.n157 DVSS.n140 4.89462
R17117 DVSS.n136 DVSS.n119 4.89462
R17118 DVSS.n2145 DVSS.n1999 4.74328
R17119 DVSS.n2040 DVSS.n2015 4.74328
R17120 DVSS.n1527 DVSS.n1381 4.74328
R17121 DVSS.n1422 DVSS.n1397 4.74328
R17122 DVSS.n914 DVSS.n768 4.74328
R17123 DVSS.n809 DVSS.n784 4.74328
R17124 DVSS.n325 DVSS.n179 4.74328
R17125 DVSS.n220 DVSS.n195 4.74328
R17126 DVSS.n2865 DVSS.n2864 4.72584
R17127 DVSS.n1751 DVSS.n1750 4.6505
R17128 DVSS.n1734 DVSS.n1733 4.6505
R17129 DVSS.n1693 DVSS.n1692 4.6505
R17130 DVSS.n2369 DVSS.n2368 4.6505
R17131 DVSS.n2352 DVSS.n2351 4.6505
R17132 DVSS.n2311 DVSS.n2310 4.6505
R17133 DVSS.n2308 DVSS.n2307 4.6505
R17134 DVSS.n2315 DVSS.n2314 4.6505
R17135 DVSS.n2319 DVSS.n2318 4.6505
R17136 DVSS.n2323 DVSS.n2322 4.6505
R17137 DVSS.n2327 DVSS.n2326 4.6505
R17138 DVSS.n2331 DVSS.n2330 4.6505
R17139 DVSS.n2335 DVSS.n2334 4.6505
R17140 DVSS.n2145 DVSS.n2144 4.6505
R17141 DVSS.n2165 DVSS.n2164 4.6505
R17142 DVSS.n2147 DVSS.n2146 4.6505
R17143 DVSS.n2150 DVSS.n1997 4.6505
R17144 DVSS.n2154 DVSS.n2153 4.6505
R17145 DVSS.n2156 DVSS.n2155 4.6505
R17146 DVSS.n1996 DVSS.n1993 4.6505
R17147 DVSS.n1981 DVSS.n1979 4.6505
R17148 DVSS.n2022 DVSS.n1958 4.6505
R17149 DVSS.n2053 DVSS.n2052 4.6505
R17150 DVSS.n2055 DVSS.n2054 4.6505
R17151 DVSS.n2039 DVSS.n2034 4.6505
R17152 DVSS.n2028 DVSS.n2024 4.6505
R17153 DVSS.n2063 DVSS.n2062 4.6505
R17154 DVSS.n2065 DVSS.n2064 4.6505
R17155 DVSS.n2041 DVSS.n2040 4.6505
R17156 DVSS.n2447 DVSS.n1831 4.6505
R17157 DVSS.n2471 DVSS.n1828 4.6505
R17158 DVSS.n2488 DVSS.n2487 4.6505
R17159 DVSS.n2504 DVSS.n2503 4.6505
R17160 DVSS.n2513 DVSS.n1827 4.6505
R17161 DVSS.n1807 DVSS.n1806 4.6505
R17162 DVSS.n1823 DVSS.n1822 4.6505
R17163 DVSS.n1823 DVSS.n1207 4.6505
R17164 DVSS.n1824 DVSS.n1823 4.6505
R17165 DVSS.n2524 DVSS.n2522 4.6505
R17166 DVSS.n2529 DVSS.n2528 4.6505
R17167 DVSS.n2534 DVSS.n2533 4.6505
R17168 DVSS.n2538 DVSS.n2537 4.6505
R17169 DVSS.n2541 DVSS.n2540 4.6505
R17170 DVSS.n2523 DVSS.n1202 4.6505
R17171 DVSS.n2530 DVSS.n1202 4.6505
R17172 DVSS.n2661 DVSS.n2660 4.6505
R17173 DVSS.n2649 DVSS.n1192 4.6505
R17174 DVSS.n2644 DVSS.n1192 4.6505
R17175 DVSS.n1193 DVSS.n1192 4.6505
R17176 DVSS.n2637 DVSS.n2636 4.6505
R17177 DVSS.n2566 DVSS.n1198 4.6505
R17178 DVSS.n2608 DVSS.n2607 4.6505
R17179 DVSS.n2591 DVSS.n2590 4.6505
R17180 DVSS.n2622 DVSS.n1195 4.6505
R17181 DVSS.n1527 DVSS.n1526 4.6505
R17182 DVSS.n1547 DVSS.n1546 4.6505
R17183 DVSS.n1529 DVSS.n1528 4.6505
R17184 DVSS.n1532 DVSS.n1379 4.6505
R17185 DVSS.n1536 DVSS.n1535 4.6505
R17186 DVSS.n1538 DVSS.n1537 4.6505
R17187 DVSS.n1378 DVSS.n1375 4.6505
R17188 DVSS.n1363 DVSS.n1361 4.6505
R17189 DVSS.n1404 DVSS.n1340 4.6505
R17190 DVSS.n1435 DVSS.n1434 4.6505
R17191 DVSS.n1437 DVSS.n1436 4.6505
R17192 DVSS.n1421 DVSS.n1416 4.6505
R17193 DVSS.n1410 DVSS.n1406 4.6505
R17194 DVSS.n1445 DVSS.n1444 4.6505
R17195 DVSS.n1447 DVSS.n1446 4.6505
R17196 DVSS.n1423 DVSS.n1422 4.6505
R17197 DVSS.n1690 DVSS.n1689 4.6505
R17198 DVSS.n1697 DVSS.n1696 4.6505
R17199 DVSS.n1701 DVSS.n1700 4.6505
R17200 DVSS.n1705 DVSS.n1704 4.6505
R17201 DVSS.n1709 DVSS.n1708 4.6505
R17202 DVSS.n1713 DVSS.n1712 4.6505
R17203 DVSS.n1717 DVSS.n1716 4.6505
R17204 DVSS.n1138 DVSS.n1137 4.6505
R17205 DVSS.n1121 DVSS.n1120 4.6505
R17206 DVSS.n1080 DVSS.n1079 4.6505
R17207 DVSS.n914 DVSS.n913 4.6505
R17208 DVSS.n934 DVSS.n933 4.6505
R17209 DVSS.n916 DVSS.n915 4.6505
R17210 DVSS.n919 DVSS.n766 4.6505
R17211 DVSS.n923 DVSS.n922 4.6505
R17212 DVSS.n925 DVSS.n924 4.6505
R17213 DVSS.n765 DVSS.n762 4.6505
R17214 DVSS.n750 DVSS.n748 4.6505
R17215 DVSS.n791 DVSS.n727 4.6505
R17216 DVSS.n822 DVSS.n821 4.6505
R17217 DVSS.n824 DVSS.n823 4.6505
R17218 DVSS.n808 DVSS.n803 4.6505
R17219 DVSS.n797 DVSS.n793 4.6505
R17220 DVSS.n832 DVSS.n831 4.6505
R17221 DVSS.n834 DVSS.n833 4.6505
R17222 DVSS.n810 DVSS.n809 4.6505
R17223 DVSS.n1077 DVSS.n1076 4.6505
R17224 DVSS.n1084 DVSS.n1083 4.6505
R17225 DVSS.n1088 DVSS.n1087 4.6505
R17226 DVSS.n1092 DVSS.n1091 4.6505
R17227 DVSS.n1096 DVSS.n1095 4.6505
R17228 DVSS.n1100 DVSS.n1099 4.6505
R17229 DVSS.n1104 DVSS.n1103 4.6505
R17230 DVSS.n1108 DVSS.n1107 4.6505
R17231 DVSS.n1113 DVSS.n1112 4.6505
R17232 DVSS.n1118 DVSS.n1117 4.6505
R17233 DVSS.n1125 DVSS.n1124 4.6505
R17234 DVSS.n1129 DVSS.n1128 4.6505
R17235 DVSS.n1134 DVSS.n1133 4.6505
R17236 DVSS.n1142 DVSS.n1141 4.6505
R17237 DVSS.n1146 DVSS.n1145 4.6505
R17238 DVSS.n1153 DVSS.n1152 4.6505
R17239 DVSS.n1161 DVSS.n1160 4.6505
R17240 DVSS.n1164 DVSS.n1163 4.6505
R17241 DVSS.n2657 DVSS.n2656 4.6505
R17242 DVSS.n2653 DVSS.n2652 4.6505
R17243 DVSS.n2648 DVSS.n2647 4.6505
R17244 DVSS.n2643 DVSS.n2642 4.6505
R17245 DVSS.n2548 DVSS.n2547 4.6505
R17246 DVSS.n2552 DVSS.n2551 4.6505
R17247 DVSS.n2556 DVSS.n2555 4.6505
R17248 DVSS.n2560 DVSS.n2559 4.6505
R17249 DVSS.n2564 DVSS.n2563 4.6505
R17250 DVSS.n2570 DVSS.n2569 4.6505
R17251 DVSS.n2575 DVSS.n2574 4.6505
R17252 DVSS.n2579 DVSS.n2578 4.6505
R17253 DVSS.n2583 DVSS.n2582 4.6505
R17254 DVSS.n2589 DVSS.n2588 4.6505
R17255 DVSS.n2595 DVSS.n2594 4.6505
R17256 DVSS.n2599 DVSS.n2598 4.6505
R17257 DVSS.n2604 DVSS.n2603 4.6505
R17258 DVSS.n2612 DVSS.n2611 4.6505
R17259 DVSS.n2616 DVSS.n2615 4.6505
R17260 DVSS.n2621 DVSS.n2620 4.6505
R17261 DVSS.n2626 DVSS.n2625 4.6505
R17262 DVSS.n2630 DVSS.n2629 4.6505
R17263 DVSS.n2634 DVSS.n2633 4.6505
R17264 DVSS.n1721 DVSS.n1720 4.6505
R17265 DVSS.n1726 DVSS.n1725 4.6505
R17266 DVSS.n1731 DVSS.n1730 4.6505
R17267 DVSS.n1738 DVSS.n1737 4.6505
R17268 DVSS.n1742 DVSS.n1741 4.6505
R17269 DVSS.n1747 DVSS.n1746 4.6505
R17270 DVSS.n1755 DVSS.n1754 4.6505
R17271 DVSS.n1759 DVSS.n1758 4.6505
R17272 DVSS.n1766 DVSS.n1765 4.6505
R17273 DVSS.n1772 DVSS.n1771 4.6505
R17274 DVSS.n1778 DVSS.n1777 4.6505
R17275 DVSS.n1812 DVSS.n1811 4.6505
R17276 DVSS.n1817 DVSS.n1816 4.6505
R17277 DVSS.n1821 DVSS.n1820 4.6505
R17278 DVSS.n1206 DVSS.n1205 4.6505
R17279 DVSS.n2516 DVSS.n2515 4.6505
R17280 DVSS.n2512 DVSS.n2511 4.6505
R17281 DVSS.n2508 DVSS.n2507 4.6505
R17282 DVSS.n2501 DVSS.n2500 4.6505
R17283 DVSS.n2496 DVSS.n2495 4.6505
R17284 DVSS.n2492 DVSS.n2491 4.6505
R17285 DVSS.n2484 DVSS.n2483 4.6505
R17286 DVSS.n2479 DVSS.n2478 4.6505
R17287 DVSS.n2475 DVSS.n2474 4.6505
R17288 DVSS.n2470 DVSS.n2469 4.6505
R17289 DVSS.n2464 DVSS.n2463 4.6505
R17290 DVSS.n2460 DVSS.n2459 4.6505
R17291 DVSS.n2456 DVSS.n2455 4.6505
R17292 DVSS.n2451 DVSS.n2450 4.6505
R17293 DVSS.n2445 DVSS.n2444 4.6505
R17294 DVSS.n2441 DVSS.n2440 4.6505
R17295 DVSS.n2437 DVSS.n2436 4.6505
R17296 DVSS.n2433 DVSS.n2430 4.6505
R17297 DVSS.n2429 DVSS.n2428 4.6505
R17298 DVSS.n2339 DVSS.n2338 4.6505
R17299 DVSS.n2344 DVSS.n2343 4.6505
R17300 DVSS.n2349 DVSS.n2348 4.6505
R17301 DVSS.n2356 DVSS.n2355 4.6505
R17302 DVSS.n2360 DVSS.n2359 4.6505
R17303 DVSS.n2365 DVSS.n2364 4.6505
R17304 DVSS.n2373 DVSS.n2372 4.6505
R17305 DVSS.n2377 DVSS.n2376 4.6505
R17306 DVSS.n2381 DVSS.n2380 4.6505
R17307 DVSS.n2387 DVSS.n2386 4.6505
R17308 DVSS.n2391 DVSS.n2390 4.6505
R17309 DVSS.n2806 DVSS.n2805 4.6505
R17310 DVSS.n2813 DVSS.n2812 4.6505
R17311 DVSS.n502 DVSS.n501 4.6505
R17312 DVSS.n2791 DVSS.n2790 4.6505
R17313 DVSS.n527 DVSS.n526 4.6505
R17314 DVSS.n518 DVSS.n517 4.6505
R17315 DVSS.n514 DVSS.n513 4.6505
R17316 DVSS.n511 DVSS.n510 4.6505
R17317 DVSS.n507 DVSS.n506 4.6505
R17318 DVSS.n504 DVSS.n503 4.6505
R17319 DVSS.n498 DVSS.n497 4.6505
R17320 DVSS.n494 DVSS.n493 4.6505
R17321 DVSS.n490 DVSS.n489 4.6505
R17322 DVSS.n487 DVSS.n486 4.6505
R17323 DVSS.n2783 DVSS.n2782 4.6505
R17324 DVSS.n2788 DVSS.n2787 4.6505
R17325 DVSS.n2836 DVSS.n2835 4.6505
R17326 DVSS.n2808 DVSS.n2807 4.6505
R17327 DVSS.n2816 DVSS.n2815 4.6505
R17328 DVSS.n2819 DVSS.n2818 4.6505
R17329 DVSS.n2823 DVSS.n2822 4.6505
R17330 DVSS.n2829 DVSS.n2828 4.6505
R17331 DVSS.n2833 DVSS.n2832 4.6505
R17332 DVSS.n2796 DVSS.n2795 4.6505
R17333 DVSS.n2800 DVSS.n2799 4.6505
R17334 DVSS.n2803 DVSS.n2802 4.6505
R17335 DVSS.n2938 DVSS.n2937 4.6505
R17336 DVSS.n2921 DVSS.n2920 4.6505
R17337 DVSS.n2880 DVSS.n2879 4.6505
R17338 DVSS.n325 DVSS.n324 4.6505
R17339 DVSS.n345 DVSS.n344 4.6505
R17340 DVSS.n327 DVSS.n326 4.6505
R17341 DVSS.n330 DVSS.n177 4.6505
R17342 DVSS.n334 DVSS.n333 4.6505
R17343 DVSS.n336 DVSS.n335 4.6505
R17344 DVSS.n176 DVSS.n173 4.6505
R17345 DVSS.n161 DVSS.n159 4.6505
R17346 DVSS.n202 DVSS.n138 4.6505
R17347 DVSS.n233 DVSS.n232 4.6505
R17348 DVSS.n235 DVSS.n234 4.6505
R17349 DVSS.n219 DVSS.n214 4.6505
R17350 DVSS.n208 DVSS.n204 4.6505
R17351 DVSS.n243 DVSS.n242 4.6505
R17352 DVSS.n245 DVSS.n244 4.6505
R17353 DVSS.n221 DVSS.n220 4.6505
R17354 DVSS.n2877 DVSS.n2876 4.6505
R17355 DVSS.n2884 DVSS.n2883 4.6505
R17356 DVSS.n2888 DVSS.n2887 4.6505
R17357 DVSS.n2892 DVSS.n2891 4.6505
R17358 DVSS.n2896 DVSS.n2895 4.6505
R17359 DVSS.n2900 DVSS.n2899 4.6505
R17360 DVSS.n2904 DVSS.n2903 4.6505
R17361 DVSS.n2908 DVSS.n2907 4.6505
R17362 DVSS.n2913 DVSS.n2912 4.6505
R17363 DVSS.n2918 DVSS.n2917 4.6505
R17364 DVSS.n2925 DVSS.n2924 4.6505
R17365 DVSS.n2929 DVSS.n2928 4.6505
R17366 DVSS.n2934 DVSS.n2933 4.6505
R17367 DVSS.n2942 DVSS.n2941 4.6505
R17368 DVSS.n2946 DVSS.n2945 4.6505
R17369 DVSS.n2950 DVSS.n2949 4.6505
R17370 DVSS.n2956 DVSS.n2955 4.6505
R17371 DVSS.n2960 DVSS.n2959 4.6505
R17372 DVSS.n3087 DVSS.n3086 4.6505
R17373 DVSS.n3072 DVSS.n7 4.6505
R17374 DVSS.n3058 DVSS.n3057 4.6505
R17375 DVSS.n3041 DVSS.n3040 4.6505
R17376 DVSS.n3016 DVSS.n3015 4.6505
R17377 DVSS.n2999 DVSS.n2996 4.6505
R17378 DVSS.n3003 DVSS.n3002 4.6505
R17379 DVSS.n3007 DVSS.n3006 4.6505
R17380 DVSS.n3011 DVSS.n3010 4.6505
R17381 DVSS.n3020 DVSS.n3019 4.6505
R17382 DVSS.n3025 DVSS.n3024 4.6505
R17383 DVSS.n3029 DVSS.n3028 4.6505
R17384 DVSS.n3033 DVSS.n3032 4.6505
R17385 DVSS.n3039 DVSS.n3038 4.6505
R17386 DVSS.n3045 DVSS.n3044 4.6505
R17387 DVSS.n3049 DVSS.n3048 4.6505
R17388 DVSS.n3054 DVSS.n3053 4.6505
R17389 DVSS.n3062 DVSS.n3061 4.6505
R17390 DVSS.n3066 DVSS.n3065 4.6505
R17391 DVSS.n3071 DVSS.n3070 4.6505
R17392 DVSS.n3076 DVSS.n3075 4.6505
R17393 DVSS.n3080 DVSS.n3079 4.6505
R17394 DVSS.n3084 DVSS.n3083 4.6505
R17395 DVSS.n2994 DVSS.n2993 4.6505
R17396 DVSS.n565 DVSS.n564 4.6505
R17397 DVSS.n570 DVSS.n569 4.6505
R17398 DVSS.n575 DVSS.n574 4.6505
R17399 DVSS.n579 DVSS.n578 4.6505
R17400 DVSS.n2754 DVSS.n2753 4.6505
R17401 DVSS.n581 DVSS.n580 4.6505
R17402 DVSS.n581 DVSS.n560 4.6505
R17403 DVSS.n2752 DVSS.n581 4.6505
R17404 DVSS.n2680 DVSS.n586 4.6505
R17405 DVSS.n2736 DVSS.n583 4.6505
R17406 DVSS.n2722 DVSS.n2721 4.6505
R17407 DVSS.n2705 DVSS.n2704 4.6505
R17408 DVSS.n2751 DVSS.n2750 4.6505
R17409 DVSS.n2748 DVSS.n2747 4.6505
R17410 DVSS.n2744 DVSS.n2743 4.6505
R17411 DVSS.n2740 DVSS.n2739 4.6505
R17412 DVSS.n2735 DVSS.n2734 4.6505
R17413 DVSS.n2730 DVSS.n2729 4.6505
R17414 DVSS.n2726 DVSS.n2725 4.6505
R17415 DVSS.n2718 DVSS.n2717 4.6505
R17416 DVSS.n2713 DVSS.n2712 4.6505
R17417 DVSS.n2709 DVSS.n2708 4.6505
R17418 DVSS.n2703 DVSS.n2702 4.6505
R17419 DVSS.n2697 DVSS.n2696 4.6505
R17420 DVSS.n2693 DVSS.n2692 4.6505
R17421 DVSS.n2689 DVSS.n2688 4.6505
R17422 DVSS.n2684 DVSS.n2683 4.6505
R17423 DVSS.n2678 DVSS.n2677 4.6505
R17424 DVSS.n2674 DVSS.n2673 4.6505
R17425 DVSS.n2670 DVSS.n2669 4.6505
R17426 DVSS.n2668 DVSS.n589 4.6505
R17427 DVSS.n592 DVSS.n591 4.6505
R17428 DVSS.n2777 DVSS.n556 4.6505
R17429 DVSS.n2775 DVSS.n2774 4.6505
R17430 DVSS.n2771 DVSS.n2770 4.6505
R17431 DVSS.n2766 DVSS.n2765 4.6505
R17432 DVSS.n2761 DVSS.n2760 4.6505
R17433 DVSS.n558 DVSS.n557 4.6505
R17434 DVSS.n2767 DVSS.n557 4.6505
R17435 DVSS.n542 DVSS.n541 4.6505
R17436 DVSS.n552 DVSS.n551 4.6505
R17437 DVSS.n548 DVSS.n547 4.6505
R17438 DVSS.n3 DVSS.n2 4.6505
R17439 DVSS.n3094 DVSS.n3093 4.6505
R17440 DVSS.n3095 DVSS.n4 4.6505
R17441 DVSS.n5 DVSS.n4 4.6505
R17442 DVSS.n2169 DVSS.n1937 4.5005
R17443 DVSS.n2399 DVSS.n2398 4.5005
R17444 DVSS.n2419 DVSS.n2418 4.5005
R17445 DVSS.n1551 DVSS.n1319 4.5005
R17446 DVSS.n1213 DVSS.n1212 4.5005
R17447 DVSS.n1785 DVSS.n1784 4.5005
R17448 DVSS.n938 DVSS.n706 4.5005
R17449 DVSS.n1171 DVSS.n1170 4.5005
R17450 DVSS.n349 DVSS.n117 4.5005
R17451 DVSS.n2968 DVSS.n2967 4.5005
R17452 DVSS.n2984 DVSS.n2983 4.5005
R17453 DVSS.n599 DVSS.n598 4.5005
R17454 DVSS.n2175 DVSS.n2174 4.40783
R17455 DVSS.n1557 DVSS.n1556 4.40783
R17456 DVSS.n944 DVSS.n943 4.40783
R17457 DVSS.n355 DVSS.n354 4.40783
R17458 DVSS.n2066 DVSS.n2022 4.31208
R17459 DVSS.n1448 DVSS.n1404 4.31208
R17460 DVSS.n835 DVSS.n791 4.31208
R17461 DVSS.n246 DVSS.n202 4.31208
R17462 DVSS.n2065 DVSS.n2023 4.04261
R17463 DVSS.n1447 DVSS.n1405 4.04261
R17464 DVSS.n834 DVSS.n792 4.04261
R17465 DVSS.n245 DVSS.n203 4.04261
R17466 DVSS.n1976 DVSS.n1961 3.93153
R17467 DVSS.n1955 DVSS.n1940 3.93153
R17468 DVSS.n1358 DVSS.n1343 3.93153
R17469 DVSS.n1337 DVSS.n1322 3.93153
R17470 DVSS.n745 DVSS.n730 3.93153
R17471 DVSS.n724 DVSS.n709 3.93153
R17472 DVSS.n156 DVSS.n141 3.93153
R17473 DVSS.n135 DVSS.n120 3.93153
R17474 DVSS.n2022 DVSS.n2009 3.8405
R17475 DVSS.n1404 DVSS.n1391 3.8405
R17476 DVSS.n791 DVSS.n778 3.8405
R17477 DVSS.n202 DVSS.n189 3.8405
R17478 DVSS.n2062 DVSS.n2061 3.77313
R17479 DVSS.n1444 DVSS.n1443 3.77313
R17480 DVSS.n831 DVSS.n830 3.77313
R17481 DVSS.n242 DVSS.n241 3.77313
R17482 DVSS.n525 DVSS.n524 3.69563
R17483 DVSS.n2303 DVSS.n2302 3.69446
R17484 DVSS.n1685 DVSS.n1682 3.69446
R17485 DVSS.n1072 DVSS.n1069 3.69446
R17486 DVSS.n2872 DVSS.n480 3.69446
R17487 DVSS.n2721 DVSS.n2720 3.68864
R17488 DVSS.n3057 DVSS.n3056 3.68864
R17489 DVSS.n1750 DVSS.n1748 3.68864
R17490 DVSS.n2607 DVSS.n2606 3.68864
R17491 DVSS.n2487 DVSS.n2486 3.68864
R17492 DVSS.n2368 DVSS.n2366 3.68864
R17493 DVSS.n1137 DVSS.n1135 3.68864
R17494 DVSS.n2937 DVSS.n2935 3.68864
R17495 DVSS.n2032 DVSS.n2028 3.50366
R17496 DVSS.n1414 DVSS.n1410 3.50366
R17497 DVSS.n801 DVSS.n797 3.50366
R17498 DVSS.n212 DVSS.n208 3.50366
R17499 DVSS.n2056 DVSS.n2034 3.23418
R17500 DVSS.n1438 DVSS.n1416 3.23418
R17501 DVSS.n825 DVSS.n803 3.23418
R17502 DVSS.n236 DVSS.n214 3.23418
R17503 DVSS.n2170 DVSS.n2168 3.20387
R17504 DVSS.n1552 DVSS.n1550 3.20387
R17505 DVSS.n939 DVSS.n937 3.20387
R17506 DVSS.n350 DVSS.n348 3.20387
R17507 DVSS.n1802 DVSS.n1801 3.03311
R17508 DVSS.n1179 DVSS.n1178 3.03311
R17509 DVSS.n1792 DVSS.n1791 3.03311
R17510 DVSS.n2415 DVSS.n2414 3.03311
R17511 DVSS.n2405 DVSS.n2404 3.03311
R17512 DVSS.n2976 DVSS.n2975 3.03311
R17513 DVSS.n12 DVSS.n11 3.03311
R17514 DVSS.n1188 DVSS.n1187 3.03311
R17515 DVSS.n2055 DVSS.n2038 2.96471
R17516 DVSS.n1437 DVSS.n1420 2.96471
R17517 DVSS.n824 DVSS.n807 2.96471
R17518 DVSS.n235 DVSS.n218 2.96471
R17519 DVSS.n586 DVSS.n585 2.84494
R17520 DVSS.n3015 DVSS.n3014 2.84494
R17521 DVSS.n1198 DVSS.n1197 2.84494
R17522 DVSS.n1831 DVSS.n1830 2.84494
R17523 DVSS.n1201 DVSS 2.78465
R17524 DVSS.n2052 DVSS.n2051 2.69524
R17525 DVSS.n1434 DVSS.n1433 2.69524
R17526 DVSS.n821 DVSS.n820 2.69524
R17527 DVSS.n232 DVSS.n231 2.69524
R17528 DVSS.n2144 DVSS.n2143 2.5605
R17529 DVSS.n1526 DVSS.n1525 2.5605
R17530 DVSS.n913 DVSS.n912 2.5605
R17531 DVSS.n324 DVSS.n323 2.5605
R17532 DVSS.n2047 DVSS.n2041 2.42576
R17533 DVSS.n2047 DVSS.n2015 2.42576
R17534 DVSS.n1429 DVSS.n1423 2.42576
R17535 DVSS.n1429 DVSS.n1397 2.42576
R17536 DVSS.n816 DVSS.n810 2.42576
R17537 DVSS.n816 DVSS.n784 2.42576
R17538 DVSS.n227 DVSS.n221 2.42576
R17539 DVSS.n227 DVSS.n195 2.42576
R17540 DVSS.n2660 DVSS.n1190 2.38846
R17541 DVSS.n1768 DVSS.n1767 2.31469
R17542 DVSS.n2383 DVSS.n2382 2.31469
R17543 DVSS.n1155 DVSS.n1154 2.31469
R17544 DVSS.n2952 DVSS.n2951 2.31469
R17545 DVSS.n2005 DVSS.n1999 2.29103
R17546 DVSS.n1387 DVSS.n1381 2.29103
R17547 DVSS.n774 DVSS.n768 2.29103
R17548 DVSS.n185 DVSS.n179 2.29103
R17549 DVSS.n2051 DVSS.n2041 2.15629
R17550 DVSS.n2109 DVSS.n2015 2.15629
R17551 DVSS.n1433 DVSS.n1423 2.15629
R17552 DVSS.n1491 DVSS.n1397 2.15629
R17553 DVSS.n820 DVSS.n810 2.15629
R17554 DVSS.n878 DVSS.n784 2.15629
R17555 DVSS.n231 DVSS.n221 2.15629
R17556 DVSS.n289 DVSS.n195 2.15629
R17557 DVSS.n2778 DVSS.n2777 2.01072
R17558 DVSS.n2540 DVSS.n1201 1.93608
R17559 DVSS.n2052 DVSS.n2038 1.88682
R17560 DVSS.n1434 DVSS.n1420 1.88682
R17561 DVSS.n821 DVSS.n807 1.88682
R17562 DVSS.n232 DVSS.n218 1.88682
R17563 DVSS.n2143 DVSS.n2141 1.68471
R17564 DVSS.n2137 DVSS.n2005 1.68471
R17565 DVSS.n1525 DVSS.n1523 1.68471
R17566 DVSS.n1519 DVSS.n1387 1.68471
R17567 DVSS.n912 DVSS.n910 1.68471
R17568 DVSS.n906 DVSS.n774 1.68471
R17569 DVSS.n323 DVSS.n321 1.68471
R17570 DVSS.n317 DVSS.n185 1.68471
R17571 DVSS.n2164 DVSS.n2163 1.64728
R17572 DVSS.n1546 DVSS.n1545 1.64728
R17573 DVSS.n933 DVSS.n932 1.64728
R17574 DVSS.n344 DVSS.n343 1.64728
R17575 DVSS.n2056 DVSS.n2055 1.61734
R17576 DVSS.n1438 DVSS.n1437 1.61734
R17577 DVSS.n825 DVSS.n824 1.61734
R17578 DVSS.n236 DVSS.n235 1.61734
R17579 DVSS.n2175 DVSS.n1908 1.59464
R17580 DVSS.n2182 DVSS.n1908 1.59464
R17581 DVSS.n2182 DVSS.n1909 1.59464
R17582 DVSS.n2178 DVSS.n1909 1.59464
R17583 DVSS.n2178 DVSS.n1875 1.59464
R17584 DVSS.n2192 DVSS.n1875 1.59464
R17585 DVSS.n2202 DVSS.n1873 1.59464
R17586 DVSS.n2197 DVSS.n1861 1.59464
R17587 DVSS.n2213 DVSS.n1861 1.59464
R17588 DVSS.n2214 DVSS.n2213 1.59464
R17589 DVSS.n2214 DVSS.n1859 1.59464
R17590 DVSS.n2220 DVSS.n2219 1.59464
R17591 DVSS.n2220 DVSS.n1856 1.59464
R17592 DVSS.n2250 DVSS.n1856 1.59464
R17593 DVSS.n2246 DVSS.n1841 1.59464
R17594 DVSS.n2284 DVSS.n1841 1.59464
R17595 DVSS.n2285 DVSS.n2284 1.59464
R17596 DVSS.n2286 DVSS.n2285 1.59464
R17597 DVSS.n2286 DVSS.n1839 1.59464
R17598 DVSS.n2290 DVSS.n1839 1.59464
R17599 DVSS.n1557 DVSS.n1290 1.59464
R17600 DVSS.n1564 DVSS.n1290 1.59464
R17601 DVSS.n1564 DVSS.n1291 1.59464
R17602 DVSS.n1560 DVSS.n1291 1.59464
R17603 DVSS.n1560 DVSS.n1257 1.59464
R17604 DVSS.n1574 DVSS.n1257 1.59464
R17605 DVSS.n1584 DVSS.n1255 1.59464
R17606 DVSS.n1579 DVSS.n1243 1.59464
R17607 DVSS.n1595 DVSS.n1243 1.59464
R17608 DVSS.n1596 DVSS.n1595 1.59464
R17609 DVSS.n1596 DVSS.n1241 1.59464
R17610 DVSS.n1602 DVSS.n1601 1.59464
R17611 DVSS.n1602 DVSS.n1238 1.59464
R17612 DVSS.n1632 DVSS.n1238 1.59464
R17613 DVSS.n1628 DVSS.n1223 1.59464
R17614 DVSS.n1666 DVSS.n1223 1.59464
R17615 DVSS.n1667 DVSS.n1666 1.59464
R17616 DVSS.n1668 DVSS.n1667 1.59464
R17617 DVSS.n1668 DVSS.n1221 1.59464
R17618 DVSS.n1672 DVSS.n1221 1.59464
R17619 DVSS.n944 DVSS.n677 1.59464
R17620 DVSS.n951 DVSS.n677 1.59464
R17621 DVSS.n951 DVSS.n678 1.59464
R17622 DVSS.n947 DVSS.n678 1.59464
R17623 DVSS.n947 DVSS.n644 1.59464
R17624 DVSS.n961 DVSS.n644 1.59464
R17625 DVSS.n971 DVSS.n642 1.59464
R17626 DVSS.n966 DVSS.n630 1.59464
R17627 DVSS.n982 DVSS.n630 1.59464
R17628 DVSS.n983 DVSS.n982 1.59464
R17629 DVSS.n983 DVSS.n628 1.59464
R17630 DVSS.n989 DVSS.n988 1.59464
R17631 DVSS.n989 DVSS.n625 1.59464
R17632 DVSS.n1019 DVSS.n625 1.59464
R17633 DVSS.n1015 DVSS.n610 1.59464
R17634 DVSS.n1053 DVSS.n610 1.59464
R17635 DVSS.n1054 DVSS.n1053 1.59464
R17636 DVSS.n1055 DVSS.n1054 1.59464
R17637 DVSS.n1055 DVSS.n608 1.59464
R17638 DVSS.n1059 DVSS.n608 1.59464
R17639 DVSS.n355 DVSS.n88 1.59464
R17640 DVSS.n362 DVSS.n88 1.59464
R17641 DVSS.n362 DVSS.n89 1.59464
R17642 DVSS.n358 DVSS.n89 1.59464
R17643 DVSS.n358 DVSS.n55 1.59464
R17644 DVSS.n372 DVSS.n55 1.59464
R17645 DVSS.n382 DVSS.n53 1.59464
R17646 DVSS.n377 DVSS.n41 1.59464
R17647 DVSS.n393 DVSS.n41 1.59464
R17648 DVSS.n394 DVSS.n393 1.59464
R17649 DVSS.n394 DVSS.n39 1.59464
R17650 DVSS.n400 DVSS.n399 1.59464
R17651 DVSS.n400 DVSS.n36 1.59464
R17652 DVSS.n430 DVSS.n36 1.59464
R17653 DVSS.n426 DVSS.n21 1.59464
R17654 DVSS.n464 DVSS.n21 1.59464
R17655 DVSS.n465 DVSS.n464 1.59464
R17656 DVSS.n466 DVSS.n465 1.59464
R17657 DVSS.n466 DVSS.n19 1.59464
R17658 DVSS.n470 DVSS.n19 1.59464
R17659 DVSS.n1992 DVSS.n1981 1.54748
R17660 DVSS.n1374 DVSS.n1363 1.54748
R17661 DVSS.n761 DVSS.n750 1.54748
R17662 DVSS.n172 DVSS.n161 1.54748
R17663 DVSS.n1962 DVSS.n1960 1.50638
R17664 DVSS.n1941 DVSS.n1939 1.50638
R17665 DVSS.n1344 DVSS.n1342 1.50638
R17666 DVSS.n1323 DVSS.n1321 1.50638
R17667 DVSS.n731 DVSS.n729 1.50638
R17668 DVSS.n710 DVSS.n708 1.50638
R17669 DVSS.n142 DVSS.n140 1.50638
R17670 DVSS.n121 DVSS.n119 1.50638
R17671 DVSS.n2219 DVSS.n2218 1.45398
R17672 DVSS.n1601 DVSS.n1600 1.45398
R17673 DVSS.n988 DVSS.n987 1.45398
R17674 DVSS.n399 DVSS.n398 1.45398
R17675 DVSS.n1969 DVSS.n1968 1.45108
R17676 DVSS.n1948 DVSS.n1947 1.45108
R17677 DVSS.n1351 DVSS.n1350 1.45108
R17678 DVSS.n1330 DVSS.n1329 1.45108
R17679 DVSS.n738 DVSS.n737 1.45108
R17680 DVSS.n717 DVSS.n716 1.45108
R17681 DVSS.n149 DVSS.n148 1.45108
R17682 DVSS.n128 DVSS.n127 1.45108
R17683 DVSS.n2157 DVSS.n1993 1.44767
R17684 DVSS.n1539 DVSS.n1375 1.44767
R17685 DVSS.n926 DVSS.n762 1.44767
R17686 DVSS.n337 DVSS.n173 1.44767
R17687 DVSS.n2804 DVSS 1.39202
R17688 DVSS DVSS.n2804 1.39044
R17689 DVSS.n2156 DVSS.n1995 1.34787
R17690 DVSS.n2034 DVSS.n2032 1.34787
R17691 DVSS.n1538 DVSS.n1377 1.34787
R17692 DVSS.n1416 DVSS.n1414 1.34787
R17693 DVSS.n925 DVSS.n764 1.34787
R17694 DVSS.n803 DVSS.n801 1.34787
R17695 DVSS.n336 DVSS.n175 1.34787
R17696 DVSS.n214 DVSS.n212 1.34787
R17697 DVSS.n2198 DVSS.n2197 1.26643
R17698 DVSS.n1580 DVSS.n1579 1.26643
R17699 DVSS.n967 DVSS.n966 1.26643
R17700 DVSS.n378 DVSS.n377 1.26643
R17701 DVSS.n2514 DVSS 1.2505
R17702 DVSS.n2153 DVSS.n2152 1.24806
R17703 DVSS.n1535 DVSS.n1534 1.24806
R17704 DVSS.n922 DVSS.n921 1.24806
R17705 DVSS.n333 DVSS.n332 1.24806
R17706 DVSS.n3085 DVSS 1.15435
R17707 DVSS.n2150 DVSS.n2149 1.14826
R17708 DVSS.n1532 DVSS.n1531 1.14826
R17709 DVSS.n919 DVSS.n918 1.14826
R17710 DVSS.n330 DVSS.n329 1.14826
R17711 DVSS.n2635 DVSS 1.13383
R17712 DVSS.n2980 DVSS.n2978 1.10812
R17713 DVSS.n2408 DVSS.n2407 1.10762
R17714 DVSS.n1796 DVSS.n1794 1.10762
R17715 DVSS.n1182 DVSS.n1181 1.10762
R17716 DVSS.n2144 DVSS.n2002 1.07839
R17717 DVSS.n2061 DVSS.n2028 1.07839
R17718 DVSS.n1526 DVSS.n1384 1.07839
R17719 DVSS.n1443 DVSS.n1410 1.07839
R17720 DVSS.n913 DVSS.n771 1.07839
R17721 DVSS.n830 DVSS.n797 1.07839
R17722 DVSS.n324 DVSS.n182 1.07839
R17723 DVSS.n241 DVSS.n208 1.07839
R17724 DVSS.n2147 DVSS.n1998 0.973599
R17725 DVSS.n1529 DVSS.n1380 0.973599
R17726 DVSS.n916 DVSS.n767 0.973599
R17727 DVSS.n327 DVSS.n178 0.973599
R17728 DVSS.n2062 DVSS.n2023 0.808921
R17729 DVSS.n1444 DVSS.n1405 0.808921
R17730 DVSS.n831 DVSS.n792 0.808921
R17731 DVSS.n242 DVSS.n203 0.808921
R17732 DVSS.n1975 DVSS.n1974 0.753441
R17733 DVSS.n1966 DVSS.n1963 0.753441
R17734 DVSS.n1954 DVSS.n1953 0.753441
R17735 DVSS.n1945 DVSS.n1942 0.753441
R17736 DVSS.n1357 DVSS.n1356 0.753441
R17737 DVSS.n1348 DVSS.n1345 0.753441
R17738 DVSS.n1336 DVSS.n1335 0.753441
R17739 DVSS.n1327 DVSS.n1324 0.753441
R17740 DVSS.n744 DVSS.n743 0.753441
R17741 DVSS.n735 DVSS.n732 0.753441
R17742 DVSS.n723 DVSS.n722 0.753441
R17743 DVSS.n714 DVSS.n711 0.753441
R17744 DVSS.n155 DVSS.n154 0.753441
R17745 DVSS.n146 DVSS.n143 0.753441
R17746 DVSS.n134 DVSS.n133 0.753441
R17747 DVSS.n125 DVSS.n122 0.753441
R17748 DVSS.n2149 DVSS.n2147 0.649233
R17749 DVSS.n1531 DVSS.n1529 0.649233
R17750 DVSS.n918 DVSS.n916 0.649233
R17751 DVSS.n329 DVSS.n327 0.649233
R17752 DVSS.n2141 DVSS.n1999 0.606816
R17753 DVSS.n1523 DVSS.n1381 0.606816
R17754 DVSS.n910 DVSS.n768 0.606816
R17755 DVSS.n321 DVSS.n179 0.606816
R17756 DVSS.n2174 DVSS.n2173 0.563137
R17757 DVSS.n1556 DVSS.n1555 0.563137
R17758 DVSS.n943 DVSS.n942 0.563137
R17759 DVSS.n354 DVSS.n353 0.563137
R17760 DVSS.n2152 DVSS.n2150 0.549428
R17761 DVSS.n1534 DVSS.n1532 0.549428
R17762 DVSS.n921 DVSS.n919 0.549428
R17763 DVSS.n332 DVSS.n330 0.549428
R17764 DVSS.n2066 DVSS.n2065 0.539447
R17765 DVSS.n1448 DVSS.n1447 0.539447
R17766 DVSS.n835 DVSS.n834 0.539447
R17767 DVSS.n246 DVSS.n245 0.539447
R17768 DVSS.n526 DVSS.n525 0.526461
R17769 DVSS.n2863 DVSS.n2862 0.526088
R17770 DVSS.n1686 DVSS.n1685 0.502212
R17771 DVSS.n2304 DVSS.n2303 0.502212
R17772 DVSS.n1073 DVSS.n1072 0.502212
R17773 DVSS.n2873 DVSS.n2872 0.502212
R17774 DVSS.n2153 DVSS.n1995 0.449623
R17775 DVSS.n1535 DVSS.n1377 0.449623
R17776 DVSS.n922 DVSS.n764 0.449623
R17777 DVSS.n333 DVSS.n175 0.449623
R17778 DVSS.n1157 DVSS.n1156 0.441318
R17779 DVSS.n2157 DVSS.n2156 0.349818
R17780 DVSS.n2002 DVSS.n2001 0.349818
R17781 DVSS.n1539 DVSS.n1538 0.349818
R17782 DVSS.n1384 DVSS.n1383 0.349818
R17783 DVSS.n926 DVSS.n925 0.349818
R17784 DVSS.n771 DVSS.n770 0.349818
R17785 DVSS.n337 DVSS.n336 0.349818
R17786 DVSS.n182 DVSS.n181 0.349818
R17787 DVSS.n2166 DVSS.n1978 0.337926
R17788 DVSS.n2168 DVSS.n1957 0.337926
R17789 DVSS.n1548 DVSS.n1360 0.337926
R17790 DVSS.n1550 DVSS.n1339 0.337926
R17791 DVSS.n935 DVSS.n747 0.337926
R17792 DVSS.n937 DVSS.n726 0.337926
R17793 DVSS.n346 DVSS.n158 0.337926
R17794 DVSS.n348 DVSS.n137 0.337926
R17795 DVSS.n2198 DVSS.n1873 0.328705
R17796 DVSS.n1580 DVSS.n1255 0.328705
R17797 DVSS.n967 DVSS.n642 0.328705
R17798 DVSS.n378 DVSS.n53 0.328705
R17799 DVSS.n1190 DVSS 0.316512
R17800 DVSS.n2780 DVSS 0.300422
R17801 DVSS.n2245 DVSS.n1857 0.281819
R17802 DVSS.n1627 DVSS.n1239 0.281819
R17803 DVSS.n1014 DVSS.n626 0.281819
R17804 DVSS.n425 DVSS.n37 0.281819
R17805 DVSS.n2778 DVSS.n553 0.256648
R17806 DVSS.n1993 DVSS.n1992 0.250013
R17807 DVSS.n1375 DVSS.n1374 0.250013
R17808 DVSS.n762 DVSS.n761 0.250013
R17809 DVSS.n173 DVSS.n172 0.250013
R17810 DVSS DVSS.n2295 0.249718
R17811 DVSS DVSS.n1677 0.249718
R17812 DVSS DVSS.n1064 0.249718
R17813 DVSS DVSS.n475 0.249718
R17814 DVSS.n1900 DVSS.n1872 0.234932
R17815 DVSS.n1282 DVSS.n1254 0.234932
R17816 DVSS.n669 DVSS.n641 0.234932
R17817 DVSS.n80 DVSS.n52 0.234932
R17818 DVSS.n2780 DVSS.n2779 0.215447
R17819 DVSS.n2658 DVSS.n1191 0.213615
R17820 DVSS.n1201 DVSS.n1191 0.211531
R17821 DVSS.n2166 DVSS.n2165 0.198603
R17822 DVSS.n1548 DVSS.n1547 0.198603
R17823 DVSS.n935 DVSS.n934 0.198603
R17824 DVSS.n346 DVSS.n345 0.198603
R17825 DVSS.n2168 DVSS.n2167 0.196998
R17826 DVSS.n1550 DVSS.n1549 0.196998
R17827 DVSS.n937 DVSS.n936 0.196998
R17828 DVSS.n348 DVSS.n347 0.196998
R17829 DVSS.n2995 DVSS 0.18712
R17830 DVSS.n2781 DVSS 0.17755
R17831 DVSS.n2865 DVSS.n2843 0.156029
R17832 DVSS.n2865 DVSS.n2850 0.156029
R17833 DVSS.n2865 DVSS.n2855 0.156029
R17834 DVSS.n2865 DVSS.n536 0.153643
R17835 DVSS.n2793 DVSS.n2792 0.153643
R17836 DVSS.n530 DVSS.n529 0.151786
R17837 DVSS.n1177 DVSS.n1176 0.151309
R17838 DVSS.n1790 DVSS.n1789 0.151309
R17839 DVSS.n1185 DVSS.n1184 0.151309
R17840 DVSS.n530 DVSS.n516 0.151294
R17841 DVSS.n530 DVSS.n509 0.151294
R17842 DVSS.n530 DVSS.n500 0.151294
R17843 DVSS.n530 DVSS.n492 0.151294
R17844 DVSS.n2785 DVSS.n530 0.151294
R17845 DVSS.n2865 DVSS.n2810 0.151294
R17846 DVSS.n2865 DVSS.n2821 0.151294
R17847 DVSS.n2865 DVSS.n2831 0.151294
R17848 DVSS.n2865 DVSS.n2838 0.151294
R17849 DVSS.n2163 DVSS.n1981 0.150208
R17850 DVSS.n1545 DVSS.n1363 0.150208
R17851 DVSS.n932 DVSS.n750 0.150208
R17852 DVSS.n343 DVSS.n161 0.150208
R17853 DVSS.n2296 DVSS 0.147302
R17854 DVSS.n1678 DVSS 0.147302
R17855 DVSS.n1065 DVSS 0.147302
R17856 DVSS.n476 DVSS 0.147302
R17857 DVSS.n1807 DVSS 0.146353
R17858 DVSS.n565 DVSS 0.143808
R17859 DVSS.n2218 DVSS.n1859 0.141159
R17860 DVSS.n1600 DVSS.n1241 0.141159
R17861 DVSS.n987 DVSS.n628 0.141159
R17862 DVSS.n398 DVSS.n39 0.141159
R17863 DVSS.n2781 DVSS.n2780 0.126683
R17864 DVSS.n2290 DVSS.n1834 0.0942729
R17865 DVSS.n1672 DVSS.n1216 0.0942729
R17866 DVSS.n1059 DVSS.n603 0.0942729
R17867 DVSS.n470 DVSS.n14 0.0942729
R17868 DVSS.n2165 DVSS.n1979 0.0932835
R17869 DVSS.n1996 DVSS.n1979 0.0932835
R17870 DVSS.n2155 DVSS.n1996 0.0932835
R17871 DVSS.n2155 DVSS.n2154 0.0932835
R17872 DVSS.n2154 DVSS.n1997 0.0932835
R17873 DVSS.n2146 DVSS.n1997 0.0932835
R17874 DVSS.n2146 DVSS.n2145 0.0932835
R17875 DVSS.n2064 DVSS.n1958 0.0932835
R17876 DVSS.n2064 DVSS.n2063 0.0932835
R17877 DVSS.n2063 DVSS.n2024 0.0932835
R17878 DVSS.n2039 DVSS.n2024 0.0932835
R17879 DVSS.n2054 DVSS.n2039 0.0932835
R17880 DVSS.n2054 DVSS.n2053 0.0932835
R17881 DVSS.n2053 DVSS.n2040 0.0932835
R17882 DVSS.n1547 DVSS.n1361 0.0932835
R17883 DVSS.n1378 DVSS.n1361 0.0932835
R17884 DVSS.n1537 DVSS.n1378 0.0932835
R17885 DVSS.n1537 DVSS.n1536 0.0932835
R17886 DVSS.n1536 DVSS.n1379 0.0932835
R17887 DVSS.n1528 DVSS.n1379 0.0932835
R17888 DVSS.n1528 DVSS.n1527 0.0932835
R17889 DVSS.n1446 DVSS.n1340 0.0932835
R17890 DVSS.n1446 DVSS.n1445 0.0932835
R17891 DVSS.n1445 DVSS.n1406 0.0932835
R17892 DVSS.n1421 DVSS.n1406 0.0932835
R17893 DVSS.n1436 DVSS.n1421 0.0932835
R17894 DVSS.n1436 DVSS.n1435 0.0932835
R17895 DVSS.n1435 DVSS.n1422 0.0932835
R17896 DVSS.n934 DVSS.n748 0.0932835
R17897 DVSS.n765 DVSS.n748 0.0932835
R17898 DVSS.n924 DVSS.n765 0.0932835
R17899 DVSS.n924 DVSS.n923 0.0932835
R17900 DVSS.n923 DVSS.n766 0.0932835
R17901 DVSS.n915 DVSS.n766 0.0932835
R17902 DVSS.n915 DVSS.n914 0.0932835
R17903 DVSS.n833 DVSS.n727 0.0932835
R17904 DVSS.n833 DVSS.n832 0.0932835
R17905 DVSS.n832 DVSS.n793 0.0932835
R17906 DVSS.n808 DVSS.n793 0.0932835
R17907 DVSS.n823 DVSS.n808 0.0932835
R17908 DVSS.n823 DVSS.n822 0.0932835
R17909 DVSS.n822 DVSS.n809 0.0932835
R17910 DVSS.n345 DVSS.n159 0.0932835
R17911 DVSS.n176 DVSS.n159 0.0932835
R17912 DVSS.n335 DVSS.n176 0.0932835
R17913 DVSS.n335 DVSS.n334 0.0932835
R17914 DVSS.n334 DVSS.n177 0.0932835
R17915 DVSS.n326 DVSS.n177 0.0932835
R17916 DVSS.n326 DVSS.n325 0.0932835
R17917 DVSS.n244 DVSS.n138 0.0932835
R17918 DVSS.n244 DVSS.n243 0.0932835
R17919 DVSS.n243 DVSS.n204 0.0932835
R17920 DVSS.n219 DVSS.n204 0.0932835
R17921 DVSS.n234 DVSS.n219 0.0932835
R17922 DVSS.n234 DVSS.n233 0.0932835
R17923 DVSS.n233 DVSS.n220 0.0932835
R17924 DVSS.n2167 DVSS.n2166 0.0870759
R17925 DVSS.n1549 DVSS.n1548 0.0870759
R17926 DVSS.n936 DVSS.n935 0.0870759
R17927 DVSS.n347 DVSS.n346 0.0870759
R17928 DVSS.n2515 DVSS 0.0854216
R17929 DVSS DVSS.n2751 0.0843846
R17930 DVSS.n3086 DVSS 0.0802544
R17931 DVSS.n1965 DVSS.n1964 0.0793691
R17932 DVSS.n1944 DVSS.n1943 0.0793691
R17933 DVSS.n1347 DVSS.n1346 0.0793691
R17934 DVSS.n1326 DVSS.n1325 0.0793691
R17935 DVSS.n734 DVSS.n733 0.0793691
R17936 DVSS.n713 DVSS.n712 0.0793691
R17937 DVSS.n145 DVSS.n144 0.0793691
R17938 DVSS.n124 DVSS.n123 0.0793691
R17939 DVSS.n2636 DVSS 0.0791394
R17940 DVSS.n2001 DVSS.n1998 0.0753538
R17941 DVSS.n1383 DVSS.n1380 0.0753538
R17942 DVSS.n770 DVSS.n767 0.0753538
R17943 DVSS.n181 DVSS.n178 0.0753538
R17944 DVSS.n2538 DVSS.n2534 0.0736707
R17945 DVSS.n2775 DVSS.n2771 0.0719286
R17946 DVSS.n2194 DVSS.n2193 0.0637979
R17947 DVSS.n2201 DVSS.n2194 0.0637979
R17948 DVSS.n2249 DVSS.n2248 0.0637979
R17949 DVSS.n2248 DVSS.n2247 0.0637979
R17950 DVSS.n1576 DVSS.n1575 0.0637979
R17951 DVSS.n1583 DVSS.n1576 0.0637979
R17952 DVSS.n1631 DVSS.n1630 0.0637979
R17953 DVSS.n1630 DVSS.n1629 0.0637979
R17954 DVSS.n963 DVSS.n962 0.0637979
R17955 DVSS.n970 DVSS.n963 0.0637979
R17956 DVSS.n1018 DVSS.n1017 0.0637979
R17957 DVSS.n1017 DVSS.n1016 0.0637979
R17958 DVSS.n374 DVSS.n373 0.0637979
R17959 DVSS.n381 DVSS.n374 0.0637979
R17960 DVSS.n429 DVSS.n428 0.0637979
R17961 DVSS.n428 DVSS.n427 0.0637979
R17962 DVSS.n2539 DVSS.n2538 0.0637622
R17963 DVSS.n2776 DVSS.n2775 0.062256
R17964 DVSS.n2513 DVSS.n2512 0.0617245
R17965 DVSS.n2512 DVSS.n2508 0.0617245
R17966 DVSS.n2496 DVSS.n2492 0.0617245
R17967 DVSS.n2479 DVSS.n2475 0.0617245
R17968 DVSS.n2464 DVSS.n2460 0.0617245
R17969 DVSS.n2460 DVSS.n2456 0.0617245
R17970 DVSS.n2445 DVSS.n2441 0.0617245
R17971 DVSS.n2441 DVSS.n2437 0.0617245
R17972 DVSS.n2430 DVSS.n2429 0.0617245
R17973 DVSS.n1701 DVSS.n1697 0.0611061
R17974 DVSS.n1705 DVSS.n1701 0.0611061
R17975 DVSS.n1709 DVSS.n1705 0.0611061
R17976 DVSS.n1713 DVSS.n1709 0.0611061
R17977 DVSS.n1717 DVSS.n1713 0.0611061
R17978 DVSS.n1721 DVSS.n1717 0.0611061
R17979 DVSS.n1726 DVSS.n1721 0.0611061
R17980 DVSS.n1742 DVSS.n1738 0.0611061
R17981 DVSS.n1759 DVSS.n1755 0.0611061
R17982 DVSS.n1766 DVSS.n1759 0.0611061
R17983 DVSS.n1778 DVSS.n1772 0.0611061
R17984 DVSS.n2319 DVSS.n2315 0.0611061
R17985 DVSS.n2323 DVSS.n2319 0.0611061
R17986 DVSS.n2327 DVSS.n2323 0.0611061
R17987 DVSS.n2331 DVSS.n2327 0.0611061
R17988 DVSS.n2335 DVSS.n2331 0.0611061
R17989 DVSS.n2339 DVSS.n2335 0.0611061
R17990 DVSS.n2344 DVSS.n2339 0.0611061
R17991 DVSS.n2360 DVSS.n2356 0.0611061
R17992 DVSS.n2377 DVSS.n2373 0.0611061
R17993 DVSS.n2381 DVSS.n2377 0.0611061
R17994 DVSS.n2391 DVSS.n2387 0.0611061
R17995 DVSS.n1088 DVSS.n1084 0.0611061
R17996 DVSS.n1092 DVSS.n1088 0.0611061
R17997 DVSS.n1096 DVSS.n1092 0.0611061
R17998 DVSS.n1100 DVSS.n1096 0.0611061
R17999 DVSS.n1104 DVSS.n1100 0.0611061
R18000 DVSS.n1108 DVSS.n1104 0.0611061
R18001 DVSS.n1113 DVSS.n1108 0.0611061
R18002 DVSS.n1129 DVSS.n1125 0.0611061
R18003 DVSS.n1146 DVSS.n1142 0.0611061
R18004 DVSS.n1153 DVSS.n1146 0.0611061
R18005 DVSS.n1164 DVSS.n1161 0.0611061
R18006 DVSS.n2888 DVSS.n2884 0.0611061
R18007 DVSS.n2892 DVSS.n2888 0.0611061
R18008 DVSS.n2896 DVSS.n2892 0.0611061
R18009 DVSS.n2900 DVSS.n2896 0.0611061
R18010 DVSS.n2904 DVSS.n2900 0.0611061
R18011 DVSS.n2908 DVSS.n2904 0.0611061
R18012 DVSS.n2913 DVSS.n2908 0.0611061
R18013 DVSS.n2929 DVSS.n2925 0.0611061
R18014 DVSS.n2946 DVSS.n2942 0.0611061
R18015 DVSS.n2950 DVSS.n2946 0.0611061
R18016 DVSS.n2960 DVSS.n2956 0.0611061
R18017 DVSS.n2475 DVSS.n2471 0.0610867
R18018 DVSS.n2429 DVSS.n2425 0.060449
R18019 DVSS.n1780 DVSS.n1778 0.0592121
R18020 DVSS.n2393 DVSS.n2391 0.0592121
R18021 DVSS.n1166 DVSS.n1164 0.0592121
R18022 DVSS.n2962 DVSS.n2960 0.0592121
R18023 DVSS.n1743 DVSS.n1742 0.0585808
R18024 DVSS.n2361 DVSS.n2360 0.0585808
R18025 DVSS.n1130 DVSS.n1129 0.0585808
R18026 DVSS.n2930 DVSS.n2929 0.0585808
R18027 DVSS.n2751 DVSS.n2748 0.0581923
R18028 DVSS.n2748 DVSS.n2744 0.0581923
R18029 DVSS.n2744 DVSS.n2740 0.0581923
R18030 DVSS.n2730 DVSS.n2726 0.0581923
R18031 DVSS.n2713 DVSS.n2709 0.0581923
R18032 DVSS.n2697 DVSS.n2693 0.0581923
R18033 DVSS.n2693 DVSS.n2689 0.0581923
R18034 DVSS.n2678 DVSS.n2674 0.0581923
R18035 DVSS.n2674 DVSS.n2670 0.0581923
R18036 DVSS.n592 DVSS.n589 0.0581923
R18037 DVSS.n2709 DVSS.n2705 0.0575913
R18038 DVSS.n594 DVSS.n592 0.0569904
R18039 DVSS.n3084 DVSS.n3080 0.056838
R18040 DVSS.n3080 DVSS.n3076 0.056838
R18041 DVSS.n3066 DVSS.n3062 0.056838
R18042 DVSS.n3049 DVSS.n3045 0.056838
R18043 DVSS.n3033 DVSS.n3029 0.056838
R18044 DVSS.n3029 DVSS.n3025 0.056838
R18045 DVSS.n3011 DVSS.n3007 0.056838
R18046 DVSS.n3007 DVSS.n3003 0.056838
R18047 DVSS.n1697 DVSS.n1693 0.0566869
R18048 DVSS.n2315 DVSS.n2311 0.0566869
R18049 DVSS.n1084 DVSS.n1080 0.0566869
R18050 DVSS.n2884 DVSS.n2880 0.0566869
R18051 DVSS.n3045 DVSS.n3041 0.0562512
R18052 DVSS.n2634 DVSS.n2630 0.0557995
R18053 DVSS.n2630 DVSS.n2626 0.0557995
R18054 DVSS.n2616 DVSS.n2612 0.0557995
R18055 DVSS.n2599 DVSS.n2595 0.0557995
R18056 DVSS.n2583 DVSS.n2579 0.0557995
R18057 DVSS.n2579 DVSS.n2575 0.0557995
R18058 DVSS.n2564 DVSS.n2560 0.0557995
R18059 DVSS.n2560 DVSS.n2556 0.0557995
R18060 DVSS.n2552 DVSS.n2548 0.0557995
R18061 DVSS.n2595 DVSS.n2591 0.0552235
R18062 DVSS.n2171 DVSS.n1937 0.0547553
R18063 DVSS.n1553 DVSS.n1319 0.0547553
R18064 DVSS.n940 DVSS.n706 0.0547553
R18065 DVSS.n351 DVSS.n117 0.0547553
R18066 DVSS.n2548 DVSS.n1200 0.0546475
R18067 DVSS.n2994 DVSS.n2990 0.0546475
R18068 DVSS.n2176 DVSS.n1910 0.0505
R18069 DVSS.n1558 DVSS.n1292 0.0505
R18070 DVSS.n945 DVSS.n679 0.0505
R18071 DVSS.n356 DVSS.n90 0.0505
R18072 DVSS.n2437 DVSS 0.0476939
R18073 DVSS.n2497 DVSS.n2496 0.0470561
R18074 DVSS.n2514 DVSS.n2513 0.0464184
R18075 DVSS.n2447 DVSS.n2446 0.0464184
R18076 DVSS.n2803 DVSS.n2800 0.0459545
R18077 DVSS.n2492 DVSS.n2488 0.0457806
R18078 DVSS.n2470 DVSS.n2465 0.0457806
R18079 DVSS.n2862 DVSS.n2861 0.0456128
R18080 DVSS.n2861 DVSS.n2860 0.0456128
R18081 DVSS.n2860 DVSS.n2859 0.0456128
R18082 DVSS.n2859 DVSS.n2858 0.0456128
R18083 DVSS.n2858 DVSS.n2857 0.0456128
R18084 DVSS.n2857 DVSS.n2856 0.0456128
R18085 DVSS.n2995 DVSS.n2994 0.0454309
R18086 DVSS.n2670 DVSS 0.0449712
R18087 DVSS.n2731 DVSS.n2730 0.0443702
R18088 DVSS.n2534 DVSS.n2530 0.0439451
R18089 DVSS.n3003 DVSS 0.0439272
R18090 DVSS.n2680 DVSS.n2679 0.0437692
R18091 DVSS.n1727 DVSS.n1726 0.0434293
R18092 DVSS.n1751 DVSS.n1747 0.0434293
R18093 DVSS.n2345 DVSS.n2344 0.0434293
R18094 DVSS.n2369 DVSS.n2365 0.0434293
R18095 DVSS.n1114 DVSS.n1113 0.0434293
R18096 DVSS.n1138 DVSS.n1134 0.0434293
R18097 DVSS.n2914 DVSS.n2913 0.0434293
R18098 DVSS.n2938 DVSS.n2934 0.0434293
R18099 DVSS.n3067 DVSS.n3066 0.0433404
R18100 DVSS.n2726 DVSS.n2722 0.0431683
R18101 DVSS.n2703 DVSS.n2698 0.0431683
R18102 DVSS.n2556 DVSS 0.0431267
R18103 DVSS.n2771 DVSS.n2767 0.0429107
R18104 DVSS.n3085 DVSS.n3084 0.0427535
R18105 DVSS.n3016 DVSS.n3012 0.0427535
R18106 DVSS.n2452 DVSS.n2451 0.0425918
R18107 DVSS.n2617 DVSS.n2616 0.0425507
R18108 DVSS.n2525 DVSS 0.0424207
R18109 DVSS.n3062 DVSS.n3058 0.0421667
R18110 DVSS.n3039 DVSS.n3034 0.0421667
R18111 DVSS.n2635 DVSS.n2634 0.0419747
R18112 DVSS.n2566 DVSS.n2565 0.0419747
R18113 DVSS.n1690 DVSS.n1686 0.0415354
R18114 DVSS.n2308 DVSS.n2304 0.0415354
R18115 DVSS.n1077 DVSS.n1073 0.0415354
R18116 DVSS.n2877 DVSS.n2873 0.0415354
R18117 DVSS.n2762 DVSS 0.0414226
R18118 DVSS.n2612 DVSS.n2608 0.0413986
R18119 DVSS.n2589 DVSS.n2584 0.0413986
R18120 DVSS.n2779 DVSS 0.0413499
R18121 DVSS.n2295 DVSS.n1833 0.0401852
R18122 DVSS.n1677 DVSS.n1215 0.0401852
R18123 DVSS.n1064 DVSS.n602 0.0401852
R18124 DVSS.n475 DVSS.n13 0.0401852
R18125 DVSS.n2685 DVSS.n2684 0.0401635
R18126 DVSS.n3021 DVSS.n3020 0.0392324
R18127 DVSS.n2571 DVSS.n2570 0.0385184
R18128 DVSS.n1768 DVSS.n1766 0.036243
R18129 DVSS.n2383 DVSS.n2381 0.036243
R18130 DVSS.n1155 DVSS.n1153 0.036243
R18131 DVSS.n2952 DVSS.n2950 0.036243
R18132 DVSS.n1738 DVSS.n1734 0.0333283
R18133 DVSS.n2356 DVSS.n2352 0.0333283
R18134 DVSS.n1125 DVSS.n1121 0.0333283
R18135 DVSS.n2925 DVSS.n2921 0.0333283
R18136 DVSS.n2504 DVSS.n2501 0.03175
R18137 DVSS.n2480 DVSS.n2479 0.03175
R18138 DVSS.n2508 DVSS.n2504 0.0304745
R18139 DVSS.n2484 DVSS.n2480 0.0304745
R18140 DVSS.n2530 DVSS.n2529 0.0302256
R18141 DVSS.n2523 DVSS 0.0302256
R18142 DVSS.n2736 DVSS.n2735 0.0299471
R18143 DVSS.n2714 DVSS.n2713 0.0299471
R18144 DVSS.n2791 DVSS.n2788 0.0298561
R18145 DVSS.n2767 DVSS.n2766 0.0295179
R18146 DVSS DVSS.n558 0.0295179
R18147 DVSS.n3072 DVSS.n3071 0.0292559
R18148 DVSS.n3050 DVSS.n3049 0.0292559
R18149 DVSS.n2740 DVSS.n2736 0.0287452
R18150 DVSS.n2718 DVSS.n2714 0.0287452
R18151 DVSS.n2622 DVSS.n2621 0.0287258
R18152 DVSS.n2600 DVSS.n2599 0.0287258
R18153 DVSS.n1937 DVSS 0.0286915
R18154 DVSS.n1319 DVSS 0.0286915
R18155 DVSS.n706 DVSS 0.0286915
R18156 DVSS.n117 DVSS 0.0286915
R18157 DVSS.n1734 DVSS.n1731 0.0282778
R18158 DVSS.n2352 DVSS.n2349 0.0282778
R18159 DVSS.n1121 DVSS.n1118 0.0282778
R18160 DVSS.n2921 DVSS.n2918 0.0282778
R18161 DVSS.n3076 DVSS.n3072 0.0280822
R18162 DVSS.n3054 DVSS.n3050 0.0280822
R18163 DVSS.n2800 DVSS.n2797 0.0279621
R18164 DVSS.n2626 DVSS.n2622 0.0275737
R18165 DVSS.n2604 DVSS.n2600 0.0275737
R18166 DVSS.n2980 DVSS.n2979 0.0275051
R18167 DVSS.n2408 DVSS.n1832 0.0271646
R18168 DVSS.n1796 DVSS.n1795 0.0271646
R18169 DVSS.n1182 DVSS.n601 0.0271646
R18170 DVSS.n1772 DVSS.n1768 0.026142
R18171 DVSS.n2387 DVSS.n2383 0.026142
R18172 DVSS.n1161 DVSS.n1155 0.026142
R18173 DVSS.n2956 DVSS.n2952 0.026142
R18174 DVSS.n2529 DVSS.n2525 0.0256524
R18175 DVSS.n2766 DVSS.n2762 0.0250536
R18176 DVSS.n1793 DVSS.n1786 0.0249644
R18177 DVSS.n2406 DVSS.n2400 0.0249644
R18178 DVSS.n1180 DVSS.n1172 0.0249644
R18179 DVSS.n2977 DVSS.n2969 0.0249644
R18180 DVSS.n1817 DVSS.n1812 0.0245
R18181 DVSS.n575 DVSS.n570 0.0245
R18182 DVSS.n2982 DVSS.n2981 0.0237334
R18183 DVSS.n1787 DVSS 0.0237145
R18184 DVSS.n2401 DVSS 0.0237145
R18185 DVSS.n1173 DVSS 0.0237145
R18186 DVSS.n2970 DVSS 0.0237145
R18187 DVSS.n552 DVSS.n548 0.0237108
R18188 DVSS.n2409 DVSS 0.0236262
R18189 DVSS.n2657 DVSS.n2653 0.0235326
R18190 DVSS DVSS.n2803 0.0232273
R18191 DVSS.n2805 DVSS 0.0230564
R18192 DVSS.n1967 DVSS.n1965 0.0228214
R18193 DVSS.n1946 DVSS.n1944 0.0228214
R18194 DVSS.n1349 DVSS.n1347 0.0228214
R18195 DVSS.n1328 DVSS.n1326 0.0228214
R18196 DVSS.n736 DVSS.n734 0.0228214
R18197 DVSS.n715 DVSS.n713 0.0228214
R18198 DVSS.n147 DVSS.n145 0.0228214
R18199 DVSS.n126 DVSS.n124 0.0228214
R18200 DVSS DVSS.n1189 0.0223216
R18201 DVSS.n486 DVSS.n485 0.0222446
R18202 DVSS DVSS.n1803 0.0214378
R18203 DVSS DVSS.n561 0.0214378
R18204 DVSS.n1812 DVSS.n1808 0.02125
R18205 DVSS.n570 DVSS.n566 0.02125
R18206 DVSS.n2419 DVSS.n2417 0.0204913
R18207 DVSS.n2407 DVSS.n2297 0.0198972
R18208 DVSS.n1794 DVSS.n1679 0.0198972
R18209 DVSS.n1181 DVSS.n1066 0.0198972
R18210 DVSS.n2978 DVSS.n477 0.0198972
R18211 DVSS.n1978 DVSS.n1959 0.0198452
R18212 DVSS.n1957 DVSS.n1938 0.0198452
R18213 DVSS.n1360 DVSS.n1341 0.0198452
R18214 DVSS.n1339 DVSS.n1320 0.0198452
R18215 DVSS.n747 DVSS.n728 0.0198452
R18216 DVSS.n726 DVSS.n707 0.0198452
R18217 DVSS.n158 DVSS.n139 0.0198452
R18218 DVSS.n137 DVSS.n118 0.0198452
R18219 DVSS.n2456 DVSS.n2452 0.0196327
R18220 DVSS.n600 DVSS.n599 0.0194094
R18221 DVSS.n2177 DVSS.n2176 0.0185851
R18222 DVSS.n2181 DVSS.n2177 0.0185851
R18223 DVSS.n2181 DVSS.n2180 0.0185851
R18224 DVSS.n2180 DVSS.n2179 0.0185851
R18225 DVSS.n2179 DVSS.n1874 0.0185851
R18226 DVSS.n2193 DVSS.n1874 0.0185851
R18227 DVSS.n2201 DVSS.n2200 0.0185851
R18228 DVSS.n2196 DVSS.n2195 0.0185851
R18229 DVSS.n2195 DVSS.n1860 0.0185851
R18230 DVSS.n2215 DVSS.n1860 0.0185851
R18231 DVSS.n2216 DVSS.n2215 0.0185851
R18232 DVSS.n2221 DVSS.n1858 0.0185851
R18233 DVSS.n2222 DVSS.n2221 0.0185851
R18234 DVSS.n2249 DVSS.n2222 0.0185851
R18235 DVSS.n2247 DVSS.n2223 0.0185851
R18236 DVSS.n2223 DVSS.n1842 0.0185851
R18237 DVSS.n1842 DVSS.n1840 0.0185851
R18238 DVSS.n2287 DVSS.n1840 0.0185851
R18239 DVSS.n2288 DVSS.n2287 0.0185851
R18240 DVSS.n2289 DVSS.n2288 0.0185851
R18241 DVSS.n1559 DVSS.n1558 0.0185851
R18242 DVSS.n1563 DVSS.n1559 0.0185851
R18243 DVSS.n1563 DVSS.n1562 0.0185851
R18244 DVSS.n1562 DVSS.n1561 0.0185851
R18245 DVSS.n1561 DVSS.n1256 0.0185851
R18246 DVSS.n1575 DVSS.n1256 0.0185851
R18247 DVSS.n1583 DVSS.n1582 0.0185851
R18248 DVSS.n1578 DVSS.n1577 0.0185851
R18249 DVSS.n1577 DVSS.n1242 0.0185851
R18250 DVSS.n1597 DVSS.n1242 0.0185851
R18251 DVSS.n1598 DVSS.n1597 0.0185851
R18252 DVSS.n1603 DVSS.n1240 0.0185851
R18253 DVSS.n1604 DVSS.n1603 0.0185851
R18254 DVSS.n1631 DVSS.n1604 0.0185851
R18255 DVSS.n1629 DVSS.n1605 0.0185851
R18256 DVSS.n1605 DVSS.n1224 0.0185851
R18257 DVSS.n1224 DVSS.n1222 0.0185851
R18258 DVSS.n1669 DVSS.n1222 0.0185851
R18259 DVSS.n1670 DVSS.n1669 0.0185851
R18260 DVSS.n1671 DVSS.n1670 0.0185851
R18261 DVSS.n946 DVSS.n945 0.0185851
R18262 DVSS.n950 DVSS.n946 0.0185851
R18263 DVSS.n950 DVSS.n949 0.0185851
R18264 DVSS.n949 DVSS.n948 0.0185851
R18265 DVSS.n948 DVSS.n643 0.0185851
R18266 DVSS.n962 DVSS.n643 0.0185851
R18267 DVSS.n970 DVSS.n969 0.0185851
R18268 DVSS.n965 DVSS.n964 0.0185851
R18269 DVSS.n964 DVSS.n629 0.0185851
R18270 DVSS.n984 DVSS.n629 0.0185851
R18271 DVSS.n985 DVSS.n984 0.0185851
R18272 DVSS.n990 DVSS.n627 0.0185851
R18273 DVSS.n991 DVSS.n990 0.0185851
R18274 DVSS.n1018 DVSS.n991 0.0185851
R18275 DVSS.n1016 DVSS.n992 0.0185851
R18276 DVSS.n992 DVSS.n611 0.0185851
R18277 DVSS.n611 DVSS.n609 0.0185851
R18278 DVSS.n1056 DVSS.n609 0.0185851
R18279 DVSS.n1057 DVSS.n1056 0.0185851
R18280 DVSS.n1058 DVSS.n1057 0.0185851
R18281 DVSS.n357 DVSS.n356 0.0185851
R18282 DVSS.n361 DVSS.n357 0.0185851
R18283 DVSS.n361 DVSS.n360 0.0185851
R18284 DVSS.n360 DVSS.n359 0.0185851
R18285 DVSS.n359 DVSS.n54 0.0185851
R18286 DVSS.n373 DVSS.n54 0.0185851
R18287 DVSS.n381 DVSS.n380 0.0185851
R18288 DVSS.n376 DVSS.n375 0.0185851
R18289 DVSS.n375 DVSS.n40 0.0185851
R18290 DVSS.n395 DVSS.n40 0.0185851
R18291 DVSS.n396 DVSS.n395 0.0185851
R18292 DVSS.n401 DVSS.n38 0.0185851
R18293 DVSS.n402 DVSS.n401 0.0185851
R18294 DVSS.n429 DVSS.n402 0.0185851
R18295 DVSS.n427 DVSS.n403 0.0185851
R18296 DVSS.n403 DVSS.n22 0.0185851
R18297 DVSS.n22 DVSS.n20 0.0185851
R18298 DVSS.n467 DVSS.n20 0.0185851
R18299 DVSS.n468 DVSS.n467 0.0185851
R18300 DVSS.n469 DVSS.n468 0.0185851
R18301 DVSS.n2689 DVSS.n2685 0.0185288
R18302 DVSS.n2797 DVSS.n2796 0.0184924
R18303 DVSS.n2815 DVSS.n2814 0.0183571
R18304 DVSS.n1214 DVSS.n1213 0.0183396
R18305 DVSS.n2828 DVSS.n2827 0.0183259
R18306 DVSS.n1731 DVSS.n1727 0.0181768
R18307 DVSS.n1755 DVSS.n1751 0.0181768
R18308 DVSS.n2349 DVSS.n2345 0.0181768
R18309 DVSS.n2373 DVSS.n2369 0.0181768
R18310 DVSS.n1118 DVSS.n1114 0.0181768
R18311 DVSS.n1142 DVSS.n1138 0.0181768
R18312 DVSS.n2918 DVSS.n2914 0.0181768
R18313 DVSS.n2942 DVSS.n2938 0.0181768
R18314 DVSS.n3025 DVSS.n3021 0.0181056
R18315 DVSS.n2417 DVSS.n2416 0.0180768
R18316 DVSS.n2297 DVSS.n2296 0.0179419
R18317 DVSS.n1679 DVSS.n1678 0.0179419
R18318 DVSS.n1066 DVSS.n1065 0.0179419
R18319 DVSS.n477 DVSS.n476 0.0179419
R18320 DVSS.n2575 DVSS.n2571 0.0177811
R18321 DVSS.n1793 DVSS.n1792 0.0175455
R18322 DVSS.n2406 DVSS.n2405 0.0175455
R18323 DVSS.n1180 DVSS.n1179 0.0175455
R18324 DVSS.n2977 DVSS.n2976 0.0175455
R18325 DVSS.n1183 DVSS.n600 0.0171144
R18326 DVSS.n2217 DVSS.n1858 0.0169894
R18327 DVSS.n1599 DVSS.n1240 0.0169894
R18328 DVSS.n986 DVSS.n627 0.0169894
R18329 DVSS.n397 DVSS.n38 0.0169894
R18330 DVSS.n1797 DVSS.n1214 0.0167984
R18331 DVSS.n2796 DVSS.n2791 0.0165985
R18332 DVSS.n2815 DVSS.n2813 0.0164774
R18333 DVSS.n2488 DVSS.n2484 0.0164439
R18334 DVSS.n2465 DVSS.n2464 0.0164439
R18335 DVSS.n2416 DVSS.n2415 0.0164439
R18336 DVSS.n497 DVSS.n496 0.016125
R18337 DVSS.n2722 DVSS.n2718 0.015524
R18338 DVSS.n2698 DVSS.n2697 0.015524
R18339 DVSS.n1188 DVSS.n1183 0.015524
R18340 DVSS.n2515 DVSS.n2514 0.0152059
R18341 DVSS.n3058 DVSS.n3054 0.0151714
R18342 DVSS.n3034 DVSS.n3033 0.0151714
R18343 DVSS.n2501 DVSS.n2497 0.0151684
R18344 DVSS.n2608 DVSS.n2604 0.0149009
R18345 DVSS.n2584 DVSS.n2583 0.0149009
R18346 DVSS.n1802 DVSS.n1797 0.0149009
R18347 DVSS.n2981 DVSS.n12 0.0149009
R18348 DVSS.n2199 DVSS.n2196 0.0148617
R18349 DVSS.n1581 DVSS.n1578 0.0148617
R18350 DVSS.n968 DVSS.n965 0.0148617
R18351 DVSS.n379 DVSS.n376 0.0148617
R18352 DVSS.n1822 DVSS.n1817 0.01475
R18353 DVSS.n580 DVSS.n575 0.01475
R18354 DVSS.n2430 DVSS 0.0145306
R18355 DVSS.n2735 DVSS.n2731 0.0143221
R18356 DVSS.n548 DVSS.n544 0.0142814
R18357 DVSS.n1207 DVSS 0.01425
R18358 DVSS.n560 DVSS 0.01425
R18359 DVSS.n2653 DVSS.n2649 0.0141756
R18360 DVSS.n3086 DVSS.n3085 0.0140747
R18361 DVSS.n3071 DVSS.n3067 0.0139977
R18362 DVSS.n2636 DVSS.n2635 0.0138333
R18363 DVSS.n553 DVSS.n543 0.0137979
R18364 DVSS.n3095 DVSS 0.0137979
R18365 DVSS.n2621 DVSS.n2617 0.0137488
R18366 DVSS.n589 DVSS 0.0137212
R18367 DVSS.n2659 DVSS.n2658 0.0136958
R18368 DVSS.n2644 DVSS 0.0136958
R18369 DVSS.n2996 DVSS 0.0134108
R18370 DVSS DVSS.n2552 0.0131728
R18371 DVSS.n2446 DVSS.n2445 0.0119796
R18372 DVSS.n2400 DVSS.n2399 0.0117068
R18373 DVSS.n1786 DVSS.n1785 0.0117068
R18374 DVSS.n1172 DVSS.n1171 0.0117068
R18375 DVSS.n2969 DVSS.n2968 0.0117068
R18376 DVSS.n2679 DVSS.n2678 0.0113173
R18377 DVSS.n3012 DVSS.n3011 0.0110634
R18378 DVSS.n2996 DVSS.n2995 0.0110634
R18379 DVSS.n2565 DVSS.n2564 0.0108687
R18380 DVSS.n2984 DVSS.n2982 0.0104846
R18381 DVSS.n2540 DVSS.n2539 0.0104085
R18382 DVSS.n1822 DVSS.n1821 0.01025
R18383 DVSS DVSS.n1824 0.01025
R18384 DVSS.n580 DVSS.n579 0.01025
R18385 DVSS.n2752 DVSS 0.01025
R18386 DVSS.n2777 DVSS.n2776 0.0101726
R18387 DVSS.n2423 DVSS.n2419 0.0100663
R18388 DVSS.n544 DVSS.n3 0.0099294
R18389 DVSS DVSS.n5 0.0099294
R18390 DVSS.n2649 DVSS.n2648 0.00985701
R18391 DVSS DVSS.n1193 0.00985701
R18392 DVSS.n599 DVSS.n597 0.00951442
R18393 DVSS.n1785 DVSS.n1783 0.00933838
R18394 DVSS.n2399 DVSS.n2397 0.00933838
R18395 DVSS.n1171 DVSS.n1169 0.00933838
R18396 DVSS.n2968 DVSS.n2966 0.00933838
R18397 DVSS.n1213 DVSS.n1211 0.00914055
R18398 DVSS.n2988 DVSS.n2984 0.00914055
R18399 DVSS.n2415 DVSS.n2409 0.00895784
R18400 DVSS.n2405 DVSS.n2401 0.00856303
R18401 DVSS.n1792 DVSS.n1787 0.00856303
R18402 DVSS.n1179 DVSS.n1173 0.00856303
R18403 DVSS.n2976 DVSS.n2970 0.00856303
R18404 DVSS.n1189 DVSS.n1188 0.0084995
R18405 DVSS.n1803 DVSS.n1802 0.00818896
R18406 DVSS.n561 DVSS.n12 0.00818896
R18407 DVSS.n1821 DVSS 0.008
R18408 DVSS.n579 DVSS 0.008
R18409 DVSS DVSS.n3 0.00775339
R18410 DVSS.n2648 DVSS 0.0076977
R18411 DVSS.n2524 DVSS.n2523 0.00735976
R18412 DVSS.n553 DVSS.n552 0.00726983
R18413 DVSS.n2658 DVSS.n2657 0.00721785
R18414 DVSS.n2761 DVSS.n558 0.00719643
R18415 DVSS.n2172 DVSS.n1910 0.00688298
R18416 DVSS.n1554 DVSS.n1292 0.00688298
R18417 DVSS.n941 DVSS.n679 0.00688298
R18418 DVSS.n352 DVSS.n90 0.00688298
R18419 DVSS DVSS.n2524 0.00659756
R18420 DVSS.n1964 DVSS.n1959 0.00645238
R18421 DVSS.n1943 DVSS.n1938 0.00645238
R18422 DVSS.n1346 DVSS.n1341 0.00645238
R18423 DVSS.n1325 DVSS.n1320 0.00645238
R18424 DVSS.n733 DVSS.n728 0.00645238
R18425 DVSS.n712 DVSS.n707 0.00645238
R18426 DVSS.n144 DVSS.n139 0.00645238
R18427 DVSS.n123 DVSS.n118 0.00645238
R18428 DVSS DVSS.n2761 0.00645238
R18429 DVSS.n2167 DVSS.n1958 0.00565464
R18430 DVSS.n1549 DVSS.n1340 0.00565464
R18431 DVSS.n936 DVSS.n727 0.00565464
R18432 DVSS.n347 DVSS.n138 0.00565464
R18433 DVSS.n1693 DVSS.n1690 0.00491919
R18434 DVSS.n2311 DVSS.n2308 0.00491919
R18435 DVSS.n1080 DVSS.n1077 0.00491919
R18436 DVSS.n2880 DVSS.n2877 0.00491919
R18437 DVSS.n503 DVSS.n502 0.00476136
R18438 DVSS.n2172 DVSS.n2171 0.00475532
R18439 DVSS.n1554 DVSS.n1553 0.00475532
R18440 DVSS.n941 DVSS.n940 0.00475532
R18441 DVSS.n352 DVSS.n351 0.00475532
R18442 DVSS.n2451 DVSS.n2447 0.00432653
R18443 DVSS.n2170 DVSS.n2169 0.00423171
R18444 DVSS.n1552 DVSS.n1551 0.00423171
R18445 DVSS.n939 DVSS.n938 0.00423171
R18446 DVSS.n350 DVSS.n349 0.00423171
R18447 DVSS.n2200 DVSS.n2199 0.0042234
R18448 DVSS.n1582 DVSS.n1581 0.0042234
R18449 DVSS.n969 DVSS.n968 0.0042234
R18450 DVSS.n380 DVSS.n379 0.0042234
R18451 DVSS.n2684 DVSS.n2680 0.00410577
R18452 DVSS.n3020 DVSS.n3016 0.00402113
R18453 DVSS.n2570 DVSS.n2566 0.00395622
R18454 DVSS.n1808 DVSS.n1807 0.00375
R18455 DVSS.n566 DVSS.n565 0.00375
R18456 DVSS.n543 DVSS.n542 0.00364313
R18457 DVSS.n2660 DVSS.n2659 0.003619
R18458 DVSS.n1968 DVSS.n1967 0.00347619
R18459 DVSS.n1947 DVSS.n1946 0.00347619
R18460 DVSS.n1350 DVSS.n1349 0.00347619
R18461 DVSS.n1329 DVSS.n1328 0.00347619
R18462 DVSS.n737 DVSS.n736 0.00347619
R18463 DVSS.n716 DVSS.n715 0.00347619
R18464 DVSS.n148 DVSS.n147 0.00347619
R18465 DVSS.n127 DVSS.n126 0.00347619
R18466 DVSS.n1747 DVSS.n1743 0.00302525
R18467 DVSS.n2365 DVSS.n2361 0.00302525
R18468 DVSS.n1134 DVSS.n1130 0.00302525
R18469 DVSS.n2934 DVSS.n2930 0.00302525
R18470 DVSS.n1824 DVSS.n1206 0.00275
R18471 DVSS.n2753 DVSS.n2752 0.00275
R18472 DVSS.n3094 DVSS.n5 0.00267602
R18473 DVSS.n2643 DVSS.n1193 0.00265931
R18474 DVSS DVSS.n1206 0.0025
R18475 DVSS.n2753 DVSS 0.0025
R18476 DVSS DVSS.n3094 0.00243424
R18477 DVSS DVSS.n2643 0.00241939
R18478 DVSS.n1783 DVSS.n1780 0.00239394
R18479 DVSS.n2397 DVSS.n2393 0.00239394
R18480 DVSS.n1169 DVSS.n1166 0.00239394
R18481 DVSS.n2966 DVSS.n2962 0.00239394
R18482 DVSS.n2217 DVSS.n2216 0.00209574
R18483 DVSS.n1599 DVSS.n1598 0.00209574
R18484 DVSS.n986 DVSS.n985 0.00209574
R18485 DVSS.n397 DVSS.n396 0.00209574
R18486 DVSS.n2425 DVSS.n2423 0.00177551
R18487 DVSS.n597 DVSS.n594 0.00170192
R18488 DVSS.n1211 DVSS.n1200 0.00165207
R18489 DVSS.n2990 DVSS.n2988 0.00165207
R18490 DVSS.n2289 DVSS.n1833 0.00156383
R18491 DVSS.n1671 DVSS.n1215 0.00156383
R18492 DVSS.n1058 DVSS.n602 0.00156383
R18493 DVSS.n469 DVSS.n13 0.00156383
R18494 DVSS.n2171 DVSS.n2170 0.00149989
R18495 DVSS.n1553 DVSS.n1552 0.00149989
R18496 DVSS.n940 DVSS.n939 0.00149989
R18497 DVSS.n351 DVSS.n350 0.00149989
R18498 DVSS.n2981 DVSS.n2980 0.00149701
R18499 DVSS DVSS.n1207 0.00125
R18500 DVSS DVSS.n560 0.00125
R18501 DVSS DVSS.n3095 0.00122534
R18502 DVSS DVSS.n2644 0.00121977
R18503 DVSS.n2471 DVSS.n2470 0.00113776
R18504 DVSS.n2705 DVSS.n2703 0.00110096
R18505 DVSS.n3041 DVSS.n3039 0.00108685
R18506 DVSS.n2591 DVSS.n2589 0.00107604
R18507 DVSS.n2407 DVSS.n2406 0.001
R18508 DVSS.n1794 DVSS.n1793 0.001
R18509 DVSS.n1181 DVSS.n1180 0.001
R18510 DVSS.n2978 DVSS.n2977 0.001
R18511 DVSS.n2416 DVSS.n2408 0.001
R18512 DVSS.n1797 DVSS.n1796 0.001
R18513 DVSS.n1183 DVSS.n1182 0.001
R18514 DVSS.n2169 DVSS.n1910 0.000500988
R18515 DVSS.n2174 DVSS.n1910 0.000500988
R18516 DVSS.n1551 DVSS.n1292 0.000500988
R18517 DVSS.n1556 DVSS.n1292 0.000500988
R18518 DVSS.n938 DVSS.n679 0.000500988
R18519 DVSS.n943 DVSS.n679 0.000500988
R18520 DVSS.n349 DVSS.n90 0.000500988
R18521 DVSS.n354 DVSS.n90 0.000500988
R18522 DVSS.n2199 DVSS.n2198 0.000500379
R18523 DVSS.n1581 DVSS.n1580 0.000500379
R18524 DVSS.n968 DVSS.n967 0.000500379
R18525 DVSS.n379 DVSS.n378 0.000500379
R18526 DVSS.n1834 DVSS.n1833 0.000500334
R18527 DVSS.n1216 DVSS.n1215 0.000500334
R18528 DVSS.n603 DVSS.n602 0.000500334
R18529 DVSS.n14 DVSS.n13 0.000500334
R18530 DVSS.n2218 DVSS.n2217 0.000500219
R18531 DVSS.n1600 DVSS.n1599 0.000500219
R18532 DVSS.n987 DVSS.n986 0.000500219
R18533 DVSS.n398 DVSS.n397 0.000500219
R18534 DVSS.n2804 DVSS.n2781 0.000500012
R18535 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 136.804
R18536 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 136.325
R18537 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 119.999
R18538 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 93.9023
R18539 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 93.3044
R18540 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 93.0848
R18541 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n4 92.5005
R18542 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 92.4623
R18543 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 69.2281
R18544 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 29.4833
R18545 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 27.6955
R18546 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 27.6955
R18547 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 15.4626
R18548 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n16 9.3005
R18549 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n8 9.3005
R18550 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n7 9.3005
R18551 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 9.3005
R18552 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 9.3005
R18553 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n15 9.3005
R18554 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n17 9.3005
R18555 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 9.02061
R18556 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 9.02061
R18557 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n34 8.28285
R18558 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n21 8.28285
R18559 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 5.64756
R18560 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 5.31864
R18561 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n42 4.14168
R18562 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n28 4.14168
R18563 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 4.06959
R18564 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n11 3.93153
R18565 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n40 3.76521
R18566 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n33 3.76521
R18567 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n24 3.76521
R18568 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n19 3.76521
R18569 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n36 3.38874
R18570 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n22 3.38874
R18571 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 3.0736
R18572 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 3.07249
R18573 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 3.07078
R18574 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 3.04338
R18575 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 3.03311
R18576 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 3.03311
R18577 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 3.03311
R18578 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n39 2.63579
R18579 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n20 2.63579
R18580 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 2.27447
R18581 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 2.25932
R18582 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 2.25932
R18583 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 1.80772
R18584 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n30 1.61433
R18585 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 1.45534
R18586 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 1.19419
R18587 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n9 0.753441
R18588 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 0.719888
R18589 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 0.22499
R18590 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 0.176176
R18591 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 2.36361
R18592 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 2.36353
R18593 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 1.14499
R18594 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 1.00043
R18595 B1.n66 B1.n65 185
R18596 B1.n64 B1.n57 185
R18597 B1.n24 B1.n15 185
R18598 B1.n23 B1.n22 185
R18599 B1.n69 B1.t2 120.037
R18600 B1.t3 B1.n14 120.037
R18601 B1.n59 B1.n57 112.831
R18602 B1.n22 B1.n21 112.831
R18603 B1.n68 B1.n67 104.172
R18604 B1.n27 B1.n26 104.172
R18605 B1.n68 B1.n56 92.5005
R18606 B1.n28 B1.n27 92.5005
R18607 B1.t2 B1.n68 66.8281
R18608 B1.n27 B1.t3 66.8281
R18609 B1.n6 B1.t4 35.2053
R18610 B1.n3 B1.t5 34.0571
R18611 B1.n67 B1.n66 29.4833
R18612 B1.n26 B1.n15 29.4833
R18613 B1.n1 B1.t1 27.6955
R18614 B1.n1 B1.t0 27.6955
R18615 B1.n45 B1.n44 19.0955
R18616 B1.n69 B1.n56 15.4558
R18617 B1.n28 B1.n14 15.4558
R18618 B1.n64 B1.n63 13.5534
R18619 B1.n23 B1.n18 13.5534
R18620 B1.n2 B1.n1 9.67857
R18621 B1.n41 B1.n34 9.30581
R18622 B1.n59 B1.n58 9.30424
R18623 B1.n21 B1.n20 9.30413
R18624 B1.n40 B1.n39 9.3005
R18625 B1.n46 B1.n45 9.3005
R18626 B1.n71 B1.n70 9.3005
R18627 B1.n55 B1.n52 9.3005
R18628 B1.n67 B1.n55 9.3005
R18629 B1.n63 B1.n62 9.3005
R18630 B1.n72 B1.n54 9.3005
R18631 B1.n29 B1.n13 9.3005
R18632 B1.n25 B1.n11 9.3005
R18633 B1.n26 B1.n25 9.3005
R18634 B1.n18 B1.n17 9.3005
R18635 B1.n31 B1.n30 9.3005
R18636 B1.n71 B1.n56 9.03579
R18637 B1.n29 B1.n28 9.03579
R18638 B1.n43 B1.n41 8.49366
R18639 B1.n43 B1.t7 8.2655
R18640 B1.n43 B1.t6 8.2655
R18641 B1.n44 B1.n43 7.97749
R18642 B1.n42 B1.n40 7.26743
R18643 B1.n43 B1.n42 6.15568
R18644 B1.n65 B1.n55 5.64756
R18645 B1.n25 B1.n24 5.64756
R18646 B1.n41 B1.n35 4.89462
R18647 B1.n60 B1.n59 4.89462
R18648 B1.n21 B1.n19 4.89462
R18649 B1.n73 B1.n55 4.51815
R18650 B1.n72 B1.n71 4.51815
R18651 B1.n25 B1.n12 4.51815
R18652 B1.n30 B1.n29 4.51815
R18653 B1.n5 B1.n4 4.5005
R18654 B1.n4 B1.n2 4.5005
R18655 B1.n51 B1.n9 4.5005
R18656 B1.n49 B1.n9 4.5005
R18657 B1.n51 B1.n50 4.5005
R18658 B1.n50 B1.n49 4.5005
R18659 B1.n74 B1.n53 4.5005
R18660 B1.n75 B1.n8 4.5005
R18661 B1.n53 B1.n8 4.5005
R18662 B1.n75 B1.n74 4.5005
R18663 B1.n48 B1.n32 4.5005
R18664 B1.n47 B1.n36 4.5005
R18665 B1.n48 B1.n47 4.5005
R18666 B1.n36 B1.n32 4.5005
R18667 B1.n38 B1.n33 4.5005
R18668 B1.n66 B1.n57 3.93153
R18669 B1.n22 B1.n15 3.93153
R18670 B1.n19 B1.n9 3.03311
R18671 B1.n50 B1.n12 3.03311
R18672 B1.n60 B1.n8 3.03311
R18673 B1.n74 B1.n73 3.03311
R18674 B1.n47 B1.n35 3.03311
R18675 B1.n3 B1.n0 2.2714
R18676 B1.n58 B1.n7 2.25261
R18677 B1.n20 B1.n10 2.25256
R18678 B1.n34 B1.n33 2.25127
R18679 B1.n37 B1.n33 2.24434
R18680 B1.n73 B1.n72 1.88285
R18681 B1.n30 B1.n12 1.88285
R18682 B1.n45 B1.n35 1.50638
R18683 B1.n63 B1.n60 1.50638
R18684 B1.n19 B1.n18 1.50638
R18685 B1.n16 B1.n10 1.49213
R18686 B1.n70 B1.n69 1.49212
R18687 B1.n61 B1.n7 1.49182
R18688 B1.n14 B1.n13 1.49166
R18689 B1.n78 B1 0.946182
R18690 B1.n65 B1.n64 0.753441
R18691 B1.n24 B1.n23 0.753441
R18692 B1.n44 B1.n40 0.521921
R18693 B1.n78 B1 0.368241
R18694 B1.n77 B1.n6 0.29767
R18695 B1.n49 B1.n48 0.238951
R18696 B1.n77 B1.n76 0.196255
R18697 B1 B1.n77 0.1855
R18698 B1.n6 B1.n5 0.149538
R18699 B1.n75 B1.n51 0.124821
R18700 B1 B1.n78 0.063
R18701 B1.n42 B1.n32 0.0579027
R18702 B1.n62 B1.n61 0.0396286
R18703 B1.n17 B1.n16 0.0383668
R18704 B1.n46 B1.n37 0.0314092
R18705 B1.n5 B1.n0 0.0281442
R18706 B1.n39 B1.n37 0.0271357
R18707 B1.n61 B1.n52 0.0202788
R18708 B1.n16 B1.n11 0.0196501
R18709 B1.n51 B1.n10 0.0168043
R18710 B1.n36 B1.n33 0.016125
R18711 B1.n74 B1.n52 0.013431
R18712 B1.n70 B1.n54 0.013431
R18713 B1.n50 B1.n11 0.013
R18714 B1.n31 B1.n13 0.013
R18715 B1.n38 B1.n32 0.0122521
R18716 B1.n58 B1.n8 0.0117689
R18717 B1.n20 B1.n9 0.0114102
R18718 B1.n47 B1.n34 0.0100704
R18719 B1.n76 B1.n7 0.0100109
R18720 B1.n74 B1.n54 0.00588793
R18721 B1.n50 B1.n31 0.00570833
R18722 B1.n62 B1.n8 0.00481034
R18723 B1.n47 B1.n46 0.0047735
R18724 B1.n17 B1.n9 0.00466667
R18725 B1.n53 B1.n7 0.00457609
R18726 B1.n76 B1.n75 0.00457609
R18727 B1.n2 B1.n0 0.00410577
R18728 B1.n39 B1.n38 0.00370513
R18729 B1.n48 B1.n33 0.00253804
R18730 B1.n4 B1.n3 0.00185919
R18731 B1.n49 B1.n10 0.0018587
R18732 a_2221_8623.n79 a_2221_8623.t9 60.2505
R18733 a_2221_8623.n57 a_2221_8623.t6 60.2505
R18734 a_2221_8623.n43 a_2221_8623.t8 60.2505
R18735 a_2221_8623.n21 a_2221_8623.t7 60.2505
R18736 a_2221_8623.n0 a_2221_8623.n131 9.3005
R18737 a_2221_8623.n0 a_2221_8623.n129 9.3005
R18738 a_2221_8623.n4 a_2221_8623.n65 9.3005
R18739 a_2221_8623.n4 a_2221_8623.n66 9.3005
R18740 a_2221_8623.n4 a_2221_8623.n64 9.3005
R18741 a_2221_8623.n64 a_2221_8623.n63 9.3005
R18742 a_2221_8623.n5 a_2221_8623.n72 9.3005
R18743 a_2221_8623.n6 a_2221_8623.n89 9.3005
R18744 a_2221_8623.n5 a_2221_8623.n78 9.3005
R18745 a_2221_8623.n78 a_2221_8623.n77 9.3005
R18746 a_2221_8623.n5 a_2221_8623.n71 9.3005
R18747 a_2221_8623.n6 a_2221_8623.n87 9.3005
R18748 a_2221_8623.n87 a_2221_8623.n86 9.3005
R18749 a_2221_8623.n6 a_2221_8623.n88 9.3005
R18750 a_2221_8623.n3 a_2221_8623.n29 9.3005
R18751 a_2221_8623.n3 a_2221_8623.n30 9.3005
R18752 a_2221_8623.n3 a_2221_8623.n28 9.3005
R18753 a_2221_8623.n28 a_2221_8623.n27 9.3005
R18754 a_2221_8623.n2 a_2221_8623.n36 9.3005
R18755 a_2221_8623.n2 a_2221_8623.n42 9.3005
R18756 a_2221_8623.n42 a_2221_8623.n41 9.3005
R18757 a_2221_8623.n2 a_2221_8623.n35 9.3005
R18758 a_2221_8623.n1 a_2221_8623.n51 9.3005
R18759 a_2221_8623.n51 a_2221_8623.n50 9.3005
R18760 a_2221_8623.n1 a_2221_8623.n53 9.3005
R18761 a_2221_8623.n1 a_2221_8623.n52 9.3005
R18762 a_2221_8623.n8 a_2221_8623.n19 9.3005
R18763 a_2221_8623.n7 a_2221_8623.n14 9.3005
R18764 a_2221_8623.n162 a_2221_8623.n159 9.3005
R18765 a_2221_8623.n162 a_2221_8623.n160 9.3005
R18766 a_2221_8623.n80 a_2221_8623.n79 8.76429
R18767 a_2221_8623.n44 a_2221_8623.n43 8.76429
R18768 a_2221_8623.n85 a_2221_8623.n84 7.45411
R18769 a_2221_8623.n76 a_2221_8623.n75 7.45411
R18770 a_2221_8623.n62 a_2221_8623.n61 7.45411
R18771 a_2221_8623.n40 a_2221_8623.n39 7.45411
R18772 a_2221_8623.n49 a_2221_8623.n48 7.45411
R18773 a_2221_8623.n26 a_2221_8623.n25 7.45411
R18774 a_2221_8623.n58 a_2221_8623.n57 6.80105
R18775 a_2221_8623.n22 a_2221_8623.n21 6.80105
R18776 a_2221_8623.n83 a_2221_8623.n82 5.64756
R18777 a_2221_8623.n74 a_2221_8623.n73 5.64756
R18778 a_2221_8623.n60 a_2221_8623.n59 5.64756
R18779 a_2221_8623.n38 a_2221_8623.n37 5.64756
R18780 a_2221_8623.n47 a_2221_8623.n46 5.64756
R18781 a_2221_8623.n24 a_2221_8623.n23 5.64756
R18782 a_2221_8623.n112 a_2221_8623.t2 5.5395
R18783 a_2221_8623.n112 a_2221_8623.t1 5.5395
R18784 a_2221_8623.t3 a_2221_8623.n162 5.5395
R18785 a_2221_8623.n162 a_2221_8623.t0 5.5395
R18786 a_2221_8623.n70 a_2221_8623.n69 4.73575
R18787 a_2221_8623.n68 a_2221_8623.n67 4.73575
R18788 a_2221_8623.n34 a_2221_8623.n33 4.73575
R18789 a_2221_8623.n32 a_2221_8623.n31 4.73575
R18790 a_2221_8623.n81 a_2221_8623.n80 4.6505
R18791 a_2221_8623.n45 a_2221_8623.n44 4.6505
R18792 a_2221_8623.n135 a_2221_8623.n134 4.51815
R18793 a_2221_8623.n17 a_2221_8623.n16 4.51815
R18794 a_2221_8623.n155 a_2221_8623.n154 4.51815
R18795 a_2221_8623.n0 a_2221_8623.n128 4.5005
R18796 a_2221_8623.n124 a_2221_8623.n133 4.5005
R18797 a_2221_8623.n125 a_2221_8623.n123 4.5005
R18798 a_2221_8623.n118 a_2221_8623.n116 4.5005
R18799 a_2221_8623.n8 a_2221_8623.n12 4.5005
R18800 a_2221_8623.n7 a_2221_8623.n17 4.5005
R18801 a_2221_8623.n102 a_2221_8623.n107 4.5005
R18802 a_2221_8623.n139 a_2221_8623.n147 4.5005
R18803 a_2221_8623.n152 a_2221_8623.n151 4.5005
R18804 a_2221_8623.n138 a_2221_8623.n141 4.5005
R18805 a_2221_8623.n162 a_2221_8623.n161 4.35791
R18806 a_2221_8623.n91 a_2221_8623.n93 4.24504
R18807 a_2221_8623.n54 a_2221_8623.n56 4.24504
R18808 a_2221_8623.n12 a_2221_8623.n11 3.76521
R18809 a_2221_8623.n4 a_2221_8623.n58 3.42768
R18810 a_2221_8623.n3 a_2221_8623.n22 3.42768
R18811 a_2221_8623.n123 a_2221_8623.n119 3.38874
R18812 a_2221_8623.n147 a_2221_8623.n144 3.38874
R18813 a_2221_8623.n131 a_2221_8623.n130 3.38537
R18814 a_2221_8623.n158 a_2221_8623.n157 3.38537
R18815 a_2221_8623.n97 a_2221_8623.t5 3.3065
R18816 a_2221_8623.n97 a_2221_8623.t4 3.3065
R18817 a_2221_8623.n107 a_2221_8623.n105 3.28194
R18818 a_2221_8623.n99 a_2221_8623.n98 3.15821
R18819 a_2221_8623.n117 a_2221_8623.n135 3.03311
R18820 a_2221_8623.n153 a_2221_8623.n155 3.03311
R18821 a_2221_8623.n107 a_2221_8623.n106 3.01226
R18822 a_2221_8623.n12 a_2221_8623.n10 2.63579
R18823 a_2221_8623.n14 a_2221_8623.n13 2.61733
R18824 a_2221_8623.n0 a_2221_8623.n126 2.57914
R18825 a_2221_8623.n122 a_2221_8623.n121 2.25932
R18826 a_2221_8623.n146 a_2221_8623.n145 2.25932
R18827 a_2221_8623.n19 a_2221_8623.n18 2.24766
R18828 a_2221_8623.n116 a_2221_8623.n114 2.22452
R18829 a_2221_8623.n151 a_2221_8623.n149 2.22452
R18830 a_2221_8623.n162 a_2221_8623.n148 1.99078
R18831 a_2221_8623.n17 a_2221_8623.n15 1.88285
R18832 a_2221_8623.n113 a_2221_8623.n112 1.72048
R18833 a_2221_8623.n99 a_2221_8623.n97 1.61799
R18834 a_2221_8623.n108 a_2221_8623.n96 1.51434
R18835 a_2221_8623.n96 a_2221_8623.n8 1.51334
R18836 a_2221_8623.n128 a_2221_8623.n127 1.50638
R18837 a_2221_8623.n159 a_2221_8623.n158 1.50638
R18838 a_2221_8623.n142 a_2221_8623.n143 1.50638
R18839 a_2221_8623.n101 a_2221_8623.n100 1.12991
R18840 a_2221_8623.n95 a_2221_8623.n94 3.28829
R18841 a_2221_8623.n86 a_2221_8623.n85 0.994314
R18842 a_2221_8623.n77 a_2221_8623.n76 0.994314
R18843 a_2221_8623.n63 a_2221_8623.n62 0.994314
R18844 a_2221_8623.n41 a_2221_8623.n40 0.994314
R18845 a_2221_8623.n50 a_2221_8623.n49 0.994314
R18846 a_2221_8623.n27 a_2221_8623.n26 0.994314
R18847 a_2221_8623.n111 a_2221_8623.n156 0.829361
R18848 a_2221_8623.n133 a_2221_8623.n132 0.753441
R18849 a_2221_8623.n87 a_2221_8623.n83 0.753441
R18850 a_2221_8623.n78 a_2221_8623.n74 0.753441
R18851 a_2221_8623.n64 a_2221_8623.n60 0.753441
R18852 a_2221_8623.n42 a_2221_8623.n38 0.753441
R18853 a_2221_8623.n51 a_2221_8623.n47 0.753441
R18854 a_2221_8623.n28 a_2221_8623.n24 0.753441
R18855 a_2221_8623.n141 a_2221_8623.n140 0.753441
R18856 a_2221_8623.n137 a_2221_8623.n136 0.754708
R18857 a_2221_8623.n93 a_2221_8623.n92 0.709906
R18858 a_2221_8623.n56 a_2221_8623.n55 0.709906
R18859 a_2221_8623.n109 a_2221_8623.n137 0.678625
R18860 a_2221_8623.n70 a_2221_8623.n68 0.458354
R18861 a_2221_8623.n34 a_2221_8623.n32 0.458354
R18862 a_2221_8623.n123 a_2221_8623.n122 0.376971
R18863 a_2221_8623.n121 a_2221_8623.n120 0.376971
R18864 a_2221_8623.n104 a_2221_8623.n103 0.376971
R18865 a_2221_8623.n147 a_2221_8623.n146 0.376971
R18866 a_2221_8623.n95 a_2221_8623.n20 0.242354
R18867 a_2221_8623.n136 a_2221_8623.n113 0.225683
R18868 a_2221_8623.n108 a_2221_8623.n99 0.224119
R18869 a_2221_8623.n6 a_2221_8623.n81 0.190717
R18870 a_2221_8623.n81 a_2221_8623.n5 0.190717
R18871 a_2221_8623.n45 a_2221_8623.n2 0.190717
R18872 a_2221_8623.n1 a_2221_8623.n45 0.190717
R18873 a_2221_8623.n94 a_2221_8623.n54 0.159981
R18874 a_2221_8623.n94 a_2221_8623.n91 0.159717
R18875 a_2221_8623.n138 a_2221_8623.n142 4.63429
R18876 a_2221_8623.n105 a_2221_8623.n104 0.0902327
R18877 a_2221_8623.n117 a_2221_8623.n125 0.0900802
R18878 a_2221_8623.n136 a_2221_8623.n118 0.0608541
R18879 a_2221_8623.n111 a_2221_8623.n110 0.0528649
R18880 a_2221_8623.n156 a_2221_8623.n153 0.0511262
R18881 a_2221_8623.n156 a_2221_8623.n139 0.040511
R18882 a_2221_8623.n114 a_2221_8623.n115 0.0303633
R18883 a_2221_8623.n149 a_2221_8623.n150 0.0303633
R18884 a_2221_8623.n102 a_2221_8623.n101 4.54542
R18885 a_2221_8623.n152 a_2221_8623.n148 0.0122188
R18886 a_2221_8623.n153 a_2221_8623.n152 0.0454219
R18887 a_2221_8623.n139 a_2221_8623.n138 0.0454219
R18888 a_2221_8623.n118 a_2221_8623.n117 0.0454219
R18889 a_2221_8623.n125 a_2221_8623.n124 0.0454219
R18890 a_2221_8623.n111 a_2221_8623.n109 0.022561
R18891 a_2221_8623.n111 a_2221_8623.n20 0.847626
R18892 a_2221_8623.n108 a_2221_8623.n102 0.0883906
R18893 a_2221_8623.n96 a_2221_8623.n95 0.905839
R18894 a_2221_8623.n91 a_2221_8623.n90 0.0410417
R18895 a_2221_8623.n8 a_2221_8623.n9 2.77239
R18896 a_2221_8623.n5 a_2221_8623.n70 0.205546
R18897 a_2221_8623.n68 a_2221_8623.n4 0.205546
R18898 a_2221_8623.n32 a_2221_8623.n3 0.205546
R18899 a_2221_8623.n2 a_2221_8623.n34 0.205546
R18900 a_2221_8623.n54 a_2221_8623.n1 0.177485
R18901 a_2221_8623.n124 a_2221_8623.n0 0.171838
R18902 a_2221_8623.n8 a_2221_8623.n7 0.167464
R18903 a_2221_8623.n90 a_2221_8623.n6 0.137941
R18904 comparator_top_0.comparator_bias_0.VBP.n29 comparator_top_0.comparator_bias_0.VBP.t3 116.841
R18905 comparator_top_0.comparator_bias_0.VBP.n56 comparator_top_0.comparator_bias_0.VBP.t2 60.2505
R18906 comparator_top_0.comparator_bias_0.VBP.n98 comparator_top_0.comparator_bias_0.VBP.t4 60.2505
R18907 comparator_top_0.comparator_bias_0.VBP.n110 comparator_top_0.comparator_bias_0.VBP.t5 60.2505
R18908 comparator_top_0.comparator_bias_0.VBP.n33 comparator_top_0.comparator_bias_0.VBP.n32 52.6902
R18909 comparator_top_0.comparator_bias_0.VBP.n41 comparator_top_0.comparator_bias_0.VBP.n40 46.104
R18910 comparator_top_0.comparator_bias_0.VBP.n89 comparator_top_0.comparator_bias_0.VBP.n88 39.5177
R18911 comparator_top_0.comparator_bias_0.VBP.n81 comparator_top_0.comparator_bias_0.VBP.n80 32.9315
R18912 comparator_top_0.comparator_bias_0.VBP.n72 comparator_top_0.comparator_bias_0.VBP.n71 29.6384
R18913 comparator_top_0.comparator_bias_0.VBP.n71 comparator_top_0.comparator_bias_0.VBP.n70 26.3453
R18914 comparator_top_0.comparator_bias_0.VBP.n82 comparator_top_0.comparator_bias_0.VBP.n81 23.0522
R18915 comparator_top_0.comparator_bias_0.VBP.n90 comparator_top_0.comparator_bias_0.VBP.n89 16.466
R18916 comparator_top_0.comparator_bias_0.VBP.n42 comparator_top_0.comparator_bias_0.VBP.n41 9.87981
R18917 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n36 9.3005
R18918 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n44 9.3005
R18919 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n43 9.3005
R18920 comparator_top_0.comparator_bias_0.VBP.n43 comparator_top_0.comparator_bias_0.VBP.n42 9.3005
R18921 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n37 9.3005
R18922 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n35 9.3005
R18923 comparator_top_0.comparator_bias_0.VBP.n35 comparator_top_0.comparator_bias_0.VBP.n34 9.3005
R18924 comparator_top_0.comparator_bias_0.VBP.n8 comparator_top_0.comparator_bias_0.VBP.n76 9.3005
R18925 comparator_top_0.comparator_bias_0.VBP.n83 comparator_top_0.comparator_bias_0.VBP.n82 9.3005
R18926 comparator_top_0.comparator_bias_0.VBP.n91 comparator_top_0.comparator_bias_0.VBP.n90 9.3005
R18927 comparator_top_0.comparator_bias_0.VBP.n8 comparator_top_0.comparator_bias_0.VBP.n73 9.3005
R18928 comparator_top_0.comparator_bias_0.VBP.n73 comparator_top_0.comparator_bias_0.VBP.n72 9.3005
R18929 comparator_top_0.comparator_bias_0.VBP.n65 comparator_top_0.comparator_bias_0.VBP.n64 9.3005
R18930 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n59 9.3005
R18931 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n48 9.3005
R18932 comparator_top_0.comparator_bias_0.VBP.n54 comparator_top_0.comparator_bias_0.VBP.n53 9.3005
R18933 comparator_top_0.comparator_bias_0.VBP.n4 comparator_top_0.comparator_bias_0.VBP.n107 9.3005
R18934 comparator_top_0.comparator_bias_0.VBP.n4 comparator_top_0.comparator_bias_0.VBP.n105 9.3005
R18935 comparator_top_0.comparator_bias_0.VBP.n105 comparator_top_0.comparator_bias_0.VBP.n104 9.3005
R18936 comparator_top_0.comparator_bias_0.VBP.n4 comparator_top_0.comparator_bias_0.VBP.n106 9.3005
R18937 comparator_top_0.comparator_bias_0.VBP.n5 comparator_top_0.comparator_bias_0.VBP.n117 9.3005
R18938 comparator_top_0.comparator_bias_0.VBP.n117 comparator_top_0.comparator_bias_0.VBP.n116 9.3005
R18939 comparator_top_0.comparator_bias_0.VBP.n5 comparator_top_0.comparator_bias_0.VBP.n119 9.3005
R18940 comparator_top_0.comparator_bias_0.VBP.n5 comparator_top_0.comparator_bias_0.VBP.n118 9.3005
R18941 comparator_top_0.comparator_bias_0.VBP.n6 comparator_top_0.comparator_bias_0.VBP.n18 9.3005
R18942 comparator_top_0.comparator_bias_0.VBP.n6 comparator_top_0.comparator_bias_0.VBP.n13 9.3005
R18943 comparator_top_0.comparator_bias_0.VBP.n57 comparator_top_0.comparator_bias_0.VBP.n56 8.76429
R18944 comparator_top_0.comparator_bias_0.VBP.n52 comparator_top_0.comparator_bias_0.VBP.n51 7.45411
R18945 comparator_top_0.comparator_bias_0.VBP.n63 comparator_top_0.comparator_bias_0.VBP.n62 7.45411
R18946 comparator_top_0.comparator_bias_0.VBP.n103 comparator_top_0.comparator_bias_0.VBP.n102 7.45411
R18947 comparator_top_0.comparator_bias_0.VBP.n115 comparator_top_0.comparator_bias_0.VBP.n114 7.45411
R18948 comparator_top_0.comparator_bias_0.VBP.n99 comparator_top_0.comparator_bias_0.VBP.n98 6.80105
R18949 comparator_top_0.comparator_bias_0.VBP.n111 comparator_top_0.comparator_bias_0.VBP.n110 6.801
R18950 comparator_top_0.comparator_bias_0.VBP.n31 comparator_top_0.comparator_bias_0.VBP.n30 6.02403
R18951 comparator_top_0.comparator_bias_0.VBP.n2 comparator_top_0.comparator_bias_0.VBP.n93 6.0005
R18952 comparator_top_0.comparator_bias_0.VBP.n2 comparator_top_0.comparator_bias_0.VBP.n86 6.0005
R18953 comparator_top_0.comparator_bias_0.VBP.n50 comparator_top_0.comparator_bias_0.VBP.n49 5.64756
R18954 comparator_top_0.comparator_bias_0.VBP.n61 comparator_top_0.comparator_bias_0.VBP.n60 5.64756
R18955 comparator_top_0.comparator_bias_0.VBP.n101 comparator_top_0.comparator_bias_0.VBP.n100 5.64756
R18956 comparator_top_0.comparator_bias_0.VBP.n113 comparator_top_0.comparator_bias_0.VBP.n112 5.64756
R18957 comparator_top_0.comparator_bias_0.VBP.n39 comparator_top_0.comparator_bias_0.VBP.n38 5.27109
R18958 comparator_top_0.comparator_bias_0.VBP.n10 comparator_top_0.comparator_bias_0.VBP.n69 5.25098
R18959 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n47 4.88281
R18960 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n58 4.88086
R18961 comparator_top_0.comparator_bias_0.VBP.n1 comparator_top_0.comparator_bias_0.VBP.n9 4.54542
R18962 comparator_top_0.comparator_bias_0.VBP.n16 comparator_top_0.comparator_bias_0.VBP.n15 4.51815
R18963 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n55 4.5005
R18964 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n66 4.5005
R18965 comparator_top_0.comparator_bias_0.VBP.n8 comparator_top_0.comparator_bias_0.VBP.n78 4.5005
R18966 comparator_top_0.comparator_bias_0.VBP.n10 comparator_top_0.comparator_bias_0.VBP.n68 4.5005
R18967 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n46 4.5005
R18968 comparator_top_0.comparator_bias_0.VBP.n6 comparator_top_0.comparator_bias_0.VBP.n16 4.5005
R18969 comparator_top_0.comparator_bias_0.VBP.n6 comparator_top_0.comparator_bias_0.VBP.n21 4.5005
R18970 comparator_top_0.comparator_bias_0.VBP.n1 comparator_top_0.comparator_bias_0.VBP.n26 4.5005
R18971 comparator_top_0.comparator_bias_0.VBP.n4 comparator_top_0.comparator_bias_0.VBP.n97 4.24504
R18972 comparator_top_0.comparator_bias_0.VBP.n5 comparator_top_0.comparator_bias_0.VBP.n109 4.24504
R18973 comparator_top_0.comparator_bias_0.VBP.n3 comparator_top_0.comparator_bias_0.VBP.n29 4.23684
R18974 comparator_top_0.comparator_bias_0.VBP.n93 comparator_top_0.comparator_bias_0.VBP.n87 4.14168
R18975 comparator_top_0.comparator_bias_0.VBP.n21 comparator_top_0.comparator_bias_0.VBP.n20 3.76521
R18976 comparator_top_0.comparator_bias_0.VBP.n5 comparator_top_0.comparator_bias_0.VBP.n111 3.42853
R18977 comparator_top_0.comparator_bias_0.VBP.n4 comparator_top_0.comparator_bias_0.VBP.n99 3.42768
R18978 comparator_top_0.comparator_bias_0.VBP.n86 comparator_top_0.comparator_bias_0.VBP.n79 3.38874
R18979 comparator_top_0.comparator_bias_0.VBP.n27 comparator_top_0.comparator_bias_0.VBP.t1 3.3065
R18980 comparator_top_0.comparator_bias_0.VBP.n27 comparator_top_0.comparator_bias_0.VBP.t0 3.3065
R18981 comparator_top_0.comparator_bias_0.VBP.n34 comparator_top_0.comparator_bias_0.VBP.n33 3.2936
R18982 comparator_top_0.comparator_bias_0.VBP.n26 comparator_top_0.comparator_bias_0.VBP.n24 3.74814
R18983 comparator_top_0.comparator_bias_0.VBP comparator_top_0.comparator_bias_0.VBP.n95 3.26842
R18984 comparator_top_0.comparator_bias_0.VBP.n1 comparator_top_0.comparator_bias_0.VBP.n28 3.15814
R18985 comparator_top_0.comparator_bias_0.VBP.n0 comparator_top_0.comparator_bias_0.VBP.n57 3.03311
R18986 comparator_top_0.comparator_bias_0.VBP.n75 comparator_top_0.comparator_bias_0.VBP.n74 3.01226
R18987 comparator_top_0.comparator_bias_0.VBP.n26 comparator_top_0.comparator_bias_0.VBP.n25 3.01226
R18988 comparator_top_0.comparator_bias_0.VBP.n6 comparator_top_0.comparator_bias_0.VBP.n11 2.77255
R18989 comparator_top_0.comparator_bias_0.VBP.n21 comparator_top_0.comparator_bias_0.VBP.n19 2.63579
R18990 comparator_top_0.comparator_bias_0.VBP.n13 comparator_top_0.comparator_bias_0.VBP.n12 2.61733
R18991 comparator_top_0.comparator_bias_0.VBP.n85 comparator_top_0.comparator_bias_0.VBP.n84 2.25932
R18992 comparator_top_0.comparator_bias_0.VBP.n18 comparator_top_0.comparator_bias_0.VBP.n17 2.24766
R18993 comparator_top_0.comparator_bias_0.VBP.n92 comparator_top_0.comparator_bias_0.VBP.n91 1.88285
R18994 comparator_top_0.comparator_bias_0.VBP.n76 comparator_top_0.comparator_bias_0.VBP.n75 1.88285
R18995 comparator_top_0.comparator_bias_0.VBP.n16 comparator_top_0.comparator_bias_0.VBP.n14 1.88285
R18996 comparator_top_0.comparator_bias_0.VBP.n7 comparator_top_0.comparator_bias_0.VBP.n0 1.85011
R18997 comparator_top_0.comparator_bias_0.VBP.n22 comparator_top_0.comparator_bias_0.VBP.n1 1.82596
R18998 comparator_top_0.comparator_bias_0.VBP.n120 comparator_top_0.comparator_bias_0.VBP.n5 1.75631
R18999 comparator_top_0.comparator_bias_0.VBP.n2 comparator_top_0.comparator_bias_0.VBP.n3 1.74716
R19000 comparator_top_0.comparator_bias_0.VBP.n22 comparator_top_0.comparator_bias_0.VBP.n6 1.6803
R19001 comparator_top_0.comparator_bias_0.VBP.n1 comparator_top_0.comparator_bias_0.VBP.n27 1.61775
R19002 comparator_top_0.comparator_bias_0.VBP.n2 comparator_top_0.comparator_bias_0.VBP.n8 1.60792
R19003 comparator_top_0.comparator_bias_0.VBP.n2 comparator_top_0.comparator_bias_0.VBP.n10 1.55128
R19004 comparator_top_0.comparator_bias_0.VBP.n68 comparator_top_0.comparator_bias_0.VBP.n67 1.50638
R19005 comparator_top_0.comparator_bias_0.VBP comparator_top_0.comparator_bias_0.VBP.n120 1.3155
R19006 comparator_top_0.comparator_bias_0.VBP.n43 comparator_top_0.comparator_bias_0.VBP.n39 1.12991
R19007 comparator_top_0.comparator_bias_0.VBP.n9 comparator_top_0.comparator_bias_0.VBP.n23 1.12991
R19008 comparator_top_0.comparator_bias_0.VBP.n95 comparator_top_0.comparator_bias_0.VBP.n22 1.04295
R19009 comparator_top_0.comparator_bias_0.VBP.n53 comparator_top_0.comparator_bias_0.VBP.n52 0.994314
R19010 comparator_top_0.comparator_bias_0.VBP.n64 comparator_top_0.comparator_bias_0.VBP.n63 0.994314
R19011 comparator_top_0.comparator_bias_0.VBP.n104 comparator_top_0.comparator_bias_0.VBP.n103 0.994314
R19012 comparator_top_0.comparator_bias_0.VBP.n116 comparator_top_0.comparator_bias_0.VBP.n115 0.994314
R19013 comparator_top_0.comparator_bias_0.VBP.n94 comparator_top_0.comparator_bias_0.VBP.n2 0.794925
R19014 comparator_top_0.comparator_bias_0.VBP.n46 comparator_top_0.comparator_bias_0.VBP.n45 0.753441
R19015 comparator_top_0.comparator_bias_0.VBP.n78 comparator_top_0.comparator_bias_0.VBP.n77 0.753441
R19016 comparator_top_0.comparator_bias_0.VBP.n55 comparator_top_0.comparator_bias_0.VBP.n54 0.753441
R19017 comparator_top_0.comparator_bias_0.VBP.n54 comparator_top_0.comparator_bias_0.VBP.n50 0.753441
R19018 comparator_top_0.comparator_bias_0.VBP.n65 comparator_top_0.comparator_bias_0.VBP.n61 0.753441
R19019 comparator_top_0.comparator_bias_0.VBP.n66 comparator_top_0.comparator_bias_0.VBP.n65 0.753441
R19020 comparator_top_0.comparator_bias_0.VBP.n105 comparator_top_0.comparator_bias_0.VBP.n101 0.753441
R19021 comparator_top_0.comparator_bias_0.VBP.n117 comparator_top_0.comparator_bias_0.VBP.n113 0.753441
R19022 comparator_top_0.comparator_bias_0.VBP.n2 comparator_top_0.comparator_bias_0.VBP.n7 0.748981
R19023 comparator_top_0.comparator_bias_0.VBP.n97 comparator_top_0.comparator_bias_0.VBP.n96 0.709906
R19024 comparator_top_0.comparator_bias_0.VBP.n109 comparator_top_0.comparator_bias_0.VBP.n108 0.709906
R19025 comparator_top_0.comparator_bias_0.VBP.n5 comparator_top_0.comparator_bias_0.VBP.n4 0.673704
R19026 comparator_top_0.comparator_bias_0.VBP.n95 comparator_top_0.comparator_bias_0.VBP.n94 0.577213
R19027 comparator_top_0.comparator_bias_0.VBP.n7 comparator_top_0.comparator_bias_0.VBP 0.538902
R19028 comparator_top_0.comparator_bias_0.VBP.n35 comparator_top_0.comparator_bias_0.VBP.n31 0.376971
R19029 comparator_top_0.comparator_bias_0.VBP.n93 comparator_top_0.comparator_bias_0.VBP.n92 0.376971
R19030 comparator_top_0.comparator_bias_0.VBP.n86 comparator_top_0.comparator_bias_0.VBP.n85 0.376971
R19031 comparator_top_0.comparator_bias_0.VBP.n84 comparator_top_0.comparator_bias_0.VBP.n83 0.376971
R19032 a_2093_3714.n47 a_2093_3714.n46 6.31679
R19033 a_2093_3714.n7 a_2093_3714.n41 6.12797
R19034 a_2093_3714.n1 a_2093_3714.n19 6.12763
R19035 a_2093_3714.n3 a_2093_3714.n25 6.12763
R19036 a_2093_3714.n17 a_2093_3714.t4 5.5395
R19037 a_2093_3714.n17 a_2093_3714.t2 5.5395
R19038 a_2093_3714.n23 a_2093_3714.t3 5.5395
R19039 a_2093_3714.n23 a_2093_3714.t1 5.5395
R19040 a_2093_3714.n29 a_2093_3714.t0 5.5395
R19041 a_2093_3714.n29 a_2093_3714.t10 5.5395
R19042 a_2093_3714.n34 a_2093_3714.t9 5.5395
R19043 a_2093_3714.n34 a_2093_3714.t8 5.5395
R19044 a_2093_3714.n36 a_2093_3714.t6 5.5395
R19045 a_2093_3714.n36 a_2093_3714.t7 5.5395
R19046 a_2093_3714.n51 a_2093_3714.t11 5.5395
R19047 a_2093_3714.t5 a_2093_3714.n51 5.5395
R19048 a_2093_3714.n49 a_2093_3714.n48 5.26941
R19049 a_2093_3714.n4 a_2093_3714.n33 4.5005
R19050 a_2093_3714.n6 a_2093_3714.n40 4.5005
R19051 a_2093_3714.n2 a_2093_3714.n22 4.5005
R19052 a_2093_3714.n5 a_2093_3714.n28 4.5005
R19053 a_2093_3714.n0 a_2093_3714.n16 4.5005
R19054 a_2093_3714.n9 a_2093_3714.n45 4.5005
R19055 a_2093_3714.n8 a_2093_3714.n43 4.5005
R19056 a_2093_3714.n51 a_2093_3714.n50 4.27411
R19057 a_2093_3714.n16 a_2093_3714.n14 3.76521
R19058 a_2093_3714.n22 a_2093_3714.n20 3.76521
R19059 a_2093_3714.n28 a_2093_3714.n26 3.76521
R19060 a_2093_3714.n33 a_2093_3714.n31 3.76521
R19061 a_2093_3714.n40 a_2093_3714.n38 3.76521
R19062 a_2093_3714.n45 a_2093_3714.n44 3.76521
R19063 a_2093_3714.n43 a_2093_3714.n42 3.01226
R19064 a_2093_3714.n16 a_2093_3714.n15 2.63579
R19065 a_2093_3714.n22 a_2093_3714.n21 2.63579
R19066 a_2093_3714.n28 a_2093_3714.n27 2.63579
R19067 a_2093_3714.n33 a_2093_3714.n32 2.63579
R19068 a_2093_3714.n40 a_2093_3714.n39 2.63579
R19069 a_2093_3714.n12 a_2093_3714.n1 2.20191
R19070 a_2093_3714.n10 a_2093_3714.n7 2.18375
R19071 a_2093_3714.n50 a_2093_3714.n49 1.8965
R19072 a_2093_3714.n8 a_2093_3714.n10 1.56196
R19073 a_2093_3714.n11 a_2093_3714.n4 1.74534
R19074 a_2093_3714.n12 a_2093_3714.n3 1.48434
R19075 a_2093_3714.n13 a_2093_3714.n5 1.745
R19076 a_2093_3714.n5 a_2093_3714.n30 1.4669
R19077 a_2093_3714.n6 a_2093_3714.n37 1.4669
R19078 a_2093_3714.n0 a_2093_3714.n18 1.46689
R19079 a_2093_3714.n2 a_2093_3714.n24 1.46689
R19080 a_2093_3714.n4 a_2093_3714.n35 1.46689
R19081 a_2093_3714.n47 a_2093_3714.n9 1.46687
R19082 a_2093_3714.n10 a_2093_3714.n11 0.753593
R19083 a_2093_3714.n11 a_2093_3714.n13 0.718062
R19084 a_2093_3714.n13 a_2093_3714.n12 0.700686
R19085 a_2093_3714.n30 a_2093_3714.n29 0.400769
R19086 a_2093_3714.n37 a_2093_3714.n36 0.400769
R19087 a_2093_3714.n18 a_2093_3714.n17 0.400768
R19088 a_2093_3714.n24 a_2093_3714.n23 0.400768
R19089 a_2093_3714.n35 a_2093_3714.n34 0.400768
R19090 a_2093_3714.n51 a_2093_3714.n47 0.40076
R19091 a_2093_3714.n1 a_2093_3714.n0 0.261498
R19092 a_2093_3714.n3 a_2093_3714.n2 0.261477
R19093 a_2093_3714.n7 a_2093_3714.n6 0.261136
R19094 a_2093_3714.n9 a_2093_3714.n8 0.183856
R19095 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 136.804
R19096 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 136.325
R19097 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 119.999
R19098 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 93.9023
R19099 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 93.3044
R19100 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 93.0848
R19101 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n4 92.5005
R19102 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 92.4623
R19103 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 69.2281
R19104 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 29.4833
R19105 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 27.6955
R19106 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 27.6955
R19107 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 15.4626
R19108 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n16 9.3005
R19109 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n8 9.3005
R19110 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n7 9.3005
R19111 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 9.3005
R19112 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 9.3005
R19113 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n15 9.3005
R19114 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n17 9.3005
R19115 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 9.02061
R19116 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 9.02061
R19117 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n34 8.28285
R19118 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n21 8.28285
R19119 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 5.64756
R19120 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 5.31864
R19121 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n42 4.14168
R19122 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n28 4.14168
R19123 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 4.06959
R19124 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n11 3.93153
R19125 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n40 3.76521
R19126 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n33 3.76521
R19127 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n24 3.76521
R19128 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n19 3.76521
R19129 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n36 3.38874
R19130 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n22 3.38874
R19131 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 3.0736
R19132 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 3.07249
R19133 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 3.07078
R19134 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 3.04338
R19135 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 3.03311
R19136 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 3.03311
R19137 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 3.03311
R19138 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n39 2.63579
R19139 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n20 2.63579
R19140 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 2.27447
R19141 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 2.25932
R19142 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 2.25932
R19143 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 1.80772
R19144 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n30 1.61433
R19145 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 1.45534
R19146 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 1.19419
R19147 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n9 0.753441
R19148 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 0.719888
R19149 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 0.22499
R19150 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 0.176176
R19151 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 2.36361
R19152 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 2.36353
R19153 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 1.14499
R19154 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 1.00043
R19155 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 120.01
R19156 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 92.9415
R19157 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n4 92.5005
R19158 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 92.4623
R19159 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 73.195
R19160 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 72.1651
R19161 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 29.4833
R19162 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 27.6955
R19163 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 27.6955
R19164 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 15.4607
R19165 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 9.3005
R19166 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 9.3005
R19167 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 9.02061
R19168 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 9.01961
R19169 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n26 8.28285
R19170 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n16 8.28285
R19171 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 5.64756
R19172 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 5.32161
R19173 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 5.31894
R19174 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n31 4.14168
R19175 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n23 4.14168
R19176 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n19 4.14168
R19177 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 4.03426
R19178 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n9 3.93153
R19179 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n33 3.76521
R19180 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n14 3.76521
R19181 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 3.20519
R19182 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 3.07304
R19183 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 3.04478
R19184 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 3.03311
R19185 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 3.03311
R19186 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 3.03311
R19187 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n27 3.01226
R19188 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n17 3.01226
R19189 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n34 2.63579
R19190 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n15 2.63579
R19191 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 2.47579
R19192 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 2.27623
R19193 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 2.25932
R19194 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 2.25932
R19195 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 1.51198
R19196 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 1.15307
R19197 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 1.04295
R19198 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n7 0.753441
R19199 a_2151_594.n7 a_2151_594.t0 60.2505
R19200 a_2151_594.n64 a_2151_594.t2 60.2505
R19201 a_2151_594.n21 a_2151_594.t9 60.2505
R19202 a_2151_594.n42 a_2151_594.t8 60.2505
R19203 a_2151_594.n4 a_2151_594.n73 9.3005
R19204 a_2151_594.n3 a_2151_594.n57 9.3005
R19205 a_2151_594.n2 a_2151_594.n51 9.3005
R19206 a_2151_594.n1 a_2151_594.n35 9.3005
R19207 a_2151_594.n1 a_2151_594.n34 9.3005
R19208 a_2151_594.n2 a_2151_594.n52 9.3005
R19209 a_2151_594.n2 a_2151_594.n50 9.3005
R19210 a_2151_594.n50 a_2151_594.n49 9.3005
R19211 a_2151_594.n1 a_2151_594.n41 9.3005
R19212 a_2151_594.n41 a_2151_594.n40 9.3005
R19213 a_2151_594.n0 a_2151_594.n29 9.3005
R19214 a_2151_594.n0 a_2151_594.n30 9.3005
R19215 a_2151_594.n0 a_2151_594.n28 9.3005
R19216 a_2151_594.n28 a_2151_594.n27 9.3005
R19217 a_2151_594.n4 a_2151_594.n74 9.3005
R19218 a_2151_594.n4 a_2151_594.n72 9.3005
R19219 a_2151_594.n72 a_2151_594.n71 9.3005
R19220 a_2151_594.n3 a_2151_594.n63 9.3005
R19221 a_2151_594.n63 a_2151_594.n62 9.3005
R19222 a_2151_594.n3 a_2151_594.n56 9.3005
R19223 a_2151_594.n5 a_2151_594.n14 9.3005
R19224 a_2151_594.n14 a_2151_594.n13 9.3005
R19225 a_2151_594.n5 a_2151_594.n16 9.3005
R19226 a_2151_594.n5 a_2151_594.n15 9.3005
R19227 a_2151_594.n43 a_2151_594.n42 8.76429
R19228 a_2151_594.n65 a_2151_594.n64 8.76429
R19229 a_2151_594.n26 a_2151_594.n25 8.21641
R19230 a_2151_594.n48 a_2151_594.n47 8.21641
R19231 a_2151_594.n39 a_2151_594.n38 8.21641
R19232 a_2151_594.n70 a_2151_594.n69 8.21641
R19233 a_2151_594.n61 a_2151_594.n60 8.21641
R19234 a_2151_594.n12 a_2151_594.n11 8.21641
R19235 a_2151_594.n22 a_2151_594.n21 6.92011
R19236 a_2151_594.n8 a_2151_594.n7 6.92007
R19237 a_2151_594.n24 a_2151_594.n23 5.64756
R19238 a_2151_594.n46 a_2151_594.n45 5.64756
R19239 a_2151_594.n37 a_2151_594.n36 5.64756
R19240 a_2151_594.n68 a_2151_594.n67 5.64756
R19241 a_2151_594.n59 a_2151_594.n58 5.64756
R19242 a_2151_594.n10 a_2151_594.n9 5.64756
R19243 a_2151_594.n97 a_2151_594.t6 5.5395
R19244 a_2151_594.n97 a_2151_594.t5 5.5395
R19245 a_2151_594.n115 a_2151_594.t4 5.5395
R19246 a_2151_594.t7 a_2151_594.n115 5.5395
R19247 a_2151_594.n78 a_2151_594.n77 5.27461
R19248 a_2151_594.n31 a_2151_594.n20 4.76425
R19249 a_2151_594.n53 a_2151_594.n19 4.76425
R19250 a_2151_594.n33 a_2151_594.n32 4.76425
R19251 a_2151_594.n75 a_2151_594.n18 4.76425
R19252 a_2151_594.n55 a_2151_594.n54 4.76425
R19253 a_2151_594.n17 a_2151_594.n6 4.76425
R19254 a_2151_594.n44 a_2151_594.n43 4.6505
R19255 a_2151_594.n66 a_2151_594.n65 4.6505
R19256 a_2151_594.n104 a_2151_594.n103 4.51815
R19257 a_2151_594.n109 a_2151_594.n108 4.51815
R19258 a_2151_594.n79 a_2151_594.n90 6.0005
R19259 a_2151_594.n80 a_2151_594.n82 4.5005
R19260 a_2151_594.n96 a_2151_594.n101 4.5005
R19261 a_2151_594.n92 a_2151_594.n112 4.5005
R19262 a_2151_594.n5 a_2151_594.n8 3.47842
R19263 a_2151_594.n0 a_2151_594.n22 3.47753
R19264 a_2151_594.n90 a_2151_594.n89 3.38238
R19265 a_2151_594.n95 a_2151_594.t1 3.3065
R19266 a_2151_594.n95 a_2151_594.t3 3.3065
R19267 a_2151_594.n84 a_2151_594.n95 3.21134
R19268 a_2151_594.n102 a_2151_594.n104 3.03311
R19269 a_2151_594.n93 a_2151_594.n109 3.03311
R19270 a_2151_594.n115 a_2151_594.n91 2.85325
R19271 a_2151_594.n94 a_2151_594.n84 2.63601
R19272 a_2151_594.n100 a_2151_594.n99 2.25932
R19273 a_2151_594.n111 a_2151_594.n110 2.25932
R19274 a_2151_594.n90 a_2151_594.n88 1.88285
R19275 a_2151_594.n115 a_2151_594.n114 1.64452
R19276 a_2151_594.n98 a_2151_594.n97 1.64446
R19277 a_2151_594.n94 a_2151_594.n106 1.62064
R19278 a_2151_594.n83 a_2151_594.n86 6.0005
R19279 a_2151_594.n86 a_2151_594.n85 1.12991
R19280 a_2151_594.n27 a_2151_594.n26 1.09595
R19281 a_2151_594.n49 a_2151_594.n48 1.09595
R19282 a_2151_594.n40 a_2151_594.n39 1.09595
R19283 a_2151_594.n71 a_2151_594.n70 1.09595
R19284 a_2151_594.n62 a_2151_594.n61 1.09595
R19285 a_2151_594.n13 a_2151_594.n12 1.09595
R19286 a_2151_594.n101 a_2151_594.n100 0.753441
R19287 a_2151_594.n28 a_2151_594.n24 0.753441
R19288 a_2151_594.n50 a_2151_594.n46 0.753441
R19289 a_2151_594.n41 a_2151_594.n37 0.753441
R19290 a_2151_594.n72 a_2151_594.n68 0.753441
R19291 a_2151_594.n63 a_2151_594.n59 0.753441
R19292 a_2151_594.n14 a_2151_594.n10 0.753441
R19293 a_2151_594.n88 a_2151_594.n87 0.753441
R19294 a_2151_594.n112 a_2151_594.n111 0.753441
R19295 a_2151_594.n107 a_2151_594.n94 0.599869
R19296 a_2151_594.n106 a_2151_594.n105 0.561382
R19297 a_2151_594.n114 a_2151_594.n113 0.462706
R19298 a_2151_594.n55 a_2151_594.n53 0.458354
R19299 a_2151_594.n33 a_2151_594.n31 0.458354
R19300 a_2151_594.n82 a_2151_594.n81 0.376971
R19301 a_2151_594.n76 a_2151_594.n17 0.229427
R19302 a_2151_594.n76 a_2151_594.n75 0.229427
R19303 a_2151_594.n78 a_2151_594.n76 0.191391
R19304 a_2151_594.n4 a_2151_594.n66 0.190717
R19305 a_2151_594.n66 a_2151_594.n3 0.190717
R19306 a_2151_594.n2 a_2151_594.n44 0.190717
R19307 a_2151_594.n44 a_2151_594.n1 0.190717
R19308 a_2151_594.n83 a_2151_594.n84 0.0960207
R19309 a_2151_594.n102 a_2151_594.n96 0.135435
R19310 a_2151_594.n92 a_2151_594.n93 0.134305
R19311 a_2151_594.n79 a_2151_594.n83 0.0765135
R19312 a_2151_594.n80 a_2151_594.n78 0.125375
R19313 a_2151_594.n106 a_2151_594.n102 0.0711242
R19314 a_2151_594.n93 a_2151_594.n107 0.0536188
R19315 a_2151_594.n113 a_2151_594.n92 0.0954783
R19316 a_2151_594.n96 a_2151_594.n98 0.55664
R19317 a_2151_594.n80 a_2151_594.n79 1.53935
R19318 a_2151_594.n17 a_2151_594.n5 0.205546
R19319 a_2151_594.n75 a_2151_594.n4 0.205546
R19320 a_2151_594.n3 a_2151_594.n55 0.205546
R19321 a_2151_594.n53 a_2151_594.n2 0.205546
R19322 a_2151_594.n1 a_2151_594.n33 0.205546
R19323 a_2151_594.n31 a_2151_594.n0 0.205546
R19324 a_2551_620.n27 a_2551_620.t6 60.2505
R19325 a_2551_620.n48 a_2551_620.t7 60.2505
R19326 a_2551_620.n70 a_2551_620.t4 60.2505
R19327 a_2551_620.n82 a_2551_620.t2 60.2505
R19328 a_2551_620.n1 a_2551_620.n90 9.3005
R19329 a_2551_620.n1 a_2551_620.n91 9.3005
R19330 a_2551_620.n1 a_2551_620.n89 9.3005
R19331 a_2551_620.n89 a_2551_620.n88 9.3005
R19332 a_2551_620.n2 a_2551_620.n79 9.3005
R19333 a_2551_620.n3 a_2551_620.n63 9.3005
R19334 a_2551_620.n3 a_2551_620.n62 9.3005
R19335 a_2551_620.n3 a_2551_620.n69 9.3005
R19336 a_2551_620.n69 a_2551_620.n68 9.3005
R19337 a_2551_620.n2 a_2551_620.n78 9.3005
R19338 a_2551_620.n78 a_2551_620.n77 9.3005
R19339 a_2551_620.n2 a_2551_620.n80 9.3005
R19340 a_2551_620.n4 a_2551_620.n57 9.3005
R19341 a_2551_620.n5 a_2551_620.n41 9.3005
R19342 a_2551_620.n5 a_2551_620.n40 9.3005
R19343 a_2551_620.n5 a_2551_620.n47 9.3005
R19344 a_2551_620.n47 a_2551_620.n46 9.3005
R19345 a_2551_620.n4 a_2551_620.n56 9.3005
R19346 a_2551_620.n56 a_2551_620.n55 9.3005
R19347 a_2551_620.n4 a_2551_620.n58 9.3005
R19348 a_2551_620.n6 a_2551_620.n35 9.3005
R19349 a_2551_620.n6 a_2551_620.n34 9.3005
R19350 a_2551_620.n34 a_2551_620.n33 9.3005
R19351 a_2551_620.n6 a_2551_620.n36 9.3005
R19352 a_2551_620.n7 a_2551_620.n98 9.3005
R19353 a_2551_620.n7 a_2551_620.n97 9.3005
R19354 a_2551_620.n100 a_2551_620.n99 9.3005
R19355 a_2551_620.n102 a_2551_620.n101 9.3005
R19356 a_2551_620.n104 a_2551_620.n103 9.3005
R19357 a_2551_620.n0 a_2551_620.n105 9.3005
R19358 a_2551_620.n125 a_2551_620.n112 9.909
R19359 a_2551_620.n125 a_2551_620.n113 11.0386
R19360 a_2551_620.n125 a_2551_620.n124 8.89115
R19361 a_2551_620.n125 a_2551_620.n121 8.88036
R19362 a_2551_620.n125 a_2551_620.n118 8.86963
R19363 a_2551_620.n125 a_2551_620.n115 8.85895
R19364 a_2551_620.n71 a_2551_620.n70 8.76429
R19365 a_2551_620.n49 a_2551_620.n48 8.76429
R19366 a_2551_620.n32 a_2551_620.n31 7.45411
R19367 a_2551_620.n45 a_2551_620.n44 7.45411
R19368 a_2551_620.n54 a_2551_620.n53 7.45411
R19369 a_2551_620.n67 a_2551_620.n66 7.45411
R19370 a_2551_620.n76 a_2551_620.n75 7.45411
R19371 a_2551_620.n87 a_2551_620.n86 7.45411
R19372 a_2551_620.n20 a_2551_620.n19 7.45281
R19373 a_2551_620.n28 a_2551_620.n27 6.80105
R19374 a_2551_620.n83 a_2551_620.n82 6.80105
R19375 a_2551_620.n0 a_2551_620.n11 6.29716
R19376 a_2551_620.n30 a_2551_620.n29 5.64756
R19377 a_2551_620.n43 a_2551_620.n42 5.64756
R19378 a_2551_620.n52 a_2551_620.n51 5.64756
R19379 a_2551_620.n65 a_2551_620.n64 5.64756
R19380 a_2551_620.n74 a_2551_620.n73 5.64756
R19381 a_2551_620.n85 a_2551_620.n84 5.64756
R19382 a_2551_620.n125 a_2551_620.t5 5.5395
R19383 a_2551_620.t3 a_2551_620.n125 5.5395
R19384 a_2551_620.n96 a_2551_620.n95 4.95534
R19385 a_2551_620.n37 a_2551_620.n26 4.73575
R19386 a_2551_620.n39 a_2551_620.n38 4.73575
R19387 a_2551_620.n59 a_2551_620.n25 4.73575
R19388 a_2551_620.n61 a_2551_620.n60 4.73575
R19389 a_2551_620.n81 a_2551_620.n24 4.73575
R19390 a_2551_620.n93 a_2551_620.n92 4.73575
R19391 a_2551_620.n72 a_2551_620.n71 4.6505
R19392 a_2551_620.n50 a_2551_620.n49 4.6505
R19393 a_2551_620.n8 a_2551_620.n21 4.5005
R19394 a_2551_620.n9 a_2551_620.n20 4.5005
R19395 a_2551_620.n8 a_2551_620.n108 4.5005
R19396 a_2551_620.n0 a_2551_620.n23 4.5005
R19397 a_2551_620.n9 a_2551_620.n110 4.5005
R19398 a_2551_620.n6 a_2551_620.n28 3.42768
R19399 a_2551_620.n1 a_2551_620.n83 3.42768
R19400 a_2551_620.n110 a_2551_620.n109 3.38874
R19401 a_2551_620.n117 a_2551_620.n116 3.38874
R19402 a_2551_620.n17 a_2551_620.n16 3.38238
R19403 a_2551_620.n106 a_2551_620.t1 3.3065
R19404 a_2551_620.n106 a_2551_620.t0 3.3065
R19405 a_2551_620.n11 a_2551_620.n106 3.21133
R19406 a_2551_620.n20 a_2551_620.n18 2.63579
R19407 a_2551_620.n120 a_2551_620.n119 2.63579
R19408 a_2551_620.n17 a_2551_620.n15 1.88285
R19409 a_2551_620.n23 a_2551_620.n22 1.88285
R19410 a_2551_620.n123 a_2551_620.n122 1.88285
R19411 a_2551_620.n125 a_2551_620.n111 1.67004
R19412 a_2551_620.n108 a_2551_620.n107 1.50638
R19413 a_2551_620.n10 a_2551_620.n13 6.0005
R19414 a_2551_620.n13 a_2551_620.n12 1.12991
R19415 a_2551_620.n33 a_2551_620.n32 0.994314
R19416 a_2551_620.n46 a_2551_620.n45 0.994314
R19417 a_2551_620.n55 a_2551_620.n54 0.994314
R19418 a_2551_620.n68 a_2551_620.n67 0.994314
R19419 a_2551_620.n77 a_2551_620.n76 0.994314
R19420 a_2551_620.n88 a_2551_620.n87 0.994314
R19421 a_2551_620.n111 a_2551_620.n9 0.944917
R19422 a_2551_620.n15 a_2551_620.n14 0.753441
R19423 a_2551_620.n34 a_2551_620.n30 0.753441
R19424 a_2551_620.n47 a_2551_620.n43 0.753441
R19425 a_2551_620.n56 a_2551_620.n52 0.753441
R19426 a_2551_620.n69 a_2551_620.n65 0.753441
R19427 a_2551_620.n78 a_2551_620.n74 0.753441
R19428 a_2551_620.n89 a_2551_620.n85 0.753441
R19429 a_2551_620.n39 a_2551_620.n37 0.458354
R19430 a_2551_620.n61 a_2551_620.n59 0.458354
R19431 a_2551_620.n94 a_2551_620.n81 0.229427
R19432 a_2551_620.n94 a_2551_620.n93 0.229427
R19433 a_2551_620.n96 a_2551_620.n94 0.215848
R19434 a_2551_620.n104 a_2551_620.n102 0.190717
R19435 a_2551_620.n50 a_2551_620.n5 0.190717
R19436 a_2551_620.n4 a_2551_620.n50 0.190717
R19437 a_2551_620.n72 a_2551_620.n3 0.190717
R19438 a_2551_620.n2 a_2551_620.n72 0.190717
R19439 a_2551_620.n0 a_2551_620.n104 0.190717
R19440 a_2551_620.n102 a_2551_620.n100 0.190717
R19441 a_2551_620.n7 a_2551_620.n96 0.164777
R19442 a_2551_620.n115 a_2551_620.n114 0.160869
R19443 a_2551_620.n118 a_2551_620.n117 0.14967
R19444 a_2551_620.n121 a_2551_620.n120 0.138414
R19445 a_2551_620.n124 a_2551_620.n123 0.127101
R19446 a_2551_620.n10 a_2551_620.n11 0.0960207
R19447 a_2551_620.n17 a_2551_620.n10 6.07651
R19448 a_2551_620.n8 a_2551_620.n0 0.208476
R19449 a_2551_620.n37 a_2551_620.n6 0.205546
R19450 a_2551_620.n5 a_2551_620.n39 0.205546
R19451 a_2551_620.n59 a_2551_620.n4 0.205546
R19452 a_2551_620.n3 a_2551_620.n61 0.205546
R19453 a_2551_620.n81 a_2551_620.n2 0.205546
R19454 a_2551_620.n93 a_2551_620.n1 0.205546
R19455 a_2551_620.n100 a_2551_620.n7 0.190717
R19456 a_2551_620.n9 a_2551_620.n8 0.135431
R19457 a_5299_3714.n53 a_5299_3714.t2 60.2505
R19458 a_5299_3714.n31 a_5299_3714.t9 60.2505
R19459 a_5299_3714.n9 a_5299_3714.t8 60.2505
R19460 a_5299_3714.n66 a_5299_3714.t0 60.2505
R19461 a_5299_3714.n0 a_5299_3714.n74 9.3005
R19462 a_5299_3714.n0 a_5299_3714.n75 9.3005
R19463 a_5299_3714.n0 a_5299_3714.n73 9.3005
R19464 a_5299_3714.n73 a_5299_3714.n72 9.3005
R19465 a_5299_3714.n3 a_5299_3714.n41 9.3005
R19466 a_5299_3714.n4 a_5299_3714.n23 9.3005
R19467 a_5299_3714.n5 a_5299_3714.n18 9.3005
R19468 a_5299_3714.n5 a_5299_3714.n17 9.3005
R19469 a_5299_3714.n5 a_5299_3714.n16 9.3005
R19470 a_5299_3714.n16 a_5299_3714.n15 9.3005
R19471 a_5299_3714.n4 a_5299_3714.n24 9.3005
R19472 a_5299_3714.n4 a_5299_3714.n30 9.3005
R19473 a_5299_3714.n30 a_5299_3714.n29 9.3005
R19474 a_5299_3714.n3 a_5299_3714.n40 9.3005
R19475 a_5299_3714.n3 a_5299_3714.n39 9.3005
R19476 a_5299_3714.n39 a_5299_3714.n38 9.3005
R19477 a_5299_3714.n2 a_5299_3714.n45 9.3005
R19478 a_5299_3714.n2 a_5299_3714.n52 9.3005
R19479 a_5299_3714.n52 a_5299_3714.n51 9.3005
R19480 a_5299_3714.n2 a_5299_3714.n46 9.3005
R19481 a_5299_3714.n1 a_5299_3714.n61 9.3005
R19482 a_5299_3714.n61 a_5299_3714.n60 9.3005
R19483 a_5299_3714.n1 a_5299_3714.n63 9.3005
R19484 a_5299_3714.n1 a_5299_3714.n62 9.3005
R19485 a_5299_3714.n32 a_5299_3714.n31 8.76429
R19486 a_5299_3714.n54 a_5299_3714.n53 8.76429
R19487 a_5299_3714.n14 a_5299_3714.n13 8.21641
R19488 a_5299_3714.n28 a_5299_3714.n27 8.21641
R19489 a_5299_3714.n37 a_5299_3714.n36 8.21641
R19490 a_5299_3714.n71 a_5299_3714.n70 8.21641
R19491 a_5299_3714.n50 a_5299_3714.n49 8.21641
R19492 a_5299_3714.n59 a_5299_3714.n58 8.21641
R19493 a_5299_3714.n10 a_5299_3714.n9 6.92242
R19494 a_5299_3714.n67 a_5299_3714.n66 6.92012
R19495 a_5299_3714.n12 a_5299_3714.n11 5.64756
R19496 a_5299_3714.n26 a_5299_3714.n25 5.64756
R19497 a_5299_3714.n35 a_5299_3714.n34 5.64756
R19498 a_5299_3714.n69 a_5299_3714.n68 5.64756
R19499 a_5299_3714.n48 a_5299_3714.n47 5.64756
R19500 a_5299_3714.n57 a_5299_3714.n56 5.64756
R19501 a_5299_3714.n98 a_5299_3714.t5 5.5395
R19502 a_5299_3714.n98 a_5299_3714.t4 5.5395
R19503 a_5299_3714.n115 a_5299_3714.t6 5.5395
R19504 a_5299_3714.t7 a_5299_3714.n115 5.5395
R19505 a_5299_3714.n79 a_5299_3714.n78 5.27461
R19506 a_5299_3714.n20 a_5299_3714.n19 4.76425
R19507 a_5299_3714.n22 a_5299_3714.n21 4.76425
R19508 a_5299_3714.n43 a_5299_3714.n42 4.76425
R19509 a_5299_3714.n76 a_5299_3714.n65 4.76425
R19510 a_5299_3714.n44 a_5299_3714.n8 4.76425
R19511 a_5299_3714.n64 a_5299_3714.n7 4.76425
R19512 a_5299_3714.n33 a_5299_3714.n32 4.6505
R19513 a_5299_3714.n55 a_5299_3714.n54 4.6505
R19514 a_5299_3714.n105 a_5299_3714.n104 4.51815
R19515 a_5299_3714.n110 a_5299_3714.n109 4.51815
R19516 a_5299_3714.n80 a_5299_3714.n91 6.0005
R19517 a_5299_3714.n81 a_5299_3714.n83 4.5005
R19518 a_5299_3714.n97 a_5299_3714.n102 4.5005
R19519 a_5299_3714.n93 a_5299_3714.n113 4.5005
R19520 a_5299_3714.n0 a_5299_3714.n67 3.47756
R19521 a_5299_3714.n5 a_5299_3714.n10 3.4767
R19522 a_5299_3714.n91 a_5299_3714.n90 3.38238
R19523 a_5299_3714.n95 a_5299_3714.t3 3.3065
R19524 a_5299_3714.n95 a_5299_3714.t1 3.3065
R19525 a_5299_3714.n85 a_5299_3714.n95 3.21134
R19526 a_5299_3714.n103 a_5299_3714.n105 3.03311
R19527 a_5299_3714.n94 a_5299_3714.n110 3.03311
R19528 a_5299_3714.n115 a_5299_3714.n92 2.85325
R19529 a_5299_3714.n6 a_5299_3714.n85 2.81636
R19530 a_5299_3714.n101 a_5299_3714.n100 2.25932
R19531 a_5299_3714.n112 a_5299_3714.n111 2.25932
R19532 a_5299_3714.n91 a_5299_3714.n89 1.88285
R19533 a_5299_3714.n99 a_5299_3714.n98 1.64453
R19534 a_5299_3714.n115 a_5299_3714.n114 1.64449
R19535 a_5299_3714.n84 a_5299_3714.n87 6.0005
R19536 a_5299_3714.n87 a_5299_3714.n86 1.12991
R19537 a_5299_3714.n15 a_5299_3714.n14 1.09595
R19538 a_5299_3714.n29 a_5299_3714.n28 1.09595
R19539 a_5299_3714.n38 a_5299_3714.n37 1.09595
R19540 a_5299_3714.n72 a_5299_3714.n71 1.09595
R19541 a_5299_3714.n51 a_5299_3714.n50 1.09595
R19542 a_5299_3714.n60 a_5299_3714.n59 1.09595
R19543 a_5299_3714.n107 a_5299_3714.n106 0.760382
R19544 a_5299_3714.n16 a_5299_3714.n12 0.753441
R19545 a_5299_3714.n30 a_5299_3714.n26 0.753441
R19546 a_5299_3714.n39 a_5299_3714.n35 0.753441
R19547 a_5299_3714.n73 a_5299_3714.n69 0.753441
R19548 a_5299_3714.n52 a_5299_3714.n48 0.753441
R19549 a_5299_3714.n61 a_5299_3714.n57 0.753441
R19550 a_5299_3714.n89 a_5299_3714.n88 0.753441
R19551 a_5299_3714.n102 a_5299_3714.n101 0.753441
R19552 a_5299_3714.n113 a_5299_3714.n112 0.753441
R19553 a_5299_3714.n6 a_5299_3714.n107 0.678625
R19554 a_5299_3714.n106 a_5299_3714.n96 0.573452
R19555 a_5299_3714.n22 a_5299_3714.n20 0.458354
R19556 a_5299_3714.n44 a_5299_3714.n43 0.458354
R19557 a_5299_3714.n83 a_5299_3714.n82 0.376971
R19558 a_5299_3714.n77 a_5299_3714.n64 0.229427
R19559 a_5299_3714.n77 a_5299_3714.n76 0.229427
R19560 a_5299_3714.n79 a_5299_3714.n77 0.191391
R19561 a_5299_3714.n33 a_5299_3714.n4 0.190717
R19562 a_5299_3714.n3 a_5299_3714.n33 0.190717
R19563 a_5299_3714.n55 a_5299_3714.n2 0.190717
R19564 a_5299_3714.n1 a_5299_3714.n55 0.190717
R19565 a_5299_3714.n84 a_5299_3714.n85 0.0960207
R19566 a_5299_3714.n93 a_5299_3714.n94 0.135434
R19567 a_5299_3714.n103 a_5299_3714.n97 0.13503
R19568 a_5299_3714.n80 a_5299_3714.n84 0.0765135
R19569 a_5299_3714.n81 a_5299_3714.n79 0.125375
R19570 a_5299_3714.n106 a_5299_3714.n103 0.0591603
R19571 a_5299_3714.n94 a_5299_3714.n108 0.0540944
R19572 a_5299_3714.n114 a_5299_3714.n93 0.556715
R19573 a_5299_3714.n97 a_5299_3714.n99 0.556623
R19574 a_5299_3714.n81 a_5299_3714.n80 1.53935
R19575 a_5299_3714.n108 a_5299_3714.n6 0.620875
R19576 a_5299_3714.n20 a_5299_3714.n5 0.205546
R19577 a_5299_3714.n4 a_5299_3714.n22 0.205546
R19578 a_5299_3714.n43 a_5299_3714.n3 0.205546
R19579 a_5299_3714.n2 a_5299_3714.n44 0.205546
R19580 a_5299_3714.n64 a_5299_3714.n1 0.205546
R19581 a_5299_3714.n76 a_5299_3714.n0 0.205546
R19582 a_2093_1782.n88 a_2093_1782.n86 8.05594
R19583 a_2093_1782.n88 a_2093_1782.n87 8.02969
R19584 a_2093_1782.n84 a_2093_1782.n83 6.13632
R19585 a_2093_1782.n46 a_2093_1782.n45 5.61041
R19586 a_2093_1782.n58 a_2093_1782.n57 5.61041
R19587 a_2093_1782.n82 a_2093_1782.n81 5.61041
R19588 a_2093_1782.n26 a_2093_1782.n25 5.61037
R19589 a_2093_1782.n72 a_2093_1782.n71 5.61037
R19590 a_2093_1782.n69 a_2093_1782.n68 5.61037
R19591 a_2093_1782.n48 a_2093_1782.n51 4.5005
R19592 a_2093_1782.n6 a_2093_1782.n66 4.5005
R19593 a_2093_1782.n15 a_2093_1782.n80 4.5005
R19594 a_2093_1782.n8 a_2093_1782.n76 4.5005
R19595 a_2093_1782.n4 a_2093_1782.n55 4.5005
R19596 a_2093_1782.n36 a_2093_1782.n39 4.5005
R19597 a_2093_1782.n13 a_2093_1782.n34 4.5005
R19598 a_2093_1782.n0 a_2093_1782.n30 4.5005
R19599 a_2093_1782.n2 a_2093_1782.n43 4.5005
R19600 a_2093_1782.n14 a_2093_1782.n62 4.5005
R19601 a_2093_1782.n20 a_2093_1782.n23 4.5005
R19602 a_2093_1782.n21 a_2093_1782.n19 4.5005
R19603 a_2093_1782.n34 a_2093_1782.n33 3.76521
R19604 a_2093_1782.n39 a_2093_1782.n38 3.76521
R19605 a_2093_1782.n80 a_2093_1782.n79 3.76521
R19606 a_2093_1782.n51 a_2093_1782.n50 3.76521
R19607 a_2093_1782.n62 a_2093_1782.n61 3.76521
R19608 a_2093_1782.n19 a_2093_1782.n18 3.76521
R19609 a_2093_1782.n30 a_2093_1782.n28 3.38874
R19610 a_2093_1782.n43 a_2093_1782.n41 3.38874
R19611 a_2093_1782.n76 a_2093_1782.n74 3.38874
R19612 a_2093_1782.n55 a_2093_1782.n53 3.38874
R19613 a_2093_1782.n66 a_2093_1782.n64 3.38874
R19614 a_2093_1782.n31 a_2093_1782.t4 3.3065
R19615 a_2093_1782.n31 a_2093_1782.t3 3.3065
R19616 a_2093_1782.n35 a_2093_1782.t0 3.3065
R19617 a_2093_1782.n35 a_2093_1782.t2 3.3065
R19618 a_2093_1782.n77 a_2093_1782.t9 3.3065
R19619 a_2093_1782.n77 a_2093_1782.t8 3.3065
R19620 a_2093_1782.n47 a_2093_1782.t11 3.3065
R19621 a_2093_1782.n47 a_2093_1782.t5 3.3065
R19622 a_2093_1782.n59 a_2093_1782.t7 3.3065
R19623 a_2093_1782.n59 a_2093_1782.t6 3.3065
R19624 a_2093_1782.n88 a_2093_1782.t1 3.3065
R19625 a_2093_1782.t10 a_2093_1782.n88 3.3065
R19626 a_2093_1782.n30 a_2093_1782.n29 3.01226
R19627 a_2093_1782.n43 a_2093_1782.n42 3.01226
R19628 a_2093_1782.n76 a_2093_1782.n75 3.01226
R19629 a_2093_1782.n55 a_2093_1782.n54 3.01226
R19630 a_2093_1782.n66 a_2093_1782.n65 3.01226
R19631 a_2093_1782.n23 a_2093_1782.n22 3.01226
R19632 a_2093_1782.n34 a_2093_1782.n32 2.63579
R19633 a_2093_1782.n39 a_2093_1782.n37 2.63579
R19634 a_2093_1782.n80 a_2093_1782.n78 2.63579
R19635 a_2093_1782.n51 a_2093_1782.n49 2.63579
R19636 a_2093_1782.n62 a_2093_1782.n60 2.63579
R19637 a_2093_1782.n16 a_2093_1782.n7 2.2019
R19638 a_2093_1782.n11 a_2093_1782.n1 2.18356
R19639 a_2093_1782.n36 a_2093_1782.n35 1.85087
R19640 a_2093_1782.n48 a_2093_1782.n47 1.85087
R19641 a_2093_1782.n13 a_2093_1782.n31 1.85087
R19642 a_2093_1782.n15 a_2093_1782.n77 1.85087
R19643 a_2093_1782.n14 a_2093_1782.n59 1.85087
R19644 a_2093_1782.n84 a_2093_1782.n21 1.48738
R19645 a_2093_1782.n11 a_2093_1782.n3 1.48434
R19646 a_2093_1782.n17 a_2093_1782.n9 1.48434
R19647 a_2093_1782.n16 a_2093_1782.n5 1.48434
R19648 a_2093_1782.n10 a_2093_1782.n12 1.48434
R19649 a_2093_1782.n12 a_2093_1782.n17 0.734472
R19650 a_2093_1782.n17 a_2093_1782.n16 0.718062
R19651 a_2093_1782.n12 a_2093_1782.n11 0.718062
R19652 a_2093_1782.n25 a_2093_1782.n24 0.461175
R19653 a_2093_1782.n45 a_2093_1782.n44 0.461175
R19654 a_2093_1782.n71 a_2093_1782.n70 0.461175
R19655 a_2093_1782.n57 a_2093_1782.n56 0.461175
R19656 a_2093_1782.n68 a_2093_1782.n67 0.461175
R19657 a_2093_1782.n28 a_2093_1782.n27 0.430121
R19658 a_2093_1782.n41 a_2093_1782.n40 0.430121
R19659 a_2093_1782.n74 a_2093_1782.n73 0.430121
R19660 a_2093_1782.n53 a_2093_1782.n52 0.430121
R19661 a_2093_1782.n64 a_2093_1782.n63 0.430121
R19662 a_2093_1782.n86 a_2093_1782.n85 0.429625
R19663 a_2093_1782.n88 a_2093_1782.n84 0.363994
R19664 a_2093_1782.n7 a_2093_1782.n69 0.297864
R19665 a_2093_1782.n1 a_2093_1782.n26 0.297864
R19666 a_2093_1782.n9 a_2093_1782.n72 0.297864
R19667 a_2093_1782.n5 a_2093_1782.n58 0.297822
R19668 a_2093_1782.n3 a_2093_1782.n46 0.297822
R19669 a_2093_1782.n10 a_2093_1782.n82 0.297822
R19670 a_2093_1782.n21 a_2093_1782.n20 0.14384
R19671 a_2093_1782.n0 a_2093_1782.n13 0.14384
R19672 a_2093_1782.n2 a_2093_1782.n36 0.142841
R19673 a_2093_1782.n4 a_2093_1782.n48 0.142841
R19674 a_2093_1782.n8 a_2093_1782.n15 0.142841
R19675 a_2093_1782.n6 a_2093_1782.n14 0.141862
R19676 a_2093_1782.n20 a_2093_1782.n10 0.136602
R19677 a_2093_1782.n9 a_2093_1782.n8 0.136602
R19678 a_2093_1782.n7 a_2093_1782.n6 0.136602
R19679 a_2093_1782.n5 a_2093_1782.n4 0.136602
R19680 a_2093_1782.n3 a_2093_1782.n2 0.136602
R19681 a_2093_1782.n1 a_2093_1782.n0 0.136602
R19682 VO.n8 VO.n7 148.663
R19683 VO.n16 VO.t1 122.728
R19684 VO.n5 VO.t0 22.4191
R19685 VO.n9 VO.n8 10.5541
R19686 VO.n7 VO 9.62836
R19687 VO.n10 VO.n9 9.3005
R19688 VO VO.n12 7.00682
R19689 VO VO.n11 6.32867
R19690 VO.n15 VO.n14 5.92892
R19691 VO.n15 VO.n3 4.72813
R19692 VO.n16 VO 4.69453
R19693 VO.n12 VO.n2 4.6505
R19694 VO.n19 VO.n18 4.6505
R19695 VO VO.n21 3.37933
R19696 VO.n12 VO 2.96471
R19697 VO VO.n15 2.42576
R19698 VO.n8 VO.n5 2.19143
R19699 VO.n13 VO 2.15629
R19700 VO.n11 VO.n2 2.04091
R19701 VO VO.n1 1.95259
R19702 VO.n18 VO.n17 1.75208
R19703 VO.n6 VO.n4 1.61734
R19704 VO.n14 VO 1.61734
R19705 VO.n11 VO.n10 0.816947
R19706 VO.n17 VO.n16 0.795743
R19707 VO.n10 VO.n4 0.674184
R19708 VO.n18 VO.n13 0.539447
R19709 VO.n7 VO 0.343399
R19710 VO VO.n6 0.269974
R19711 VO.n1 VO.n0 0.202535
R19712 VO.n21 VO.n20 0.0807632
R19713 VO.n1 VO 0.0730901
R19714 VO.n19 VO.n3 0.0176053
R19715 VO.n21 VO.n2 0.00971053
R19716 VO.n20 VO.n19 0.00576316
R19717 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 136.804
R19718 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 136.325
R19719 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 119.999
R19720 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 93.9023
R19721 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 93.3044
R19722 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 93.0848
R19723 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n4 92.5005
R19724 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 92.4623
R19725 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 69.2281
R19726 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 29.4833
R19727 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 27.6955
R19728 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 27.6955
R19729 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 15.4626
R19730 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n16 9.3005
R19731 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n8 9.3005
R19732 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n7 9.3005
R19733 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 9.3005
R19734 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 9.3005
R19735 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n15 9.3005
R19736 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n17 9.3005
R19737 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 9.02061
R19738 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 9.02061
R19739 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n34 8.28285
R19740 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n21 8.28285
R19741 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 5.64756
R19742 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 5.31864
R19743 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n42 4.14168
R19744 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n28 4.14168
R19745 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 4.06959
R19746 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n11 3.93153
R19747 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n40 3.76521
R19748 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n33 3.76521
R19749 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n24 3.76521
R19750 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n19 3.76521
R19751 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n36 3.38874
R19752 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n22 3.38874
R19753 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 3.0736
R19754 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 3.07249
R19755 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 3.07078
R19756 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 3.04338
R19757 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 3.03311
R19758 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 3.03311
R19759 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 3.03311
R19760 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n39 2.63579
R19761 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n20 2.63579
R19762 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 2.27447
R19763 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 2.25932
R19764 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 2.25932
R19765 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 1.80772
R19766 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n30 1.61433
R19767 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 1.45534
R19768 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 1.19419
R19769 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n9 0.753441
R19770 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 0.719888
R19771 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 0.22499
R19772 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 0.176176
R19773 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 2.36361
R19774 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 2.36353
R19775 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 1.14499
R19776 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 1.00043
R19777 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 120.01
R19778 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 92.9415
R19779 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n4 92.5005
R19780 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 92.4623
R19781 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 73.195
R19782 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 72.1651
R19783 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 29.4833
R19784 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 27.6955
R19785 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 27.6955
R19786 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 15.4607
R19787 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 9.3005
R19788 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 9.3005
R19789 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n33 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 9.02061
R19790 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 9.01961
R19791 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n15 8.28285
R19792 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 8.28285
R19793 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 5.64756
R19794 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 5.31894
R19795 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n23 4.14168
R19796 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 4.14168
R19797 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n34 4.14168
R19798 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n27 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n26 4.14168
R19799 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 4.03426
R19800 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n9 3.93153
R19801 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n19 3.76521
R19802 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n36 3.76521
R19803 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 3.20519
R19804 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 3.07304
R19805 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 3.07194
R19806 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n27 3.07027
R19807 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n39 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n38 3.04478
R19808 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 3.03311
R19809 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n14 3.03311
R19810 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 3.03311
R19811 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n16 3.01226
R19812 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n29 3.01226
R19813 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n20 2.63579
R19814 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n37 2.63579
R19815 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 2.47579
R19816 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n39 2.27091
R19817 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 2.25932
R19818 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n33 2.25932
R19819 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 2.25549
R19820 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 1.51198
R19821 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 1.15307
R19822 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 1.04295
R19823 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n7 0.753441
R19824 SELA.n1 SELA.t2 186.374
R19825 SELA.n1 SELA.t3 170.308
R19826 SELA.n2 SELA.n1 139.876
R19827 SELA.n5 SELA.t4 84.8325
R19828 SELA.n6 SELA.t0 84.8325
R19829 SELA.n6 SELA.n5 60.1541
R19830 SELA.n7 SELA.n6 50.1642
R19831 SELA.n5 SELA.t5 48.6825
R19832 SELA.n6 SELA.t1 48.6825
R19833 SELA.n0 SELA 42.9181
R19834 SELA.n9 SELA 17.169
R19835 SELA.n8 SELA.n7 15.2731
R19836 SELA.n0 SELA 12.8005
R19837 SELA.n9 SELA.n8 4.77356
R19838 SELA.n3 SELA 2.73914
R19839 SELA.n10 SELA 2.70667
R19840 SELA SELA.n8 2.13383
R19841 SELA SELA.n2 1.61978
R19842 SELA.n4 SELA.n3 1.31185
R19843 SELA.n7 SELA 1.1768
R19844 SELA.n2 SELA.n0 0.925801
R19845 SELA.n12 SELA.n11 0.659992
R19846 SELA.n11 SELA 0.559032
R19847 SELA.n13 SELA 0.34425
R19848 SELA.n10 SELA 0.321549
R19849 SELA SELA.n14 0.0255
R19850 SELA.n14 SELA.n13 0.0194024
R19851 SELA SELA.n9 0.0180439
R19852 SELA SELA.n12 0.0151341
R19853 SELA.n3 SELA 0.00770734
R19854 SELA.n12 SELA 0.00415854
R19855 SELA.n13 SELA 0.00171951
R19856 SELA.n12 SELA.n4 0.000502048
R19857 SELA.n11 SELA.n10 0.000500307
R19858 DVDD.n282 DVDD.t22 591.327
R19859 DVDD.n284 DVDD.t26 591.327
R19860 DVDD.n293 DVDD.n292 585
R19861 DVDD.n166 DVDD.n153 321.882
R19862 DVDD.n200 DVDD.n153 321.882
R19863 DVDD.n200 DVDD.n151 321.882
R19864 DVDD.n26 DVDD.n13 321.882
R19865 DVDD.n60 DVDD.n13 321.882
R19866 DVDD.n60 DVDD.n11 321.882
R19867 DVDD.n201 DVDD.n152 175.386
R19868 DVDD.n61 DVDD.n12 175.386
R19869 DVDD.n166 DVDD.t2 171.452
R19870 DVDD.n26 DVDD.t18 171.452
R19871 DVDD.n316 DVDD.n315 161.37
R19872 DVDD.n82 DVDD.n75 161.37
R19873 DVDD.n229 DVDD.n228 161.37
R19874 DVDD.n130 DVDD.n129 161.37
R19875 DVDD.n173 DVDD.t3 160.743
R19876 DVDD.n33 DVDD.t19 160.743
R19877 DVDD.n185 DVDD.t7 158.225
R19878 DVDD.n45 DVDD.t9 158.225
R19879 DVDD.n287 DVDD.t23 148.294
R19880 DVDD.t10 DVDD.n77 129.546
R19881 DVDD.t24 DVDD.n224 129.546
R19882 DVDD.t12 DVDD.n125 129.546
R19883 DVDD.n203 DVDD.n202 124.013
R19884 DVDD.n63 DVDD.n62 124.013
R19885 DVDD.n291 DVDD.n288 107.746
R19886 DVDD.n310 DVDD.t16 100.874
R19887 DVDD.n78 DVDD.t10 100.874
R19888 DVDD.n225 DVDD.t24 100.874
R19889 DVDD.n126 DVDD.t12 100.874
R19890 DVDD.t6 DVDD.n201 96.8274
R19891 DVDD.t8 DVDD.n61 96.8274
R19892 DVDD.n284 DVDD.n279 92.5005
R19893 DVDD.n311 DVDD.n309 92.5005
R19894 DVDD.n79 DVDD.n77 92.5005
R19895 DVDD.n77 DVDD.n76 92.5005
R19896 DVDD.n226 DVDD.n224 92.5005
R19897 DVDD.n224 DVDD.n223 92.5005
R19898 DVDD.n127 DVDD.n125 92.5005
R19899 DVDD.n125 DVDD.n124 92.5005
R19900 DVDD.n284 DVDD.n283 81.7536
R19901 DVDD.n202 DVDD.t6 81.7266
R19902 DVDD.n62 DVDD.t8 81.7266
R19903 DVDD.n312 DVDD.n308 55.3934
R19904 DVDD.n80 DVDD.n76 55.3934
R19905 DVDD.n227 DVDD.n223 55.3934
R19906 DVDD.n128 DVDD.n124 55.3934
R19907 DVDD.n287 DVDD.n280 52.9371
R19908 DVDD.n294 DVDD.n279 49.5938
R19909 DVDD.n285 DVDD.n284 47.5553
R19910 DVDD.n309 DVDD.t20 47.2949
R19911 DVDD.n77 DVDD.t0 47.2949
R19912 DVDD.n224 DVDD.t14 47.2949
R19913 DVDD.n125 DVDD.t4 47.2949
R19914 DVDD.n287 DVDD.n286 46.2505
R19915 DVDD.n312 DVDD.n311 46.2505
R19916 DVDD.n80 DVDD.n79 46.2505
R19917 DVDD.n227 DVDD.n226 46.2505
R19918 DVDD.n128 DVDD.n127 46.2505
R19919 DVDD.n285 DVDD.n280 42.3392
R19920 DVDD.n283 DVDD.n282 40.8773
R19921 DVDD.n167 DVDD.n154 36.1417
R19922 DVDD.n199 DVDD.n154 36.1417
R19923 DVDD.n199 DVDD.n150 36.1417
R19924 DVDD.n203 DVDD.n150 36.1417
R19925 DVDD.n27 DVDD.n14 36.1417
R19926 DVDD.n59 DVDD.n14 36.1417
R19927 DVDD.n59 DVDD.n10 36.1417
R19928 DVDD.n63 DVDD.n10 36.1417
R19929 DVDD.n283 DVDD.n280 34.4168
R19930 DVDD.n315 DVDD.t17 32.8338
R19931 DVDD.n315 DVDD.t21 32.8338
R19932 DVDD.n75 DVDD.t11 32.8338
R19933 DVDD.n75 DVDD.t1 32.8338
R19934 DVDD.n228 DVDD.t25 32.8338
R19935 DVDD.n228 DVDD.t15 32.8338
R19936 DVDD.n129 DVDD.t13 32.8338
R19937 DVDD.n129 DVDD.t5 32.8338
R19938 DVDD.n282 DVDD.n281 32.0046
R19939 DVDD.n286 DVDD.n281 28.4938
R19940 DVDD.n281 DVDD.n279 28.4938
R19941 DVDD.n311 DVDD.n310 26.4697
R19942 DVDD.n78 DVDD.n76 26.4697
R19943 DVDD.n79 DVDD.n78 26.4697
R19944 DVDD.n225 DVDD.n223 26.4697
R19945 DVDD.n226 DVDD.n225 26.4697
R19946 DVDD.n126 DVDD.n124 26.4697
R19947 DVDD.n127 DVDD.n126 26.4697
R19948 DVDD.n290 DVDD.t27 22.8666
R19949 DVDD.n286 DVDD.n285 21.17
R19950 DVDD.n314 DVDD.n313 17.8772
R19951 DVDD.n81 DVDD.n74 17.8772
R19952 DVDD.n231 DVDD.n230 17.8772
R19953 DVDD.n132 DVDD.n131 17.8772
R19954 DVDD.n82 DVDD.n81 17.4938
R19955 DVDD.n230 DVDD.n229 17.4938
R19956 DVDD.n131 DVDD.n130 17.4938
R19957 DVDD.n292 DVDD.n291 13.514
R19958 DVDD.t2 DVDD.n152 12.789
R19959 DVDD.t18 DVDD.n12 12.789
R19960 DVDD.n292 DVDD.t28 11.4335
R19961 DVDD.n295 DVDD.n294 10.8623
R19962 DVDD.n290 DVDD.n289 9.3005
R19963 DVDD.n173 DVDD.n172 9.3005
R19964 DVDD.n173 DVDD.n162 9.3005
R19965 DVDD.n173 DVDD.n161 9.3005
R19966 DVDD.n33 DVDD.n32 9.3005
R19967 DVDD.n33 DVDD.n22 9.3005
R19968 DVDD.n33 DVDD.n21 9.3005
R19969 DVDD.n167 DVDD.n166 8.85536
R19970 DVDD.n154 DVDD.n153 8.85536
R19971 DVDD.n153 DVDD.n152 8.85536
R19972 DVDD.n200 DVDD.n199 8.85536
R19973 DVDD.n201 DVDD.n200 8.85536
R19974 DVDD.n151 DVDD.n150 8.85536
R19975 DVDD.n27 DVDD.n26 8.85536
R19976 DVDD.n14 DVDD.n13 8.85536
R19977 DVDD.n13 DVDD.n12 8.85536
R19978 DVDD.n60 DVDD.n59 8.85536
R19979 DVDD.n61 DVDD.n60 8.85536
R19980 DVDD.n11 DVDD.n10 8.85536
R19981 DVDD.n202 DVDD.n151 5.53567
R19982 DVDD.n62 DVDD.n11 5.53567
R19983 DVDD.n317 DVDD.n316 4.6505
R19984 DVDD.n83 DVDD.n82 4.6505
R19985 DVDD.n229 DVDD.n222 4.6505
R19986 DVDD.n130 DVDD.n123 4.6505
R19987 DVDD.n185 DVDD.n149 4.6505
R19988 DVDD.n192 DVDD.n185 4.6505
R19989 DVDD.n174 DVDD.n173 4.6505
R19990 DVDD.n45 DVDD.n9 4.6505
R19991 DVDD.n52 DVDD.n45 4.6505
R19992 DVDD.n34 DVDD.n33 4.6505
R19993 DVDD.n256 DVDD.n70 4.5005
R19994 DVDD.n240 DVDD.n88 4.5005
R19995 DVDD.n251 DVDD.n250 4.5005
R19996 DVDD.n235 DVDD.n234 4.5005
R19997 DVDD.n93 DVDD.n92 4.5005
R19998 DVDD.n212 DVDD.n211 4.5005
R19999 DVDD.n136 DVDD.n135 4.5005
R20000 DVDD.n104 DVDD.n103 4.5005
R20001 DVDD.n112 DVDD.n108 4.5005
R20002 DVDD.n169 DVDD.n168 4.5005
R20003 DVDD.n171 DVDD.n170 4.5005
R20004 DVDD.n176 DVDD.n175 4.5005
R20005 DVDD.n179 DVDD.n178 4.5005
R20006 DVDD.n182 DVDD.n181 4.5005
R20007 DVDD.n198 DVDD.n197 4.5005
R20008 DVDD.n195 DVDD.n194 4.5005
R20009 DVDD.n190 DVDD.n189 4.5005
R20010 DVDD.n146 DVDD.n144 4.5005
R20011 DVDD DVDD.n145 4.5005
R20012 DVDD.n177 DVDD.n158 4.5005
R20013 DVDD.n183 DVDD.n155 4.5005
R20014 DVDD.n193 DVDD.n184 4.5005
R20015 DVDD.n188 DVDD.n187 4.5005
R20016 DVDD.n148 DVDD.n147 4.5005
R20017 DVDD.n29 DVDD.n28 4.5005
R20018 DVDD.n31 DVDD.n30 4.5005
R20019 DVDD.n36 DVDD.n35 4.5005
R20020 DVDD.n39 DVDD.n38 4.5005
R20021 DVDD.n42 DVDD.n41 4.5005
R20022 DVDD.n58 DVDD.n57 4.5005
R20023 DVDD.n55 DVDD.n54 4.5005
R20024 DVDD.n50 DVDD.n49 4.5005
R20025 DVDD.n6 DVDD.n4 4.5005
R20026 DVDD DVDD.n5 4.5005
R20027 DVDD.n37 DVDD.n18 4.5005
R20028 DVDD.n43 DVDD.n15 4.5005
R20029 DVDD.n53 DVDD.n44 4.5005
R20030 DVDD.n48 DVDD.n47 4.5005
R20031 DVDD.n8 DVDD.n7 4.5005
R20032 DVDD.n313 DVDD.n312 4.32258
R20033 DVDD.n81 DVDD.n80 4.32258
R20034 DVDD.n230 DVDD.n227 4.32258
R20035 DVDD.n131 DVDD.n128 4.32258
R20036 DVDD.n294 DVDD.n293 3.76521
R20037 DVDD.n294 DVDD.n287 3.34378
R20038 DVDD.n298 DVDD.n297 3.18888
R20039 DVDD.n186 DVDD.n185 3.09891
R20040 DVDD.n46 DVDD.n45 3.09891
R20041 DVDD.n171 DVDD.n167 3.03311
R20042 DVDD.n179 DVDD.n154 3.03311
R20043 DVDD.n199 DVDD.n198 3.03311
R20044 DVDD.n190 DVDD.n150 3.03311
R20045 DVDD DVDD.n203 3.03311
R20046 DVDD.n31 DVDD.n27 3.03311
R20047 DVDD.n39 DVDD.n14 3.03311
R20048 DVDD.n59 DVDD.n58 3.03311
R20049 DVDD.n50 DVDD.n10 3.03311
R20050 DVDD DVDD.n63 3.03311
R20051 DVDD.n293 DVDD.n288 2.82403
R20052 DVDD DVDD.n295 2.78431
R20053 DVDD.n289 DVDD.n278 2.54327
R20054 DVDD DVDD.n307 1.93032
R20055 DVDD DVDD.n73 1.93032
R20056 DVDD.n232 DVDD 1.93032
R20057 DVDD.n133 DVDD 1.93032
R20058 DVDD.n278 DVDD 1.8288
R20059 DVDD DVDD.n141 1.75727
R20060 DVDD DVDD.n1 1.75727
R20061 DVDD.n307 DVDD 1.61911
R20062 DVDD.n73 DVDD 1.61911
R20063 DVDD.n232 DVDD 1.61911
R20064 DVDD.n133 DVDD 1.61911
R20065 DVDD.n291 DVDD.n290 1.43457
R20066 DVDD.n318 DVDD 1.11892
R20067 DVDD.n84 DVDD 1.11892
R20068 DVDD.n221 DVDD 1.11892
R20069 DVDD.n122 DVDD 1.11892
R20070 DVDD.n244 DVDD.n239 0.433917
R20071 DVDD.n318 DVDD.n317 0.417167
R20072 DVDD.n84 DVDD.n83 0.417167
R20073 DVDD.n222 DVDD.n221 0.417167
R20074 DVDD.n123 DVDD.n122 0.417167
R20075 DVDD.n297 DVDD.n296 0.397498
R20076 DVDD.n262 DVDD 0.377693
R20077 DVDD.n241 DVDD 0.377693
R20078 DVDD.n98 DVDD 0.377693
R20079 DVDD.n109 DVDD 0.377693
R20080 DVDD.n289 DVDD.n288 0.376971
R20081 DVDD.n261 DVDD.n260 0.312991
R20082 DVDD.n208 DVDD.n140 0.296735
R20083 DVDD DVDD.n94 0.272089
R20084 DVDD.n314 DVDD 0.268044
R20085 DVDD.n74 DVDD 0.268044
R20086 DVDD DVDD.n231 0.268044
R20087 DVDD DVDD.n132 0.268044
R20088 DVDD DVDD.n105 0.243821
R20089 DVDD DVDD.n0 0.238894
R20090 DVDD.n254 DVDD 0.234986
R20091 DVDD DVDD.n207 0.206256
R20092 DVDD.n261 DVDD.n67 0.185367
R20093 DVDD.n295 DVDD.n278 0.163151
R20094 DVDD.n317 DVDD.n314 0.158395
R20095 DVDD.n83 DVDD.n74 0.158395
R20096 DVDD.n231 DVDD.n222 0.158395
R20097 DVDD.n132 DVDD.n123 0.158395
R20098 DVDD.n262 DVDD 0.15085
R20099 DVDD.n241 DVDD 0.15085
R20100 DVDD.n98 DVDD 0.15085
R20101 DVDD.n109 DVDD 0.15085
R20102 DVDD.n119 DVDD 0.14163
R20103 DVDD.n218 DVDD 0.14163
R20104 DVDD DVDD.n322 0.124528
R20105 DVDD DVDD.n253 0.12237
R20106 DVDD.n265 DVDD 0.112517
R20107 DVDD.n209 DVDD.n208 0.110693
R20108 DVDD.n307 DVDD.n306 0.0728282
R20109 DVDD.n73 DVDD.n71 0.0728282
R20110 DVDD.n233 DVDD.n232 0.0728282
R20111 DVDD.n134 DVDD.n133 0.0728282
R20112 DVDD.n263 DVDD.n262 0.0471653
R20113 DVDD.n242 DVDD.n241 0.0471653
R20114 DVDD.n99 DVDD.n98 0.0471653
R20115 DVDD.n110 DVDD.n109 0.0471653
R20116 DVDD.n319 DVDD.n318 0.0401723
R20117 DVDD.n85 DVDD.n84 0.0401723
R20118 DVDD.n221 DVDD.n220 0.0401723
R20119 DVDD.n122 DVDD.n121 0.0401723
R20120 DVDD.n260 DVDD.n259 0.0390074
R20121 DVDD.n239 DVDD.n238 0.0390074
R20122 DVDD.n140 DVDD.n139 0.0390074
R20123 DVDD.n305 DVDD.n304 0.0378134
R20124 DVDD.n256 DVDD.n255 0.0378134
R20125 DVDD.n235 DVDD.n91 0.0378134
R20126 DVDD.n136 DVDD.n102 0.0378134
R20127 DVDD.n319 DVDD.n276 0.0359671
R20128 DVDD.n250 DVDD.n85 0.0359671
R20129 DVDD.n242 DVDD.n240 0.0359671
R20130 DVDD.n220 DVDD.n92 0.0359671
R20131 DVDD.n212 DVDD.n99 0.0359671
R20132 DVDD.n121 DVDD.n103 0.0359671
R20133 DVDD.n110 DVDD.n108 0.0359671
R20134 DVDD.n321 DVDD.n320 0.0357113
R20135 DVDD.n269 DVDD.n268 0.0357113
R20136 DVDD.n252 DVDD.n251 0.0357113
R20137 DVDD.n251 DVDD.n86 0.0357113
R20138 DVDD.n247 DVDD.n86 0.0357113
R20139 DVDD.n247 DVDD.n246 0.0357113
R20140 DVDD.n246 DVDD.n88 0.0357113
R20141 DVDD.n243 DVDD.n88 0.0357113
R20142 DVDD.n219 DVDD.n93 0.0357113
R20143 DVDD.n216 DVDD.n93 0.0357113
R20144 DVDD.n216 DVDD.n215 0.0357113
R20145 DVDD.n215 DVDD.n97 0.0357113
R20146 DVDD.n211 DVDD.n97 0.0357113
R20147 DVDD.n211 DVDD.n210 0.0357113
R20148 DVDD.n120 DVDD.n104 0.0357113
R20149 DVDD.n117 DVDD.n104 0.0357113
R20150 DVDD.n117 DVDD.n107 0.0357113
R20151 DVDD.n113 DVDD.n107 0.0357113
R20152 DVDD.n113 DVDD.n112 0.0357113
R20153 DVDD.n112 DVDD.n111 0.0357113
R20154 DVDD.n273 DVDD.n272 0.035465
R20155 DVDD.n267 DVDD.n266 0.035465
R20156 DVDD.n250 DVDD.n249 0.035465
R20157 DVDD.n249 DVDD.n248 0.035465
R20158 DVDD.n248 DVDD.n87 0.035465
R20159 DVDD.n240 DVDD.n87 0.035465
R20160 DVDD.n96 DVDD.n92 0.035465
R20161 DVDD.n214 DVDD.n96 0.035465
R20162 DVDD.n214 DVDD.n213 0.035465
R20163 DVDD.n213 DVDD.n212 0.035465
R20164 DVDD.n116 DVDD.n103 0.035465
R20165 DVDD.n116 DVDD.n115 0.035465
R20166 DVDD.n115 DVDD.n114 0.035465
R20167 DVDD.n114 DVDD.n108 0.035465
R20168 DVDD.n257 DVDD.n256 0.0340821
R20169 DVDD.n236 DVDD.n235 0.0340821
R20170 DVDD.n137 DVDD.n136 0.0340821
R20171 DVDD.n169 DVDD.n159 0.0333947
R20172 DVDD.n184 DVDD.n143 0.0333947
R20173 DVDD.n147 DVDD.n141 0.0333947
R20174 DVDD.n29 DVDD.n19 0.0333947
R20175 DVDD.n44 DVDD.n3 0.0333947
R20176 DVDD.n7 DVDD.n1 0.0333947
R20177 DVDD.n303 DVDD.n302 0.0333467
R20178 DVDD.n258 DVDD.n70 0.0333467
R20179 DVDD.n234 DVDD.n90 0.0333467
R20180 DVDD.n135 DVDD.n101 0.0333467
R20181 DVDD.n170 DVDD.n165 0.03175
R20182 DVDD.n196 DVDD.n195 0.03175
R20183 DVDD.n30 DVDD.n25 0.03175
R20184 DVDD.n56 DVDD.n55 0.03175
R20185 DVDD.n177 DVDD.n176 0.0284605
R20186 DVDD.n189 DVDD.n188 0.0284605
R20187 DVDD.n37 DVDD.n36 0.0284605
R20188 DVDD.n49 DVDD.n48 0.0284605
R20189 DVDD.n306 DVDD 0.0274625
R20190 DVDD.n71 DVDD 0.0274625
R20191 DVDD DVDD.n233 0.0274625
R20192 DVDD DVDD.n134 0.0274625
R20193 DVDD.n296 DVDD 0.0264901
R20194 DVDD.n296 DVDD 0.0262353
R20195 DVDD.n165 DVDD.n164 0.0255919
R20196 DVDD.n25 DVDD.n24 0.0255919
R20197 DVDD.n164 DVDD.n163 0.0252368
R20198 DVDD.n163 DVDD.n142 0.0252368
R20199 DVDD.n24 DVDD.n23 0.0252368
R20200 DVDD.n23 DVDD.n2 0.0252368
R20201 DVDD.n197 DVDD.n183 0.0251711
R20202 DVDD.n57 DVDD.n43 0.0251711
R20203 DVDD.n111 DVDD.n106 0.024355
R20204 DVDD.n239 DVDD.n89 0.0242975
R20205 DVDD.n94 DVDD.n89 0.0242975
R20206 DVDD.n119 DVDD.n118 0.024
R20207 DVDD.n118 DVDD.n106 0.024
R20208 DVDD.n218 DVDD.n217 0.024
R20209 DVDD.n217 DVDD.n95 0.024
R20210 DVDD.n209 DVDD.n95 0.024
R20211 DVDD.n192 DVDD.n191 0.0232804
R20212 DVDD.n52 DVDD.n51 0.0232804
R20213 DVDD.n194 DVDD.n156 0.0226963
R20214 DVDD.n54 DVDD.n16 0.0226963
R20215 DVDD.n178 DVDD.n157 0.0218816
R20216 DVDD.n205 DVDD.n144 0.0218816
R20217 DVDD.n38 DVDD.n17 0.0218816
R20218 DVDD.n65 DVDD.n4 0.0218816
R20219 DVDD.n162 DVDD.n160 0.021528
R20220 DVDD.n22 DVDD.n20 0.021528
R20221 DVDD.n140 DVDD.n100 0.0215056
R20222 DVDD.n105 DVDD.n100 0.0215056
R20223 DVDD.n299 DVDD.n298 0.0213889
R20224 DVDD.n299 DVDD.n0 0.0213889
R20225 DVDD.n322 DVDD.n275 0.0213889
R20226 DVDD.n275 DVDD.n270 0.0213889
R20227 DVDD.n270 DVDD.n265 0.0213889
R20228 DVDD.n260 DVDD.n68 0.0210464
R20229 DVDD.n254 DVDD.n68 0.0210464
R20230 DVDD.n253 DVDD.n72 0.0208243
R20231 DVDD.n245 DVDD.n72 0.0208243
R20232 DVDD.n245 DVDD.n244 0.0208243
R20233 DVDD.n182 DVDD.n157 0.0185921
R20234 DVDD.n205 DVDD.n145 0.0185921
R20235 DVDD.n42 DVDD.n17 0.0185921
R20236 DVDD.n65 DVDD.n5 0.0185921
R20237 DVDD.n198 DVDD.n155 0.0180234
R20238 DVDD.n148 DVDD 0.0180234
R20239 DVDD.n58 DVDD.n15 0.0180234
R20240 DVDD.n8 DVDD 0.0180234
R20241 DVDD.n172 DVDD.n165 0.016626
R20242 DVDD.n32 DVDD.n25 0.016626
R20243 DVDD.n180 DVDD.n179 0.0156869
R20244 DVDD.n204 DVDD.n146 0.0156869
R20245 DVDD.n40 DVDD.n39 0.0156869
R20246 DVDD.n64 DVDD.n6 0.0156869
R20247 DVDD.n190 DVDD.n186 0.0153479
R20248 DVDD.n50 DVDD.n46 0.0153479
R20249 DVDD.n183 DVDD.n182 0.0153026
R20250 DVDD.n147 DVDD.n145 0.0153026
R20251 DVDD.n43 DVDD.n42 0.0153026
R20252 DVDD.n7 DVDD.n5 0.0153026
R20253 DVDD.n175 DVDD.n174 0.0151028
R20254 DVDD.n35 DVDD.n34 0.0151028
R20255 DVDD.n297 DVDD 0.0143584
R20256 DVDD.n181 DVDD.n180 0.0133505
R20257 DVDD.n204 DVDD 0.0133505
R20258 DVDD.n41 DVDD.n40 0.0133505
R20259 DVDD.n64 DVDD 0.0133505
R20260 DVDD.n178 DVDD.n177 0.0120132
R20261 DVDD.n188 DVDD.n144 0.0120132
R20262 DVDD.n38 DVDD.n37 0.0120132
R20263 DVDD.n48 DVDD.n4 0.0120132
R20264 DVDD.n181 DVDD.n155 0.011014
R20265 DVDD.n41 DVDD.n15 0.011014
R20266 DVDD DVDD.n303 0.0105365
R20267 DVDD DVDD.n70 0.0105365
R20268 DVDD.n234 DVDD 0.0105365
R20269 DVDD.n135 DVDD 0.0105365
R20270 DVDD.n207 DVDD.n142 0.0103947
R20271 DVDD.n67 DVDD.n2 0.0103947
R20272 DVDD.n207 DVDD.n141 0.00951292
R20273 DVDD.n67 DVDD.n1 0.00951292
R20274 DVDD.n149 DVDD.n148 0.00926168
R20275 DVDD.n9 DVDD.n8 0.00926168
R20276 DVDD DVDD.n261 0.00885556
R20277 DVDD.n197 DVDD.n196 0.00872368
R20278 DVDD.n57 DVDD.n56 0.00872368
R20279 DVDD.n179 DVDD.n158 0.00867757
R20280 DVDD.n187 DVDD.n146 0.00867757
R20281 DVDD.n39 DVDD.n18 0.00867757
R20282 DVDD.n47 DVDD.n6 0.00867757
R20283 DVDD.n187 DVDD.n186 0.00750551
R20284 DVDD.n47 DVDD.n46 0.00750551
R20285 DVDD.n172 DVDD.n171 0.00692523
R20286 DVDD.n32 DVDD.n31 0.00692523
R20287 DVDD.n198 DVDD.n156 0.00634112
R20288 DVDD.n58 DVDD.n16 0.00634112
R20289 DVDD.n174 DVDD.n158 0.00575701
R20290 DVDD.n34 DVDD.n18 0.00575701
R20291 DVDD.n176 DVDD.n159 0.00543421
R20292 DVDD.n189 DVDD.n143 0.00543421
R20293 DVDD.n36 DVDD.n19 0.00543421
R20294 DVDD.n49 DVDD.n3 0.00543421
R20295 DVDD.n208 DVDD 0.00493889
R20296 DVDD.n259 DVDD.n258 0.00482522
R20297 DVDD.n238 DVDD.n90 0.00482522
R20298 DVDD.n139 DVDD.n101 0.00482522
R20299 DVDD.n301 DVDD.n300 0.00423134
R20300 DVDD.n257 DVDD.n69 0.00423134
R20301 DVDD.n237 DVDD.n236 0.00423134
R20302 DVDD.n138 DVDD.n137 0.00423134
R20303 DVDD.n175 DVDD.n160 0.00400467
R20304 DVDD.n191 DVDD.n190 0.00400467
R20305 DVDD.n35 DVDD.n20 0.00400467
R20306 DVDD.n51 DVDD.n50 0.00400467
R20307 DVDD.n168 DVDD.n162 0.00283645
R20308 DVDD.n28 DVDD.n22 0.00283645
R20309 DVDD.n207 DVDD.n206 0.00258889
R20310 DVDD.n67 DVDD.n66 0.00258889
R20311 DVDD DVDD.n149 0.00225234
R20312 DVDD DVDD.n9 0.00225234
R20313 DVDD.n170 DVDD.n169 0.00214474
R20314 DVDD.n195 DVDD.n184 0.00214474
R20315 DVDD.n30 DVDD.n29 0.00214474
R20316 DVDD.n55 DVDD.n44 0.00214474
R20317 DVDD.n194 DVDD.n193 0.00166822
R20318 DVDD.n54 DVDD.n53 0.00166822
R20319 DVDD.n321 DVDD.n319 0.00135292
R20320 DVDD.n264 DVDD.n263 0.00135292
R20321 DVDD.n252 DVDD.n85 0.00135292
R20322 DVDD.n243 DVDD.n242 0.00135292
R20323 DVDD.n220 DVDD.n219 0.00135292
R20324 DVDD.n210 DVDD.n99 0.00135292
R20325 DVDD.n121 DVDD.n120 0.00135292
R20326 DVDD.n111 DVDD.n110 0.00135292
R20327 DVDD.n306 DVDD.n305 0.00135241
R20328 DVDD.n255 DVDD.n71 0.00135241
R20329 DVDD.n233 DVDD.n91 0.00135241
R20330 DVDD.n134 DVDD.n102 0.00135241
R20331 DVDD.n238 DVDD.n237 0.00117863
R20332 DVDD.n139 DVDD.n138 0.00117863
R20333 DVDD.n259 DVDD.n69 0.00117863
R20334 DVDD.n300 DVDD.n277 0.00117863
R20335 DVDD.n171 DVDD.n161 0.00108411
R20336 DVDD.n168 DVDD.n161 0.00108411
R20337 DVDD.n193 DVDD.n192 0.00108411
R20338 DVDD.n31 DVDD.n21 0.00108411
R20339 DVDD.n28 DVDD.n21 0.00108411
R20340 DVDD.n53 DVDD.n52 0.00108411
R20341 DVDD.n117 DVDD.n116 0.00085506
R20342 DVDD.n114 DVDD.n113 0.00085506
R20343 DVDD.n160 DVDD.n159 0.00085506
R20344 DVDD.n180 DVDD.n157 0.00085506
R20345 DVDD.n191 DVDD.n143 0.00085506
R20346 DVDD.n205 DVDD.n204 0.00085506
R20347 DVDD.n216 DVDD.n96 0.00085506
R20348 DVDD.n213 DVDD.n97 0.00085506
R20349 DVDD.n246 DVDD.n87 0.00085506
R20350 DVDD.n249 DVDD.n86 0.00085506
R20351 DVDD.n20 DVDD.n19 0.00085506
R20352 DVDD.n40 DVDD.n17 0.00085506
R20353 DVDD.n51 DVDD.n3 0.00085506
R20354 DVDD.n65 DVDD.n64 0.00085506
R20355 DVDD.n269 DVDD.n267 0.00085506
R20356 DVDD.n274 DVDD.n273 0.00085506
R20357 DVDD.n120 DVDD.n119 0.000855023
R20358 DVDD.n118 DVDD.n117 0.000855023
R20359 DVDD.n113 DVDD.n106 0.000855023
R20360 DVDD.n138 DVDD.n100 0.000855023
R20361 DVDD.n105 DVDD.n102 0.000855023
R20362 DVDD.n164 DVDD.n159 0.000855023
R20363 DVDD.n163 DVDD.n157 0.000855023
R20364 DVDD.n196 DVDD.n142 0.000855023
R20365 DVDD.n206 DVDD.n143 0.000855023
R20366 DVDD.n206 DVDD.n205 0.000855023
R20367 DVDD.n219 DVDD.n218 0.000855023
R20368 DVDD.n217 DVDD.n216 0.000855023
R20369 DVDD.n97 DVDD.n95 0.000855023
R20370 DVDD.n210 DVDD.n209 0.000855023
R20371 DVDD.n237 DVDD.n89 0.000855023
R20372 DVDD.n94 DVDD.n91 0.000855023
R20373 DVDD.n246 DVDD.n245 0.000855023
R20374 DVDD.n86 DVDD.n72 0.000855023
R20375 DVDD.n253 DVDD.n252 0.000855023
R20376 DVDD.n244 DVDD.n243 0.000855023
R20377 DVDD.n69 DVDD.n68 0.000855023
R20378 DVDD.n255 DVDD.n254 0.000855023
R20379 DVDD.n24 DVDD.n19 0.000855023
R20380 DVDD.n23 DVDD.n17 0.000855023
R20381 DVDD.n56 DVDD.n2 0.000855023
R20382 DVDD.n66 DVDD.n3 0.000855023
R20383 DVDD.n66 DVDD.n65 0.000855023
R20384 DVDD.n270 DVDD.n269 0.000855023
R20385 DVDD.n275 DVDD.n274 0.000855023
R20386 DVDD.n322 DVDD.n321 0.000855023
R20387 DVDD.n300 DVDD.n299 0.000855023
R20388 DVDD.n305 DVDD.n0 0.000855023
R20389 DVDD.n265 DVDD.n264 0.000855023
R20390 DVDD.n196 DVDD.n156 0.000854948
R20391 DVDD.n56 DVDD.n16 0.000854948
R20392 DVDD.n236 DVDD.n90 0.000500614
R20393 DVDD.n137 DVDD.n101 0.000500614
R20394 DVDD.n302 DVDD.n301 0.000500614
R20395 DVDD.n258 DVDD.n257 0.000500614
R20396 DVDD.n215 DVDD.n214 0.000500461
R20397 DVDD.n115 DVDD.n107 0.000500461
R20398 DVDD.n272 DVDD.n271 0.000500461
R20399 DVDD.n248 DVDD.n247 0.000500461
R20400 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 120.01
R20401 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 92.9415
R20402 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n4 92.5005
R20403 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 92.4623
R20404 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 73.195
R20405 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 72.1651
R20406 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 29.4833
R20407 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 27.6955
R20408 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 27.6955
R20409 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 15.4607
R20410 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 9.3005
R20411 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 9.3005
R20412 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 9.02061
R20413 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 9.01961
R20414 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n26 8.28285
R20415 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n16 8.28285
R20416 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 5.64756
R20417 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 5.32161
R20418 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 5.31894
R20419 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n31 4.14168
R20420 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n23 4.14168
R20421 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n19 4.14168
R20422 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 4.03426
R20423 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n9 3.93153
R20424 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n33 3.76521
R20425 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n14 3.76521
R20426 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 3.20519
R20427 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 3.07304
R20428 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 3.04478
R20429 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 3.03311
R20430 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 3.03311
R20431 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 3.03311
R20432 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n27 3.01226
R20433 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n17 3.01226
R20434 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n34 2.63579
R20435 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n15 2.63579
R20436 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 2.47579
R20437 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 2.27623
R20438 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 2.25932
R20439 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 2.25932
R20440 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 1.51198
R20441 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 1.15307
R20442 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 1.04295
R20443 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n7 0.753441
R20444 a_5299_620.n27 a_5299_620.t9 129.037
R20445 a_5299_620.n27 a_5299_620.t8 68.9672
R20446 a_5299_620.n42 a_5299_620.n40 8.0439
R20447 a_5299_620.n3 a_5299_620.n20 7.45281
R20448 a_5299_620.n35 a_5299_620.n33 5.63
R20449 a_5299_620.n36 a_5299_620.t0 5.5395
R20450 a_5299_620.n36 a_5299_620.t7 5.5395
R20451 a_5299_620.n24 a_5299_620.t4 5.5395
R20452 a_5299_620.n24 a_5299_620.t3 5.5395
R20453 a_5299_620.n2 a_5299_620.n1 4.54542
R20454 a_5299_620.n6 a_5299_620.n39 4.5005
R20455 a_5299_620.n5 a_5299_620.n31 4.5005
R20456 a_5299_620.n0 a_5299_620.n42 4.5005
R20457 a_5299_620.n0 a_5299_620.n46 4.5005
R20458 a_5299_620.n4 a_5299_620.n23 4.5005
R20459 a_5299_620.n2 a_5299_620.n17 4.5005
R20460 a_5299_620.n2 a_5299_620.n12 4.5005
R20461 a_5299_620.n2 a_5299_620.n14 4.5005
R20462 a_5299_620.n47 a_5299_620.n0 4.3695
R20463 a_5299_620.n23 a_5299_620.n21 4.14168
R20464 a_5299_620.n7 a_5299_620.n26 3.82535
R20465 a_5299_620.n39 a_5299_620.n38 3.76521
R20466 a_5299_620.n46 a_5299_620.n45 3.76521
R20467 a_5299_620.n31 a_5299_620.n28 3.38874
R20468 a_5299_620.n42 a_5299_620.n41 3.38874
R20469 a_5299_620.n12 a_5299_620.n11 3.38238
R20470 a_5299_620.n44 a_5299_620.t6 3.3065
R20471 a_5299_620.n44 a_5299_620.t5 3.3065
R20472 a_5299_620.t2 a_5299_620.n50 3.3065
R20473 a_5299_620.n50 a_5299_620.t1 3.3065
R20474 a_5299_620.n31 a_5299_620.n30 3.01226
R20475 a_5299_620.n16 a_5299_620.n15 3.01226
R20476 a_5299_620.n39 a_5299_620.n37 2.63579
R20477 a_5299_620.n3 a_5299_620.n19 2.63579
R20478 a_5299_620.n7 a_5299_620.n27 2.423
R20479 a_5299_620.n18 a_5299_620.n48 2.2208
R20480 a_5299_620.n25 a_5299_620.n24 2.12431
R20481 a_5299_620.n47 a_5299_620.n6 3.11985
R20482 a_5299_620.n6 a_5299_620.n36 1.90815
R20483 a_5299_620.n12 a_5299_620.n10 1.88285
R20484 a_5299_620.n0 a_5299_620.n44 2.5496
R20485 a_5299_620.n23 a_5299_620.n22 1.50638
R20486 a_5299_620.n50 a_5299_620.n49 1.33804
R20487 a_5299_620.n14 a_5299_620.n13 1.12991
R20488 a_5299_620.n17 a_5299_620.n16 1.12991
R20489 a_5299_620.n26 a_5299_620.n4 0.922158
R20490 a_5299_620.n48 a_5299_620.n7 0.824928
R20491 a_5299_620.n10 a_5299_620.n9 0.753441
R20492 a_5299_620.n7 a_5299_620.n47 0.504252
R20493 a_5299_620.n1 a_5299_620.n8 0.376971
R20494 a_5299_620.n49 a_5299_620.n18 0.352626
R20495 a_5299_620.n32 a_5299_620.n35 0.278788
R20496 a_5299_620.n33 a_5299_620.n34 0.161367
R20497 a_5299_620.n28 a_5299_620.n29 0.150167
R20498 a_5299_620.n6 a_5299_620.n5 0.143833
R20499 a_5299_620.n5 a_5299_620.n32 0.1366
R20500 a_5299_620.n4 a_5299_620.n3 4.63501
R20501 a_5299_620.n0 a_5299_620.n43 1.11727
R20502 a_5299_620.n4 a_5299_620.n25 0.422157
R20503 a_5299_620.n18 a_5299_620.n2 0.221203
R20504 A1.n66 A1.n65 185
R20505 A1.n64 A1.n57 185
R20506 A1.n24 A1.n15 185
R20507 A1.n23 A1.n22 185
R20508 A1.n69 A1.t4 120.037
R20509 A1.t5 A1.n14 120.037
R20510 A1.n59 A1.n57 112.831
R20511 A1.n22 A1.n21 112.831
R20512 A1.n68 A1.n67 104.172
R20513 A1.n27 A1.n26 104.172
R20514 A1.n68 A1.n56 92.5005
R20515 A1.n28 A1.n27 92.5005
R20516 A1.t4 A1.n68 66.8281
R20517 A1.n27 A1.t5 66.8281
R20518 A1.n6 A1.t0 35.2053
R20519 A1.n3 A1.t1 34.0571
R20520 A1.n67 A1.n66 29.4833
R20521 A1.n26 A1.n15 29.4833
R20522 A1.n1 A1.t6 27.6955
R20523 A1.n1 A1.t7 27.6955
R20524 A1.n45 A1.n44 19.0955
R20525 A1.n69 A1.n56 15.4558
R20526 A1.n28 A1.n14 15.4558
R20527 A1.n64 A1.n63 13.5534
R20528 A1.n23 A1.n18 13.5534
R20529 A1.n2 A1.n1 9.67857
R20530 A1.n41 A1.n34 9.30581
R20531 A1.n59 A1.n58 9.30424
R20532 A1.n21 A1.n20 9.30413
R20533 A1.n40 A1.n39 9.3005
R20534 A1.n46 A1.n45 9.3005
R20535 A1.n71 A1.n70 9.3005
R20536 A1.n55 A1.n52 9.3005
R20537 A1.n67 A1.n55 9.3005
R20538 A1.n63 A1.n62 9.3005
R20539 A1.n72 A1.n54 9.3005
R20540 A1.n29 A1.n13 9.3005
R20541 A1.n25 A1.n11 9.3005
R20542 A1.n26 A1.n25 9.3005
R20543 A1.n18 A1.n17 9.3005
R20544 A1.n31 A1.n30 9.3005
R20545 A1.n71 A1.n56 9.03579
R20546 A1.n29 A1.n28 9.03579
R20547 A1.n43 A1.n41 8.49366
R20548 A1.n43 A1.t2 8.2655
R20549 A1.n43 A1.t3 8.2655
R20550 A1.n44 A1.n43 7.97749
R20551 A1.n42 A1.n40 7.26743
R20552 A1.n43 A1.n42 6.15568
R20553 A1.n65 A1.n55 5.64756
R20554 A1.n25 A1.n24 5.64756
R20555 A1.n41 A1.n35 4.89462
R20556 A1.n60 A1.n59 4.89462
R20557 A1.n21 A1.n19 4.89462
R20558 A1.n73 A1.n55 4.51815
R20559 A1.n72 A1.n71 4.51815
R20560 A1.n25 A1.n12 4.51815
R20561 A1.n30 A1.n29 4.51815
R20562 A1.n5 A1.n4 4.5005
R20563 A1.n4 A1.n2 4.5005
R20564 A1.n51 A1.n9 4.5005
R20565 A1.n49 A1.n9 4.5005
R20566 A1.n51 A1.n50 4.5005
R20567 A1.n50 A1.n49 4.5005
R20568 A1.n74 A1.n53 4.5005
R20569 A1.n75 A1.n8 4.5005
R20570 A1.n53 A1.n8 4.5005
R20571 A1.n75 A1.n74 4.5005
R20572 A1.n48 A1.n32 4.5005
R20573 A1.n47 A1.n36 4.5005
R20574 A1.n48 A1.n47 4.5005
R20575 A1.n36 A1.n32 4.5005
R20576 A1.n38 A1.n33 4.5005
R20577 A1.n66 A1.n57 3.93153
R20578 A1.n22 A1.n15 3.93153
R20579 A1.n19 A1.n9 3.03311
R20580 A1.n50 A1.n12 3.03311
R20581 A1.n60 A1.n8 3.03311
R20582 A1.n74 A1.n73 3.03311
R20583 A1.n47 A1.n35 3.03311
R20584 A1.n3 A1.n0 2.2714
R20585 A1.n58 A1.n7 2.25261
R20586 A1.n20 A1.n10 2.25256
R20587 A1.n34 A1.n33 2.25127
R20588 A1.n37 A1.n33 2.24434
R20589 A1.n73 A1.n72 1.88285
R20590 A1.n30 A1.n12 1.88285
R20591 A1.n45 A1.n35 1.50638
R20592 A1.n63 A1.n60 1.50638
R20593 A1.n19 A1.n18 1.50638
R20594 A1.n16 A1.n10 1.49213
R20595 A1.n70 A1.n69 1.49212
R20596 A1.n61 A1.n7 1.49182
R20597 A1.n14 A1.n13 1.49166
R20598 A1.n78 A1 0.830453
R20599 A1.n65 A1.n64 0.753441
R20600 A1.n24 A1.n23 0.753441
R20601 A1.n44 A1.n40 0.521921
R20602 A1.n78 A1 0.377842
R20603 A1.n77 A1.n6 0.29767
R20604 A1.n49 A1.n48 0.238951
R20605 A1.n77 A1.n76 0.196255
R20606 A1 A1.n77 0.1855
R20607 A1.n6 A1.n5 0.149538
R20608 A1.n75 A1.n51 0.124821
R20609 A1.n42 A1.n32 0.0579027
R20610 A1 A1.n78 0.0478131
R20611 A1.n62 A1.n61 0.0396286
R20612 A1.n17 A1.n16 0.0383668
R20613 A1.n46 A1.n37 0.0314092
R20614 A1.n5 A1.n0 0.0281442
R20615 A1.n39 A1.n37 0.0271357
R20616 A1.n61 A1.n52 0.0202788
R20617 A1.n16 A1.n11 0.0196501
R20618 A1.n51 A1.n10 0.0168043
R20619 A1.n36 A1.n33 0.016125
R20620 A1.n74 A1.n52 0.013431
R20621 A1.n70 A1.n54 0.013431
R20622 A1.n50 A1.n11 0.013
R20623 A1.n31 A1.n13 0.013
R20624 A1.n38 A1.n32 0.0122521
R20625 A1.n58 A1.n8 0.0117689
R20626 A1.n20 A1.n9 0.0114102
R20627 A1.n47 A1.n34 0.0100704
R20628 A1.n76 A1.n7 0.0100109
R20629 A1.n74 A1.n54 0.00588793
R20630 A1.n50 A1.n31 0.00570833
R20631 A1.n62 A1.n8 0.00481034
R20632 A1.n47 A1.n46 0.0047735
R20633 A1.n17 A1.n9 0.00466667
R20634 A1.n53 A1.n7 0.00457609
R20635 A1.n76 A1.n75 0.00457609
R20636 A1.n2 A1.n0 0.00410577
R20637 A1.n39 A1.n38 0.00370513
R20638 A1.n48 A1.n33 0.00253804
R20639 A1.n4 A1.n3 0.00185919
R20640 A1.n49 A1.n10 0.0018587
R20641 a_5299_1782.n21 a_5299_1782.t8 60.2505
R20642 a_5299_1782.n42 a_5299_1782.t9 60.2505
R20643 a_5299_1782.n64 a_5299_1782.t4 60.2505
R20644 a_5299_1782.n76 a_5299_1782.t6 60.2505
R20645 a_5299_1782.n2 a_5299_1782.n84 9.3005
R20646 a_5299_1782.n2 a_5299_1782.n85 9.3005
R20647 a_5299_1782.n2 a_5299_1782.n83 9.3005
R20648 a_5299_1782.n83 a_5299_1782.n82 9.3005
R20649 a_5299_1782.n3 a_5299_1782.n73 9.3005
R20650 a_5299_1782.n4 a_5299_1782.n57 9.3005
R20651 a_5299_1782.n4 a_5299_1782.n56 9.3005
R20652 a_5299_1782.n4 a_5299_1782.n63 9.3005
R20653 a_5299_1782.n63 a_5299_1782.n62 9.3005
R20654 a_5299_1782.n3 a_5299_1782.n72 9.3005
R20655 a_5299_1782.n72 a_5299_1782.n71 9.3005
R20656 a_5299_1782.n3 a_5299_1782.n74 9.3005
R20657 a_5299_1782.n5 a_5299_1782.n51 9.3005
R20658 a_5299_1782.n6 a_5299_1782.n35 9.3005
R20659 a_5299_1782.n6 a_5299_1782.n34 9.3005
R20660 a_5299_1782.n6 a_5299_1782.n41 9.3005
R20661 a_5299_1782.n41 a_5299_1782.n40 9.3005
R20662 a_5299_1782.n5 a_5299_1782.n50 9.3005
R20663 a_5299_1782.n50 a_5299_1782.n49 9.3005
R20664 a_5299_1782.n5 a_5299_1782.n52 9.3005
R20665 a_5299_1782.n7 a_5299_1782.n29 9.3005
R20666 a_5299_1782.n7 a_5299_1782.n28 9.3005
R20667 a_5299_1782.n28 a_5299_1782.n27 9.3005
R20668 a_5299_1782.n7 a_5299_1782.n30 9.3005
R20669 a_5299_1782.n1 a_5299_1782.n91 9.3005
R20670 a_5299_1782.n119 a_5299_1782.n118 10.743
R20671 a_5299_1782.n65 a_5299_1782.n64 8.76429
R20672 a_5299_1782.n43 a_5299_1782.n42 8.76429
R20673 a_5299_1782.n26 a_5299_1782.n25 7.45411
R20674 a_5299_1782.n39 a_5299_1782.n38 7.45411
R20675 a_5299_1782.n48 a_5299_1782.n47 7.45411
R20676 a_5299_1782.n61 a_5299_1782.n60 7.45411
R20677 a_5299_1782.n70 a_5299_1782.n69 7.45411
R20678 a_5299_1782.n81 a_5299_1782.n80 7.45411
R20679 a_5299_1782.n22 a_5299_1782.n21 6.80105
R20680 a_5299_1782.n77 a_5299_1782.n76 6.80105
R20681 a_5299_1782.n24 a_5299_1782.n23 5.64756
R20682 a_5299_1782.n37 a_5299_1782.n36 5.64756
R20683 a_5299_1782.n46 a_5299_1782.n45 5.64756
R20684 a_5299_1782.n59 a_5299_1782.n58 5.64756
R20685 a_5299_1782.n68 a_5299_1782.n67 5.64756
R20686 a_5299_1782.n79 a_5299_1782.n78 5.64756
R20687 a_5299_1782.n96 a_5299_1782.t5 5.5395
R20688 a_5299_1782.n96 a_5299_1782.t7 5.5395
R20689 a_5299_1782.n90 a_5299_1782.n89 4.95584
R20690 a_5299_1782.n31 a_5299_1782.n20 4.73575
R20691 a_5299_1782.n33 a_5299_1782.n32 4.73575
R20692 a_5299_1782.n53 a_5299_1782.n19 4.73575
R20693 a_5299_1782.n55 a_5299_1782.n54 4.73575
R20694 a_5299_1782.n75 a_5299_1782.n18 4.73575
R20695 a_5299_1782.n87 a_5299_1782.n86 4.73575
R20696 a_5299_1782.n11 a_5299_1782.n13 4.66695
R20697 a_5299_1782.n66 a_5299_1782.n65 4.6505
R20698 a_5299_1782.n44 a_5299_1782.n43 4.6505
R20699 a_5299_1782.n1 a_5299_1782.n17 4.5005
R20700 a_5299_1782.n13 a_5299_1782.n99 4.5005
R20701 a_5299_1782.n12 a_5299_1782.n95 4.5005
R20702 a_5299_1782.n0 a_5299_1782.n110 4.5005
R20703 a_5299_1782.n0 a_5299_1782.n105 4.5005
R20704 a_5299_1782.n10 a_5299_1782.n117 4.5005
R20705 a_5299_1782.n9 a_5299_1782.n114 4.5005
R20706 a_5299_1782.n9 a_5299_1782.n112 4.5005
R20707 a_5299_1782.n110 a_5299_1782.n109 4.14168
R20708 a_5299_1782.n99 a_5299_1782.n98 3.76521
R20709 a_5299_1782.n114 a_5299_1782.n113 3.76521
R20710 a_5299_1782.n7 a_5299_1782.n22 3.42768
R20711 a_5299_1782.n2 a_5299_1782.n77 3.42768
R20712 a_5299_1782.n95 a_5299_1782.n93 3.38874
R20713 a_5299_1782.n17 a_5299_1782.n16 3.38874
R20714 a_5299_1782.n106 a_5299_1782.t1 3.3065
R20715 a_5299_1782.n106 a_5299_1782.t0 3.3065
R20716 a_5299_1782.n119 a_5299_1782.t2 3.3065
R20717 a_5299_1782.t3 a_5299_1782.n119 3.3065
R20718 a_5299_1782.n95 a_5299_1782.n94 3.01226
R20719 a_5299_1782.n17 a_5299_1782.n15 3.01226
R20720 a_5299_1782.n119 a_5299_1782.n100 2.66355
R20721 a_5299_1782.n99 a_5299_1782.n97 2.63579
R20722 a_5299_1782.n104 a_5299_1782.n103 2.25932
R20723 a_5299_1782.n116 a_5299_1782.n115 2.25932
R20724 a_5299_1782.n9 a_5299_1782.n11 1.68471
R20725 a_5299_1782.n107 a_5299_1782.n106 1.46875
R20726 a_5299_1782.n27 a_5299_1782.n26 0.994314
R20727 a_5299_1782.n40 a_5299_1782.n39 0.994314
R20728 a_5299_1782.n49 a_5299_1782.n48 0.994314
R20729 a_5299_1782.n62 a_5299_1782.n61 0.994314
R20730 a_5299_1782.n71 a_5299_1782.n70 0.994314
R20731 a_5299_1782.n82 a_5299_1782.n81 0.994314
R20732 a_5299_1782.n28 a_5299_1782.n24 0.753441
R20733 a_5299_1782.n41 a_5299_1782.n37 0.753441
R20734 a_5299_1782.n50 a_5299_1782.n46 0.753441
R20735 a_5299_1782.n63 a_5299_1782.n59 0.753441
R20736 a_5299_1782.n72 a_5299_1782.n68 0.753441
R20737 a_5299_1782.n83 a_5299_1782.n79 0.753441
R20738 a_5299_1782.n102 a_5299_1782.n101 0.603501
R20739 a_5299_1782.n119 a_5299_1782.n10 2.11613
R20740 a_5299_1782.n8 a_5299_1782.n107 0.555049
R20741 a_5299_1782.n33 a_5299_1782.n31 0.458354
R20742 a_5299_1782.n55 a_5299_1782.n53 0.458354
R20743 a_5299_1782.n13 a_5299_1782.n96 1.90913
R20744 a_5299_1782.n11 a_5299_1782.n102 0.710352
R20745 a_5299_1782.n110 a_5299_1782.n108 0.376971
R20746 a_5299_1782.n105 a_5299_1782.n104 0.376971
R20747 a_5299_1782.n112 a_5299_1782.n111 0.376971
R20748 a_5299_1782.n117 a_5299_1782.n116 0.376971
R20749 a_5299_1782.n88 a_5299_1782.n75 0.229427
R20750 a_5299_1782.n88 a_5299_1782.n87 0.229427
R20751 a_5299_1782.n90 a_5299_1782.n88 0.215848
R20752 a_5299_1782.n31 a_5299_1782.n7 0.205546
R20753 a_5299_1782.n6 a_5299_1782.n33 0.205546
R20754 a_5299_1782.n53 a_5299_1782.n5 0.205546
R20755 a_5299_1782.n4 a_5299_1782.n55 0.205546
R20756 a_5299_1782.n75 a_5299_1782.n3 0.205546
R20757 a_5299_1782.n87 a_5299_1782.n2 0.205546
R20758 a_5299_1782.n44 a_5299_1782.n6 0.190717
R20759 a_5299_1782.n5 a_5299_1782.n44 0.190717
R20760 a_5299_1782.n66 a_5299_1782.n4 0.190717
R20761 a_5299_1782.n3 a_5299_1782.n66 0.190717
R20762 a_5299_1782.n0 a_5299_1782.n8 0.183965
R20763 a_5299_1782.n12 a_5299_1782.n1 0.169804
R20764 a_5299_1782.n15 a_5299_1782.n14 0.161367
R20765 a_5299_1782.n93 a_5299_1782.n92 0.150167
R20766 a_5299_1782.n1 a_5299_1782.n90 0.140745
R20767 a_5299_1782.n13 a_5299_1782.n12 0.14187
R20768 a_5299_1782.n10 a_5299_1782.n9 0.135427
R20769 a_5299_1782.n102 a_5299_1782.n0 0.107619
R20770 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 136.804
R20771 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 136.325
R20772 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 119.999
R20773 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 93.9023
R20774 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 93.3044
R20775 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 93.0848
R20776 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n4 92.5005
R20777 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 92.4623
R20778 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 69.2281
R20779 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 29.4833
R20780 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 27.6955
R20781 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 27.6955
R20782 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 15.4626
R20783 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n16 9.3005
R20784 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n8 9.3005
R20785 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n7 9.3005
R20786 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 9.3005
R20787 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 9.3005
R20788 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n15 9.3005
R20789 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n17 9.3005
R20790 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 9.02061
R20791 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 9.02061
R20792 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n34 8.28285
R20793 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n21 8.28285
R20794 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 5.64756
R20795 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 5.31864
R20796 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n42 4.14168
R20797 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n28 4.14168
R20798 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 4.06959
R20799 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n11 3.93153
R20800 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n40 3.76521
R20801 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n33 3.76521
R20802 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n24 3.76521
R20803 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n19 3.76521
R20804 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n36 3.38874
R20805 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n22 3.38874
R20806 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 3.0736
R20807 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 3.07249
R20808 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 3.07078
R20809 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 3.04338
R20810 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 3.03311
R20811 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 3.03311
R20812 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 3.03311
R20813 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n39 2.63579
R20814 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n20 2.63579
R20815 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 2.27447
R20816 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 2.25932
R20817 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 2.25932
R20818 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 1.80772
R20819 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n30 1.61433
R20820 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 1.45534
R20821 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 1.19419
R20822 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n9 0.753441
R20823 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 0.719888
R20824 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 0.22499
R20825 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 0.176176
R20826 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 2.36361
R20827 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 2.36353
R20828 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 1.14499
R20829 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 1.00043
R20830 B2.n66 B2.n65 185
R20831 B2.n64 B2.n57 185
R20832 B2.n24 B2.n15 185
R20833 B2.n23 B2.n22 185
R20834 B2.n69 B2.t0 120.037
R20835 B2.t1 B2.n14 120.037
R20836 B2.n59 B2.n57 112.831
R20837 B2.n22 B2.n21 112.831
R20838 B2.n68 B2.n67 104.172
R20839 B2.n27 B2.n26 104.172
R20840 B2.n68 B2.n56 92.5005
R20841 B2.n28 B2.n27 92.5005
R20842 B2.t0 B2.n68 66.8281
R20843 B2.n27 B2.t1 66.8281
R20844 B2.n6 B2.t4 35.2053
R20845 B2.n3 B2.t5 34.0571
R20846 B2.n67 B2.n66 29.4833
R20847 B2.n26 B2.n15 29.4833
R20848 B2.n1 B2.t3 27.6955
R20849 B2.n1 B2.t2 27.6955
R20850 B2.n45 B2.n44 19.0955
R20851 B2.n69 B2.n56 15.4558
R20852 B2.n28 B2.n14 15.4558
R20853 B2.n64 B2.n63 13.5534
R20854 B2.n23 B2.n18 13.5534
R20855 B2.n2 B2.n1 9.67857
R20856 B2.n41 B2.n34 9.30581
R20857 B2.n59 B2.n58 9.30424
R20858 B2.n21 B2.n20 9.30413
R20859 B2.n40 B2.n39 9.3005
R20860 B2.n46 B2.n45 9.3005
R20861 B2.n71 B2.n70 9.3005
R20862 B2.n55 B2.n52 9.3005
R20863 B2.n67 B2.n55 9.3005
R20864 B2.n63 B2.n62 9.3005
R20865 B2.n72 B2.n54 9.3005
R20866 B2.n29 B2.n13 9.3005
R20867 B2.n25 B2.n11 9.3005
R20868 B2.n26 B2.n25 9.3005
R20869 B2.n18 B2.n17 9.3005
R20870 B2.n31 B2.n30 9.3005
R20871 B2.n71 B2.n56 9.03579
R20872 B2.n29 B2.n28 9.03579
R20873 B2.n43 B2.n41 8.49366
R20874 B2.n43 B2.t7 8.2655
R20875 B2.n43 B2.t6 8.2655
R20876 B2.n44 B2.n43 7.97749
R20877 B2.n42 B2.n40 7.26743
R20878 B2.n43 B2.n42 6.15568
R20879 B2.n65 B2.n55 5.64756
R20880 B2.n25 B2.n24 5.64756
R20881 B2.n41 B2.n35 4.89462
R20882 B2.n60 B2.n59 4.89462
R20883 B2.n21 B2.n19 4.89462
R20884 B2.n73 B2.n55 4.51815
R20885 B2.n72 B2.n71 4.51815
R20886 B2.n25 B2.n12 4.51815
R20887 B2.n30 B2.n29 4.51815
R20888 B2.n5 B2.n4 4.5005
R20889 B2.n4 B2.n2 4.5005
R20890 B2.n51 B2.n9 4.5005
R20891 B2.n49 B2.n9 4.5005
R20892 B2.n51 B2.n50 4.5005
R20893 B2.n50 B2.n49 4.5005
R20894 B2.n74 B2.n53 4.5005
R20895 B2.n75 B2.n8 4.5005
R20896 B2.n53 B2.n8 4.5005
R20897 B2.n75 B2.n74 4.5005
R20898 B2.n48 B2.n32 4.5005
R20899 B2.n47 B2.n36 4.5005
R20900 B2.n48 B2.n47 4.5005
R20901 B2.n36 B2.n32 4.5005
R20902 B2.n38 B2.n33 4.5005
R20903 B2.n66 B2.n57 3.93153
R20904 B2.n22 B2.n15 3.93153
R20905 B2.n19 B2.n9 3.03311
R20906 B2.n50 B2.n12 3.03311
R20907 B2.n60 B2.n8 3.03311
R20908 B2.n74 B2.n73 3.03311
R20909 B2.n47 B2.n35 3.03311
R20910 B2.n3 B2.n0 2.2714
R20911 B2.n58 B2.n7 2.25261
R20912 B2.n20 B2.n10 2.25256
R20913 B2.n34 B2.n33 2.25127
R20914 B2.n37 B2.n33 2.24434
R20915 B2.n73 B2.n72 1.88285
R20916 B2.n30 B2.n12 1.88285
R20917 B2.n45 B2.n35 1.50638
R20918 B2.n63 B2.n60 1.50638
R20919 B2.n19 B2.n18 1.50638
R20920 B2.n16 B2.n10 1.49213
R20921 B2.n70 B2.n69 1.49212
R20922 B2.n61 B2.n7 1.49182
R20923 B2.n14 B2.n13 1.49166
R20924 B2.n78 B2 0.90653
R20925 B2.n65 B2.n64 0.753441
R20926 B2.n24 B2.n23 0.753441
R20927 B2.n44 B2.n40 0.521921
R20928 B2.n78 B2 0.384338
R20929 B2.n77 B2.n6 0.29767
R20930 B2.n49 B2.n48 0.238951
R20931 B2.n77 B2.n76 0.196255
R20932 B2 B2.n77 0.1855
R20933 B2.n6 B2.n5 0.149538
R20934 B2 B2.n78 0.135601
R20935 B2.n75 B2.n51 0.124821
R20936 B2.n42 B2.n32 0.0579027
R20937 B2.n62 B2.n61 0.0396286
R20938 B2.n17 B2.n16 0.0383668
R20939 B2.n46 B2.n37 0.0314092
R20940 B2.n5 B2.n0 0.0281442
R20941 B2.n39 B2.n37 0.0271357
R20942 B2.n61 B2.n52 0.0202788
R20943 B2.n16 B2.n11 0.0196501
R20944 B2.n51 B2.n10 0.0168043
R20945 B2.n36 B2.n33 0.016125
R20946 B2.n74 B2.n52 0.013431
R20947 B2.n70 B2.n54 0.013431
R20948 B2.n50 B2.n11 0.013
R20949 B2.n31 B2.n13 0.013
R20950 B2.n38 B2.n32 0.0122521
R20951 B2.n58 B2.n8 0.0117689
R20952 B2.n20 B2.n9 0.0114102
R20953 B2.n47 B2.n34 0.0100704
R20954 B2.n76 B2.n7 0.0100109
R20955 B2.n74 B2.n54 0.00588793
R20956 B2.n50 B2.n31 0.00570833
R20957 B2.n62 B2.n8 0.00481034
R20958 B2.n47 B2.n46 0.0047735
R20959 B2.n17 B2.n9 0.00466667
R20960 B2.n53 B2.n7 0.00457609
R20961 B2.n76 B2.n75 0.00457609
R20962 B2.n2 B2.n0 0.00410577
R20963 B2.n39 B2.n38 0.00370513
R20964 B2.n48 B2.n33 0.00253804
R20965 B2.n4 B2.n3 0.00185919
R20966 B2.n49 B2.n10 0.0018587
R20967 SELB.n1 SELB.t4 186.374
R20968 SELB.n1 SELB.t5 170.308
R20969 SELB.n2 SELB.n1 139.876
R20970 SELB.n5 SELB.t1 84.8325
R20971 SELB.n6 SELB.t0 84.8325
R20972 SELB.n6 SELB.n5 60.1541
R20973 SELB.n7 SELB.n6 50.1642
R20974 SELB.n5 SELB.t3 48.6825
R20975 SELB.n6 SELB.t2 48.6825
R20976 SELB.n0 SELB 42.9181
R20977 SELB.n9 SELB 17.169
R20978 SELB.n8 SELB.n7 15.2731
R20979 SELB.n0 SELB 12.8005
R20980 SELB.n9 SELB.n8 4.77356
R20981 SELB.n10 SELB 2.74121
R20982 SELB.n3 SELB 2.73914
R20983 SELB SELB.n8 2.13383
R20984 SELB SELB.n2 1.61978
R20985 SELB.n4 SELB.n3 1.31185
R20986 SELB.n7 SELB 1.1768
R20987 SELB.n2 SELB.n0 0.925801
R20988 SELB.n12 SELB.n11 0.661383
R20989 SELB.n11 SELB 0.563656
R20990 SELB.n13 SELB 0.34425
R20991 SELB.n10 SELB 0.321549
R20992 SELB SELB.n14 0.0255
R20993 SELB.n14 SELB.n13 0.0194024
R20994 SELB SELB.n9 0.0180439
R20995 SELB SELB.n12 0.0151341
R20996 SELB.n3 SELB 0.00770734
R20997 SELB.n12 SELB 0.00415854
R20998 SELB.n13 SELB 0.00171951
R20999 SELB.n12 SELB.n4 0.000502048
R21000 SELB.n11 SELB.n10 0.000500307
R21001 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 120.01
R21002 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 92.9415
R21003 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n4 92.5005
R21004 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 92.4623
R21005 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 73.195
R21006 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 72.1651
R21007 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 29.4833
R21008 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 27.6955
R21009 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 27.6955
R21010 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 15.4607
R21011 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 9.3005
R21012 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 9.3005
R21013 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 9.02061
R21014 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n29 9.01961
R21015 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n26 8.28285
R21016 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n16 8.28285
R21017 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 5.64756
R21018 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 5.32161
R21019 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 5.31894
R21020 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 4.14168
R21021 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n23 4.14168
R21022 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n20 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n19 4.14168
R21023 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 4.03426
R21024 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n9 3.93153
R21025 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n33 3.76521
R21026 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n14 3.76521
R21027 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 3.20519
R21028 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 3.07304
R21029 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n36 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 3.04478
R21030 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 3.03311
R21031 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n20 3.03311
R21032 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 3.03311
R21033 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n27 3.01226
R21034 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 3.01226
R21035 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n34 2.63579
R21036 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n15 2.63579
R21037 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 2.47579
R21038 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n36 2.27623
R21039 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 2.25932
R21040 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 2.25932
R21041 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 1.51198
R21042 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 1.15307
R21043 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 1.04295
R21044 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n7 0.753441
R21045 A2.n66 A2.n65 185
R21046 A2.n64 A2.n57 185
R21047 A2.n24 A2.n15 185
R21048 A2.n23 A2.n22 185
R21049 A2.n69 A2.t6 120.037
R21050 A2.t7 A2.n14 120.037
R21051 A2.n59 A2.n57 112.831
R21052 A2.n22 A2.n21 112.831
R21053 A2.n68 A2.n67 104.172
R21054 A2.n27 A2.n26 104.172
R21055 A2.n68 A2.n56 92.5005
R21056 A2.n28 A2.n27 92.5005
R21057 A2.t6 A2.n68 66.8281
R21058 A2.n27 A2.t7 66.8281
R21059 A2.n6 A2.t2 35.2053
R21060 A2.n3 A2.t3 34.0571
R21061 A2.n67 A2.n66 29.4833
R21062 A2.n26 A2.n15 29.4833
R21063 A2.n1 A2.t4 27.6955
R21064 A2.n1 A2.t5 27.6955
R21065 A2.n45 A2.n44 19.0955
R21066 A2.n69 A2.n56 15.4558
R21067 A2.n28 A2.n14 15.4558
R21068 A2.n64 A2.n63 13.5534
R21069 A2.n23 A2.n18 13.5534
R21070 A2.n2 A2.n1 9.67857
R21071 A2.n41 A2.n34 9.30581
R21072 A2.n59 A2.n58 9.30424
R21073 A2.n21 A2.n20 9.30413
R21074 A2.n40 A2.n39 9.3005
R21075 A2.n46 A2.n45 9.3005
R21076 A2.n71 A2.n70 9.3005
R21077 A2.n55 A2.n52 9.3005
R21078 A2.n67 A2.n55 9.3005
R21079 A2.n63 A2.n62 9.3005
R21080 A2.n72 A2.n54 9.3005
R21081 A2.n29 A2.n13 9.3005
R21082 A2.n25 A2.n11 9.3005
R21083 A2.n26 A2.n25 9.3005
R21084 A2.n18 A2.n17 9.3005
R21085 A2.n31 A2.n30 9.3005
R21086 A2.n71 A2.n56 9.03579
R21087 A2.n29 A2.n28 9.03579
R21088 A2.n43 A2.n41 8.49366
R21089 A2.n43 A2.t0 8.2655
R21090 A2.n43 A2.t1 8.2655
R21091 A2.n44 A2.n43 7.97749
R21092 A2.n42 A2.n40 7.26743
R21093 A2.n43 A2.n42 6.15568
R21094 A2.n65 A2.n55 5.64756
R21095 A2.n25 A2.n24 5.64756
R21096 A2.n41 A2.n35 4.89462
R21097 A2.n60 A2.n59 4.89462
R21098 A2.n21 A2.n19 4.89462
R21099 A2.n73 A2.n55 4.51815
R21100 A2.n72 A2.n71 4.51815
R21101 A2.n25 A2.n12 4.51815
R21102 A2.n30 A2.n29 4.51815
R21103 A2.n5 A2.n4 4.5005
R21104 A2.n4 A2.n2 4.5005
R21105 A2.n51 A2.n9 4.5005
R21106 A2.n49 A2.n9 4.5005
R21107 A2.n51 A2.n50 4.5005
R21108 A2.n50 A2.n49 4.5005
R21109 A2.n74 A2.n53 4.5005
R21110 A2.n75 A2.n8 4.5005
R21111 A2.n53 A2.n8 4.5005
R21112 A2.n75 A2.n74 4.5005
R21113 A2.n48 A2.n32 4.5005
R21114 A2.n47 A2.n36 4.5005
R21115 A2.n48 A2.n47 4.5005
R21116 A2.n36 A2.n32 4.5005
R21117 A2.n38 A2.n33 4.5005
R21118 A2.n66 A2.n57 3.93153
R21119 A2.n22 A2.n15 3.93153
R21120 A2.n19 A2.n9 3.03311
R21121 A2.n50 A2.n12 3.03311
R21122 A2.n60 A2.n8 3.03311
R21123 A2.n74 A2.n73 3.03311
R21124 A2.n47 A2.n35 3.03311
R21125 A2.n3 A2.n0 2.2714
R21126 A2.n58 A2.n7 2.25261
R21127 A2.n20 A2.n10 2.25256
R21128 A2.n34 A2.n33 2.25127
R21129 A2.n37 A2.n33 2.24434
R21130 A2.n73 A2.n72 1.88285
R21131 A2.n30 A2.n12 1.88285
R21132 A2.n45 A2.n35 1.50638
R21133 A2.n63 A2.n60 1.50638
R21134 A2.n19 A2.n18 1.50638
R21135 A2.n16 A2.n10 1.49213
R21136 A2.n70 A2.n69 1.49212
R21137 A2.n61 A2.n7 1.49182
R21138 A2.n14 A2.n13 1.49166
R21139 A2.n78 A2 1.01398
R21140 A2.n65 A2.n64 0.753441
R21141 A2.n24 A2.n23 0.753441
R21142 A2.n44 A2.n40 0.521921
R21143 A2.n78 A2 0.399268
R21144 A2.n77 A2.n6 0.29767
R21145 A2.n49 A2.n48 0.238951
R21146 A2.n77 A2.n76 0.196255
R21147 A2 A2.n77 0.1855
R21148 A2.n6 A2.n5 0.149538
R21149 A2 A2.n78 0.129964
R21150 A2.n75 A2.n51 0.124821
R21151 A2.n42 A2.n32 0.0579027
R21152 A2.n62 A2.n61 0.0396286
R21153 A2.n17 A2.n16 0.0383668
R21154 A2.n46 A2.n37 0.0314092
R21155 A2.n5 A2.n0 0.0281442
R21156 A2.n39 A2.n37 0.0271357
R21157 A2.n61 A2.n52 0.0202788
R21158 A2.n16 A2.n11 0.0196501
R21159 A2.n51 A2.n10 0.0168043
R21160 A2.n36 A2.n33 0.016125
R21161 A2.n74 A2.n52 0.013431
R21162 A2.n70 A2.n54 0.013431
R21163 A2.n50 A2.n11 0.013
R21164 A2.n31 A2.n13 0.013
R21165 A2.n38 A2.n32 0.0122521
R21166 A2.n58 A2.n8 0.0117689
R21167 A2.n20 A2.n9 0.0114102
R21168 A2.n47 A2.n34 0.0100704
R21169 A2.n76 A2.n7 0.0100109
R21170 A2.n74 A2.n54 0.00588793
R21171 A2.n50 A2.n31 0.00570833
R21172 A2.n62 A2.n8 0.00481034
R21173 A2.n47 A2.n46 0.0047735
R21174 A2.n17 A2.n9 0.00466667
R21175 A2.n53 A2.n7 0.00457609
R21176 A2.n76 A2.n75 0.00457609
R21177 A2.n2 A2.n0 0.00410577
R21178 A2.n39 A2.n38 0.00370513
R21179 A2.n48 A2.n33 0.00253804
R21180 A2.n4 A2.n3 0.00185919
R21181 A2.n49 A2.n10 0.0018587
C0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVDD 0.0946f
C1 a_10442_n5795# VDD 0.335f
C2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_11235_n6821# 0.00288f
C3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00684f
C4 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 DVDD 0.126f
C5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp A1 2.59e-19
C6 a_10542_n5707# B2 0.00545f
C7 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.00152f
C8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_0.l0 8.17e-19
C9 a_4184_n6773# DVDD 0.24f
C10 a_10809_9307# a_10811_8247# 0.139f
C11 a_7889_n6842# SELB 0.0046f
C12 a_7196_n5728# DVDD 0.117f
C13 EF_AMUX21m_1.array_1ls_1tgm_0.l0 a_4184_n6773# 0.0217f
C14 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.282f
C15 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp VDD 2.65f
C16 a_10442_n5795# a_10810_n6777# 0.139f
C17 a_8403_n6064# a_7889_n6842# 2.63e-19
C18 a_3816_n5791# a_4184_n6773# 0.139f
C19 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_7889_n6842# 7.05e-21
C20 comparator_top_0.comparator_bias_0.VBP comparator_top_0.VINM 0.0131f
C21 a_11749_n6043# VDD 0.489f
C22 a_10542_n5707# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.0154f
C23 A1 A2 6.92e-20
C24 a_6351_6657# VDD 0.684f
C25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 B1 2.1e-19
C26 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_11235_n6821# 7.05e-21
C27 VSS A1 9e-20
C28 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.34f
C29 A2 B1 7.46e-20
C30 a_5123_n6039# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.145f
C31 a_11271_4224# VO 0.0548f
C32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 VDD 2.18f
C33 a_7464_n6798# DVDD 0.236f
C34 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.124f
C35 a_6349_9307# a_6351_7717# 0.14f
C36 B1 B2 6.81e-20
C37 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.668f
C38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_10442_n5795# 0.00188f
C39 a_10442_n5795# DVDD 0.437f
C40 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 a_4609_n6817# 3.13e-19
C41 VDD A2 2.45f
C42 VSS SELA 0.032f
C43 a_11749_n6043# a_10810_n6777# 6.24e-19
C44 VDD VSS 0.152p
C45 a_4609_n6817# A2 0.00722f
C46 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X B1 0.0285f
C47 comparator_top_0.VINM comparator_top_0.VINP 3.44f
C48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 a_11749_n6043# 0.00121f
C49 VDD B2 2.31f
C50 a_5123_n6039# a_4184_n6773# 6.24e-19
C51 a_470_n5812# a_1263_n6838# 8.36e-19
C52 a_470_n5812# A1 3.15e-19
C53 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_7196_n5728# 4.56e-19
C54 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD 1.2f
C55 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 0.839f
C56 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 1.54e-19
C57 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb A2 1.01f
C58 a_470_n5812# SELA 0.235f
C59 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_10542_n5707# 0.00139f
C60 a_11031_3400# VO 0.0102f
C61 a_470_n5812# VDD 0.326f
C62 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_4184_n6773# 7.03e-19
C63 a_838_n6794# VSS 0.0013f
C64 a_10809_9307# a_10811_7187# 4.42e-21
C65 a_10810_n6777# B2 0.00652f
C66 a_11749_n6043# DVDD 0.0136f
C67 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 B2 0.892f
C68 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_7196_n5728# 8.72e-21
C69 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_11749_n6043# 0.00108f
C70 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD 1.2f
C71 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 a_7196_n5728# 6.2e-19
C72 a_570_n5724# VSS 0.00169f
C73 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_3816_n5791# 0.00188f
C74 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_10810_n6777# 4.53e-21
C75 m2_2600_n8446# A1 0.0196f
C76 comparator_top_0.comparator_bias_0.VBN VSS 11.2f
C77 a_7889_n6842# B1 0.007f
C78 a_7096_n5816# SELB 0.235f
C79 a_11271_4224# VDD 0.17f
C80 a_1777_n6060# a_1263_n6838# 2.63e-19
C81 a_1777_n6060# A1 0.00748f
C82 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 DVDD 0.11f
C83 m2_2600_n8446# SELA 0.00706f
C84 a_7096_n5816# a_8403_n6064# 3.88e-20
C85 DVDD A2 0.252f
C86 a_470_n5812# a_838_n6794# 0.139f
C87 comparator_top_0.comparator_bias_0.VBP VDD 10.8f
C88 a_7889_n6842# VDD 0.607f
C89 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp A1 1.51f
C90 VSS DVDD 0.00708f
C91 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_10810_n6777# 7.03e-19
C92 comparator_top_0.VINM a_7096_n5816# 0.00115f
C93 a_1777_n6060# SELA 5.58e-20
C94 DVDD B2 0.305f
C95 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp B2 1.51f
C96 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.282f
C97 a_470_n5812# a_570_n5724# 0.405f
C98 a_1777_n6060# VDD 0.489f
C99 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_7464_n6798# 1.96e-19
C100 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 a_7464_n6798# 1.09e-19
C101 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVDD 0.102f
C102 a_3816_n5791# A2 3.15e-19
C103 comparator_top_0.VINP A1 2.88f
C104 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VDD 2.64f
C105 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 a_10442_n5795# 0.0085f
C106 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_5123_n6039# 0.00108f
C107 a_10809_9307# VDD 0.697f
C108 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD 3.43f
C109 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 a_1263_n6838# 3.13e-19
C110 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 A1 0.965f
C111 comparator_top_0.comparator_0.VOUT VSS 0.872f
C112 a_8403_n6064# SELB 5.62e-20
C113 a_11031_3400# VDD 0.51f
C114 a_3916_n5703# A1 0.00179f
C115 a_470_n5812# DVDD 0.428f
C116 a_7196_n5728# a_7464_n6798# 0.0272f
C117 a_6349_9307# VSS 3.54e-19
C118 comparator_top_0.VINP VDD 12.7f
C119 a_1777_n6060# a_838_n6794# 6.24e-19
C120 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVDD 0.0982f
C121 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 SELA 1.27e-19
C122 comparator_top_0.VINM a_8403_n6064# 0.00136f
C123 comparator_top_0.comparator_bias_0.VBN comparator_top_0.comparator_bias_0.VBP 1.78f
C124 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 VDD 2.16f
C125 a_570_n5724# a_1777_n6060# 0.289f
C126 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 a_5123_n6039# 0.00121f
C127 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.00724f
C128 a_3916_n5703# VDD 1.12f
C129 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.682f
C130 a_11271_4224# a_10975_4108# 0.136f
C131 a_10811_8247# a_10811_7187# 0.14f
C132 a_11271_4224# DVDD 0.449f
C133 a_3916_n5703# a_4609_n6817# 0.265f
C134 a_5123_n6039# A2 0.00717f
C135 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp A2 2.99e-19
C136 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 0.839f
C137 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_570_n5724# 4.56e-19
C138 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.668f
C139 m2_2600_n8446# DVDD 2.22e-19
C140 a_7889_n6842# DVDD 0.188f
C141 EF_AMUX21m_2.array_1ls_1tgm_0.l0 SELB 0.241f
C142 m2_2600_n8446# m3_2600_n8446# 0.262f
C143 a_11235_n6821# EF_AMUX21m_2.array_1ls_1tgm_0.l0 0.00503f
C144 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 2.72e-19
C145 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_1263_n6838# 0.00288f
C146 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X A1 0.0306f
C147 a_1777_n6060# DVDD 0.0139f
C148 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.282f
C149 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_3916_n5703# 0.00139f
C150 a_10542_n5707# a_11235_n6821# 0.265f
C151 comparator_top_0.VINP a_570_n5724# 0.0032f
C152 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 a_838_n6794# 1.09e-19
C153 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 3.11e-19
C154 comparator_top_0.comparator_0.VOUT a_11271_4224# 0.00564f
C155 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X A2 0.028f
C156 comparator_top_0.comparator_bias_0.VBN comparator_top_0.VINP 0.09f
C157 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VSS 8.77e-20
C158 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 a_570_n5724# 6.2e-19
C159 comparator_top_0.VINM a_10542_n5707# 0.0032f
C160 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X SELA 3.51e-19
C161 a_7096_n5816# B1 3.15e-19
C162 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.34f
C163 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD 1.2f
C164 a_11271_4224# a_10965_3602# 7.97e-19
C165 a_10975_4108# a_11031_3400# 0.166f
C166 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 a_4184_n6773# 1.09e-19
C167 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 B2 1.85e-19
C168 a_6351_7717# a_6351_6657# 0.14f
C169 a_11031_3400# DVDD 0.0693f
C170 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 a_7196_n5728# 0.00196f
C171 a_7096_n5816# VDD 0.336f
C172 a_4184_n6773# A2 0.00632f
C173 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.282f
C174 a_7196_n5728# A2 0.00174f
C175 a_10811_8247# VDD 0.508f
C176 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 DVDD 0.124f
C177 a_3916_n5703# DVDD 0.115f
C178 a_10542_n5707# EF_AMUX21m_2.array_1ls_1tgm_0.l0 0.00242f
C179 comparator_top_0.VINP a_3816_n5791# 0.00115f
C180 a_6351_7717# VSS 3.36e-19
C181 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 m3_2600_n8446# 3.28e-19
C182 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.l0 1.69e-19
C183 B1 SELB 0.0643f
C184 comparator_top_0.comparator_0.VOUT a_11031_3400# 0.225f
C185 a_3916_n5703# EF_AMUX21m_1.array_1ls_1tgm_0.l0 0.00242f
C186 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_838_n6794# 7.03e-19
C187 a_7196_n5728# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.0154f
C188 a_10442_n5795# a_11749_n6043# 3.88e-20
C189 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 a_3816_n5791# 0.0085f
C190 a_8403_n6064# B1 0.0072f
C191 a_570_n5724# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.0154f
C192 VDD SELB 0.0248f
C193 a_3816_n5791# a_3916_n5703# 0.405f
C194 a_11031_3400# a_10965_3602# 0.17f
C195 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb B1 1.01f
C196 a_11235_n6821# VDD 0.607f
C197 comparator_top_0.VINM B1 2.88f
C198 a_8403_n6064# VDD 0.489f
C199 a_7464_n6798# A2 0.0018f
C200 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD 3.43f
C201 comparator_top_0.VINM VDD 14.1f
C202 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 a_7889_n6842# 3.13e-19
C203 a_10442_n5795# B2 3.15e-19
C204 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVDD 0.101f
C205 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_7464_n6798# 7.03e-19
C206 comparator_top_0.VINP a_5123_n6039# 0.00136f
C207 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.34f
C208 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X m3_2600_n8446# 2.65e-19
C209 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 5.32e-19
C210 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_0.l0 8.17e-19
C211 a_7096_n5816# DVDD 0.431f
C212 a_11235_n6821# a_10810_n6777# 0.461f
C213 EF_AMUX21m_2.array_1ls_1tgm_0.l0 B1 0.0202f
C214 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 a_11235_n6821# 3.13e-19
C215 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.124f
C216 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.00181f
C217 a_10542_n5707# B1 0.00174f
C218 a_7196_n5728# a_7889_n6842# 0.265f
C219 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 5.32e-19
C220 a_3916_n5703# a_5123_n6039# 0.289f
C221 EF_AMUX21m_2.array_1ls_1tgm_0.l0 VDD 0.0233f
C222 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp A2 1.51f
C223 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 2.72e-19
C224 VDD VO 0.268f
C225 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 0.0365f
C226 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.683f
C227 a_10542_n5707# VDD 1.12f
C228 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.00152f
C229 a_10811_7187# VDD 0.512f
C230 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 0.839f
C231 comparator_top_0.comparator_bias_0.VBN comparator_top_0.VINM 0.494f
C232 a_11749_n6043# B2 0.00734f
C233 DVDD SELB 0.921f
C234 a_3916_n5703# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.0154f
C235 a_6351_6657# VSS 0.0236f
C236 a_11235_n6821# DVDD 0.19f
C237 a_1263_n6838# A1 0.00735f
C238 a_8403_n6064# DVDD 0.0139f
C239 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 A2 0.895f
C240 EF_AMUX21m_2.array_1ls_1tgm_0.l0 a_10810_n6777# 0.0217f
C241 a_7889_n6842# a_7464_n6798# 0.461f
C242 a_10542_n5707# a_10810_n6777# 0.0272f
C243 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.07f
C244 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 a_10542_n5707# 6.2e-19
C245 a_3916_n5703# a_4184_n6773# 0.0272f
C246 a_1263_n6838# SELA 0.00469f
C247 A1 SELA 0.0517f
C248 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_7096_n5816# 0.00188f
C249 a_1263_n6838# VDD 0.607f
C250 VDD A1 2.49f
C251 a_11749_n6043# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.145f
C252 VDD B1 2.45f
C253 VDD SELA 0.0304f
C254 a_10975_4108# VO 0.169f
C255 EF_AMUX21m_2.array_1ls_1tgm_0.l0 DVDD 0.958f
C256 DVDD VO 0.78f
C257 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_7096_n5816# 5.3e-19
C258 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_10542_n5707# 4.56e-19
C259 a_10542_n5707# DVDD 0.116f
C260 a_4609_n6817# VDD 0.607f
C261 a_470_n5812# VSS 0.00701f
C262 a_1263_n6838# a_838_n6794# 0.461f
C263 a_838_n6794# A1 0.0067f
C264 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_4184_n6773# 4.53e-21
C265 a_10810_n6777# B1 0.00151f
C266 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X B2 0.0289f
C267 a_570_n5724# a_1263_n6838# 0.265f
C268 a_570_n5724# A1 0.00546f
C269 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_8403_n6064# 0.00108f
C270 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD 3.43f
C271 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.34f
C272 comparator_top_0.comparator_0.VOUT VO 0.0406f
C273 a_838_n6794# SELA 0.0224f
C274 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.08f
C275 a_7096_n5816# a_7196_n5728# 0.405f
C276 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_4609_n6817# 7.05e-21
C277 a_10810_n6777# VDD 0.154f
C278 a_838_n6794# VDD 0.154f
C279 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 VDD 2.05f
C280 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X SELB 5.01e-19
C281 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.07f
C282 a_570_n5724# SELA 0.00244f
C283 a_10965_3602# VO 0.0178f
C284 a_570_n5724# VDD 1.12f
C285 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 SELB 1.27e-19
C286 comparator_top_0.comparator_bias_0.VBP VSS 2.22f
C287 a_1263_n6838# DVDD 0.189f
C288 DVDD A1 0.372f
C289 comparator_top_0.comparator_bias_0.VBN VDD 9.88f
C290 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00684f
C291 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 1.54e-19
C292 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 a_8403_n6064# 0.00121f
C293 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_3916_n5703# 4.56e-19
C294 m3_2600_n8446# A1 0.308f
C295 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_7889_n6842# 0.00288f
C296 EF_AMUX21m_1.array_1ls_1tgm_0.l0 A1 0.0211f
C297 DVDD B1 0.351f
C298 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp B1 2.53e-19
C299 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 0.839f
C300 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 0.301f
C301 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VSS 3.09e-19
C302 a_7196_n5728# SELB 0.00244f
C303 a_10975_4108# VDD 0.248f
C304 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 a_10810_n6777# 1.09e-19
C305 DVDD SELA 0.921f
C306 a_3816_n5791# A1 0.00526f
C307 VDD DVDD 11.6f
C308 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp VDD 2.65f
C309 a_7096_n5816# a_7464_n6798# 0.139f
C310 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 0.0365f
C311 m3_2600_n8446# SELA 0.00883f
C312 EF_AMUX21m_1.array_1ls_1tgm_0.l0 SELA 0.241f
C313 a_4609_n6817# DVDD 0.186f
C314 a_570_n5724# a_838_n6794# 0.0272f
C315 a_7196_n5728# a_8403_n6064# 0.289f
C316 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb B2 1.01f
C317 EF_AMUX21m_1.array_1ls_1tgm_0.l0 VDD 0.0233f
C318 comparator_top_0.VINP A2 2.83f
C319 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_7196_n5728# 0.00139f
C320 a_4609_n6817# EF_AMUX21m_1.array_1ls_1tgm_0.l0 0.00503f
C321 comparator_top_0.VINM a_7196_n5728# 0.0032f
C322 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 2.6e-19
C323 comparator_top_0.VINP VSS 4.62f
C324 a_470_n5812# a_1777_n6060# 3.88e-20
C325 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 a_3916_n5703# 6.2e-19
C326 a_3816_n5791# VDD 0.335f
C327 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 A2 1.85e-19
C328 a_3916_n5703# A2 0.0054f
C329 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.l0 1.69e-19
C330 a_3816_n5791# a_4609_n6817# 8.36e-19
C331 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_470_n5812# 0.00188f
C332 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 VSS 9.51e-19
C333 comparator_top_0.comparator_0.VOUT VDD 2.93f
C334 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 a_10542_n5707# 0.00162f
C335 a_10810_n6777# DVDD 0.243f
C336 a_838_n6794# DVDD 0.238f
C337 a_6349_9307# VDD 0.701f
C338 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 DVDD 0.147f
C339 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.124f
C340 a_7464_n6798# SELB 0.0221f
C341 a_10965_3602# VDD 0.0939f
C342 a_570_n5724# DVDD 0.116f
C343 comparator_top_0.VINP a_470_n5812# 0.00115f
C344 a_10442_n5795# a_11235_n6821# 8.36e-19
C345 a_8403_n6064# a_7464_n6798# 6.24e-19
C346 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp B1 1.51f
C347 comparator_top_0.VINM a_10442_n5795# 0.00115f
C348 a_5123_n6039# VDD 0.489f
C349 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VDD 2.65f
C350 a_11271_4224# a_11031_3400# 0.25f
C351 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_1263_n6838# 7.05e-21
C352 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb A1 1.01f
C353 a_10975_4108# DVDD 0.466f
C354 a_5123_n6039# a_4609_n6817# 2.63e-19
C355 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 a_7096_n5816# 0.00935f
C356 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_1777_n6060# 0.00108f
C357 m3_2600_n8446# DVDD 0.00989f
C358 EF_AMUX21m_1.array_1ls_1tgm_0.l0 DVDD 0.946f
C359 a_7096_n5816# A2 0.0053f
C360 comparator_top_0.comparator_bias_0.VBP comparator_top_0.VINP 0.355f
C361 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 B1 0.901f
C362 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD 3.42f
C363 a_3816_n5791# DVDD 0.435f
C364 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD 1.21f
C365 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_0.l0 0.235f
C366 comparator_top_0.VINP a_1777_n6060# 0.00136f
C367 a_4184_n6773# A1 0.00161f
C368 a_11749_n6043# a_11235_n6821# 2.63e-19
C369 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 3.05e-19
C370 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 m2_2600_n8446# 4.22e-19
C371 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 VDD 2.16f
C372 comparator_top_0.comparator_0.VOUT a_10975_4108# 0.0135f
C373 a_10442_n5795# a_10542_n5707# 0.405f
C374 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_4609_n6817# 0.00288f
C375 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_0.l0 0.235f
C376 a_7096_n5816# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.00152f
C377 comparator_top_0.comparator_0.VOUT DVDD 0.0256f
C378 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.08f
C379 comparator_top_0.VINM a_11749_n6043# 0.00136f
C380 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 a_1777_n6060# 0.00121f
C381 a_7196_n5728# B1 0.00533f
C382 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 SELB 1.12e-20
C383 a_470_n5812# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.00152f
C384 a_10975_4108# a_10965_3602# 0.249f
C385 a_4184_n6773# VDD 0.154f
C386 a_10965_3602# DVDD 0.033f
C387 A2 SELB 0.0606f
C388 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.124f
C389 a_7196_n5728# VDD 1.12f
C390 a_4609_n6817# a_4184_n6773# 0.461f
C391 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 3.37e-19
C392 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.s0 0.207f
C393 a_6351_7717# VDD 0.522f
C394 a_11235_n6821# B2 0.00724f
C395 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.s0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.s0 2.6e-19
C396 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_570_n5724# 0.00139f
C397 comparator_top_0.VINM A2 0.0517f
C398 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X SELB 3.51e-19
C399 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 0.303f
C400 a_5123_n6039# DVDD 0.0134f
C401 comparator_top_0.VINM VSS 4.14f
C402 comparator_top_0.VINP a_3916_n5703# 0.0032f
C403 comparator_top_0.VINM B2 2.83f
C404 comparator_top_0.comparator_0.VOUT a_10965_3602# 0.0309f
C405 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X m2_2600_n8446# 2.82e-19
C406 a_10542_n5707# a_11749_n6043# 0.289f
C407 a_8403_n6064# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.145f
C408 a_7464_n6798# B1 0.00613f
C409 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.s0 a_3916_n5703# 0.00162f
C410 a_7096_n5816# a_7889_n6842# 8.36e-19
C411 a_10442_n5795# B1 0.00501f
C412 a_1777_n6060# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.145f
C413 a_3816_n5791# a_5123_n6039# 3.88e-20
C414 a_7464_n6798# VDD 0.153f
.ends

