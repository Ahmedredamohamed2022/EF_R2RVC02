magic
tech sky130A
magscale 1 2
timestamp 1699954036
<< locali >>
rect 3345 479 3607 520
rect 2409 455 2855 468
rect 2409 421 2433 455
rect 2467 421 2505 455
rect 2539 421 2577 455
rect 2611 421 2649 455
rect 2683 421 2721 455
rect 2755 421 2793 455
rect 2827 421 2855 455
rect 2409 412 2855 421
rect 3345 445 3390 479
rect 3424 445 3462 479
rect 3496 445 3534 479
rect 3568 445 3607 479
rect 3345 412 3607 445
<< viali >>
rect 2433 421 2467 455
rect 2505 421 2539 455
rect 2577 421 2611 455
rect 2649 421 2683 455
rect 2721 421 2755 455
rect 2793 421 2827 455
rect 3390 445 3424 479
rect 3462 445 3496 479
rect 3534 445 3568 479
<< metal1 >>
rect 325 12170 3827 12274
rect 325 11934 429 12170
rect 2735 3104 2839 3218
rect 6139 3094 6239 3310
rect 349 1791 601 1822
rect 349 1675 382 1791
rect 562 1675 601 1791
rect 349 1632 601 1675
rect 3747 1792 4009 1816
rect 3747 1676 3790 1792
rect 3970 1676 4009 1792
rect 3747 1646 4009 1676
rect 2631 1198 3683 1496
rect 2603 957 3601 1022
rect 2603 841 2675 957
rect 3559 841 3601 957
rect 2603 788 3601 841
rect 1 576 209 582
rect 357 576 609 578
rect 2283 576 2495 578
rect 0 553 2495 576
rect 0 501 390 553
rect 442 501 454 553
rect 506 501 518 553
rect 570 501 2495 553
rect 3763 526 4001 530
rect 3357 520 4011 526
rect 0 486 2495 501
rect 1 484 209 486
rect 357 484 609 486
rect 2283 476 2495 486
rect 3345 498 4011 520
rect 3345 479 3792 498
rect 2283 474 2649 476
rect 2283 455 2865 474
rect 2283 421 2433 455
rect 2467 421 2505 455
rect 2539 421 2577 455
rect 2611 421 2649 455
rect 2683 421 2721 455
rect 2755 421 2793 455
rect 2827 421 2865 455
rect 2283 386 2865 421
rect 3345 445 3390 479
rect 3424 445 3462 479
rect 3496 445 3534 479
rect 3568 446 3792 479
rect 3844 446 3856 498
rect 3908 446 3920 498
rect 3972 446 4011 498
rect 3568 445 4011 446
rect 3345 412 4011 445
rect 3357 410 4011 412
rect 5978 326 6204 1413
rect 4111 226 6204 326
rect 2603 100 6204 226
rect 2603 0 6200 100
<< via1 >>
rect 382 1675 562 1791
rect 3790 1676 3970 1792
rect 2675 841 3559 957
rect 390 501 442 553
rect 454 501 506 553
rect 518 501 570 553
rect 3792 446 3844 498
rect 3856 446 3908 498
rect 3920 446 3972 498
<< metal2 >>
rect 349 1791 601 1822
rect 349 1675 382 1791
rect 562 1675 601 1791
rect 349 1632 601 1675
rect 3747 1792 4009 1816
rect 3747 1676 3790 1792
rect 3970 1676 4009 1792
rect 3747 1646 4009 1676
rect 405 578 535 1632
rect 3801 1258 3939 1646
rect 3799 1128 3939 1258
rect 2603 967 3601 1022
rect 2603 957 2689 967
rect 3545 957 3601 967
rect 2603 841 2675 957
rect 3559 841 3601 957
rect 2603 831 2689 841
rect 3545 831 3601 841
rect 2603 788 3601 831
rect 357 553 609 578
rect 357 501 390 553
rect 442 501 454 553
rect 506 501 518 553
rect 570 501 609 553
rect 3801 530 3939 1128
rect 357 484 609 501
rect 3763 498 4001 530
rect 3763 446 3792 498
rect 3844 446 3856 498
rect 3908 446 3920 498
rect 3972 446 4001 498
rect 3763 410 4001 446
<< via2 >>
rect 2689 957 3545 967
rect 2689 841 3545 957
rect 2689 831 3545 841
<< metal3 >>
rect 3097 8142 3297 8146
rect 693 7942 4289 8142
rect 3023 2022 3165 2026
rect 1001 1890 4671 2022
rect 3021 1022 3153 1890
rect 2603 967 3601 1022
rect 2603 831 2689 967
rect 3545 831 3601 967
rect 2603 788 3601 831
use single_ls_2tgwd_sw  single_ls_2tgwd_sw_0
timestamp 1699954036
transform 1 0 3403 0 1 1296
box 0 -100 2973 10946
use single_ls_2tgwd_sw  single_ls_2tgwd_sw_1
timestamp 1699954036
transform 1 0 3 0 1 1296
box 0 -100 2973 10946
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_0
timestamp 1699954036
transform 1 0 2711 0 1 99
box -66 -43 834 897
<< labels >>
flabel metal1 s 3041 1350 3153 1436 0 FreeSans 976 0 0 0 DVSS
port 1 nsew
flabel metal3 s 3097 7946 3297 8146 0 FreeSans 976 0 0 0 VDD
port 2 nsew
flabel metal1 s 3069 12170 3173 12274 0 FreeSans 976 0 0 0 VO
port 3 nsew
flabel metal3 s 3023 1900 3165 2026 0 FreeSans 195 0 0 0 DVDD
port 4 nsew
flabel metal1 s 1 484 209 582 0 FreeSans 195 0 0 0 SEL
port 5 nsew
flabel metal1 s 2735 3104 2839 3218 0 FreeSans 195 0 0 0 VIN1
port 6 nsew
flabel metal1 s 6139 3094 6239 3310 0 FreeSans 195 0 0 0 VIN2
port 7 nsew
<< end >>
