magic
tech sky130A
magscale 1 2
timestamp 1699286160
<< checkpaint >>
rect -1260 -1260 17674 28088
<< metal1 >>
rect 4516 12957 5316 12986
rect 4516 12905 4539 12957
rect 4591 12905 4603 12957
rect 4655 12905 4667 12957
rect 4719 12905 4731 12957
rect 4783 12905 4795 12957
rect 4847 12905 4859 12957
rect 4911 12905 4923 12957
rect 4975 12905 4987 12957
rect 5039 12905 5051 12957
rect 5103 12905 5115 12957
rect 5167 12905 5179 12957
rect 5231 12905 5243 12957
rect 5295 12905 5316 12957
rect 4516 12876 5316 12905
rect 10992 12960 11812 12990
rect 10992 12908 11033 12960
rect 11085 12908 11097 12960
rect 11149 12908 11161 12960
rect 11213 12908 11225 12960
rect 11277 12908 11289 12960
rect 11341 12908 11353 12960
rect 11405 12908 11417 12960
rect 11469 12908 11481 12960
rect 11533 12908 11545 12960
rect 11597 12908 11609 12960
rect 11661 12908 11673 12960
rect 11725 12908 11737 12960
rect 11789 12908 11812 12960
rect 10992 12880 11812 12908
rect 4542 4375 4648 4418
rect 4542 4323 4570 4375
rect 4622 4323 4648 4375
rect 4542 4311 4648 4323
rect 4542 4259 4570 4311
rect 4622 4259 4648 4311
rect 4542 4247 4648 4259
rect 4542 4195 4570 4247
rect 4622 4195 4648 4247
rect 4542 4183 4648 4195
rect 4542 4131 4570 4183
rect 4622 4131 4648 4183
rect 4542 4119 4648 4131
rect 4542 4067 4570 4119
rect 4622 4067 4648 4119
rect 4542 4055 4648 4067
rect 4542 4003 4570 4055
rect 4622 4003 4648 4055
rect 4542 3991 4648 4003
rect 4542 3939 4570 3991
rect 4622 3939 4648 3991
rect 4542 3927 4648 3939
rect 4542 3875 4570 3927
rect 4622 3875 4648 3927
rect 4542 3820 4648 3875
rect 7940 4359 8046 4406
rect 7940 4307 7966 4359
rect 8018 4307 8046 4359
rect 7940 4295 8046 4307
rect 7940 4243 7966 4295
rect 8018 4243 8046 4295
rect 7940 4231 8046 4243
rect 7940 4179 7966 4231
rect 8018 4179 8046 4231
rect 7940 4167 8046 4179
rect 7940 4115 7966 4167
rect 8018 4115 8046 4167
rect 7940 4103 8046 4115
rect 7940 4051 7966 4103
rect 8018 4051 8046 4103
rect 7940 4039 8046 4051
rect 7940 3987 7966 4039
rect 8018 3987 8046 4039
rect 7940 3975 8046 3987
rect 7940 3923 7966 3975
rect 8018 3923 8046 3975
rect 7940 3911 8046 3923
rect 7940 3859 7966 3911
rect 8018 3859 8046 3911
rect 7940 3808 8046 3859
rect 11136 4365 11242 4414
rect 11136 4313 11162 4365
rect 11214 4313 11242 4365
rect 11136 4301 11242 4313
rect 11136 4249 11162 4301
rect 11214 4249 11242 4301
rect 11136 4237 11242 4249
rect 11136 4185 11162 4237
rect 11214 4185 11242 4237
rect 11136 4173 11242 4185
rect 11136 4121 11162 4173
rect 11214 4121 11242 4173
rect 11136 4109 11242 4121
rect 11136 4057 11162 4109
rect 11214 4057 11242 4109
rect 11136 4045 11242 4057
rect 11136 3993 11162 4045
rect 11214 3993 11242 4045
rect 11136 3981 11242 3993
rect 11136 3929 11162 3981
rect 11214 3929 11242 3981
rect 11136 3917 11242 3929
rect 11136 3865 11162 3917
rect 11214 3865 11242 3917
rect 11136 3816 11242 3865
rect 14538 4363 14644 4412
rect 14538 4311 14568 4363
rect 14620 4311 14644 4363
rect 14538 4299 14644 4311
rect 14538 4247 14568 4299
rect 14620 4247 14644 4299
rect 14538 4235 14644 4247
rect 14538 4183 14568 4235
rect 14620 4183 14644 4235
rect 14538 4171 14644 4183
rect 14538 4119 14568 4171
rect 14620 4119 14644 4171
rect 14538 4107 14644 4119
rect 14538 4055 14568 4107
rect 14620 4055 14644 4107
rect 14538 4043 14644 4055
rect 14538 3991 14568 4043
rect 14620 3991 14644 4043
rect 14538 3979 14644 3991
rect 14538 3927 14568 3979
rect 14620 3927 14644 3979
rect 14538 3915 14644 3927
rect 14538 3863 14568 3915
rect 14620 3863 14644 3915
rect 14538 3814 14644 3863
rect 1799 808 5997 1034
rect 7563 1014 15203 1038
rect 7563 834 15049 1014
rect 15165 834 15203 1014
rect 7563 812 15203 834
<< via1 >>
rect 4539 12905 4591 12957
rect 4603 12905 4655 12957
rect 4667 12905 4719 12957
rect 4731 12905 4783 12957
rect 4795 12905 4847 12957
rect 4859 12905 4911 12957
rect 4923 12905 4975 12957
rect 4987 12905 5039 12957
rect 5051 12905 5103 12957
rect 5115 12905 5167 12957
rect 5179 12905 5231 12957
rect 5243 12905 5295 12957
rect 11033 12908 11085 12960
rect 11097 12908 11149 12960
rect 11161 12908 11213 12960
rect 11225 12908 11277 12960
rect 11289 12908 11341 12960
rect 11353 12908 11405 12960
rect 11417 12908 11469 12960
rect 11481 12908 11533 12960
rect 11545 12908 11597 12960
rect 11609 12908 11661 12960
rect 11673 12908 11725 12960
rect 11737 12908 11789 12960
rect 4570 4323 4622 4375
rect 4570 4259 4622 4311
rect 4570 4195 4622 4247
rect 4570 4131 4622 4183
rect 4570 4067 4622 4119
rect 4570 4003 4622 4055
rect 4570 3939 4622 3991
rect 4570 3875 4622 3927
rect 7966 4307 8018 4359
rect 7966 4243 8018 4295
rect 7966 4179 8018 4231
rect 7966 4115 8018 4167
rect 7966 4051 8018 4103
rect 7966 3987 8018 4039
rect 7966 3923 8018 3975
rect 7966 3859 8018 3911
rect 11162 4313 11214 4365
rect 11162 4249 11214 4301
rect 11162 4185 11214 4237
rect 11162 4121 11214 4173
rect 11162 4057 11214 4109
rect 11162 3993 11214 4045
rect 11162 3929 11214 3981
rect 11162 3865 11214 3917
rect 14568 4311 14620 4363
rect 14568 4247 14620 4299
rect 14568 4183 14620 4235
rect 14568 4119 14620 4171
rect 14568 4055 14620 4107
rect 14568 3991 14620 4043
rect 14568 3927 14620 3979
rect 14568 3863 14620 3915
rect 15049 834 15165 1014
<< metal2 >>
rect 1204 14757 1404 14812
rect 1204 14461 1226 14757
rect 1362 14707 1404 14757
rect 1362 14547 7248 14707
rect 1362 14461 1404 14547
rect 1204 14408 1404 14461
rect 4516 12959 5316 12986
rect 4516 12957 4569 12959
rect 4625 12957 4649 12959
rect 4705 12957 4729 12959
rect 4785 12957 4809 12959
rect 4865 12957 4889 12959
rect 4945 12957 4969 12959
rect 5025 12957 5049 12959
rect 5105 12957 5129 12959
rect 5185 12957 5209 12959
rect 5265 12957 5316 12959
rect 4516 12905 4539 12957
rect 4719 12905 4729 12957
rect 4785 12905 4795 12957
rect 5039 12905 5049 12957
rect 5105 12905 5115 12957
rect 5295 12905 5316 12957
rect 4516 12903 4569 12905
rect 4625 12903 4649 12905
rect 4705 12903 4729 12905
rect 4785 12903 4809 12905
rect 4865 12903 4889 12905
rect 4945 12903 4969 12905
rect 5025 12903 5049 12905
rect 5105 12903 5129 12905
rect 5185 12903 5209 12905
rect 5265 12903 5316 12905
rect 4516 12876 5316 12903
rect 10992 12962 11812 12990
rect 10992 12906 11023 12962
rect 11079 12960 11103 12962
rect 11159 12960 11183 12962
rect 11239 12960 11263 12962
rect 11319 12960 11343 12962
rect 11399 12960 11423 12962
rect 11479 12960 11503 12962
rect 11559 12960 11583 12962
rect 11639 12960 11663 12962
rect 11719 12960 11743 12962
rect 11085 12908 11097 12960
rect 11159 12908 11161 12960
rect 11341 12908 11343 12960
rect 11405 12908 11417 12960
rect 11479 12908 11481 12960
rect 11661 12908 11663 12960
rect 11725 12908 11737 12960
rect 11079 12906 11103 12908
rect 11159 12906 11183 12908
rect 11239 12906 11263 12908
rect 11319 12906 11343 12908
rect 11399 12906 11423 12908
rect 11479 12906 11503 12908
rect 11559 12906 11583 12908
rect 11639 12906 11663 12908
rect 11719 12906 11743 12908
rect 11799 12906 11812 12962
rect 10992 12880 11812 12906
rect 4542 4393 4648 4418
rect 4542 4337 4568 4393
rect 4624 4337 4648 4393
rect 4542 4323 4570 4337
rect 4622 4323 4648 4337
rect 4542 4313 4648 4323
rect 4542 4257 4568 4313
rect 4624 4257 4648 4313
rect 4542 4247 4648 4257
rect 4542 4233 4570 4247
rect 4622 4233 4648 4247
rect 4542 4177 4568 4233
rect 4624 4177 4648 4233
rect 4542 4153 4570 4177
rect 4622 4153 4648 4177
rect 4542 4097 4568 4153
rect 4624 4097 4648 4153
rect 4542 4073 4570 4097
rect 4622 4073 4648 4097
rect 4542 4017 4568 4073
rect 4624 4017 4648 4073
rect 4542 4003 4570 4017
rect 4622 4003 4648 4017
rect 4542 3993 4648 4003
rect 4542 3937 4568 3993
rect 4624 3937 4648 3993
rect 4542 3927 4648 3937
rect 4542 3913 4570 3927
rect 4622 3913 4648 3927
rect 4542 3857 4568 3913
rect 4624 3857 4648 3913
rect 4542 3820 4648 3857
rect 7940 4377 8046 4406
rect 7940 4321 7964 4377
rect 8020 4321 8046 4377
rect 7940 4307 7966 4321
rect 8018 4307 8046 4321
rect 7940 4297 8046 4307
rect 7940 4241 7964 4297
rect 8020 4241 8046 4297
rect 7940 4231 8046 4241
rect 7940 4217 7966 4231
rect 8018 4217 8046 4231
rect 7940 4161 7964 4217
rect 8020 4161 8046 4217
rect 7940 4137 7966 4161
rect 8018 4137 8046 4161
rect 7940 4081 7964 4137
rect 8020 4081 8046 4137
rect 7940 4057 7966 4081
rect 8018 4057 8046 4081
rect 7940 4001 7964 4057
rect 8020 4001 8046 4057
rect 7940 3987 7966 4001
rect 8018 3987 8046 4001
rect 7940 3977 8046 3987
rect 7940 3921 7964 3977
rect 8020 3921 8046 3977
rect 7940 3911 8046 3921
rect 7940 3897 7966 3911
rect 8018 3897 8046 3911
rect 7940 3841 7964 3897
rect 8020 3841 8046 3897
rect 7940 3808 8046 3841
rect 11136 4383 11242 4414
rect 11136 4327 11160 4383
rect 11216 4327 11242 4383
rect 11136 4313 11162 4327
rect 11214 4313 11242 4327
rect 11136 4303 11242 4313
rect 11136 4247 11160 4303
rect 11216 4247 11242 4303
rect 11136 4237 11242 4247
rect 11136 4223 11162 4237
rect 11214 4223 11242 4237
rect 11136 4167 11160 4223
rect 11216 4167 11242 4223
rect 11136 4143 11162 4167
rect 11214 4143 11242 4167
rect 11136 4087 11160 4143
rect 11216 4087 11242 4143
rect 11136 4063 11162 4087
rect 11214 4063 11242 4087
rect 11136 4007 11160 4063
rect 11216 4007 11242 4063
rect 11136 3993 11162 4007
rect 11214 3993 11242 4007
rect 11136 3983 11242 3993
rect 11136 3927 11160 3983
rect 11216 3927 11242 3983
rect 11136 3917 11242 3927
rect 11136 3903 11162 3917
rect 11214 3903 11242 3917
rect 11136 3847 11160 3903
rect 11216 3847 11242 3903
rect 11136 3816 11242 3847
rect 14538 4381 14644 4412
rect 14538 4325 14566 4381
rect 14622 4325 14644 4381
rect 14538 4311 14568 4325
rect 14620 4311 14644 4325
rect 14538 4301 14644 4311
rect 14538 4245 14566 4301
rect 14622 4245 14644 4301
rect 14538 4235 14644 4245
rect 14538 4221 14568 4235
rect 14620 4221 14644 4235
rect 14538 4165 14566 4221
rect 14622 4165 14644 4221
rect 14538 4141 14568 4165
rect 14620 4141 14644 4165
rect 14538 4085 14566 4141
rect 14622 4085 14644 4141
rect 14538 4061 14568 4085
rect 14620 4061 14644 4085
rect 14538 4005 14566 4061
rect 14622 4005 14644 4061
rect 14538 3991 14568 4005
rect 14620 3991 14644 4005
rect 14538 3981 14644 3991
rect 14538 3925 14566 3981
rect 14622 3925 14644 3981
rect 14538 3915 14644 3925
rect 14538 3901 14568 3915
rect 14620 3901 14644 3915
rect 14538 3845 14566 3901
rect 14622 3845 14644 3901
rect 14538 3814 14644 3845
rect 2213 624 2343 1627
rect 2208 20 2344 624
rect 7942 610 8054 616
rect 4540 578 4652 610
rect 4540 522 4561 578
rect 4617 522 4652 578
rect 4540 498 4652 522
rect 4540 442 4561 498
rect 4617 442 4652 498
rect 4540 418 4652 442
rect 4540 362 4561 418
rect 4617 362 4652 418
rect 4540 338 4652 362
rect 4540 282 4561 338
rect 4617 282 4652 338
rect 4540 258 4652 282
rect 4540 202 4561 258
rect 4617 202 4652 258
rect 4540 178 4652 202
rect 4540 122 4561 178
rect 4617 122 4652 178
rect 4540 98 4652 122
rect 4540 42 4561 98
rect 4617 42 4652 98
rect 2213 7 2343 20
rect 4540 4 4652 42
rect 7940 574 8054 610
rect 8811 608 8941 1575
rect 15002 1014 15208 1042
rect 15002 992 15049 1014
rect 15165 992 15208 1014
rect 15002 856 15039 992
rect 15175 856 15208 992
rect 15002 834 15049 856
rect 15165 834 15208 856
rect 15002 812 15208 834
rect 7940 518 7963 574
rect 8019 518 8054 574
rect 7940 494 8054 518
rect 7940 438 7963 494
rect 8019 438 8054 494
rect 7940 414 8054 438
rect 7940 358 7963 414
rect 8019 358 8054 414
rect 7940 334 8054 358
rect 7940 278 7963 334
rect 8019 278 8054 334
rect 7940 254 8054 278
rect 7940 198 7963 254
rect 8019 198 8054 254
rect 7940 174 8054 198
rect 7940 118 7963 174
rect 8019 118 8054 174
rect 7940 94 8054 118
rect 7940 38 7963 94
rect 8019 38 8054 94
rect 7940 8 8054 38
rect 7942 6 8054 8
rect 8808 0 8946 608
rect 11134 578 11244 618
rect 11134 522 11161 578
rect 11217 522 11244 578
rect 11134 498 11244 522
rect 11134 442 11161 498
rect 11217 442 11244 498
rect 11134 418 11244 442
rect 11134 362 11161 418
rect 11217 362 11244 418
rect 11134 338 11244 362
rect 11134 282 11161 338
rect 11217 282 11244 338
rect 11134 258 11244 282
rect 11134 202 11161 258
rect 11217 202 11244 258
rect 11134 178 11244 202
rect 11134 122 11161 178
rect 11217 122 11244 178
rect 11134 98 11244 122
rect 11134 42 11161 98
rect 11217 42 11244 98
rect 11134 10 11244 42
rect 14540 584 14646 612
rect 14540 528 14570 584
rect 14626 528 14646 584
rect 14540 504 14646 528
rect 14540 448 14570 504
rect 14626 448 14646 504
rect 14540 424 14646 448
rect 14540 368 14570 424
rect 14626 368 14646 424
rect 14540 344 14646 368
rect 14540 288 14570 344
rect 14626 288 14646 344
rect 14540 264 14646 288
rect 14540 208 14570 264
rect 14626 208 14646 264
rect 14540 184 14646 208
rect 14540 128 14570 184
rect 14626 128 14646 184
rect 14540 104 14646 128
rect 14540 48 14570 104
rect 14626 48 14646 104
rect 14540 10 14646 48
rect 14546 8 14640 10
<< via2 >>
rect 1226 14461 1362 14757
rect 4569 12957 4625 12959
rect 4649 12957 4705 12959
rect 4729 12957 4785 12959
rect 4809 12957 4865 12959
rect 4889 12957 4945 12959
rect 4969 12957 5025 12959
rect 5049 12957 5105 12959
rect 5129 12957 5185 12959
rect 5209 12957 5265 12959
rect 4569 12905 4591 12957
rect 4591 12905 4603 12957
rect 4603 12905 4625 12957
rect 4649 12905 4655 12957
rect 4655 12905 4667 12957
rect 4667 12905 4705 12957
rect 4729 12905 4731 12957
rect 4731 12905 4783 12957
rect 4783 12905 4785 12957
rect 4809 12905 4847 12957
rect 4847 12905 4859 12957
rect 4859 12905 4865 12957
rect 4889 12905 4911 12957
rect 4911 12905 4923 12957
rect 4923 12905 4945 12957
rect 4969 12905 4975 12957
rect 4975 12905 4987 12957
rect 4987 12905 5025 12957
rect 5049 12905 5051 12957
rect 5051 12905 5103 12957
rect 5103 12905 5105 12957
rect 5129 12905 5167 12957
rect 5167 12905 5179 12957
rect 5179 12905 5185 12957
rect 5209 12905 5231 12957
rect 5231 12905 5243 12957
rect 5243 12905 5265 12957
rect 4569 12903 4625 12905
rect 4649 12903 4705 12905
rect 4729 12903 4785 12905
rect 4809 12903 4865 12905
rect 4889 12903 4945 12905
rect 4969 12903 5025 12905
rect 5049 12903 5105 12905
rect 5129 12903 5185 12905
rect 5209 12903 5265 12905
rect 11023 12960 11079 12962
rect 11103 12960 11159 12962
rect 11183 12960 11239 12962
rect 11263 12960 11319 12962
rect 11343 12960 11399 12962
rect 11423 12960 11479 12962
rect 11503 12960 11559 12962
rect 11583 12960 11639 12962
rect 11663 12960 11719 12962
rect 11743 12960 11799 12962
rect 11023 12908 11033 12960
rect 11033 12908 11079 12960
rect 11103 12908 11149 12960
rect 11149 12908 11159 12960
rect 11183 12908 11213 12960
rect 11213 12908 11225 12960
rect 11225 12908 11239 12960
rect 11263 12908 11277 12960
rect 11277 12908 11289 12960
rect 11289 12908 11319 12960
rect 11343 12908 11353 12960
rect 11353 12908 11399 12960
rect 11423 12908 11469 12960
rect 11469 12908 11479 12960
rect 11503 12908 11533 12960
rect 11533 12908 11545 12960
rect 11545 12908 11559 12960
rect 11583 12908 11597 12960
rect 11597 12908 11609 12960
rect 11609 12908 11639 12960
rect 11663 12908 11673 12960
rect 11673 12908 11719 12960
rect 11743 12908 11789 12960
rect 11789 12908 11799 12960
rect 11023 12906 11079 12908
rect 11103 12906 11159 12908
rect 11183 12906 11239 12908
rect 11263 12906 11319 12908
rect 11343 12906 11399 12908
rect 11423 12906 11479 12908
rect 11503 12906 11559 12908
rect 11583 12906 11639 12908
rect 11663 12906 11719 12908
rect 11743 12906 11799 12908
rect 4568 4375 4624 4393
rect 4568 4337 4570 4375
rect 4570 4337 4622 4375
rect 4622 4337 4624 4375
rect 4568 4311 4624 4313
rect 4568 4259 4570 4311
rect 4570 4259 4622 4311
rect 4622 4259 4624 4311
rect 4568 4257 4624 4259
rect 4568 4195 4570 4233
rect 4570 4195 4622 4233
rect 4622 4195 4624 4233
rect 4568 4183 4624 4195
rect 4568 4177 4570 4183
rect 4570 4177 4622 4183
rect 4622 4177 4624 4183
rect 4568 4131 4570 4153
rect 4570 4131 4622 4153
rect 4622 4131 4624 4153
rect 4568 4119 4624 4131
rect 4568 4097 4570 4119
rect 4570 4097 4622 4119
rect 4622 4097 4624 4119
rect 4568 4067 4570 4073
rect 4570 4067 4622 4073
rect 4622 4067 4624 4073
rect 4568 4055 4624 4067
rect 4568 4017 4570 4055
rect 4570 4017 4622 4055
rect 4622 4017 4624 4055
rect 4568 3991 4624 3993
rect 4568 3939 4570 3991
rect 4570 3939 4622 3991
rect 4622 3939 4624 3991
rect 4568 3937 4624 3939
rect 4568 3875 4570 3913
rect 4570 3875 4622 3913
rect 4622 3875 4624 3913
rect 4568 3857 4624 3875
rect 7964 4359 8020 4377
rect 7964 4321 7966 4359
rect 7966 4321 8018 4359
rect 8018 4321 8020 4359
rect 7964 4295 8020 4297
rect 7964 4243 7966 4295
rect 7966 4243 8018 4295
rect 8018 4243 8020 4295
rect 7964 4241 8020 4243
rect 7964 4179 7966 4217
rect 7966 4179 8018 4217
rect 8018 4179 8020 4217
rect 7964 4167 8020 4179
rect 7964 4161 7966 4167
rect 7966 4161 8018 4167
rect 8018 4161 8020 4167
rect 7964 4115 7966 4137
rect 7966 4115 8018 4137
rect 8018 4115 8020 4137
rect 7964 4103 8020 4115
rect 7964 4081 7966 4103
rect 7966 4081 8018 4103
rect 8018 4081 8020 4103
rect 7964 4051 7966 4057
rect 7966 4051 8018 4057
rect 8018 4051 8020 4057
rect 7964 4039 8020 4051
rect 7964 4001 7966 4039
rect 7966 4001 8018 4039
rect 8018 4001 8020 4039
rect 7964 3975 8020 3977
rect 7964 3923 7966 3975
rect 7966 3923 8018 3975
rect 8018 3923 8020 3975
rect 7964 3921 8020 3923
rect 7964 3859 7966 3897
rect 7966 3859 8018 3897
rect 8018 3859 8020 3897
rect 7964 3841 8020 3859
rect 11160 4365 11216 4383
rect 11160 4327 11162 4365
rect 11162 4327 11214 4365
rect 11214 4327 11216 4365
rect 11160 4301 11216 4303
rect 11160 4249 11162 4301
rect 11162 4249 11214 4301
rect 11214 4249 11216 4301
rect 11160 4247 11216 4249
rect 11160 4185 11162 4223
rect 11162 4185 11214 4223
rect 11214 4185 11216 4223
rect 11160 4173 11216 4185
rect 11160 4167 11162 4173
rect 11162 4167 11214 4173
rect 11214 4167 11216 4173
rect 11160 4121 11162 4143
rect 11162 4121 11214 4143
rect 11214 4121 11216 4143
rect 11160 4109 11216 4121
rect 11160 4087 11162 4109
rect 11162 4087 11214 4109
rect 11214 4087 11216 4109
rect 11160 4057 11162 4063
rect 11162 4057 11214 4063
rect 11214 4057 11216 4063
rect 11160 4045 11216 4057
rect 11160 4007 11162 4045
rect 11162 4007 11214 4045
rect 11214 4007 11216 4045
rect 11160 3981 11216 3983
rect 11160 3929 11162 3981
rect 11162 3929 11214 3981
rect 11214 3929 11216 3981
rect 11160 3927 11216 3929
rect 11160 3865 11162 3903
rect 11162 3865 11214 3903
rect 11214 3865 11216 3903
rect 11160 3847 11216 3865
rect 14566 4363 14622 4381
rect 14566 4325 14568 4363
rect 14568 4325 14620 4363
rect 14620 4325 14622 4363
rect 14566 4299 14622 4301
rect 14566 4247 14568 4299
rect 14568 4247 14620 4299
rect 14620 4247 14622 4299
rect 14566 4245 14622 4247
rect 14566 4183 14568 4221
rect 14568 4183 14620 4221
rect 14620 4183 14622 4221
rect 14566 4171 14622 4183
rect 14566 4165 14568 4171
rect 14568 4165 14620 4171
rect 14620 4165 14622 4171
rect 14566 4119 14568 4141
rect 14568 4119 14620 4141
rect 14620 4119 14622 4141
rect 14566 4107 14622 4119
rect 14566 4085 14568 4107
rect 14568 4085 14620 4107
rect 14620 4085 14622 4107
rect 14566 4055 14568 4061
rect 14568 4055 14620 4061
rect 14620 4055 14622 4061
rect 14566 4043 14622 4055
rect 14566 4005 14568 4043
rect 14568 4005 14620 4043
rect 14620 4005 14622 4043
rect 14566 3979 14622 3981
rect 14566 3927 14568 3979
rect 14568 3927 14620 3979
rect 14620 3927 14622 3979
rect 14566 3925 14622 3927
rect 14566 3863 14568 3901
rect 14568 3863 14620 3901
rect 14620 3863 14622 3901
rect 14566 3845 14622 3863
rect 4561 522 4617 578
rect 4561 442 4617 498
rect 4561 362 4617 418
rect 4561 282 4617 338
rect 4561 202 4617 258
rect 4561 122 4617 178
rect 4561 42 4617 98
rect 15039 856 15049 992
rect 15049 856 15165 992
rect 15165 856 15175 992
rect 7963 518 8019 574
rect 7963 438 8019 494
rect 7963 358 8019 414
rect 7963 278 8019 334
rect 7963 198 8019 254
rect 7963 118 8019 174
rect 7963 38 8019 94
rect 11161 522 11217 578
rect 11161 442 11217 498
rect 11161 362 11217 418
rect 11161 282 11217 338
rect 11161 202 11217 258
rect 11161 122 11217 178
rect 11161 42 11217 98
rect 14570 528 14626 584
rect 14570 448 14626 504
rect 14570 368 14626 424
rect 14570 288 14626 344
rect 14570 208 14626 264
rect 14570 128 14626 184
rect 14570 48 14626 104
<< metal3 >>
rect 930 25291 1980 25312
rect 930 25067 954 25291
rect 1098 25067 1980 25291
rect 930 25048 1980 25067
rect 14110 20655 16414 20696
rect 14110 20191 15315 20655
rect 15459 20191 16414 20655
rect 14110 20168 16414 20191
rect 15804 19578 16410 19582
rect 14010 19404 16410 19578
rect 1498 18274 2030 18496
rect 1204 14761 1404 14812
rect 0 14714 612 14722
rect 1204 14714 1222 14761
rect 0 14508 1222 14714
rect 1204 14457 1222 14508
rect 1366 14457 1404 14761
rect 1204 14408 1404 14457
rect 1498 13427 1720 18274
rect 1805 18196 2195 18213
rect 1805 17996 2404 18196
rect 1805 17991 2195 17996
rect 1805 13753 2027 17991
rect 15794 17660 16404 17662
rect 14372 17588 16408 17660
rect 13704 14120 16414 14146
rect 13704 13896 15037 14120
rect 15181 13896 16414 14120
rect 13704 13866 16414 13896
rect 1805 13531 11409 13753
rect 1498 13205 5009 13427
rect 4787 12986 5009 13205
rect 11187 12990 11409 13531
rect 4516 12959 5316 12986
rect 4516 12903 4569 12959
rect 4625 12903 4649 12959
rect 4705 12903 4729 12959
rect 4785 12903 4809 12959
rect 4865 12903 4889 12959
rect 4945 12903 4969 12959
rect 5025 12903 5049 12959
rect 5105 12903 5129 12959
rect 5185 12903 5209 12959
rect 5265 12903 5316 12959
rect 4516 12876 5316 12903
rect 10992 12962 11812 12990
rect 10992 12906 11023 12962
rect 11079 12906 11103 12962
rect 11159 12906 11183 12962
rect 11239 12906 11263 12962
rect 11319 12906 11343 12962
rect 11399 12906 11423 12962
rect 11479 12906 11503 12962
rect 11559 12906 11583 12962
rect 11639 12906 11663 12962
rect 11719 12906 11743 12962
rect 11799 12906 11812 12962
rect 10992 12880 11812 12906
rect 11187 12875 11409 12880
rect 0 8854 822 8860
rect 0 8828 11680 8854
rect 0 8684 962 8828
rect 1106 8684 11680 8828
rect 0 8660 11680 8684
rect 14 8654 11680 8660
rect 14 8650 5096 8654
rect 4542 4397 4648 4418
rect 4542 4333 4564 4397
rect 4628 4333 4648 4397
rect 4542 4317 4648 4333
rect 4542 4253 4564 4317
rect 4628 4253 4648 4317
rect 4542 4237 4648 4253
rect 4542 4173 4564 4237
rect 4628 4173 4648 4237
rect 4542 4157 4648 4173
rect 4542 4093 4564 4157
rect 4628 4093 4648 4157
rect 4542 4077 4648 4093
rect 4542 4013 4564 4077
rect 4628 4013 4648 4077
rect 4542 3997 4648 4013
rect 4542 3933 4564 3997
rect 4628 3933 4648 3997
rect 4542 3917 4648 3933
rect 4542 3853 4564 3917
rect 4628 3853 4648 3917
rect 4542 3820 4648 3853
rect 7940 4381 8046 4406
rect 7940 4317 7960 4381
rect 8024 4317 8046 4381
rect 7940 4301 8046 4317
rect 7940 4237 7960 4301
rect 8024 4237 8046 4301
rect 7940 4221 8046 4237
rect 7940 4157 7960 4221
rect 8024 4157 8046 4221
rect 7940 4141 8046 4157
rect 7940 4077 7960 4141
rect 8024 4077 8046 4141
rect 7940 4061 8046 4077
rect 7940 3997 7960 4061
rect 8024 3997 8046 4061
rect 7940 3981 8046 3997
rect 7940 3917 7960 3981
rect 8024 3917 8046 3981
rect 7940 3901 8046 3917
rect 7940 3837 7960 3901
rect 8024 3837 8046 3901
rect 7940 3808 8046 3837
rect 11136 4387 11242 4414
rect 11136 4323 11156 4387
rect 11220 4323 11242 4387
rect 11136 4307 11242 4323
rect 11136 4243 11156 4307
rect 11220 4243 11242 4307
rect 11136 4227 11242 4243
rect 11136 4163 11156 4227
rect 11220 4163 11242 4227
rect 11136 4147 11242 4163
rect 11136 4083 11156 4147
rect 11220 4083 11242 4147
rect 11136 4067 11242 4083
rect 11136 4003 11156 4067
rect 11220 4003 11242 4067
rect 11136 3987 11242 4003
rect 11136 3923 11156 3987
rect 11220 3923 11242 3987
rect 11136 3907 11242 3923
rect 11136 3843 11156 3907
rect 11220 3843 11242 3907
rect 11136 3816 11242 3843
rect 14538 4385 14644 4412
rect 14538 4321 14562 4385
rect 14626 4321 14644 4385
rect 14538 4305 14644 4321
rect 14538 4241 14562 4305
rect 14626 4241 14644 4305
rect 14538 4225 14644 4241
rect 14538 4161 14562 4225
rect 14626 4161 14644 4225
rect 14538 4145 14644 4161
rect 14538 4081 14562 4145
rect 14626 4081 14644 4145
rect 14538 4065 14644 4081
rect 14538 4001 14562 4065
rect 14626 4001 14644 4065
rect 14538 3985 14644 4001
rect 14538 3921 14562 3985
rect 14626 3921 14644 3985
rect 14538 3905 14644 3921
rect 14538 3841 14562 3905
rect 14626 3841 14644 3905
rect 14538 3814 14644 3841
rect 4926 2699 15506 2734
rect 4926 2635 15321 2699
rect 15385 2635 15401 2699
rect 15465 2635 15506 2699
rect 4926 2602 15506 2635
rect 15002 996 15208 1042
rect 15002 852 15035 996
rect 15179 852 15208 996
rect 15002 812 15208 852
rect 4534 582 4640 610
rect 4534 518 4557 582
rect 4621 518 4640 582
rect 4534 502 4640 518
rect 4534 438 4557 502
rect 4621 438 4640 502
rect 4534 422 4640 438
rect 4534 358 4557 422
rect 4621 358 4640 422
rect 4534 342 4640 358
rect 4534 278 4557 342
rect 4621 278 4640 342
rect 4534 262 4640 278
rect 4534 198 4557 262
rect 4621 198 4640 262
rect 4534 182 4640 198
rect 4534 118 4557 182
rect 4621 118 4640 182
rect 4534 102 4640 118
rect 4534 38 4557 102
rect 4621 38 4640 102
rect 4534 8 4640 38
rect 7940 578 8046 610
rect 7940 514 7959 578
rect 8023 514 8046 578
rect 7940 498 8046 514
rect 7940 434 7959 498
rect 8023 434 8046 498
rect 7940 418 8046 434
rect 7940 354 7959 418
rect 8023 354 8046 418
rect 7940 338 8046 354
rect 7940 274 7959 338
rect 8023 274 8046 338
rect 7940 258 8046 274
rect 7940 194 7959 258
rect 8023 194 8046 258
rect 7940 178 8046 194
rect 7940 114 7959 178
rect 8023 114 8046 178
rect 7940 98 8046 114
rect 7940 34 7959 98
rect 8023 34 8046 98
rect 7940 8 8046 34
rect 11134 582 11240 612
rect 11134 518 11157 582
rect 11221 518 11240 582
rect 11134 502 11240 518
rect 11134 438 11157 502
rect 11221 438 11240 502
rect 11134 422 11240 438
rect 11134 358 11157 422
rect 11221 358 11240 422
rect 11134 342 11240 358
rect 11134 278 11157 342
rect 11221 278 11240 342
rect 11134 262 11240 278
rect 11134 198 11157 262
rect 11221 198 11240 262
rect 11134 182 11240 198
rect 11134 118 11157 182
rect 11221 118 11240 182
rect 11134 102 11240 118
rect 11134 38 11157 102
rect 11221 38 11240 102
rect 11134 10 11240 38
rect 14546 588 14648 612
rect 14546 524 14566 588
rect 14630 524 14648 588
rect 14546 508 14648 524
rect 14546 444 14566 508
rect 14630 444 14648 508
rect 14546 428 14648 444
rect 14546 364 14566 428
rect 14630 364 14648 428
rect 14546 348 14648 364
rect 14546 284 14566 348
rect 14630 284 14648 348
rect 14546 268 14648 284
rect 14546 204 14566 268
rect 14630 204 14648 268
rect 14546 188 14648 204
rect 14546 124 14566 188
rect 14630 124 14648 188
rect 14546 108 14648 124
rect 14546 44 14566 108
rect 14630 44 14648 108
rect 14546 12 14648 44
<< via3 >>
rect 954 25067 1098 25291
rect 15315 20191 15459 20655
rect 1222 14757 1366 14761
rect 1222 14461 1226 14757
rect 1226 14461 1362 14757
rect 1362 14461 1366 14757
rect 1222 14457 1366 14461
rect 15037 13896 15181 14120
rect 962 8684 1106 8828
rect 4564 4393 4628 4397
rect 4564 4337 4568 4393
rect 4568 4337 4624 4393
rect 4624 4337 4628 4393
rect 4564 4333 4628 4337
rect 4564 4313 4628 4317
rect 4564 4257 4568 4313
rect 4568 4257 4624 4313
rect 4624 4257 4628 4313
rect 4564 4253 4628 4257
rect 4564 4233 4628 4237
rect 4564 4177 4568 4233
rect 4568 4177 4624 4233
rect 4624 4177 4628 4233
rect 4564 4173 4628 4177
rect 4564 4153 4628 4157
rect 4564 4097 4568 4153
rect 4568 4097 4624 4153
rect 4624 4097 4628 4153
rect 4564 4093 4628 4097
rect 4564 4073 4628 4077
rect 4564 4017 4568 4073
rect 4568 4017 4624 4073
rect 4624 4017 4628 4073
rect 4564 4013 4628 4017
rect 4564 3993 4628 3997
rect 4564 3937 4568 3993
rect 4568 3937 4624 3993
rect 4624 3937 4628 3993
rect 4564 3933 4628 3937
rect 4564 3913 4628 3917
rect 4564 3857 4568 3913
rect 4568 3857 4624 3913
rect 4624 3857 4628 3913
rect 4564 3853 4628 3857
rect 7960 4377 8024 4381
rect 7960 4321 7964 4377
rect 7964 4321 8020 4377
rect 8020 4321 8024 4377
rect 7960 4317 8024 4321
rect 7960 4297 8024 4301
rect 7960 4241 7964 4297
rect 7964 4241 8020 4297
rect 8020 4241 8024 4297
rect 7960 4237 8024 4241
rect 7960 4217 8024 4221
rect 7960 4161 7964 4217
rect 7964 4161 8020 4217
rect 8020 4161 8024 4217
rect 7960 4157 8024 4161
rect 7960 4137 8024 4141
rect 7960 4081 7964 4137
rect 7964 4081 8020 4137
rect 8020 4081 8024 4137
rect 7960 4077 8024 4081
rect 7960 4057 8024 4061
rect 7960 4001 7964 4057
rect 7964 4001 8020 4057
rect 8020 4001 8024 4057
rect 7960 3997 8024 4001
rect 7960 3977 8024 3981
rect 7960 3921 7964 3977
rect 7964 3921 8020 3977
rect 8020 3921 8024 3977
rect 7960 3917 8024 3921
rect 7960 3897 8024 3901
rect 7960 3841 7964 3897
rect 7964 3841 8020 3897
rect 8020 3841 8024 3897
rect 7960 3837 8024 3841
rect 11156 4383 11220 4387
rect 11156 4327 11160 4383
rect 11160 4327 11216 4383
rect 11216 4327 11220 4383
rect 11156 4323 11220 4327
rect 11156 4303 11220 4307
rect 11156 4247 11160 4303
rect 11160 4247 11216 4303
rect 11216 4247 11220 4303
rect 11156 4243 11220 4247
rect 11156 4223 11220 4227
rect 11156 4167 11160 4223
rect 11160 4167 11216 4223
rect 11216 4167 11220 4223
rect 11156 4163 11220 4167
rect 11156 4143 11220 4147
rect 11156 4087 11160 4143
rect 11160 4087 11216 4143
rect 11216 4087 11220 4143
rect 11156 4083 11220 4087
rect 11156 4063 11220 4067
rect 11156 4007 11160 4063
rect 11160 4007 11216 4063
rect 11216 4007 11220 4063
rect 11156 4003 11220 4007
rect 11156 3983 11220 3987
rect 11156 3927 11160 3983
rect 11160 3927 11216 3983
rect 11216 3927 11220 3983
rect 11156 3923 11220 3927
rect 11156 3903 11220 3907
rect 11156 3847 11160 3903
rect 11160 3847 11216 3903
rect 11216 3847 11220 3903
rect 11156 3843 11220 3847
rect 14562 4381 14626 4385
rect 14562 4325 14566 4381
rect 14566 4325 14622 4381
rect 14622 4325 14626 4381
rect 14562 4321 14626 4325
rect 14562 4301 14626 4305
rect 14562 4245 14566 4301
rect 14566 4245 14622 4301
rect 14622 4245 14626 4301
rect 14562 4241 14626 4245
rect 14562 4221 14626 4225
rect 14562 4165 14566 4221
rect 14566 4165 14622 4221
rect 14622 4165 14626 4221
rect 14562 4161 14626 4165
rect 14562 4141 14626 4145
rect 14562 4085 14566 4141
rect 14566 4085 14622 4141
rect 14622 4085 14626 4141
rect 14562 4081 14626 4085
rect 14562 4061 14626 4065
rect 14562 4005 14566 4061
rect 14566 4005 14622 4061
rect 14622 4005 14626 4061
rect 14562 4001 14626 4005
rect 14562 3981 14626 3985
rect 14562 3925 14566 3981
rect 14566 3925 14622 3981
rect 14622 3925 14626 3981
rect 14562 3921 14626 3925
rect 14562 3901 14626 3905
rect 14562 3845 14566 3901
rect 14566 3845 14622 3901
rect 14622 3845 14626 3901
rect 14562 3841 14626 3845
rect 15321 2635 15385 2699
rect 15401 2635 15465 2699
rect 15035 992 15179 996
rect 15035 856 15039 992
rect 15039 856 15175 992
rect 15175 856 15179 992
rect 15035 852 15179 856
rect 4557 578 4621 582
rect 4557 522 4561 578
rect 4561 522 4617 578
rect 4617 522 4621 578
rect 4557 518 4621 522
rect 4557 498 4621 502
rect 4557 442 4561 498
rect 4561 442 4617 498
rect 4617 442 4621 498
rect 4557 438 4621 442
rect 4557 418 4621 422
rect 4557 362 4561 418
rect 4561 362 4617 418
rect 4617 362 4621 418
rect 4557 358 4621 362
rect 4557 338 4621 342
rect 4557 282 4561 338
rect 4561 282 4617 338
rect 4617 282 4621 338
rect 4557 278 4621 282
rect 4557 258 4621 262
rect 4557 202 4561 258
rect 4561 202 4617 258
rect 4617 202 4621 258
rect 4557 198 4621 202
rect 4557 178 4621 182
rect 4557 122 4561 178
rect 4561 122 4617 178
rect 4617 122 4621 178
rect 4557 118 4621 122
rect 4557 98 4621 102
rect 4557 42 4561 98
rect 4561 42 4617 98
rect 4617 42 4621 98
rect 4557 38 4621 42
rect 7959 574 8023 578
rect 7959 518 7963 574
rect 7963 518 8019 574
rect 8019 518 8023 574
rect 7959 514 8023 518
rect 7959 494 8023 498
rect 7959 438 7963 494
rect 7963 438 8019 494
rect 8019 438 8023 494
rect 7959 434 8023 438
rect 7959 414 8023 418
rect 7959 358 7963 414
rect 7963 358 8019 414
rect 8019 358 8023 414
rect 7959 354 8023 358
rect 7959 334 8023 338
rect 7959 278 7963 334
rect 7963 278 8019 334
rect 8019 278 8023 334
rect 7959 274 8023 278
rect 7959 254 8023 258
rect 7959 198 7963 254
rect 7963 198 8019 254
rect 8019 198 8023 254
rect 7959 194 8023 198
rect 7959 174 8023 178
rect 7959 118 7963 174
rect 7963 118 8019 174
rect 8019 118 8023 174
rect 7959 114 8023 118
rect 7959 94 8023 98
rect 7959 38 7963 94
rect 7963 38 8019 94
rect 8019 38 8023 94
rect 7959 34 8023 38
rect 11157 578 11221 582
rect 11157 522 11161 578
rect 11161 522 11217 578
rect 11217 522 11221 578
rect 11157 518 11221 522
rect 11157 498 11221 502
rect 11157 442 11161 498
rect 11161 442 11217 498
rect 11217 442 11221 498
rect 11157 438 11221 442
rect 11157 418 11221 422
rect 11157 362 11161 418
rect 11161 362 11217 418
rect 11217 362 11221 418
rect 11157 358 11221 362
rect 11157 338 11221 342
rect 11157 282 11161 338
rect 11161 282 11217 338
rect 11217 282 11221 338
rect 11157 278 11221 282
rect 11157 258 11221 262
rect 11157 202 11161 258
rect 11161 202 11217 258
rect 11217 202 11221 258
rect 11157 198 11221 202
rect 11157 178 11221 182
rect 11157 122 11161 178
rect 11161 122 11217 178
rect 11217 122 11221 178
rect 11157 118 11221 122
rect 11157 98 11221 102
rect 11157 42 11161 98
rect 11161 42 11217 98
rect 11217 42 11221 98
rect 11157 38 11221 42
rect 14566 584 14630 588
rect 14566 528 14570 584
rect 14570 528 14626 584
rect 14626 528 14630 584
rect 14566 524 14630 528
rect 14566 504 14630 508
rect 14566 448 14570 504
rect 14570 448 14626 504
rect 14626 448 14630 504
rect 14566 444 14630 448
rect 14566 424 14630 428
rect 14566 368 14570 424
rect 14570 368 14626 424
rect 14626 368 14630 424
rect 14566 364 14630 368
rect 14566 344 14630 348
rect 14566 288 14570 344
rect 14570 288 14626 344
rect 14626 288 14630 344
rect 14566 284 14630 288
rect 14566 264 14630 268
rect 14566 208 14570 264
rect 14570 208 14626 264
rect 14626 208 14630 264
rect 14566 204 14630 208
rect 14566 184 14630 188
rect 14566 128 14570 184
rect 14570 128 14626 184
rect 14626 128 14630 184
rect 14566 124 14630 128
rect 14566 104 14630 108
rect 14566 48 14570 104
rect 14570 48 14626 104
rect 14626 48 14630 104
rect 14566 44 14630 48
<< metal4 >>
rect 932 25291 1132 26826
rect 932 25067 954 25291
rect 1098 25067 1132 25291
rect 932 8828 1132 25067
rect 932 8684 962 8828
rect 1106 8684 1132 8828
rect 932 1010 1132 8684
rect 1206 14761 1406 26828
rect 1206 14457 1222 14761
rect 1366 14457 1406 14761
rect 1206 1012 1406 14457
rect 15006 14120 15206 26624
rect 15006 13896 15037 14120
rect 15181 13896 15206 14120
rect 4542 4397 4648 4418
rect 4542 4333 4564 4397
rect 4628 4333 4648 4397
rect 4542 4317 4648 4333
rect 4542 4253 4564 4317
rect 4628 4253 4648 4317
rect 4542 4237 4648 4253
rect 4542 4173 4564 4237
rect 4628 4173 4648 4237
rect 4542 4157 4648 4173
rect 4542 4093 4564 4157
rect 4628 4093 4648 4157
rect 4542 4077 4648 4093
rect 4542 4013 4564 4077
rect 4628 4013 4648 4077
rect 4542 3997 4648 4013
rect 4542 3933 4564 3997
rect 4628 3933 4648 3997
rect 4542 3917 4648 3933
rect 4542 3853 4564 3917
rect 4628 3853 4648 3917
rect 4542 3820 4648 3853
rect 7940 4381 8046 4406
rect 7940 4317 7960 4381
rect 8024 4317 8046 4381
rect 7940 4301 8046 4317
rect 7940 4237 7960 4301
rect 8024 4237 8046 4301
rect 7940 4221 8046 4237
rect 7940 4157 7960 4221
rect 8024 4157 8046 4221
rect 7940 4141 8046 4157
rect 7940 4077 7960 4141
rect 8024 4077 8046 4141
rect 7940 4061 8046 4077
rect 7940 3997 7960 4061
rect 8024 3997 8046 4061
rect 7940 3981 8046 3997
rect 7940 3917 7960 3981
rect 8024 3917 8046 3981
rect 7940 3901 8046 3917
rect 7940 3837 7960 3901
rect 8024 3858 8046 3901
rect 11136 4387 11242 4414
rect 11136 4323 11156 4387
rect 11220 4323 11242 4387
rect 11136 4307 11242 4323
rect 11136 4243 11156 4307
rect 11220 4243 11242 4307
rect 11136 4227 11242 4243
rect 11136 4163 11156 4227
rect 11220 4163 11242 4227
rect 11136 4147 11242 4163
rect 11136 4083 11156 4147
rect 11220 4083 11242 4147
rect 11136 4067 11242 4083
rect 11136 4003 11156 4067
rect 11220 4003 11242 4067
rect 11136 3987 11242 4003
rect 11136 3923 11156 3987
rect 11220 3923 11242 3987
rect 11136 3907 11242 3923
rect 8024 3837 8048 3858
rect 4542 610 4644 3820
rect 7940 3782 8048 3837
rect 11136 3843 11156 3907
rect 11220 3843 11242 3907
rect 11136 3800 11242 3843
rect 14538 4385 14644 4412
rect 14538 4321 14562 4385
rect 14626 4321 14644 4385
rect 14538 4305 14644 4321
rect 14538 4241 14562 4305
rect 14626 4241 14644 4305
rect 14538 4225 14644 4241
rect 14538 4161 14562 4225
rect 14626 4161 14644 4225
rect 14538 4145 14644 4161
rect 14538 4081 14562 4145
rect 14626 4081 14644 4145
rect 14538 4065 14644 4081
rect 14538 4001 14562 4065
rect 14626 4001 14644 4065
rect 14538 3985 14644 4001
rect 14538 3921 14562 3985
rect 14626 3921 14644 3985
rect 14538 3905 14644 3921
rect 14538 3841 14562 3905
rect 14626 3841 14644 3905
rect 14538 3814 14644 3841
rect 7948 610 8048 3782
rect 11138 612 11238 3800
rect 4534 582 4644 610
rect 4534 518 4557 582
rect 4621 518 4644 582
rect 4534 502 4644 518
rect 4534 438 4557 502
rect 4621 438 4644 502
rect 4534 422 4644 438
rect 4534 358 4557 422
rect 4621 358 4644 422
rect 4534 342 4644 358
rect 4534 278 4557 342
rect 4621 278 4644 342
rect 4534 262 4644 278
rect 4534 198 4557 262
rect 4621 198 4644 262
rect 4534 182 4644 198
rect 4534 118 4557 182
rect 4621 118 4644 182
rect 4534 102 4644 118
rect 4534 38 4557 102
rect 4621 38 4644 102
rect 4534 9 4644 38
rect 7940 578 8048 610
rect 7940 514 7959 578
rect 8023 514 8048 578
rect 7940 498 8048 514
rect 7940 434 7959 498
rect 8023 434 8048 498
rect 7940 418 8048 434
rect 7940 354 7959 418
rect 8023 354 8048 418
rect 7940 338 8048 354
rect 7940 274 7959 338
rect 8023 274 8048 338
rect 7940 258 8048 274
rect 7940 194 7959 258
rect 8023 194 8048 258
rect 7940 178 8048 194
rect 7940 114 7959 178
rect 8023 114 8048 178
rect 7940 98 8048 114
rect 7940 34 7959 98
rect 8023 34 8048 98
rect 7940 12 8048 34
rect 11134 582 11240 612
rect 11134 518 11157 582
rect 11221 518 11240 582
rect 11134 502 11240 518
rect 11134 438 11157 502
rect 11221 438 11240 502
rect 11134 422 11240 438
rect 11134 358 11157 422
rect 11221 358 11240 422
rect 11134 342 11240 358
rect 11134 278 11157 342
rect 11221 278 11240 342
rect 11134 262 11240 278
rect 11134 198 11157 262
rect 11221 198 11240 262
rect 11134 182 11240 198
rect 11134 118 11157 182
rect 11221 118 11240 182
rect 11134 102 11240 118
rect 11134 38 11157 102
rect 11221 38 11240 102
rect 4534 8 4640 9
rect 7940 8 8046 12
rect 11134 10 11240 38
rect 14544 588 14644 3814
rect 15006 996 15206 13896
rect 15006 852 15035 996
rect 15179 852 15206 996
rect 15006 808 15206 852
rect 15298 20655 15498 26626
rect 15298 20191 15315 20655
rect 15459 20191 15498 20655
rect 15298 2699 15498 20191
rect 15298 2635 15321 2699
rect 15385 2635 15401 2699
rect 15465 2635 15498 2699
rect 15298 810 15498 2635
rect 14544 524 14566 588
rect 14630 524 14644 588
rect 14544 508 14644 524
rect 14544 444 14566 508
rect 14630 444 14644 508
rect 14544 428 14644 444
rect 14544 364 14566 428
rect 14630 364 14644 428
rect 14544 348 14644 364
rect 14544 284 14566 348
rect 14630 284 14644 348
rect 14544 268 14644 284
rect 14544 204 14566 268
rect 14630 204 14644 268
rect 14544 188 14644 204
rect 14544 124 14566 188
rect 14630 124 14644 188
rect 14544 108 14644 124
rect 14544 44 14566 108
rect 14630 44 14644 108
rect 14544 6 14644 44
use EF_AMUX2to1ISO  EF_AMUX2to1ISO_0
timestamp 1699022965
transform 1 0 1811 0 1 2004
box -3 -1196 6373 10978
use EF_AMUX2to1ISO  EF_AMUX2to1ISO_1
timestamp 1699022965
transform 1 0 8409 0 1 2008
box -3 -1196 6373 10978
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699022965
transform 1 0 2612 0 1 15273
box -804 -1465 11921 11144
<< labels >>
flabel metal2 s 2208 20 2344 624 0 FreeSans 1563 0 0 0 SELA
port 1 nsew
flabel metal2 s 8808 0 8946 608 0 FreeSans 1563 0 0 0 SELB
port 2 nsew
flabel metal2 s 4540 4 4652 610 0 FreeSans 1563 0 0 0 A1
port 3 nsew
flabel metal2 s 7942 6 8054 616 0 FreeSans 1563 0 0 0 A2
port 4 nsew
flabel metal2 s 11134 10 11244 618 0 FreeSans 1563 0 0 0 B1
port 5 nsew
flabel metal2 s 14540 10 14646 612 0 FreeSans 1563 0 0 0 B2
port 6 nsew
flabel metal3 s 0 8660 822 8860 0 FreeSans 1563 0 0 0 VDD
port 7 nsew
flabel metal3 s 0 14508 612 14722 0 FreeSans 1563 0 0 0 VSS
port 8 nsew
flabel metal3 s 15654 13874 16408 14144 0 FreeSans 1563 0 0 0 DVSS
port 9 nsew
flabel metal3 s 15792 20178 16408 20694 0 FreeSans 1563 0 0 0 DVDD
port 10 nsew
flabel metal3 s 15804 19406 16410 19582 0 FreeSans 1563 0 0 0 VO
port 11 nsew
flabel metal3 s 15794 17590 16404 17662 0 FreeSans 1563 0 0 0 EN
port 12 nsew
<< end >>
