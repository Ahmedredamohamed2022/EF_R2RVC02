magic
tech sky130A
magscale 1 2
timestamp 1689934956
<< checkpaint >>
rect -2527 -9292 15212 12428
<< metal1 >>
rect 518 -833 3398 -806
rect 518 -949 524 -833
rect 3392 -949 3398 -833
rect 518 -976 3398 -949
rect 7128 -828 10212 -806
rect 7128 -944 7140 -828
rect 10200 -944 10212 -828
rect 7128 -966 10212 -944
rect 2600 -4620 2796 -4086
rect 5978 -4602 6146 -4226
rect 9246 -4516 9438 -4022
rect 12586 -4546 12768 -4100
rect 2834 -7003 12762 -6799
rect 1216 -7670 1734 -7558
rect 8114 -7684 8640 -7570
rect 13236 -7834 13452 -7822
rect -26 -7863 13456 -7834
rect -26 -7979 13254 -7863
rect 13434 -7979 13456 -7863
rect -26 -7998 13456 -7979
rect 11192 -8002 13456 -7998
rect 13236 -8010 13452 -8002
<< via1 >>
rect 524 -949 3392 -833
rect 7140 -944 10200 -828
rect 13254 -7979 13434 -7863
<< metal2 >>
rect 12182 5615 13904 5678
rect 12182 5239 13731 5615
rect 13867 5239 13904 5615
rect 12182 5168 13904 5239
rect 11862 4416 11988 4494
rect -216 3590 238 3596
rect -216 3572 244 3590
rect -216 3356 -179 3572
rect 197 3362 244 3572
rect 197 3356 238 3362
rect -216 3324 238 3356
rect 178 3107 410 3176
rect 178 2658 212 3107
rect 182 2571 212 2658
rect 348 2658 410 3107
rect 348 2571 404 2658
rect 182 2486 404 2571
rect 12248 672 13438 710
rect 12248 136 13278 672
rect 13414 136 13438 672
rect 12248 70 13438 136
rect 488 -823 3470 -784
rect 488 -833 530 -823
rect 3386 -833 3470 -823
rect 488 -949 524 -833
rect 3392 -949 3470 -833
rect 488 -959 530 -949
rect 3386 -959 3470 -949
rect 488 -996 3470 -959
rect 7026 -818 10310 -780
rect 7026 -828 7162 -818
rect 10178 -828 10310 -818
rect 7026 -944 7140 -828
rect 10200 -944 10310 -828
rect 7026 -954 7162 -944
rect 10178 -954 10310 -944
rect 7026 -976 10310 -954
rect 13236 -7853 13452 -7822
rect 13236 -7863 13276 -7853
rect 13412 -7863 13452 -7853
rect 13236 -7979 13254 -7863
rect 13434 -7979 13452 -7863
rect 13236 -7989 13276 -7979
rect 13412 -7989 13452 -7979
rect 13236 -8010 13452 -7989
<< via2 >>
rect 13731 5239 13867 5615
rect -179 3356 197 3572
rect 212 2571 348 3107
rect 13278 136 13414 672
rect 530 -833 3386 -823
rect 530 -949 3386 -833
rect 530 -959 3386 -949
rect 7162 -828 10178 -818
rect 7162 -944 10178 -828
rect 7162 -954 10178 -944
rect 13276 -7863 13412 -7853
rect 13276 -7979 13412 -7863
rect 13276 -7989 13412 -7979
<< metal3 >>
rect -820 10866 -586 10872
rect -346 10866 4754 10876
rect -820 10804 4754 10866
rect -820 10180 -772 10804
rect -628 10799 4754 10804
rect -628 10575 3677 10799
rect 4701 10575 4754 10799
rect -628 10448 4754 10575
rect -628 10180 -586 10448
rect -820 10112 -586 10180
rect 13690 5619 13916 5674
rect 13690 5235 13727 5619
rect 13871 5235 13916 5619
rect 13690 5182 13916 5235
rect -216 3572 238 3596
rect -216 3356 -179 3572
rect 197 3356 238 3572
rect -216 3324 238 3356
rect -206 -370 6 3324
rect 182 3107 394 3176
rect 182 2571 212 3107
rect 348 2571 394 3107
rect 182 2 394 2571
rect 12248 676 13438 710
rect 12248 132 13274 676
rect 13418 132 13438 676
rect 12248 70 13438 132
rect 182 -210 8618 2
rect -206 -582 2008 -370
rect 1450 -784 1998 -582
rect 8212 -780 8618 -210
rect 488 -823 3470 -784
rect 488 -959 530 -823
rect 3386 -959 3470 -823
rect 488 -996 3470 -959
rect 7026 -818 10310 -780
rect 7026 -954 7162 -818
rect 10178 -954 10310 -818
rect 7026 -976 10310 -954
rect -1266 -2687 -1042 -2628
rect -1266 -2915 -1235 -2687
rect -1267 -3141 -1235 -2915
rect -1266 -3471 -1235 -3141
rect -1091 -2915 -1042 -2687
rect -1091 -3141 10085 -2915
rect -1091 -3471 -1042 -3141
rect -1266 -3536 -1042 -3471
rect 13672 -6216 13952 -6138
rect 13672 -6246 13728 -6216
rect 3211 -6404 13728 -6246
rect 9726 -6426 13728 -6404
rect 13672 -6520 13728 -6426
rect 13872 -6520 13952 -6216
rect 13672 -6614 13952 -6520
rect 13236 -7849 13452 -7822
rect 13236 -7993 13272 -7849
rect 13416 -7993 13452 -7849
rect 13236 -8010 13452 -7993
<< via3 >>
rect -772 10180 -628 10804
rect 3677 10575 4701 10799
rect 13727 5615 13871 5619
rect 13727 5239 13731 5615
rect 13731 5239 13867 5615
rect 13867 5239 13871 5615
rect 13727 5235 13871 5239
rect 13274 672 13418 676
rect 13274 136 13278 672
rect 13278 136 13414 672
rect 13414 136 13418 672
rect 13274 132 13418 136
rect -1235 -3471 -1091 -2687
rect 13728 -6520 13872 -6216
rect 13272 -7853 13416 -7849
rect 13272 -7989 13276 -7853
rect 13276 -7989 13412 -7853
rect 13412 -7989 13416 -7853
rect 13272 -7993 13416 -7989
<< metal4 >>
rect -920 11162 2472 11168
rect -1262 10944 2472 11162
rect -1262 -2687 -1038 10944
rect 1216 10932 2472 10944
rect -1262 -3471 -1235 -2687
rect -1091 -3471 -1038 -2687
rect -1262 -8030 -1038 -3471
rect -814 10804 -590 10866
rect 1216 10842 2478 10932
rect -814 10180 -772 10804
rect -628 10180 -590 10804
rect -814 -8006 -590 10180
rect 1284 9978 2478 10842
rect 3570 10799 4764 10866
rect 3570 10575 3677 10799
rect 4701 10575 4764 10799
rect 3570 9912 4764 10575
rect 13246 676 13446 10132
rect 13246 132 13274 676
rect 13418 132 13446 676
rect 13246 -7822 13446 132
rect 13700 5619 13900 10132
rect 13700 5235 13727 5619
rect 13871 5235 13900 5619
rect 13700 -6138 13900 5235
rect 13672 -6216 13952 -6138
rect 13672 -6520 13728 -6216
rect 13872 -6520 13952 -6216
rect 13672 -6614 13952 -6520
rect 13236 -7849 13452 -7822
rect 13236 -7993 13272 -7849
rect 13416 -7993 13452 -7849
rect 13700 -7974 13900 -6614
rect 13236 -8010 13452 -7993
rect 13246 -8012 13446 -8010
use EF_AMUX21m  EF_AMUX21m_1
timestamp 1689843535
transform 1 0 -3364 0 1 -7208
box 2505 -820 10000 6424
use EF_AMUX21m  EF_AMUX21m_2
timestamp 1689843535
transform 1 0 3262 0 1 -7212
box 2505 -820 10000 6424
use comparator_top  comparator_top_0
timestamp 1689839963
transform 1 0 800 0 1 265
box -802 -265 11765 10234
<< labels >>
flabel metal1 s 2682 -4524 2770 -4372 0 FreeSans 200 0 0 0 a1
port 1 nsew
flabel metal1 s 2652 -4450 2712 -4352 0 FreeSans 1000 0 0 0 a1
port 1 nsew
flabel metal1 s 6022 -4482 6090 -4352 0 FreeSans 1000 0 0 0 a2
port 2 nsew
flabel metal1 s 9268 -4352 9326 -4238 0 FreeSans 1000 0 0 0 b1
port 3 nsew
flabel metal1 s 12654 -4386 12680 -4316 0 FreeSans 1000 0 0 0 b2
port 4 nsew
flabel metal4 s 13298 -7084 13358 -6862 0 FreeSans 1000 0 0 0 dvss
port 5 nsew
flabel metal4 s -1166 11022 -1070 11100 0 FreeSans 1000 0 0 0 vdd3p3
port 6 nsew
flabel metal3 s -244 10608 -148 10686 0 FreeSans 1000 0 0 0 vss
port 7 nsew
flabel metal2 s 11896 4438 11940 4464 0 FreeSans 1000 0 0 0 vo
port 8 nsew
flabel metal1 s 1388 -7634 1464 -7584 0 FreeSans 1000 0 0 0 sela
port 9 nsew
flabel metal1 s 8280 -7624 8392 -7584 0 FreeSans 1000 0 0 0 selb
port 10 nsew
flabel metal4 s 13732 -7434 13790 -7284 0 FreeSans 1000 0 0 0 vdd1p8
port 11 nsew
<< end >>
