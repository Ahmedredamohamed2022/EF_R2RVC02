.subckt EF_R2RVC02 VSS A1 A2 SELB VO B2 B1 SELA VDD DVSS DVDD EN
*.PININFO DVDD:I VSS:I SELA:I SELB:I VDD:I DVSS:I A1:I A2:I B1:I B2:I VO:I EN:I
x1 VO EN DVDD VDD vinp VSS DVSS vinm EF_R2RVCE1x
x4 VDD DVDD DVSS vinp A1 A2 SELA EF_AMUX2to1ISOp
x5 VDD DVDD DVSS vinm B1 B2 SELB EF_AMUX2to1ISOp
.ends

* expanding   symbol:  Project/AR_SAR_ADC/comparator_top_up/spice/xschem/EF_R2RVCE1x.sym # of pins=8
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_up/spice/xschem/EF_R2RVCE1x.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_up/spice/xschem/EF_R2RVCE1x.sch
.subckt EF_R2RVCE1x VOUT EN DVDD VDD VINP VSS DVSS VINM
*.PININFO VOUT:O VINP:I VINM:I VDD:B VSS:B DVSS:B DVDD:B EN:I
x4 net1 DVDD DVSS DVSS VDD VDD VOUT sky130_fd_sc_hvl__lsbufhv2lv_1
x1 VDD VSS up down VBP VBN BIASE
x3 VDD VBP VBN VSS VINP net1 VINM AVOUT COMPARATOR
XM4 down ENB_C up VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM27 AVOUT ENB_C VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
x2 EN DVDD DVSS DVSS VDD VDD net2 sky130_fd_sc_hvl__lsbuflv2hv_1
x11 net2 DVSS DVSS VDD VDD ENB_C sky130_fd_sc_hvl__inv_4
.ends


* expanding   symbol:  Project/AR_SAR_ADC/comparator_top_02ch _up/spice/xschem/EF_AMUX2to1ISOp.sym #
*+ of pins=7
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_02ch
*+ _up/spice/xschem/EF_AMUX2to1ISOp.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_02ch
*+ _up/spice/xschem/EF_AMUX2to1ISOp.sch
.subckt EF_AMUX2to1ISOp VDD DVDD DVSS VO VIN1 VIN2 SEL
*.PININFO DVDD:I VDD:I DVSS:I SEL:I VO:I VIN1:I VIN2:I
x1 VO VDD DVDD DVSS SEL VIN1 single_ls_2tg_sw
x4 VO VDD DVDD DVSS SELB VIN2 single_ls_2tg_sw
x11 SEL DVSS DVSS DVDD DVDD SELB sky130_fd_sc_hvl__inv_4
.ends


* expanding   symbol:  Project/AR_SAR_ADC/comparator_top_up/spice/xschem/BIASE.sym # of pins=6
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_up/spice/xschem/BIASE.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_up/spice/xschem/BIASE.sch
.subckt BIASE VDD VSS up down VBP VBN
*.PININFO VBP:O VBN:O VDD:B VSS:B up:B down:B
XR1 up VDD VSS sky130_fd_pr__res_high_po W=1.41 L=141 mult=1 m=1
XM3 net1 down VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM4 VBN net1 down VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=20 nf=1 m=1
XM5 VBN VBN down VDD sky130_fd_pr__pfet_g5v0d10v5 L=15 W=1 nf=1 m=1
XM7 VBP VBP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM1 VBN VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM2 net1 VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM6 VBP VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM8 VBN VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM9 net1 VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM10 VBP VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
.ends


* expanding   symbol:  Project/AR_SAR_ADC/comparator_top_up/spice/xschem/COMPARATOR.sym # of pins=8
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_up/spice/xschem/COMPARATOR.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_up/spice/xschem/COMPARATOR.sch
.subckt COMPARATOR VDD VBP VBN VSS VINP VOUT VINM VOUTANALOG
*.PININFO VINP:I VINM:I VBN:I VBP:I VDD:B VSS:B VOUT:O VOUTANALOG:O
XM1 net3 VINM net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=4
XM2 net2 VINP net1 VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=4
XM3 net1 VBN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM4 net4 net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM5 VOUTANALOG net4 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM6 net3 net3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM7 net2 net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM8 net4 net3 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM9 VOUTANALOG net2 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM10 net6 VINM net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=4
XM11 net7 VINP net5 VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=4
XM12 net5 VBP VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM13 net8 net8 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM14 VOUTANALOG net8 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM15 net6 net6 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM16 net7 net7 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM17 net8 net6 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM18 VOUTANALOG net7 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM19 voinv1 VOUTANALOG VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 m=1
XM20 voinv1 VOUTANALOG VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM21 VOUT voinv1 VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=10 nf=1 m=1
XM22 VOUT voinv1 VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=1
XM23 net1 VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM24 net5 VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=2
XM25 VSS VSS VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=2 W=5 nf=1 m=8
XM26 VDD VDD VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=2 W=5 nf=1 m=8
.ends


* expanding   symbol:  Project/AR_SAR_ADC/comparator_top_02ch _up/spice/xschem/single_ls_2tg_sw.sym
*+ # of pins=6
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_02ch
*+ _up/spice/xschem/single_ls_2tg_sw.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_02ch
*+ _up/spice/xschem/single_ls_2tg_sw.sch
.subckt single_ls_2tg_sw VOUT VDD DVDD DVSS DINL VIN
*.PININFO DVDD:I VDD:I DVSS:I DINL:I VOUT:O VIN:I
x2 DOHB DOH VDD DVDD DVSS DINL single_lsp
x1 DOHB DVSS VOUT1 VIN VDD single_tgp
XM2 VOUT1 DOH DVSS DVSS sky130_fd_pr__nfet_g5v0d10v5 L=8 W=0.5 nf=1 m=1
x3 DOHB DVSS VOUT VOUT1 VDD single_tgp
.ends


* expanding   symbol:  Project/AR_SAR_ADC/analog_mux_up/spice/xschem/single_lsp.sym # of pins=6
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/analog_mux_up/spice/xschem/single_lsp.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/analog_mux_up/spice/xschem/single_lsp.sch
.subckt single_lsp DOHB DOH VDD DVDD DVSS DINL
*.PININFO DVDD:I VDD:I DVSS:I DINL:I DOH:O DOHB:O
x5 DINL DVDD DVSS DVSS VDD VDD DOH sky130_fd_sc_hvl__lsbuflv2hv_1
x11 DOH DVSS DVSS VDD VDD DOHB sky130_fd_sc_hvl__inv_2
.ends


* expanding   symbol:  Project/AR_SAR_ADC/analog_mux_up/spice/xschem/single_tgp.sym # of pins=5
** sym_path: /home/ahmedreda/Project/AR_SAR_ADC/analog_mux_up/spice/xschem/single_tgp.sym
** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/analog_mux_up/spice/xschem/single_tgp.sch
.subckt single_tgp SEL VSS VOUT VIN VDD
*.PININFO VIN:I VOUT:O VSS:I VDD:I SEL:I
XM1 VIN SELN VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=4 nf=2 m=1
XM2 VIN SELP VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=2 m=1
XM3 VOUT SELP VOUT VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM4 VOUT SELN VOUT VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM5 VIN SELP VIN VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM6 VIN SELN VIN VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=1 nf=1 m=1
XM7 SELN SEL VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM8 SELN SEL VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM9 SELP SELN VDD VDD sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
XM10 SELP SELN VSS VSS sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=2 nf=1 m=1
D1 VSS SEL sky130_fd_pr__diode_pw2nd_05v5
.ends

.end
