magic
tech sky130A
magscale 1 2
timestamp 1694943448
<< metal1 >>
rect 1896 2794 2621 2986
rect 1896 14 2088 2794
rect 4120 2183 4442 2190
rect 4120 2003 4127 2183
rect 4435 2003 4442 2183
rect 4120 1996 4442 2003
rect 4604 1732 4796 4114
rect 4418 1540 4796 1732
rect 2156 1148 2603 1340
rect 2156 4 2348 1148
rect 3846 420 4488 422
rect 3846 240 3853 420
rect 4481 240 4488 420
rect 3846 238 4488 240
<< via1 >>
rect 4127 2003 4435 2183
rect 3853 240 4481 420
<< metal2 >>
rect 4108 2212 4466 2214
rect 4108 2183 4886 2212
rect 4108 2003 4127 2183
rect 4435 2003 4886 2183
rect 4108 1984 4886 2003
rect 4108 1980 4466 1984
rect 3790 438 4886 450
rect 3788 420 4886 438
rect 3788 240 3853 420
rect 4481 240 4886 420
rect 3788 218 4886 240
rect 3788 214 4602 218
use tg4dm  tg4dm_1
timestamp 1694943448
transform 1 0 2091 0 1 2311
box 301 -2311 2543 1830
<< labels >>
flabel metal2 s 4744 238 4812 390 0 FreeSans 355 0 0 0 vss3p3
port 1 nsew
flabel metal2 s 4836 2020 4874 2114 0 FreeSans 355 0 0 0 vdd3p3
port 2 nsew
flabel metal1 s 1926 68 1964 162 0 FreeSans 355 0 0 0 s0
port 3 nsew
flabel metal1 s 2210 58 2248 152 0 FreeSans 355 0 0 0 in0
port 4 nsew
flabel metal1 s 4698 3594 4722 3660 0 FreeSans 30 0 0 0 vo
port 5 nsew
<< end >>
