** NOTE: ngspice DOES NOT handle environment variables used in the test benches. the Makefile handles that for you, if you wish to use your own command make sure you manually update the spice files

V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
C1 VOUT VSS 1p m=1
V5 DVDD VSS 1.8
.save i(v5)



x1 VSS VO SELB A2 B2 B1 SELA DVSS A1 DVDD VDD EF_R2RVC02



V10 DVSS GND 0
.save i(v10)
V8 SELB VSS 1.8
.save i(v8)
V9 SELA VSS 1.8
.save i(v9)
V3 A1 VSS 1.65
.save i(v3)
V4 B1 VSS 1.65
.save i(v4)
V6 B2 VSS 1.65
.save i(v6)
V7 A2 VSS 1.65
.save i(v7)
**** begin user architecture code


.include /home/ahmedreda/PDK/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /home/ahmedreda/PDK/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl__lsbuflv2hv_1.spice


.lib $PDK_ROOT/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include ../../spice/$SIM/EF_R2RVC02.spice



.option wnflag=1
.option TEMP=27
.option TNOM=27
.option wnflag=1
.control
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
save all
run
op
dc V3 0 3.3 0.01
let icom=abs(v2#branch)
let ibuf=abs(v5#branch)
let itot=icom+ibuf
let voutdigital=vout
plot vinp voutdigital vinm
meas dc offset1 WHEN vinp=1.65
meas dc offset2 FIND vout AT=1.65

plot itot
meas dc itot_1.65 FIND itot AT=1.65
meas dc itot_0 FIND itot AT=0.01
meas dc itot_3.3 FIND itot AT=3.29
meas dc offset_actual WHEN voutdigital=0.9

print (offset_actual-1.65)*1000

plot A1 B2 vout
.endc






.GLOBAL GND
.end
