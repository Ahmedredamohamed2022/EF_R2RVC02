magic
tech sky130A
magscale 1 2
timestamp 1692726716
<< pwell >>
rect -268 -448 268 448
<< mvnmos >>
rect -50 -200 50 200
<< mvndiff >>
rect -108 187 -50 200
rect -108 153 -96 187
rect -62 153 -50 187
rect -108 119 -50 153
rect -108 85 -96 119
rect -62 85 -50 119
rect -108 51 -50 85
rect -108 17 -96 51
rect -62 17 -50 51
rect -108 -17 -50 17
rect -108 -51 -96 -17
rect -62 -51 -50 -17
rect -108 -85 -50 -51
rect -108 -119 -96 -85
rect -62 -119 -50 -85
rect -108 -153 -50 -119
rect -108 -187 -96 -153
rect -62 -187 -50 -153
rect -108 -200 -50 -187
rect 50 187 108 200
rect 50 153 62 187
rect 96 153 108 187
rect 50 119 108 153
rect 50 85 62 119
rect 96 85 108 119
rect 50 51 108 85
rect 50 17 62 51
rect 96 17 108 51
rect 50 -17 108 17
rect 50 -51 62 -17
rect 96 -51 108 -17
rect 50 -85 108 -51
rect 50 -119 62 -85
rect 96 -119 108 -85
rect 50 -153 108 -119
rect 50 -187 62 -153
rect 96 -187 108 -153
rect 50 -200 108 -187
<< mvndiffc >>
rect -96 153 -62 187
rect -96 85 -62 119
rect -96 17 -62 51
rect -96 -51 -62 -17
rect -96 -119 -62 -85
rect -96 -187 -62 -153
rect 62 153 96 187
rect 62 85 96 119
rect 62 17 96 51
rect 62 -51 96 -17
rect 62 -119 96 -85
rect 62 -187 96 -153
<< mvpsubdiff >>
rect -242 410 242 422
rect -242 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 242 410
rect -242 364 242 376
rect -242 289 -184 364
rect -242 255 -230 289
rect -196 255 -184 289
rect 184 289 242 364
rect -242 221 -184 255
rect -242 187 -230 221
rect -196 187 -184 221
rect 184 255 196 289
rect 230 255 242 289
rect 184 221 242 255
rect -242 153 -184 187
rect -242 119 -230 153
rect -196 119 -184 153
rect -242 85 -184 119
rect -242 51 -230 85
rect -196 51 -184 85
rect -242 17 -184 51
rect -242 -17 -230 17
rect -196 -17 -184 17
rect -242 -51 -184 -17
rect -242 -85 -230 -51
rect -196 -85 -184 -51
rect -242 -119 -184 -85
rect -242 -153 -230 -119
rect -196 -153 -184 -119
rect -242 -187 -184 -153
rect -242 -221 -230 -187
rect -196 -221 -184 -187
rect 184 187 196 221
rect 230 187 242 221
rect 184 153 242 187
rect 184 119 196 153
rect 230 119 242 153
rect 184 85 242 119
rect 184 51 196 85
rect 230 51 242 85
rect 184 17 242 51
rect 184 -17 196 17
rect 230 -17 242 17
rect 184 -51 242 -17
rect 184 -85 196 -51
rect 230 -85 242 -51
rect 184 -119 242 -85
rect 184 -153 196 -119
rect 230 -153 242 -119
rect 184 -187 242 -153
rect -242 -255 -184 -221
rect -242 -289 -230 -255
rect -196 -289 -184 -255
rect 184 -221 196 -187
rect 230 -221 242 -187
rect 184 -255 242 -221
rect -242 -364 -184 -289
rect 184 -289 196 -255
rect 230 -289 242 -255
rect 184 -364 242 -289
rect -242 -376 242 -364
rect -242 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 242 -376
rect -242 -422 242 -410
<< mvpsubdiffcont >>
rect -119 376 -85 410
rect -51 376 -17 410
rect 17 376 51 410
rect 85 376 119 410
rect -230 255 -196 289
rect -230 187 -196 221
rect 196 255 230 289
rect -230 119 -196 153
rect -230 51 -196 85
rect -230 -17 -196 17
rect -230 -85 -196 -51
rect -230 -153 -196 -119
rect -230 -221 -196 -187
rect 196 187 230 221
rect 196 119 230 153
rect 196 51 230 85
rect 196 -17 230 17
rect 196 -85 230 -51
rect 196 -153 230 -119
rect -230 -289 -196 -255
rect 196 -221 230 -187
rect 196 -289 230 -255
rect -119 -410 -85 -376
rect -51 -410 -17 -376
rect 17 -410 51 -376
rect 85 -410 119 -376
<< poly >>
rect -50 272 50 288
rect -50 238 -17 272
rect 17 238 50 272
rect -50 200 50 238
rect -50 -238 50 -200
rect -50 -272 -17 -238
rect 17 -272 50 -238
rect -50 -288 50 -272
<< polycont >>
rect -17 238 17 272
rect -17 -272 17 -238
<< locali >>
rect -230 376 -119 410
rect -85 376 -51 410
rect -17 376 17 410
rect 51 376 85 410
rect 119 376 230 410
rect -230 289 -196 376
rect 196 289 230 376
rect -230 221 -196 255
rect -50 238 -17 272
rect 17 238 50 272
rect 196 221 230 255
rect -230 153 -196 187
rect -230 85 -196 119
rect -230 17 -196 51
rect -230 -51 -196 -17
rect -230 -119 -196 -85
rect -230 -187 -196 -153
rect -96 187 -62 204
rect -96 119 -62 127
rect -96 51 -62 55
rect -96 -55 -62 -51
rect -96 -127 -62 -119
rect -96 -204 -62 -187
rect 62 187 96 204
rect 62 119 96 127
rect 62 51 96 55
rect 62 -55 96 -51
rect 62 -127 96 -119
rect 62 -204 96 -187
rect 196 153 230 187
rect 196 85 230 119
rect 196 17 230 51
rect 196 -51 230 -17
rect 196 -119 230 -85
rect 196 -187 230 -153
rect -230 -255 -196 -221
rect -50 -272 -17 -238
rect 17 -272 50 -238
rect 196 -255 230 -221
rect -230 -376 -196 -289
rect 196 -376 230 -289
rect -230 -410 -119 -376
rect -85 -410 -51 -376
rect -17 -410 17 -376
rect 51 -410 85 -376
rect 119 -410 230 -376
<< viali >>
rect -17 238 17 272
rect -96 153 -62 161
rect -96 127 -62 153
rect -96 85 -62 89
rect -96 55 -62 85
rect -96 -17 -62 17
rect -96 -85 -62 -55
rect -96 -89 -62 -85
rect -96 -153 -62 -127
rect -96 -161 -62 -153
rect 62 153 96 161
rect 62 127 96 153
rect 62 85 96 89
rect 62 55 96 85
rect 62 -17 96 17
rect 62 -85 96 -55
rect 62 -89 96 -85
rect 62 -153 96 -127
rect 62 -161 96 -153
rect -17 -272 17 -238
<< metal1 >>
rect -46 272 46 278
rect -46 238 -17 272
rect 17 238 46 272
rect -46 232 46 238
rect -102 161 -56 200
rect -102 127 -96 161
rect -62 127 -56 161
rect -102 89 -56 127
rect -102 55 -96 89
rect -62 55 -56 89
rect -102 17 -56 55
rect -102 -17 -96 17
rect -62 -17 -56 17
rect -102 -55 -56 -17
rect -102 -89 -96 -55
rect -62 -89 -56 -55
rect -102 -127 -56 -89
rect -102 -161 -96 -127
rect -62 -161 -56 -127
rect -102 -200 -56 -161
rect 56 161 102 200
rect 56 127 62 161
rect 96 127 102 161
rect 56 89 102 127
rect 56 55 62 89
rect 96 55 102 89
rect 56 17 102 55
rect 56 -17 62 17
rect 96 -17 102 17
rect 56 -55 102 -17
rect 56 -89 62 -55
rect 96 -89 102 -55
rect 56 -127 102 -89
rect 56 -161 62 -127
rect 96 -161 102 -127
rect 56 -200 102 -161
rect -46 -238 46 -232
rect -46 -272 -17 -238
rect 17 -272 46 -238
rect -46 -278 46 -272
<< properties >>
string FIXED_BBOX -212 -392 212 392
<< end >>
