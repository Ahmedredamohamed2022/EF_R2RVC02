* NGSPICE file created from EF_R2RVC02.ext - technology: sky130A

.subckt EF_R2RVC02 VSS VO SELB A2 B2 B1 SELA DVSS A1 DVDD VDD
X0 a_1821_8526.t3 comparator_top_0.comparator_0.VBN.t3 comparator_top_0.comparator_0.VBN.t4 VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=15
X1 VSS.t66 VSS.t65 VSS.t66 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X2 VSS.t64 VSS.t62 VSS.t63 VSS.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X3 a_2551_4880.t5 a_2151_4783.t8 VDD.t137 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X4 comparator_top_0.comparator_0.VOUT a_8881_1782.t2 VDD.t47 VDD.t46 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=2
X5 a_570_n5724# a_470_n5812# DVSS.t139 DVSS.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X6 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb B1.t7 DVSS.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X7 DVSS.t77 a_570_n5724# a_1777_n6060# DVSS.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X8 VDD.t55 a_1821_8526.t6 a_2221_8623.t3 VDD.t54 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X9 a_2093_3714.t1 comparator_top_0.comparator_0.VBP VDD.t9 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X10 VDD.t29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VDD.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
D0 DVSS.t8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X11 a_6351_6657# a_10811_7187# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X12 VSS.t25 a_2151_594.t8 a_2551_620.t1 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X13 a_5299_3714.t7 comparator_top_0.VINP a_2093_3714.t10 VDD.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X14 DVSS.t38 a_3916_n5703# a_5123_n6039# DVSS.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X15 VSS.t19 comparator_top_0.comparator_0.VBN.t9 a_2093_1782.t1 VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X16 a_10542_n5707# a_10442_n5795# DVSS.t127 DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X17 a_2093_3714.t7 VDD.t125 VDD.t127 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X18 DVSS.t36 a_10965_3602# a_10975_4108# DVSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X19 a_7889_n6842# a_7464_n6798# DVSS.t103 DVSS.t102 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X20 VDD.t124 VDD.t123 VDD.t124 VDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X21 DVSS.t5 a_10975_4108# VO.t0 DVSS.t4 sky130_fd_pr__nfet_01v8 ad=0.196 pd=2.01 as=0.196 ps=2.01 w=0.74 l=0.15
X22 DVSS.t42 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp DVSS.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X23 VDD.t3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD.t62 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X25 EF_AMUX21m_1.invm_0.Y SELA.t0 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X26 DVSS.t101 a_7464_n6798# a_7889_n6842# DVSS.t100 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X27 DVDD.t16 EF_AMUX21m_2.invm_0.Y a_10442_n5795# DVDD.t15 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X28 a_7464_n6798# a_7096_n5816# DVDD.t12 DVDD.t11 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_5123_n6039# DVSS.t89 DVSS.t88 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X30 a_4184_n6773# a_3816_n5791# DVDD.t22 DVDD.t21 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X31 VSS.t61 VSS.t59 comparator_top_0.comparator_0.VBN.t2 VSS.t60 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X32 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINM DVSS.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=0.5
X33 a_2093_3714.t9 comparator_top_0.VINP a_5299_3714.t6 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X34 VSS.t31 a_5299_620.t8 a_8881_1782.t0 VSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
D1 DVSS.t13 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X35 DVSS.t65 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp DVSS.t64 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X36 a_4609_n6817# a_4184_n6773# DVSS.t190 DVSS.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X37 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_1777_n6060# VDD.t97 VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X38 A1.t7 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINP VDD.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X39 a_838_n6794# a_470_n5812# DVDD.t26 DVDD.t25 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X40 DVSS.t59 comparator_top_0.comparator_0.VOUT a_11031_3400# DVSS.t58 sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X41 VSS.t58 VSS.t57 VSS.t58 VSS.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X42 VDD.t135 a_11235_n6821# a_10542_n5707# VDD.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X43 VDD.t122 VDD.t121 VDD.t122 VDD.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X44 a_2151_594.t7 comparator_top_0.VINM a_2093_3714.t5 VDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
D2 DVSS.t180 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X45 comparator_top_0.comparator_0.VBN.t0 a_2221_8623.t6 a_1821_8526.t1 VDD.t40 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X46 a_7464_n6798# a_7096_n5816# DVSS.t29 DVSS.t28 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVSS.t163 DVSS.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_11749_n6043# VDD.t154 VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X49 VDD.t76 a_570_n5724# a_1777_n6060# VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X50 a_5299_1782.t3 a_5299_1782.t2 VDD.t143 VDD.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X51 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp A1.t6 VDD.t72 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X52 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINP VDD.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.32 ps=20.6 w=1 l=0.5
X53 a_7889_n6842# a_7464_n6798# DVSS.t99 DVSS.t98 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X54 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD.t17 VDD.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X55 comparator_top_0.comparator_0.VOUT a_8881_1782.t3 VSS.t7 VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X56 EF_AMUX21m_1.invm_0.Y SELA.t1 DVSS.t3 DVSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X57 DVSS.t12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb DVSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X58 DVDD.t14 a_11271_4224# a_10975_4108# DVDD.t13 sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.297 ps=2.77 w=1.12 l=0.15
X59 a_11271_4224# a_11031_3400# DVSS.t171 DVSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X60 B1.t5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb B1.t4 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X61 VDD.t92 a_10542_n5707# a_11749_n6043# VDD.t91 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X62 VDD.t138 a_2151_4783.t9 a_2551_4880.t4 VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X63 a_2093_1782.t0 comparator_top_0.comparator_0.VBN.t10 VSS.t17 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X64 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp B2.t7 VDD.t139 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X65 a_838_n6794# a_470_n5812# DVSS.t137 DVSS.t136 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X66 a_2093_3714.t4 comparator_top_0.VINM a_2151_594.t6 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X67 a_11271_4224# a_10975_4108# DVDD.t10 DVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.157 ps=1.4 w=1.12 l=0.15
X68 EF_AMUX21m_2.invm_0.Y SELB.t0 DVDD.t20 DVDD.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X69 VDD.t21 a_3916_n5703# a_5123_n6039# VDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X70 a_3916_n5703# a_3816_n5791# DVSS.t115 DVSS.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X71 a_5299_1782.t7 comparator_top_0.VINP a_2093_1782.t9 VSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X72 VSS.t9 a_5299_3714.t8 a_5299_620.t1 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X73 DVSS.t113 a_3816_n5791# a_3916_n5703# DVSS.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X74 VDD.t120 VDD.t118 VDD.t119 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X75 VDD.t152 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp VDD.t151 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X76 VDD.t78 a_5299_1782.t0 a_5299_1782.t1 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X77 comparator_top_0.comparator_0.VBN.t6 comparator_top_0.comparator_0.VBN.t5 VSS.t15 VSS.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X78 DVSS.t34 a_10965_3602# a_10975_4108# DVSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X79 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_5123_n6039# VDD.t93 VDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X80 DVSS.t57 a_7196_n5728# a_8403_n6064# DVSS.t56 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X81 a_2093_1782.t7 VSS.t55 VSS.t56 VSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X82 a_570_n5724# a_470_n5812# DVSS.t135 DVSS.t134 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X83 a_10810_n6777# a_10442_n5795# DVSS.t125 DVSS.t124 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X84 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVSS.t17 DVSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X85 a_6349_9307# a_10809_9307# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X86 A2.t3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINP VDD.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X87 a_2151_4783.t7 a_2151_4783.t6 VDD.t136 VDD.t99 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X88 DVDD.t28 SELB.t1 EF_AMUX21m_2.invm_0.Y DVDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X89 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD.t147 VDD.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X90 a_6351_7717# a_10811_7187# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X91 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD.t150 VDD.t86 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X92 DVSS.t52 a_10810_n6777# a_11235_n6821# DVSS.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X93 DVSS.t97 a_7464_n6798# a_7889_n6842# DVSS.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X94 a_1821_8526.t2 a_2221_8623.t7 comparator_top_0.comparator_0.VBN.t1 VDD.t41 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X95 a_7889_n6842# a_7464_n6798# DVSS.t95 DVSS.t94 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X96 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_8403_n6064# DVSS.t141 DVSS.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X97 B2.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb B2.t0 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X98 a_2093_1782.t8 comparator_top_0.VINP a_5299_1782.t6 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X99 DVSS.t175 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp DVSS.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X100 EF_AMUX21m_2.invm_0.Y SELB.t2 DVSS.t10 DVSS.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X101 VSS.t54 VSS.t52 VSS.t54 VSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X102 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb B2.t3 DVSS.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X103 DVDD.t9 a_10975_4108# VO.t1 DVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.4 as=0.297 ps=2.77 w=1.12 l=0.15
X104 a_2151_4783.t0 comparator_top_0.VINM a_2093_1782.t5 VSS.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X105 A2.t1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp A2.t0 DVSS.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X106 VDD.t84 a_2551_620.t4 a_2551_620.t5 VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X107 DVSS.t170 a_11031_3400# a_10965_3602# DVSS.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X108 VSS.t1 a_5299_3714.t2 a_5299_3714.t3 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X109 a_2151_594.t5 comparator_top_0.VINM a_2093_3714.t3 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X110 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD.t27 VDD.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X111 a_1263_n6838# a_838_n6794# DVSS.t155 DVSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X112 VDD.t117 VDD.t114 VDD.t116 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X113 DVSS.t168 a_11031_3400# a_11271_4224# DVSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X114 a_570_n5724# a_470_n5812# DVSS.t133 DVSS.t132 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X115 DVSS.t91 SELB.t3 EF_AMUX21m_2.invm_0.Y DVSS.t90 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X116 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD.t71 VDD.t70 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X117 VDD.t31 a_1263_n6838# a_570_n5724# VDD.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X118 VSS.t51 VSS.t49 VSS.t51 VSS.t50 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X119 DVSS.t179 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb DVSS.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X120 VDD.t53 a_1821_8526.t7 a_2221_8623.t2 VDD.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X121 a_6351_6657# a_1821_8526.t0 DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X122 a_11235_n6821# a_10810_n6777# DVSS.t50 DVSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X123 a_6349_9307# a_10811_8247# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X124 VDD.t113 VDD.t112 VDD.t113 VDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X125 a_2093_1782.t4 comparator_top_0.VINM a_2151_4783.t3 VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X126 comparator_top_0.comparator_0.VBP comparator_top_0.comparator_0.VBP VDD.t7 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=2
X127 VDD.t133 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VDD.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X128 a_10810_n6777# a_10442_n5795# DVDD.t24 DVDD.t23 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X129 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 VDD.t1 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X130 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINM DVSS.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X131 a_7196_n5728# a_7096_n5816# DVSS.t27 DVSS.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X132 VSS.t48 VSS.t45 VSS.t47 VSS.t46 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
D3 DVSS.t55 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X133 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINM VDD.t131 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.32 ps=20.6 w=1 l=0.5
X134 DVSS.t111 a_3816_n5791# a_3916_n5703# DVSS.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X135 A2.t7 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINP DVSS.t173 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X136 DVSS.t25 a_7096_n5816# a_7196_n5728# DVSS.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X137 comparator_top_0.comparator_0.VBN.t7 a_2221_8623.t8 a_1821_8526.t4 VDD.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X138 VDD.t157 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X139 DVSS.t153 a_838_n6794# a_1263_n6838# DVSS.t152 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X140 a_1263_n6838# a_838_n6794# DVSS.t151 DVSS.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X141 DVSS.t131 a_470_n5812# a_570_n5724# DVSS.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X142 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVSS.t73 DVSS.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X143 VSS.t13 comparator_top_0.comparator_0.VBN.t11 a_2221_8623.t4 VSS.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X144 VDD.t13 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X145 DVSS.t48 a_10810_n6777# a_11235_n6821# DVSS.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X146 a_2551_620.t3 a_2551_620.t2 VDD.t128 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X147 a_2093_3714.t11 comparator_top_0.VINP a_5299_3714.t5 VDD.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X148 a_4609_n6817# a_4184_n6773# DVSS.t188 DVSS.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X149 DVDD.t5 SELA.t2 a_470_n5812# DVDD.t4 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X150 a_11235_n6821# a_10810_n6777# DVSS.t46 DVSS.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X151 VSS.t69 a_2551_4880.t6 a_5299_620.t3 VSS.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X152 a_5299_620.t0 a_5299_3714.t9 VSS.t67 VSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X153 VDD.t35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X154 A1.t5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp A1.t4 DVSS.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X155 DVSS.t54 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb DVSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X156 A1.t3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINP DVSS.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X157 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 VDD.t11 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X158 VDD.t82 a_5299_1782.t8 a_5299_620.t4 VDD.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X159 B1.t3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINM VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X160 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINM VDD.t60 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X161 DVSS.t83 EF_AMUX21m_1.invm_0.Y a_3816_n5791# DVSS.t82 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X162 DVSS.t23 a_7096_n5816# a_7196_n5728# DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X163 B1.t1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp B1.t0 DVSS.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X164 a_3916_n5703# a_3816_n5791# DVSS.t109 DVSS.t108 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X165 a_2221_8623.t1 a_1821_8526.t8 VDD.t51 VDD.t50 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X166 VDD.t111 VDD.t110 a_2093_3714.t6 VDD.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X167 a_2151_4783.t2 comparator_top_0.VINM a_2093_1782.t3 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X168 a_7196_n5728# a_7096_n5816# DVSS.t21 DVSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X169 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb A1.t2 DVSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X170 DVSS.t61 SELA.t3 a_470_n5812# DVSS.t60 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X171 VDD.t74 a_570_n5724# a_1263_n6838# VDD.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X172 a_5299_620.t2 a_2551_4880.t7 VSS.t23 VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X173 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINP VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X174 A1.t1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb A1.t0 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X175 a_1263_n6838# a_838_n6794# DVSS.t149 DVSS.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X176 DVSS.t129 a_470_n5812# a_570_n5724# DVSS.t128 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X177 a_2093_3714.t2 comparator_top_0.VINM a_2151_594.t4 VDD.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X178 VDD.t69 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 VDD.t68 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X179 VDD.t90 a_10542_n5707# a_11235_n6821# VDD.t89 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X180 VSS.t44 VSS.t43 VSS.t44 VSS.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X181 a_11271_4224# a_11031_3400# DVSS.t167 DVSS.t166 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X182 a_11235_n6821# a_10810_n6777# DVSS.t44 DVSS.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X183 DVSS.t186 a_4184_n6773# a_4609_n6817# DVSS.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X184 a_2151_594.t3 a_2151_594.t2 VSS.t70 VSS.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X185 VSS.t21 a_2551_4880.t2 a_2551_4880.t3 VSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X186 a_10975_4108# a_10965_3602# DVSS.t32 DVSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X187 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp A2.t2 VDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X188 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_11749_n6043# DVSS.t177 DVSS.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X189 a_2221_8623.t5 VSS.t40 VSS.t42 VSS.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X190 VDD.t158 a_2551_620.t6 a_5299_620.t7 VDD.t141 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X191 VDD.t23 a_7889_n6842# a_7196_n5728# VDD.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X192 a_5299_3714.t4 comparator_top_0.VINP a_2093_3714.t8 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X193 B1.t6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINM DVSS.t144 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X194 comparator_top_0.comparator_0.VBP VSS.t37 VSS.t39 VSS.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X195 a_5299_3714.t1 a_5299_3714.t0 VSS.t28 VSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X196 a_10542_n5707# a_10442_n5795# DVSS.t123 DVSS.t122 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X197 DVSS.t87 a_10542_n5707# a_11749_n6043# DVSS.t86 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X198 DVDD.t3 SELA.t4 EF_AMUX21m_1.invm_0.Y DVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X199 DVDD.t1 SELB.t4 a_7096_n5816# DVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X200 a_1821_8526.t5 a_2221_8623.t9 comparator_top_0.comparator_0.VBN.t8 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X201 a_10965_3602# a_11031_3400# VDD.t149 VDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X202 a_11031_3400# comparator_top_0.comparator_0.VOUT VDD.t43 VDD.t42 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X203 a_2093_1782.t11 comparator_top_0.VINP a_5299_1782.t5 VSS.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X204 a_2551_4880.t1 a_2551_4880.t0 VSS.t5 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X205 DVSS.t7 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb DVSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X206 DVSS.t71 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 DVSS.t70 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X207 DVDD.t18 EF_AMUX21m_1.invm_0.Y a_3816_n5791# DVDD.t17 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X208 a_5299_620.t5 a_5299_1782.t9 VDD.t95 VDD.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X209 VDD.t109 VDD.t108 VDD.t109 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X210 VDD.t39 a_7196_n5728# a_8403_n6064# VDD.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X211 a_4609_n6817# a_4184_n6773# DVSS.t184 DVSS.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X212 DVSS.t182 a_4184_n6773# a_4609_n6817# DVSS.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X213 DVSS.t69 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 DVSS.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X214 VDD.t59 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp VDD.t58 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X215 VDD.t45 a_2151_4783.t4 a_2151_4783.t5 VDD.t44 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X216 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVSS.t67 DVSS.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X217 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_8403_n6064# VDD.t129 VDD.t38 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X218 a_2551_620.t0 a_2151_594.t9 VSS.t26 VSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X219 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINP DVSS.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=0.5
X220 DVSS.t161 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 DVSS.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X221 VSS.t36 VSS.t34 a_2093_1782.t6 VSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X222 a_3916_n5703# a_3816_n5791# DVSS.t107 DVSS.t106 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X223 DVSS.t159 SELB.t5 a_7096_n5816# DVSS.t158 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X224 VDD.t96 a_10809_9307# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X225 VDD.t5 comparator_top_0.comparator_0.VBP a_2093_3714.t0 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X226 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD.t130 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X227 B2.t6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINM VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X228 VDD.t15 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X229 a_7196_n5728# a_7096_n5816# DVSS.t19 DVSS.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X230 DVSS.t1 SELA.t5 EF_AMUX21m_1.invm_0.Y DVSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X231 DVSS.t165 a_11031_3400# a_11271_4224# DVSS.t164 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X232 VSS.t3 a_2151_594.t0 a_2151_594.t1 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X233 a_5299_620.t6 a_2551_620.t7 VDD.t159 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X234 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp B1.t2 VDD.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X235 a_2093_1782.t2 comparator_top_0.VINM a_2151_4783.t1 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X236 DVSS.t143 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp DVSS.t142 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X237 DVSS.t147 a_838_n6794# a_1263_n6838# DVSS.t146 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X238 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp comparator_top_0.VINP DVSS.t80 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X239 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb A2.t6 DVSS.t172 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X240 VDD.t19 a_3916_n5703# a_4609_n6817# VDD.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X241 DVSS.t31 a_10965_3602# a_10975_4108# DVSS.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X242 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 VDD.t155 VDD.t24 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X243 VSS.t33 VSS.t32 VSS.t33 VSS.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X244 a_6351_7717# a_10811_8247# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X245 VDD.t101 a_5299_620.t9 a_8881_1782.t1 VDD.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=2
X246 VDD.t107 VDD.t105 VDD.t107 VDD.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X247 VDD.t57 a_4609_n6817# a_3916_n5703# VDD.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X248 VDD.t66 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X249 a_2221_8623.t0 a_1821_8526.t9 VDD.t49 VDD.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X250 VDD.t104 VDD.t102 VDD.t104 VDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X251 a_5299_1782.t4 comparator_top_0.VINP a_2093_1782.t10 VSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X252 A2.t5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb A2.t4 VDD.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X253 DVSS.t121 a_10442_n5795# a_10542_n5707# DVSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X254 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD.t64 VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X255 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 VDD.t33 VDD.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X256 DVSS.t79 EF_AMUX21m_2.invm_0.Y a_10442_n5795# DVSS.t78 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X257 DVSS.t15 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 DVSS.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X258 a_4184_n6773# a_3816_n5791# DVSS.t105 DVSS.t104 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X259 a_10542_n5707# a_10442_n5795# DVSS.t119 DVSS.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X260 VSS.t11 comparator_top_0.comparator_0.VBN.t12 comparator_top_0.comparator_0.VBP VSS.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X261 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_1777_n6060# DVSS.t93 DVSS.t92 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X262 VDD.t145 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 VDD.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X263 VDD.t37 a_7196_n5728# a_7889_n6842# VDD.t36 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X264 B2.t2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb comparator_top_0.VINM DVSS.t62 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X265 B2.t5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp B2.t4 DVSS.t156 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X266 DVSS.t117 a_10442_n5795# a_10542_n5707# DVSS.t116 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
R0 comparator_top_0.comparator_0.VBN.n263 comparator_top_0.comparator_0.VBN.t5 60.2505
R1 comparator_top_0.comparator_0.VBN.n284 comparator_top_0.comparator_0.VBN.t11 60.2505
R2 comparator_top_0.comparator_0.VBN.n304 comparator_top_0.comparator_0.VBN.t12 60.2505
R3 comparator_top_0.comparator_0.VBN.n306 comparator_top_0.comparator_0.VBN.t10 60.2505
R4 comparator_top_0.comparator_0.VBN.n318 comparator_top_0.comparator_0.VBN.t9 60.2505
R5 comparator_top_0.comparator_0.VBN.n97 comparator_top_0.comparator_0.VBN.n95 41.8847
R6 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.t4 35.1154
R7 comparator_top_0.comparator_0.VBN.n105 comparator_top_0.comparator_0.VBN.n102 26.3366
R8 comparator_top_0.comparator_0.VBN.n52 comparator_top_0.comparator_0.VBN.n51 26.3366
R9 comparator_top_0.comparator_0.VBN.n38 comparator_top_0.comparator_0.VBN.n35 26.3366
R10 comparator_top_0.comparator_0.VBN.n97 comparator_top_0.comparator_0.VBN.n96 15.9528
R11 comparator_top_0.comparator_0.VBN.n44 comparator_top_0.comparator_0.VBN.n42 12.8005
R12 comparator_top_0.comparator_0.VBN.n44 comparator_top_0.comparator_0.VBN.n43 12.8005
R13 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n267 9.3005
R14 comparator_top_0.comparator_0.VBN.n273 comparator_top_0.comparator_0.VBN.n272 9.3005
R15 comparator_top_0.comparator_0.VBN.n282 comparator_top_0.comparator_0.VBN.n281 9.3005
R16 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n276 9.3005
R17 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n287 9.3005
R18 comparator_top_0.comparator_0.VBN.n302 comparator_top_0.comparator_0.VBN.n301 9.3005
R19 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n296 9.3005
R20 comparator_top_0.comparator_0.VBN.n293 comparator_top_0.comparator_0.VBN.n292 9.3005
R21 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n23 9.3005
R22 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n31 9.3005
R23 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n40 9.3005
R24 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n46 9.3005
R25 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n55 9.3005
R26 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n63 9.3005
R27 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n71 9.3005
R28 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n79 9.3005
R29 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n87 9.3005
R30 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n86 9.3005
R31 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n85 9.3005
R32 comparator_top_0.comparator_0.VBN.n85 comparator_top_0.comparator_0.VBN.n84 9.3005
R33 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n78 9.3005
R34 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n77 9.3005
R35 comparator_top_0.comparator_0.VBN.n77 comparator_top_0.comparator_0.VBN.n76 9.3005
R36 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n70 9.3005
R37 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n69 9.3005
R38 comparator_top_0.comparator_0.VBN.n69 comparator_top_0.comparator_0.VBN.n68 9.3005
R39 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n62 9.3005
R40 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n61 9.3005
R41 comparator_top_0.comparator_0.VBN.n61 comparator_top_0.comparator_0.VBN.n60 9.3005
R42 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n54 9.3005
R43 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n53 9.3005
R44 comparator_top_0.comparator_0.VBN.n53 comparator_top_0.comparator_0.VBN.n52 9.3005
R45 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n45 9.3005
R46 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n41 9.3005
R47 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n39 9.3005
R48 comparator_top_0.comparator_0.VBN.n39 comparator_top_0.comparator_0.VBN.n38 9.3005
R49 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n32 9.3005
R50 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n30 9.3005
R51 comparator_top_0.comparator_0.VBN.n30 comparator_top_0.comparator_0.VBN.n29 9.3005
R52 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n24 9.3005
R53 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n22 9.3005
R54 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n155 9.3005
R55 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n147 9.3005
R56 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n139 9.3005
R57 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n131 9.3005
R58 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n123 9.3005
R59 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n115 9.3005
R60 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n107 9.3005
R61 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n98 9.3005
R62 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n106 9.3005
R63 comparator_top_0.comparator_0.VBN.n106 comparator_top_0.comparator_0.VBN.n105 9.3005
R64 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n99 9.3005
R65 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n108 9.3005
R66 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n114 9.3005
R67 comparator_top_0.comparator_0.VBN.n114 comparator_top_0.comparator_0.VBN.n113 9.3005
R68 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n122 9.3005
R69 comparator_top_0.comparator_0.VBN.n122 comparator_top_0.comparator_0.VBN.n121 9.3005
R70 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n116 9.3005
R71 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n124 9.3005
R72 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n130 9.3005
R73 comparator_top_0.comparator_0.VBN.n130 comparator_top_0.comparator_0.VBN.n129 9.3005
R74 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n138 9.3005
R75 comparator_top_0.comparator_0.VBN.n138 comparator_top_0.comparator_0.VBN.n137 9.3005
R76 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n132 9.3005
R77 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n140 9.3005
R78 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n146 9.3005
R79 comparator_top_0.comparator_0.VBN.n146 comparator_top_0.comparator_0.VBN.n145 9.3005
R80 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n154 9.3005
R81 comparator_top_0.comparator_0.VBN.n154 comparator_top_0.comparator_0.VBN.n153 9.3005
R82 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n148 9.3005
R83 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n156 9.3005
R84 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n162 9.3005
R85 comparator_top_0.comparator_0.VBN.n162 comparator_top_0.comparator_0.VBN.n161 9.3005
R86 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n170 9.3005
R87 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n171 9.3005
R88 comparator_top_0.comparator_0.VBN.n177 comparator_top_0.comparator_0.VBN.n176 9.3005
R89 comparator_top_0.comparator_0.VBN.n92 comparator_top_0.comparator_0.VBN.n91 9.3005
R90 comparator_top_0.comparator_0.VBN.n167 comparator_top_0.comparator_0.VBN.n166 9.3005
R91 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n315 9.3005
R92 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n313 9.3005
R93 comparator_top_0.comparator_0.VBN.n313 comparator_top_0.comparator_0.VBN.n312 9.3005
R94 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n314 9.3005
R95 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n327 9.3005
R96 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n326 9.3005
R97 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n325 9.3005
R98 comparator_top_0.comparator_0.VBN.n325 comparator_top_0.comparator_0.VBN.n324 9.3005
R99 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n246 9.3005
R100 comparator_top_0.comparator_0.VBN.n252 comparator_top_0.comparator_0.VBN.n251 9.3005
R101 comparator_top_0.comparator_0.VBN.n261 comparator_top_0.comparator_0.VBN.n260 9.3005
R102 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n255 9.3005
R103 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n242 9.3005
R104 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n241 9.3005
R105 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n243 9.3005
R106 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n197 9.3005
R107 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n192 9.3005
R108 comparator_top_0.comparator_0.VBN.n285 comparator_top_0.comparator_0.VBN.n284 8.76429
R109 comparator_top_0.comparator_0.VBN.n305 comparator_top_0.comparator_0.VBN.n304 8.76429
R110 comparator_top_0.comparator_0.VBN.n264 comparator_top_0.comparator_0.VBN.n263 8.76429
R111 comparator_top_0.comparator_0.VBN.n271 comparator_top_0.comparator_0.VBN.n270 8.21641
R112 comparator_top_0.comparator_0.VBN.n280 comparator_top_0.comparator_0.VBN.n279 8.21641
R113 comparator_top_0.comparator_0.VBN.n291 comparator_top_0.comparator_0.VBN.n290 8.21641
R114 comparator_top_0.comparator_0.VBN.n300 comparator_top_0.comparator_0.VBN.n299 8.21641
R115 comparator_top_0.comparator_0.VBN.n311 comparator_top_0.comparator_0.VBN.n310 8.21641
R116 comparator_top_0.comparator_0.VBN.n323 comparator_top_0.comparator_0.VBN.n322 8.21641
R117 comparator_top_0.comparator_0.VBN.n250 comparator_top_0.comparator_0.VBN.n249 8.21641
R118 comparator_top_0.comparator_0.VBN.n259 comparator_top_0.comparator_0.VBN.n258 8.21641
R119 comparator_top_0.comparator_0.VBN.n160 comparator_top_0.comparator_0.VBN.n159 7.95102
R120 comparator_top_0.comparator_0.VBN.n165 comparator_top_0.comparator_0.VBN.n164 7.95102
R121 comparator_top_0.comparator_0.VBN.n105 comparator_top_0.comparator_0.VBN.n104 7.45411
R122 comparator_top_0.comparator_0.VBN.n52 comparator_top_0.comparator_0.VBN.n50 7.45411
R123 comparator_top_0.comparator_0.VBN.n38 comparator_top_0.comparator_0.VBN.n37 7.45411
R124 comparator_top_0.comparator_0.VBN.n152 comparator_top_0.comparator_0.VBN.n151 6.9572
R125 comparator_top_0.comparator_0.VBN.n175 comparator_top_0.comparator_0.VBN.n174 6.9572
R126 comparator_top_0.comparator_0.VBN.n319 comparator_top_0.comparator_0.VBN.n318 6.92242
R127 comparator_top_0.comparator_0.VBN.n307 comparator_top_0.comparator_0.VBN.n306 6.92012
R128 comparator_top_0.comparator_0.VBN.n113 comparator_top_0.comparator_0.VBN.n112 6.46029
R129 comparator_top_0.comparator_0.VBN.n60 comparator_top_0.comparator_0.VBN.n59 6.46029
R130 comparator_top_0.comparator_0.VBN.n29 comparator_top_0.comparator_0.VBN.n28 6.46029
R131 comparator_top_0.comparator_0.VBN.n158 comparator_top_0.comparator_0.VBN.n157 6.02403
R132 comparator_top_0.comparator_0.VBN.n144 comparator_top_0.comparator_0.VBN.n143 5.96339
R133 comparator_top_0.comparator_0.VBN.n90 comparator_top_0.comparator_0.VBN.n89 5.96339
R134 comparator_top_0.comparator_0.VBN.n269 comparator_top_0.comparator_0.VBN.n268 5.64756
R135 comparator_top_0.comparator_0.VBN.n278 comparator_top_0.comparator_0.VBN.n277 5.64756
R136 comparator_top_0.comparator_0.VBN.n289 comparator_top_0.comparator_0.VBN.n288 5.64756
R137 comparator_top_0.comparator_0.VBN.n298 comparator_top_0.comparator_0.VBN.n297 5.64756
R138 comparator_top_0.comparator_0.VBN.n106 comparator_top_0.comparator_0.VBN.n101 5.64756
R139 comparator_top_0.comparator_0.VBN.n53 comparator_top_0.comparator_0.VBN.n48 5.64756
R140 comparator_top_0.comparator_0.VBN.n39 comparator_top_0.comparator_0.VBN.n34 5.64756
R141 comparator_top_0.comparator_0.VBN.n309 comparator_top_0.comparator_0.VBN.n308 5.64756
R142 comparator_top_0.comparator_0.VBN.n321 comparator_top_0.comparator_0.VBN.n320 5.64756
R143 comparator_top_0.comparator_0.VBN.n248 comparator_top_0.comparator_0.VBN.n247 5.64756
R144 comparator_top_0.comparator_0.VBN.n257 comparator_top_0.comparator_0.VBN.n256 5.64756
R145 comparator_top_0.comparator_0.VBN.n210 comparator_top_0.comparator_0.VBN.t1 5.5395
R146 comparator_top_0.comparator_0.VBN.n210 comparator_top_0.comparator_0.VBN.t7 5.5395
R147 comparator_top_0.comparator_0.VBN.n227 comparator_top_0.comparator_0.VBN.t8 5.5395
R148 comparator_top_0.comparator_0.VBN.n227 comparator_top_0.comparator_0.VBN.t0 5.5395
R149 comparator_top_0.comparator_0.VBN.n121 comparator_top_0.comparator_0.VBN.n120 5.46648
R150 comparator_top_0.comparator_0.VBN.n68 comparator_top_0.comparator_0.VBN.n67 5.46648
R151 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n244 5.28563
R152 comparator_top_0.comparator_0.VBN.n150 comparator_top_0.comparator_0.VBN.n149 5.27109
R153 comparator_top_0.comparator_0.VBN.n136 comparator_top_0.comparator_0.VBN.n135 4.96957
R154 comparator_top_0.comparator_0.VBN.n83 comparator_top_0.comparator_0.VBN.n82 4.96957
R155 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n266 4.911
R156 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n286 4.911
R157 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n275 4.91005
R158 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n254 4.91005
R159 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n295 4.90905
R160 comparator_top_0.comparator_0.VBN.n114 comparator_top_0.comparator_0.VBN.n110 4.89462
R161 comparator_top_0.comparator_0.VBN.n61 comparator_top_0.comparator_0.VBN.n57 4.89462
R162 comparator_top_0.comparator_0.VBN.n30 comparator_top_0.comparator_0.VBN.n26 4.89462
R163 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n245 4.76425
R164 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n44 4.6505
R165 comparator_top_0.comparator_0.VBN.n142 comparator_top_0.comparator_0.VBN.n141 4.51815
R166 comparator_top_0.comparator_0.VBN.n169 comparator_top_0.comparator_0.VBN.n163 4.51815
R167 comparator_top_0.comparator_0.VBN.n195 comparator_top_0.comparator_0.VBN.n194 4.51815
R168 comparator_top_0.comparator_0.VBN.n206 comparator_top_0.comparator_0.VBN.n205 4.51815
R169 comparator_top_0.comparator_0.VBN.n236 comparator_top_0.comparator_0.VBN.n235 4.51815
R170 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n94 4.5005
R171 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n182 4.5005
R172 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n179 4.5005
R173 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n169 4.5005
R174 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n274 4.5005
R175 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n283 4.5005
R176 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n303 4.5005
R177 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n294 4.5005
R178 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n253 4.5005
R179 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n262 4.5005
R180 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n195 4.5005
R181 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n190 4.5005
R182 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n185 4.5005
R183 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n239 4.5005
R184 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n200 4.5005
R185 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n216 4.5005
R186 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n204 4.5005
R187 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n213 4.5005
R188 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n209 4.5005
R189 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n226 4.5005
R190 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n231 4.5005
R191 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n234 4.5005
R192 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n220 4.5005
R193 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n224 4.5005
R194 comparator_top_0.comparator_0.VBN.n129 comparator_top_0.comparator_0.VBN.n128 4.47267
R195 comparator_top_0.comparator_0.VBN.n76 comparator_top_0.comparator_0.VBN.n75 4.47267
R196 comparator_top_0.comparator_0.VBN.n21 comparator_top_0.comparator_0.VBN.n7 4.44875
R197 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n316 7.3305
R198 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n329 4.24504
R199 comparator_top_0.comparator_0.VBN.n122 comparator_top_0.comparator_0.VBN.n118 4.14168
R200 comparator_top_0.comparator_0.VBN.n69 comparator_top_0.comparator_0.VBN.n65 4.14168
R201 comparator_top_0.comparator_0.VBN.n128 comparator_top_0.comparator_0.VBN.n127 3.97576
R202 comparator_top_0.comparator_0.VBN.n75 comparator_top_0.comparator_0.VBN.n74 3.97576
R203 comparator_top_0.comparator_0.VBN.n134 comparator_top_0.comparator_0.VBN.n133 3.76521
R204 comparator_top_0.comparator_0.VBN.n179 comparator_top_0.comparator_0.VBN.n173 3.76521
R205 comparator_top_0.comparator_0.VBN.n182 comparator_top_0.comparator_0.VBN.n180 3.76521
R206 comparator_top_0.comparator_0.VBN.n81 comparator_top_0.comparator_0.VBN.n80 3.76521
R207 comparator_top_0.comparator_0.VBN.n239 comparator_top_0.comparator_0.VBN.n238 3.76521
R208 comparator_top_0.comparator_0.VBN.n137 comparator_top_0.comparator_0.VBN.n136 3.47885
R209 comparator_top_0.comparator_0.VBN.n84 comparator_top_0.comparator_0.VBN.n83 3.47885
R210 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n307 3.47756
R211 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n319 3.4767
R212 comparator_top_0.comparator_0.VBN.n130 comparator_top_0.comparator_0.VBN.n126 3.38874
R213 comparator_top_0.comparator_0.VBN.n77 comparator_top_0.comparator_0.VBN.n73 3.38874
R214 comparator_top_0.comparator_0.VBN.n186 comparator_top_0.comparator_0.VBN.t2 3.3065
R215 comparator_top_0.comparator_0.VBN.n186 comparator_top_0.comparator_0.VBN.t6 3.3065
R216 comparator_top_0.comparator_0.VBN.n190 comparator_top_0.comparator_0.VBN.n188 3.74814
R217 comparator_top_0.comparator_0.VBN.n15 comparator_top_0.comparator_0.VBN.n187 3.15814
R218 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n285 3.03311
R219 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n305 3.03311
R220 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n264 3.03311
R221 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n206 3.03311
R222 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n236 3.03311
R223 comparator_top_0.comparator_0.VBN.n126 comparator_top_0.comparator_0.VBN.n125 3.01226
R224 comparator_top_0.comparator_0.VBN.n94 comparator_top_0.comparator_0.VBN.n88 3.01226
R225 comparator_top_0.comparator_0.VBN.n73 comparator_top_0.comparator_0.VBN.n72 3.01226
R226 comparator_top_0.comparator_0.VBN.n190 comparator_top_0.comparator_0.VBN.n189 3.01226
R227 comparator_top_0.comparator_0.VBN.n120 comparator_top_0.comparator_0.VBN.n119 2.98194
R228 comparator_top_0.comparator_0.VBN.n67 comparator_top_0.comparator_0.VBN.n66 2.98194
R229 comparator_top_0.comparator_0.VBN.n138 comparator_top_0.comparator_0.VBN.n134 2.63579
R230 comparator_top_0.comparator_0.VBN.n85 comparator_top_0.comparator_0.VBN.n81 2.63579
R231 comparator_top_0.comparator_0.VBN.n239 comparator_top_0.comparator_0.VBN.n237 2.63579
R232 comparator_top_0.comparator_0.VBN.n204 comparator_top_0.comparator_0.VBN.n202 2.63579
R233 comparator_top_0.comparator_0.VBN.n224 comparator_top_0.comparator_0.VBN.n222 2.63579
R234 comparator_top_0.comparator_0.VBN.n192 comparator_top_0.comparator_0.VBN.n191 2.61733
R235 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n198 2.60826
R236 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n218 2.60817
R237 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n183 2.53421
R238 comparator_top_0.comparator_0.VBN.n145 comparator_top_0.comparator_0.VBN.n144 2.48504
R239 comparator_top_0.comparator_0.VBN.n91 comparator_top_0.comparator_0.VBN.n90 2.48504
R240 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n17 2.42663
R241 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n20 2.39724
R242 comparator_top_0.comparator_0.VBN.n118 comparator_top_0.comparator_0.VBN.n117 2.25932
R243 comparator_top_0.comparator_0.VBN.n65 comparator_top_0.comparator_0.VBN.n64 2.25932
R244 comparator_top_0.comparator_0.VBN.n216 comparator_top_0.comparator_0.VBN.n214 2.25932
R245 comparator_top_0.comparator_0.VBN.n208 comparator_top_0.comparator_0.VBN.n207 2.25932
R246 comparator_top_0.comparator_0.VBN.n234 comparator_top_0.comparator_0.VBN.n232 2.25932
R247 comparator_top_0.comparator_0.VBN.n230 comparator_top_0.comparator_0.VBN.n229 2.25932
R248 comparator_top_0.comparator_0.VBN.n216 comparator_top_0.comparator_0.VBN.n215 2.25379
R249 comparator_top_0.comparator_0.VBN.n234 comparator_top_0.comparator_0.VBN.n233 2.25379
R250 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n317 2.2505
R251 comparator_top_0.comparator_0.VBN.n197 comparator_top_0.comparator_0.VBN.n196 2.24766
R252 comparator_top_0.comparator_0.VBN.n265 comparator_top_0.comparator_0.VBN.n18 2.073
R253 comparator_top_0.comparator_0.VBN comparator_top_0.comparator_0.VBN.n19 2.06925
R254 comparator_top_0.comparator_0.VBN.n112 comparator_top_0.comparator_0.VBN.n111 1.98813
R255 comparator_top_0.comparator_0.VBN.n59 comparator_top_0.comparator_0.VBN.n58 1.98813
R256 comparator_top_0.comparator_0.VBN.n28 comparator_top_0.comparator_0.VBN.n27 1.98813
R257 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n172 1.94045
R258 comparator_top_0.comparator_0.VBN.n146 comparator_top_0.comparator_0.VBN.n142 1.88285
R259 comparator_top_0.comparator_0.VBN.n93 comparator_top_0.comparator_0.VBN.n92 1.88285
R260 comparator_top_0.comparator_0.VBN.n195 comparator_top_0.comparator_0.VBN.n193 1.88285
R261 comparator_top_0.comparator_0.VBN.n204 comparator_top_0.comparator_0.VBN.n203 1.87949
R262 comparator_top_0.comparator_0.VBN.n224 comparator_top_0.comparator_0.VBN.n223 1.87949
R263 comparator_top_0.comparator_0.VBN.n265 comparator_top_0.comparator_0.VBN.n3 1.85011
R264 comparator_top_0.comparator_0.VBN.n217 comparator_top_0.comparator_0.VBN.n1 1.73899
R265 comparator_top_0.comparator_0.VBN.n21 comparator_top_0.comparator_0.VBN.n172 1.70776
R266 comparator_top_0.comparator_0.VBN.n19 comparator_top_0.comparator_0.VBN.n2 1.70567
R267 comparator_top_0.comparator_0.VBN.n15 comparator_top_0.comparator_0.VBN.n186 1.61779
R268 comparator_top_0.comparator_0.VBN.n95 comparator_top_0.comparator_0.VBN.t3 1.60717
R269 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN 1.60425
R270 comparator_top_0.comparator_0.VBN.n110 comparator_top_0.comparator_0.VBN.n109 1.50638
R271 comparator_top_0.comparator_0.VBN.n169 comparator_top_0.comparator_0.VBN.n168 1.50638
R272 comparator_top_0.comparator_0.VBN.n179 comparator_top_0.comparator_0.VBN.n178 1.50638
R273 comparator_top_0.comparator_0.VBN.n94 comparator_top_0.comparator_0.VBN.n93 1.50638
R274 comparator_top_0.comparator_0.VBN.n57 comparator_top_0.comparator_0.VBN.n56 1.50638
R275 comparator_top_0.comparator_0.VBN.n26 comparator_top_0.comparator_0.VBN.n25 1.50638
R276 comparator_top_0.comparator_0.VBN.n213 comparator_top_0.comparator_0.VBN.n212 1.50638
R277 comparator_top_0.comparator_0.VBN.n226 comparator_top_0.comparator_0.VBN.n225 1.50638
R278 comparator_top_0.comparator_0.VBN.n228 comparator_top_0.comparator_0.VBN.n227 1.50151
R279 comparator_top_0.comparator_0.VBN.n211 comparator_top_0.comparator_0.VBN.n210 1.50148
R280 comparator_top_0.comparator_0.VBN.n153 comparator_top_0.comparator_0.VBN.n152 1.49122
R281 comparator_top_0.comparator_0.VBN.n176 comparator_top_0.comparator_0.VBN.n175 1.49122
R282 comparator_top_0.comparator_0.VBN.n19 comparator_top_0.comparator_0.VBN.n265 1.26925
R283 comparator_top_0.comparator_0.VBN.n217 comparator_top_0.comparator_0.VBN.n0 1.1968
R284 comparator_top_0.comparator_0.VBN.n19 comparator_top_0.comparator_0.VBN.n21 1.1545
R285 comparator_top_0.comparator_0.VBN.n154 comparator_top_0.comparator_0.VBN.n150 1.12991
R286 comparator_top_0.comparator_0.VBN.n178 comparator_top_0.comparator_0.VBN.n177 1.12991
R287 comparator_top_0.comparator_0.VBN.n185 comparator_top_0.comparator_0.VBN.n184 1.12991
R288 comparator_top_0.comparator_0.VBN.n272 comparator_top_0.comparator_0.VBN.n271 1.09595
R289 comparator_top_0.comparator_0.VBN.n281 comparator_top_0.comparator_0.VBN.n280 1.09595
R290 comparator_top_0.comparator_0.VBN.n292 comparator_top_0.comparator_0.VBN.n291 1.09595
R291 comparator_top_0.comparator_0.VBN.n301 comparator_top_0.comparator_0.VBN.n300 1.09595
R292 comparator_top_0.comparator_0.VBN.n312 comparator_top_0.comparator_0.VBN.n311 1.09595
R293 comparator_top_0.comparator_0.VBN.n324 comparator_top_0.comparator_0.VBN.n323 1.09595
R294 comparator_top_0.comparator_0.VBN.n251 comparator_top_0.comparator_0.VBN.n250 1.09595
R295 comparator_top_0.comparator_0.VBN.n260 comparator_top_0.comparator_0.VBN.n259 1.09595
R296 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n97 1.03132
R297 comparator_top_0.comparator_0.VBN.n104 comparator_top_0.comparator_0.VBN.n103 0.994314
R298 comparator_top_0.comparator_0.VBN.n50 comparator_top_0.comparator_0.VBN.n49 0.994314
R299 comparator_top_0.comparator_0.VBN.n37 comparator_top_0.comparator_0.VBN.n36 0.994314
R300 comparator_top_0.comparator_0.VBN.n183 comparator_top_0.comparator_0.VBN.n217 0.890264
R301 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n228 0.833627
R302 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n211 0.833623
R303 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n16 0.766876
R304 comparator_top_0.comparator_0.VBN.n274 comparator_top_0.comparator_0.VBN.n273 0.753441
R305 comparator_top_0.comparator_0.VBN.n273 comparator_top_0.comparator_0.VBN.n269 0.753441
R306 comparator_top_0.comparator_0.VBN.n282 comparator_top_0.comparator_0.VBN.n278 0.753441
R307 comparator_top_0.comparator_0.VBN.n283 comparator_top_0.comparator_0.VBN.n282 0.753441
R308 comparator_top_0.comparator_0.VBN.n294 comparator_top_0.comparator_0.VBN.n293 0.753441
R309 comparator_top_0.comparator_0.VBN.n293 comparator_top_0.comparator_0.VBN.n289 0.753441
R310 comparator_top_0.comparator_0.VBN.n302 comparator_top_0.comparator_0.VBN.n298 0.753441
R311 comparator_top_0.comparator_0.VBN.n303 comparator_top_0.comparator_0.VBN.n302 0.753441
R312 comparator_top_0.comparator_0.VBN.n101 comparator_top_0.comparator_0.VBN.n100 0.753441
R313 comparator_top_0.comparator_0.VBN.n48 comparator_top_0.comparator_0.VBN.n47 0.753441
R314 comparator_top_0.comparator_0.VBN.n34 comparator_top_0.comparator_0.VBN.n33 0.753441
R315 comparator_top_0.comparator_0.VBN.n313 comparator_top_0.comparator_0.VBN.n309 0.753441
R316 comparator_top_0.comparator_0.VBN.n325 comparator_top_0.comparator_0.VBN.n321 0.753441
R317 comparator_top_0.comparator_0.VBN.n253 comparator_top_0.comparator_0.VBN.n252 0.753441
R318 comparator_top_0.comparator_0.VBN.n252 comparator_top_0.comparator_0.VBN.n248 0.753441
R319 comparator_top_0.comparator_0.VBN.n261 comparator_top_0.comparator_0.VBN.n257 0.753441
R320 comparator_top_0.comparator_0.VBN.n262 comparator_top_0.comparator_0.VBN.n261 0.753441
R321 comparator_top_0.comparator_0.VBN.n200 comparator_top_0.comparator_0.VBN.n199 0.753441
R322 comparator_top_0.comparator_0.VBN.n209 comparator_top_0.comparator_0.VBN.n208 0.753441
R323 comparator_top_0.comparator_0.VBN.n220 comparator_top_0.comparator_0.VBN.n219 0.753441
R324 comparator_top_0.comparator_0.VBN.n231 comparator_top_0.comparator_0.VBN.n230 0.753441
R325 comparator_top_0.comparator_0.VBN.n329 comparator_top_0.comparator_0.VBN.n328 0.738413
R326 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n4 0.700653
R327 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n10 0.571152
R328 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n6 0.498175
R329 comparator_top_0.comparator_0.VBN.n161 comparator_top_0.comparator_0.VBN.n160 0.497407
R330 comparator_top_0.comparator_0.VBN.n166 comparator_top_0.comparator_0.VBN.n165 0.497407
R331 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n15 0.48986
R332 comparator_top_0.comparator_0.VBN.n241 comparator_top_0.comparator_0.VBN.n240 0.461175
R333 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n11 0.42713
R334 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n5 0.387304
R335 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n14 0.380935
R336 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n8 0.380935
R337 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n13 0.380935
R338 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n12 0.380935
R339 comparator_top_0.comparator_0.VBN.n162 comparator_top_0.comparator_0.VBN.n158 0.376971
R340 comparator_top_0.comparator_0.VBN.n168 comparator_top_0.comparator_0.VBN.n167 0.376971
R341 comparator_top_0.comparator_0.VBN.n182 comparator_top_0.comparator_0.VBN.n181 0.376971
R342 comparator_top_0.comparator_0.VBN.n202 comparator_top_0.comparator_0.VBN.n201 0.376971
R343 comparator_top_0.comparator_0.VBN.n222 comparator_top_0.comparator_0.VBN.n221 0.376971
R344 a_1821_8526.t1 a_1821_8526.n12 121.124
R345 a_1821_8526.n171 a_1821_8526.t2 116.841
R346 a_1821_8526.n109 a_1821_8526.t6 60.2505
R347 a_1821_8526.n88 a_1821_8526.t9 60.2505
R348 a_1821_8526.n68 a_1821_8526.t7 60.2505
R349 a_1821_8526.n48 a_1821_8526.t8 60.2505
R350 a_1821_8526.n175 a_1821_8526.n174 52.6902
R351 a_1821_8526.n183 a_1821_8526.n182 46.104
R352 a_1821_8526.n199 a_1821_8526.n198 46.104
R353 a_1821_8526.n144 a_1821_8526.n143 39.5177
R354 a_1821_8526.n40 a_1821_8526.n39 39.5177
R355 a_1821_8526.n151 a_1821_8526.n150 32.9315
R356 a_1821_8526.n30 a_1821_8526.n29 32.9315
R357 a_1821_8526.n162 a_1821_8526.n161 29.6384
R358 a_1821_8526.n23 a_1821_8526.n22 29.6384
R359 a_1821_8526.n140 a_1821_8526.t3 27.6955
R360 a_1821_8526.n161 a_1821_8526.n160 26.3453
R361 a_1821_8526.n22 a_1821_8526.n21 26.3453
R362 a_1821_8526.n152 a_1821_8526.n151 23.0522
R363 a_1821_8526.n31 a_1821_8526.n30 23.0522
R364 a_1821_8526.n145 a_1821_8526.n144 16.466
R365 a_1821_8526.n41 a_1821_8526.n40 16.466
R366 a_1821_8526.n138 a_1821_8526.n137 13.177
R367 a_1821_8526.n184 a_1821_8526.n183 9.87981
R368 a_1821_8526.n200 a_1821_8526.n199 9.87981
R369 a_1821_8526.n10 a_1821_8526.n134 9.31646
R370 a_1821_8526.n3 a_1821_8526.n130 9.3005
R371 a_1821_8526.n3 a_1821_8526.n132 9.3005
R372 a_1821_8526.n11 a_1821_8526.n178 9.3005
R373 a_1821_8526.n1 a_1821_8526.n186 9.3005
R374 a_1821_8526.n11 a_1821_8526.n177 9.3005
R375 a_1821_8526.n177 a_1821_8526.n176 9.3005
R376 a_1821_8526.n11 a_1821_8526.n179 9.3005
R377 a_1821_8526.n1 a_1821_8526.n185 9.3005
R378 a_1821_8526.n185 a_1821_8526.n184 9.3005
R379 a_1821_8526.n1 a_1821_8526.n163 9.3005
R380 a_1821_8526.n163 a_1821_8526.n162 9.3005
R381 a_1821_8526.n1 a_1821_8526.n166 9.3005
R382 a_1821_8526.n153 a_1821_8526.n152 9.3005
R383 a_1821_8526.n146 a_1821_8526.n145 9.3005
R384 a_1821_8526.n10 a_1821_8526.n141 9.3005
R385 a_1821_8526.n9 a_1821_8526.n56 9.3005
R386 a_1821_8526.n9 a_1821_8526.n57 9.3005
R387 a_1821_8526.n9 a_1821_8526.n55 9.3005
R388 a_1821_8526.n55 a_1821_8526.n54 9.3005
R389 a_1821_8526.n7 a_1821_8526.n61 9.3005
R390 a_1821_8526.n8 a_1821_8526.n76 9.3005
R391 a_1821_8526.n8 a_1821_8526.n77 9.3005
R392 a_1821_8526.n8 a_1821_8526.n75 9.3005
R393 a_1821_8526.n75 a_1821_8526.n74 9.3005
R394 a_1821_8526.n7 a_1821_8526.n67 9.3005
R395 a_1821_8526.n67 a_1821_8526.n66 9.3005
R396 a_1821_8526.n7 a_1821_8526.n60 9.3005
R397 a_1821_8526.n5 a_1821_8526.n81 9.3005
R398 a_1821_8526.n6 a_1821_8526.n96 9.3005
R399 a_1821_8526.n6 a_1821_8526.n97 9.3005
R400 a_1821_8526.n6 a_1821_8526.n95 9.3005
R401 a_1821_8526.n95 a_1821_8526.n94 9.3005
R402 a_1821_8526.n5 a_1821_8526.n87 9.3005
R403 a_1821_8526.n87 a_1821_8526.n86 9.3005
R404 a_1821_8526.n5 a_1821_8526.n80 9.3005
R405 a_1821_8526.n4 a_1821_8526.n101 9.3005
R406 a_1821_8526.n13 a_1821_8526.n108 9.3005
R407 a_1821_8526.n13 a_1821_8526.n110 9.3005
R408 a_1821_8526.n4 a_1821_8526.n107 9.3005
R409 a_1821_8526.n107 a_1821_8526.n106 9.3005
R410 a_1821_8526.n4 a_1821_8526.n100 9.3005
R411 a_1821_8526.n117 a_1821_8526.n116 9.3005
R412 a_1821_8526.n12 a_1821_8526.n195 9.3005
R413 a_1821_8526.n12 a_1821_8526.n202 9.3005
R414 a_1821_8526.n2 a_1821_8526.n27 9.3005
R415 a_1821_8526.n12 a_1821_8526.n201 9.3005
R416 a_1821_8526.n201 a_1821_8526.n200 9.3005
R417 a_1821_8526.n42 a_1821_8526.n41 9.3005
R418 a_1821_8526.n2 a_1821_8526.n24 9.3005
R419 a_1821_8526.n24 a_1821_8526.n23 9.3005
R420 a_1821_8526.n32 a_1821_8526.n31 9.3005
R421 a_1821_8526.n141 a_1821_8526.n140 9.0206
R422 a_1821_8526.n69 a_1821_8526.n68 8.76429
R423 a_1821_8526.n89 a_1821_8526.n88 8.76429
R424 a_1821_8526.n110 a_1821_8526.n109 8.76429
R425 a_1821_8526.n14 a_1821_8526.t0 7.50197
R426 a_1821_8526.n115 a_1821_8526.n114 7.45411
R427 a_1821_8526.n105 a_1821_8526.n104 7.45411
R428 a_1821_8526.n93 a_1821_8526.n92 7.45411
R429 a_1821_8526.n85 a_1821_8526.n84 7.45411
R430 a_1821_8526.n73 a_1821_8526.n72 7.45411
R431 a_1821_8526.n65 a_1821_8526.n64 7.45411
R432 a_1821_8526.n53 a_1821_8526.n52 7.45411
R433 a_1821_8526.n49 a_1821_8526.n48 6.80105
R434 a_1821_8526.n173 a_1821_8526.n172 6.02403
R435 a_1821_8526.n103 a_1821_8526.n102 5.64756
R436 a_1821_8526.n91 a_1821_8526.n90 5.64756
R437 a_1821_8526.n83 a_1821_8526.n82 5.64756
R438 a_1821_8526.n71 a_1821_8526.n70 5.64756
R439 a_1821_8526.n63 a_1821_8526.n62 5.64756
R440 a_1821_8526.n51 a_1821_8526.n50 5.64756
R441 a_1821_8526.n192 a_1821_8526.t4 5.5395
R442 a_1821_8526.n192 a_1821_8526.t5 5.5395
R443 a_1821_8526.n181 a_1821_8526.n180 5.27109
R444 a_1821_8526.n197 a_1821_8526.n196 5.27109
R445 a_1821_8526.n2 a_1821_8526.n18 5.266
R446 a_1821_8526.n1 a_1821_8526.n159 5.266
R447 a_1821_8526.n4 a_1821_8526.n99 4.73575
R448 a_1821_8526.n6 a_1821_8526.n98 4.73575
R449 a_1821_8526.n5 a_1821_8526.n79 4.73575
R450 a_1821_8526.n8 a_1821_8526.n78 4.73575
R451 a_1821_8526.n7 a_1821_8526.n59 4.73575
R452 a_1821_8526.n9 a_1821_8526.n58 4.73575
R453 a_1821_8526.n7 a_1821_8526.n69 4.6505
R454 a_1821_8526.n5 a_1821_8526.n89 4.6505
R455 a_1821_8526.n15 a_1821_8526.n47 6.76219
R456 a_1821_8526.n191 a_1821_8526.n190 4.51815
R457 a_1821_8526.n170 a_1821_8526.n169 4.51815
R458 a_1821_8526.n37 a_1821_8526.n36 4.51815
R459 a_1821_8526.n3 a_1821_8526.n128 4.5005
R460 a_1821_8526.n1 a_1821_8526.n158 4.5005
R461 a_1821_8526.n1 a_1821_8526.n188 4.5005
R462 a_1821_8526.n10 a_1821_8526.n136 4.5005
R463 a_1821_8526.n10 a_1821_8526.n139 4.5005
R464 a_1821_8526.n13 a_1821_8526.n111 4.5005
R465 a_1821_8526.n112 a_1821_8526.n118 4.5005
R466 a_1821_8526.n3 a_1821_8526.n126 4.5005
R467 a_1821_8526.n3 a_1821_8526.n124 4.5005
R468 a_1821_8526.n1 a_1821_8526.n168 4.5005
R469 a_1821_8526.n1 a_1821_8526.n156 4.5005
R470 a_1821_8526.n1 a_1821_8526.n148 4.5005
R471 a_1821_8526.n2 a_1821_8526.n17 4.5005
R472 a_1821_8526.n2 a_1821_8526.n35 4.5005
R473 a_1821_8526.n2 a_1821_8526.n44 4.5005
R474 a_1821_8526.n12 a_1821_8526.n194 4.5005
R475 a_1821_8526.n2 a_1821_8526.n20 4.5005
R476 a_1821_8526.n11 a_1821_8526.n171 4.23684
R477 a_1821_8526.n148 a_1821_8526.n142 4.14168
R478 a_1821_8526.n118 a_1821_8526.n117 4.14168
R479 a_1821_8526.n44 a_1821_8526.n38 4.14168
R480 a_1821_8526.n47 a_1821_8526.n45 3.76521
R481 a_1821_8526.n9 a_1821_8526.n49 3.42768
R482 a_1821_8526.n124 a_1821_8526.n120 3.38874
R483 a_1821_8526.n156 a_1821_8526.n149 3.38874
R484 a_1821_8526.n35 a_1821_8526.n28 3.38874
R485 a_1821_8526.n132 a_1821_8526.n131 3.38537
R486 a_1821_8526.n176 a_1821_8526.n175 3.2936
R487 a_1821_8526.n0 a_1821_8526.n191 3.03311
R488 a_1821_8526.n1 a_1821_8526.n170 3.03311
R489 a_1821_8526.n2 a_1821_8526.n37 3.03311
R490 a_1821_8526.n165 a_1821_8526.n164 3.01226
R491 a_1821_8526.n26 a_1821_8526.n25 3.01226
R492 a_1821_8526.n3 a_1821_8526.n129 2.57905
R493 a_1821_8526.n123 a_1821_8526.n122 2.25932
R494 a_1821_8526.n155 a_1821_8526.n154 2.25932
R495 a_1821_8526.n118 a_1821_8526.n113 2.25932
R496 a_1821_8526.n34 a_1821_8526.n33 2.25932
R497 a_1821_8526.n15 a_1821_8526.n13 2.25727
R498 a_1821_8526.n15 a_1821_8526.n112 2.29192
R499 a_1821_8526.n189 a_1821_8526.n133 1.90999
R500 a_1821_8526.n147 a_1821_8526.n146 1.88285
R501 a_1821_8526.n166 a_1821_8526.n165 1.88285
R502 a_1821_8526.n47 a_1821_8526.n46 1.88285
R503 a_1821_8526.n43 a_1821_8526.n42 1.88285
R504 a_1821_8526.n27 a_1821_8526.n26 1.88285
R505 a_1821_8526.n0 a_1821_8526.n192 1.72048
R506 a_1821_8526.n133 a_1821_8526.n10 1.67144
R507 a_1821_8526.n128 a_1821_8526.n127 1.50638
R508 a_1821_8526.n158 a_1821_8526.n157 1.50638
R509 a_1821_8526.n20 a_1821_8526.n19 1.50638
R510 a_1821_8526.n14 a_1821_8526.n3 1.28885
R511 a_1821_8526.n14 a_1821_8526.n0 1.22346
R512 a_1821_8526.n185 a_1821_8526.n181 1.12991
R513 a_1821_8526.n201 a_1821_8526.n197 1.12991
R514 a_1821_8526.n189 a_1821_8526.n1 1.07918
R515 a_1821_8526.n116 a_1821_8526.n115 0.994314
R516 a_1821_8526.n106 a_1821_8526.n105 0.994314
R517 a_1821_8526.n94 a_1821_8526.n93 0.994314
R518 a_1821_8526.n86 a_1821_8526.n85 0.994314
R519 a_1821_8526.n74 a_1821_8526.n73 0.994314
R520 a_1821_8526.n66 a_1821_8526.n65 0.994314
R521 a_1821_8526.n54 a_1821_8526.n53 0.994314
R522 a_1821_8526.n126 a_1821_8526.n125 0.753441
R523 a_1821_8526.n188 a_1821_8526.n187 0.753441
R524 a_1821_8526.n168 a_1821_8526.n167 0.753441
R525 a_1821_8526.n107 a_1821_8526.n103 0.753441
R526 a_1821_8526.n95 a_1821_8526.n91 0.753441
R527 a_1821_8526.n87 a_1821_8526.n83 0.753441
R528 a_1821_8526.n75 a_1821_8526.n71 0.753441
R529 a_1821_8526.n67 a_1821_8526.n63 0.753441
R530 a_1821_8526.n55 a_1821_8526.n51 0.753441
R531 a_1821_8526.n194 a_1821_8526.n193 0.753441
R532 a_1821_8526.n17 a_1821_8526.n16 0.753441
R533 a_1821_8526.n12 a_1821_8526.n119 0.737441
R534 a_1821_8526.n119 a_1821_8526.n14 0.718062
R535 a_1821_8526.n1 a_1821_8526.n11 0.676808
R536 a_1821_8526.n7 a_1821_8526.n9 0.6634
R537 a_1821_8526.n5 a_1821_8526.n8 0.6634
R538 a_1821_8526.n4 a_1821_8526.n6 0.6634
R539 a_1821_8526.n12 a_1821_8526.n2 0.631263
R540 a_1821_8526.n8 a_1821_8526.n7 0.585981
R541 a_1821_8526.n6 a_1821_8526.n5 0.585981
R542 a_1821_8526.n14 a_1821_8526.n189 0.511626
R543 a_1821_8526.n13 a_1821_8526.n4 0.447235
R544 a_1821_8526.n119 a_1821_8526.n15 0.389962
R545 a_1821_8526.n124 a_1821_8526.n123 0.376971
R546 a_1821_8526.n122 a_1821_8526.n121 0.376971
R547 a_1821_8526.n177 a_1821_8526.n173 0.376971
R548 a_1821_8526.n148 a_1821_8526.n147 0.376971
R549 a_1821_8526.n156 a_1821_8526.n155 0.376971
R550 a_1821_8526.n154 a_1821_8526.n153 0.376971
R551 a_1821_8526.n136 a_1821_8526.n135 0.376971
R552 a_1821_8526.n139 a_1821_8526.n138 0.376971
R553 a_1821_8526.n44 a_1821_8526.n43 0.376971
R554 a_1821_8526.n35 a_1821_8526.n34 0.376971
R555 a_1821_8526.n33 a_1821_8526.n32 0.376971
R556 VDD.n4014 VDD.n2474 2851.48
R557 VDD.n2494 VDD.n2472 2851.48
R558 VDD.n2492 VDD.n2472 2851.48
R559 VDD.n4014 VDD.n2473 2823.94
R560 VDD.n4197 VDD.n4027 1758.86
R561 VDD.n4197 VDD.n4196 1758.86
R562 VDD.n4024 VDD.n2461 1758.86
R563 VDD.n2461 VDD.n2441 1758.86
R564 VDD.n2345 VDD.t42 840.188
R565 VDD.n2345 VDD.t148 840.188
R566 VDD.n2236 VDD.n2214 784.588
R567 VDD.n2613 VDD.n2609 783.936
R568 VDD.n1732 VDD.n1725 767.823
R569 VDD.n4354 VDD.n2218 737.648
R570 VDD.n1403 VDD.n1374 720.883
R571 VDD.n2622 VDD.n2601 644.766
R572 VDD.n4024 VDD.n2288 609.235
R573 VDD.n3609 VDD.n2638 585
R574 VDD.n2641 VDD.n2639 585
R575 VDD.n2656 VDD.n2655 585
R576 VDD.n3596 VDD.n2647 585
R577 VDD.n3588 VDD.n3587 585
R578 VDD.n2665 VDD.n2662 585
R579 VDD.n2651 VDD.n2650 585
R580 VDD.n2657 VDD.n2646 585
R581 VDD.n2668 VDD.n2667 585
R582 VDD.n3586 VDD.n2661 585
R583 VDD.n3595 VDD.n3594 585
R584 VDD.n3611 VDD.n3610 585
R585 VDD.n3168 VDD.n3095 585
R586 VDD.n3134 VDD.n3131 585
R587 VDD.n3144 VDD.n3143 585
R588 VDD.n3152 VDD.n3120 585
R589 VDD.n3125 VDD.n3124 585
R590 VDD.n3137 VDD.n3136 585
R591 VDD.n3142 VDD.n3130 585
R592 VDD.n3151 VDD.n3150 585
R593 VDD.n3126 VDD.n3119 585
R594 VDD.n3122 VDD.n3104 585
R595 VDD.n3100 VDD.n3096 585
R596 VDD.n3170 VDD.n3169 585
R597 VDD.n3810 VDD.n3805 585
R598 VDD.n3811 VDD.n3810 585
R599 VDD.n3926 VDD.n3925 585
R600 VDD.n3927 VDD.n3926 585
R601 VDD.n3910 VDD.n3909 585
R602 VDD.n3910 VDD.n3672 585
R603 VDD.n3787 VDD.n3786 585
R604 VDD.n3642 VDD.n3640 585
R605 VDD.n3792 VDD.n3791 585
R606 VDD.n3790 VDD.n3765 585
R607 VDD.n3781 VDD.n3780 585
R608 VDD.n3784 VDD.n3768 585
R609 VDD.n2857 VDD.n2856 585
R610 VDD.n2858 VDD.n2857 585
R611 VDD.n3024 VDD.n2875 585
R612 VDD.n2930 VDD.n2929 585
R613 VDD.n2914 VDD.n2912 585
R614 VDD.n2998 VDD.n2997 585
R615 VDD.n2938 VDD.n2937 585
R616 VDD.n2922 VDD.n2921 585
R617 VDD.n2924 VDD.n2923 585
R618 VDD.n2940 VDD.n2939 585
R619 VDD.n2989 VDD.n2951 585
R620 VDD.n2984 VDD.n2956 585
R621 VDD.n2991 VDD.n2990 585
R622 VDD.n2986 VDD.n2985 585
R623 VDD.n2917 VDD.n2915 585
R624 VDD.n77 VDD.n76 585
R625 VDD.n88 VDD.n87 585
R626 VDD.n97 VDD.n96 585
R627 VDD.n86 VDD.n85 585
R628 VDD.n95 VDD.n47 585
R629 VDD.n56 VDD.n54 585
R630 VDD.n67 VDD.n61 585
R631 VDD.n66 VDD.n65 585
R632 VDD.n63 VDD.n60 585
R633 VDD.n78 VDD.n50 585
R634 VDD.n5566 VDD.n5563 585
R635 VDD.n5594 VDD.n5593 585
R636 VDD.n5555 VDD.n5554 585
R637 VDD.n5553 VDD.n5548 585
R638 VDD.n5592 VDD.n5529 585
R639 VDD.n5581 VDD.n5564 585
R640 VDD.n5573 VDD.n5572 585
R641 VDD.n5571 VDD.n5570 585
R642 VDD.n5580 VDD.n5579 585
R643 VDD.n5562 VDD.n5531 585
R644 VDD.n223 VDD.n222 585
R645 VDD.n224 VDD.n179 585
R646 VDD.n233 VDD.n177 585
R647 VDD.n235 VDD.n234 585
R648 VDD.n213 VDD.n207 585
R649 VDD.n212 VDD.n211 585
R650 VDD.n209 VDD.n206 585
R651 VDD.n184 VDD.n182 585
R652 VDD.n196 VDD.n195 585
R653 VDD.n194 VDD.n192 585
R654 VDD.n2505 VDD.n2503 550.754
R655 VDD.n4007 VDD.n2484 550.754
R656 VDD.n2614 VDD.n2613 479.688
R657 VDD.n2614 VDD.n2494 479.688
R658 VDD.n3947 VDD.n3946 456.74
R659 VDD.n4003 VDD.n4001 456.74
R660 VDD.n2343 VDD.t43 403.574
R661 VDD.n2342 VDD.t149 403.574
R662 VDD.n8386 VDD.n8269 373.449
R663 VDD.n8292 VDD.n8266 373.449
R664 VDD.n8839 VDD.n8838 373.449
R665 VDD.n8855 VDD.n8681 373.449
R666 VDD.n7531 VDD.n7414 373.449
R667 VDD.n7437 VDD.n7411 373.449
R668 VDD.n7984 VDD.n7983 373.449
R669 VDD.n8000 VDD.n7826 373.449
R670 VDD.n6677 VDD.n6560 373.449
R671 VDD.n6583 VDD.n6557 373.449
R672 VDD.n7130 VDD.n7129 373.449
R673 VDD.n7146 VDD.n6972 373.449
R674 VDD.n5822 VDD.n5705 373.449
R675 VDD.n5728 VDD.n5702 373.449
R676 VDD.n6275 VDD.n6274 373.449
R677 VDD.n6291 VDD.n6117 373.449
R678 VDD.n4013 VDD.n4012 357.288
R679 VDD.n3988 VDD.n3987 357.288
R680 VDD.n3989 VDD.n3988 357.288
R681 VDD.n4013 VDD.n2475 354.019
R682 VDD.n8768 VDD.n8697 351.829
R683 VDD.n8789 VDD.n8788 351.829
R684 VDD.n8399 VDD.n8288 351.829
R685 VDD.n8401 VDD.n8285 351.829
R686 VDD.n7913 VDD.n7842 351.829
R687 VDD.n7934 VDD.n7933 351.829
R688 VDD.n7544 VDD.n7433 351.829
R689 VDD.n7546 VDD.n7430 351.829
R690 VDD.n7059 VDD.n6988 351.829
R691 VDD.n7080 VDD.n7079 351.829
R692 VDD.n6690 VDD.n6579 351.829
R693 VDD.n6692 VDD.n6576 351.829
R694 VDD.n6204 VDD.n6133 351.829
R695 VDD.n6225 VDD.n6224 351.829
R696 VDD.n5835 VDD.n5724 351.829
R697 VDD.n5837 VDD.n5721 351.829
R698 VDD.n5664 VDD.n5646 321.882
R699 VDD.n5650 VDD.n5645 321.882
R700 VDD.n5627 VDD.n5619 321.882
R701 VDD.n5640 VDD.n5619 321.882
R702 VDD.n5640 VDD.n5617 321.882
R703 VDD.n5669 VDD.n5617 321.882
R704 VDD.n6515 VDD.n6508 321.882
R705 VDD.n6507 VDD.n6469 321.882
R706 VDD.n6487 VDD.n6478 321.882
R707 VDD.n6490 VDD.n6478 321.882
R708 VDD.n6490 VDD.n6471 321.882
R709 VDD.n6503 VDD.n6471 321.882
R710 VDD.n7373 VDD.n7355 321.882
R711 VDD.n7359 VDD.n7354 321.882
R712 VDD.n7336 VDD.n7328 321.882
R713 VDD.n7349 VDD.n7328 321.882
R714 VDD.n7349 VDD.n7326 321.882
R715 VDD.n7378 VDD.n7326 321.882
R716 VDD.n8224 VDD.n8217 321.882
R717 VDD.n8216 VDD.n8178 321.882
R718 VDD.n8196 VDD.n8187 321.882
R719 VDD.n8199 VDD.n8187 321.882
R720 VDD.n8199 VDD.n8180 321.882
R721 VDD.n8212 VDD.n8180 321.882
R722 VDD.n2457 VDD.n2441 300.546
R723 VDD.n2577 VDD.n2518 292.5
R724 VDD.n132 VDD.n121 291.75
R725 VDD.n132 VDD.n131 291.562
R726 VDD.n5668 VDD.n5667 266.731
R727 VDD.n6505 VDD.n6504 266.731
R728 VDD.n7377 VDD.n7376 266.731
R729 VDD.n8214 VDD.n8213 266.731
R730 VDD.n2616 VDD.n2603 247.893
R731 VDD.n2616 VDD.n2473 247.893
R732 VDD.n6524 VDD.t23 240.534
R733 VDD.n8233 VDD.t31 240.534
R734 VDD.n8734 VDD.n8710 239.793
R735 VDD.n8734 VDD.n8733 239.793
R736 VDD.n8724 VDD.n8707 239.793
R737 VDD.n8729 VDD.n8724 239.793
R738 VDD.n8817 VDD.n8715 239.793
R739 VDD.n9010 VDD.n8261 239.793
R740 VDD.n8815 VDD.n8748 239.793
R741 VDD.n9012 VDD.n8257 239.793
R742 VDD.n7879 VDD.n7855 239.793
R743 VDD.n7879 VDD.n7878 239.793
R744 VDD.n7869 VDD.n7852 239.793
R745 VDD.n7874 VDD.n7869 239.793
R746 VDD.n7962 VDD.n7860 239.793
R747 VDD.n8155 VDD.n7406 239.793
R748 VDD.n7960 VDD.n7893 239.793
R749 VDD.n8157 VDD.n7402 239.793
R750 VDD.n7025 VDD.n7001 239.793
R751 VDD.n7025 VDD.n7024 239.793
R752 VDD.n7015 VDD.n6998 239.793
R753 VDD.n7020 VDD.n7015 239.793
R754 VDD.n7108 VDD.n7006 239.793
R755 VDD.n7301 VDD.n6552 239.793
R756 VDD.n7106 VDD.n7039 239.793
R757 VDD.n7303 VDD.n6548 239.793
R758 VDD.n6170 VDD.n6146 239.793
R759 VDD.n6170 VDD.n6169 239.793
R760 VDD.n6160 VDD.n6143 239.793
R761 VDD.n6165 VDD.n6160 239.793
R762 VDD.n6253 VDD.n6151 239.793
R763 VDD.n6446 VDD.n5697 239.793
R764 VDD.n6251 VDD.n6184 239.793
R765 VDD.n6448 VDD.n5693 239.793
R766 VDD.n5657 VDD.t135 239.697
R767 VDD.n7366 VDD.t57 239.697
R768 VDD.n1817 VDD.n1088 232.623
R769 VDD.n3938 VDD.n3937 231.905
R770 VDD.n98 VDD.n46 229.476
R771 VDD.n5556 VDD.n5547 229.476
R772 VDD.n197 VDD.n191 229.476
R773 VDD.n2982 VDD.n2981 228.99
R774 VDD.n1487 VDD.n1374 228
R775 VDD.n1487 VDD.n1365 228
R776 VDD.n1498 VDD.n1365 228
R777 VDD.n1499 VDD.n1498 228
R778 VDD.n1499 VDD.n1359 228
R779 VDD.n1511 VDD.n1359 228
R780 VDD.n1511 VDD.n1352 228
R781 VDD.n1519 VDD.n1352 228
R782 VDD.n1519 VDD.n1346 228
R783 VDD.n1531 VDD.n1346 228
R784 VDD.n1531 VDD.n1337 228
R785 VDD.n1542 VDD.n1337 228
R786 VDD.n1543 VDD.n1542 228
R787 VDD.n1543 VDD.n1331 228
R788 VDD.n1555 VDD.n1331 228
R789 VDD.n1555 VDD.n1324 228
R790 VDD.n1563 VDD.n1324 228
R791 VDD.n1563 VDD.n1314 228
R792 VDD.n1573 VDD.n1314 228
R793 VDD.n1574 VDD.n1573 228
R794 VDD.n1574 VDD.n1308 228
R795 VDD.n1586 VDD.n1308 228
R796 VDD.n1586 VDD.n1301 228
R797 VDD.n1594 VDD.n1301 228
R798 VDD.n1594 VDD.n1295 228
R799 VDD.n1606 VDD.n1295 228
R800 VDD.n1606 VDD.n1286 228
R801 VDD.n1618 VDD.n1286 228
R802 VDD.n1619 VDD.n1618 228
R803 VDD.n1620 VDD.n1619 228
R804 VDD.n1806 VDD.n1620 228
R805 VDD.n1806 VDD.n1621 228
R806 VDD.n1799 VDD.n1621 228
R807 VDD.n1799 VDD.n1629 228
R808 VDD.n1791 VDD.n1629 228
R809 VDD.n1791 VDD.n1636 228
R810 VDD.n1784 VDD.n1636 228
R811 VDD.n1784 VDD.n1646 228
R812 VDD.n1777 VDD.n1646 228
R813 VDD.n1777 VDD.n1652 228
R814 VDD.n1770 VDD.n1652 228
R815 VDD.n1770 VDD.n1662 228
R816 VDD.n1762 VDD.n1662 228
R817 VDD.n1762 VDD.n1669 228
R818 VDD.n1755 VDD.n1669 228
R819 VDD.n1755 VDD.n1679 228
R820 VDD.n1747 VDD.n1679 228
R821 VDD.n1747 VDD.n1686 228
R822 VDD.n1740 VDD.n1686 228
R823 VDD.n1740 VDD.n1696 228
R824 VDD.n1732 VDD.n1696 228
R825 VDD.n1457 VDD.n1456 228
R826 VDD.n1447 VDD.n1446 228
R827 VDD.n1439 VDD.n1438 228
R828 VDD.n1429 VDD.n1428 228
R829 VDD.n1416 VDD.n1386 228
R830 VDD.n1478 VDD.n1029 228
R831 VDD.n1893 VDD.n1029 228
R832 VDD.n1893 VDD.n1007 228
R833 VDD.n4572 VDD.n1007 228
R834 VDD.n4572 VDD.n4571 228
R835 VDD.n4571 VDD.n1008 228
R836 VDD.n4563 VDD.n1008 228
R837 VDD.n4563 VDD.n1020 228
R838 VDD.n4553 VDD.n1020 228
R839 VDD.n4553 VDD.n4552 228
R840 VDD.n4552 VDD.n1913 228
R841 VDD.n4544 VDD.n1913 228
R842 VDD.n4544 VDD.n1925 228
R843 VDD.n4534 VDD.n1925 228
R844 VDD.n4534 VDD.n4533 228
R845 VDD.n4533 VDD.n1944 228
R846 VDD.n4525 VDD.n1944 228
R847 VDD.n4525 VDD.n1955 228
R848 VDD.n4518 VDD.n1955 228
R849 VDD.n4518 VDD.n1965 228
R850 VDD.n4509 VDD.n1965 228
R851 VDD.n4509 VDD.n4508 228
R852 VDD.n4508 VDD.n1982 228
R853 VDD.n4500 VDD.n1982 228
R854 VDD.n4500 VDD.n1997 228
R855 VDD.n4490 VDD.n1997 228
R856 VDD.n4490 VDD.n4489 228
R857 VDD.n4489 VDD.n2017 228
R858 VDD.n4481 VDD.n2017 228
R859 VDD.n4481 VDD.n2030 228
R860 VDD.n4471 VDD.n2030 228
R861 VDD.n4471 VDD.n4470 228
R862 VDD.n4470 VDD.n2049 228
R863 VDD.n4462 VDD.n2049 228
R864 VDD.n4462 VDD.n2059 228
R865 VDD.n4455 VDD.n2059 228
R866 VDD.n4455 VDD.n2067 228
R867 VDD.n4447 VDD.n2067 228
R868 VDD.n4447 VDD.n2077 228
R869 VDD.n4437 VDD.n2077 228
R870 VDD.n4437 VDD.n4436 228
R871 VDD.n4436 VDD.n2102 228
R872 VDD.n4428 VDD.n2102 228
R873 VDD.n4428 VDD.n2114 228
R874 VDD.n4418 VDD.n2114 228
R875 VDD.n4418 VDD.n4417 228
R876 VDD.n4417 VDD.n2132 228
R877 VDD.n4409 VDD.n2132 228
R878 VDD.n4409 VDD.n2145 228
R879 VDD.n4399 VDD.n2145 228
R880 VDD.n4399 VDD.n4398 228
R881 VDD.n4398 VDD.n2164 228
R882 VDD.n4390 VDD.n2164 228
R883 VDD.n4390 VDD.n2176 228
R884 VDD.n4383 VDD.n2176 228
R885 VDD.n4383 VDD.n2186 228
R886 VDD.n4374 VDD.n2186 228
R887 VDD.n4374 VDD.n4373 228
R888 VDD.n4373 VDD.n2203 228
R889 VDD.n4365 VDD.n2203 228
R890 VDD.n4365 VDD.n2218 228
R891 VDD.n2290 VDD.n2236 228
R892 VDD.n1722 VDD.n1721 228
R893 VDD.n1718 VDD.n1717 228
R894 VDD.n1714 VDD.n1713 228
R895 VDD.n1710 VDD.n1709 228
R896 VDD.n1706 VDD.n1036 228
R897 VDD.n1886 VDD.n1033 228
R898 VDD.n1891 VDD.n1033 228
R899 VDD.n1891 VDD.n1034 228
R900 VDD.n1034 VDD.n1013 228
R901 VDD.n4569 VDD.n1013 228
R902 VDD.n4569 VDD.n1014 228
R903 VDD.n4565 VDD.n1014 228
R904 VDD.n4565 VDD.n1017 228
R905 VDD.n1912 VDD.n1017 228
R906 VDD.n4550 VDD.n1912 228
R907 VDD.n4550 VDD.n1918 228
R908 VDD.n4546 VDD.n1918 228
R909 VDD.n4546 VDD.n1921 228
R910 VDD.n1943 VDD.n1921 228
R911 VDD.n4531 VDD.n1943 228
R912 VDD.n4531 VDD.n1949 228
R913 VDD.n4527 VDD.n1949 228
R914 VDD.n4527 VDD.n1952 228
R915 VDD.n1964 VDD.n1952 228
R916 VDD.n1989 VDD.n1964 228
R917 VDD.n1989 VDD.n1981 228
R918 VDD.n4506 VDD.n1981 228
R919 VDD.n4506 VDD.n1987 228
R920 VDD.n4502 VDD.n1987 228
R921 VDD.n4502 VDD.n1993 228
R922 VDD.n2016 VDD.n1993 228
R923 VDD.n4487 VDD.n2016 228
R924 VDD.n4487 VDD.n2023 228
R925 VDD.n4483 VDD.n2023 228
R926 VDD.n4483 VDD.n2026 228
R927 VDD.n2048 VDD.n2026 228
R928 VDD.n4468 VDD.n2048 228
R929 VDD.n4468 VDD.n2053 228
R930 VDD.n4464 VDD.n2053 228
R931 VDD.n4464 VDD.n2056 228
R932 VDD.n4453 VDD.n2056 228
R933 VDD.n4453 VDD.n2071 228
R934 VDD.n4449 VDD.n2071 228
R935 VDD.n4449 VDD.n2073 228
R936 VDD.n2101 VDD.n2073 228
R937 VDD.n4434 VDD.n2101 228
R938 VDD.n4434 VDD.n2107 228
R939 VDD.n4430 VDD.n2107 228
R940 VDD.n4430 VDD.n2110 228
R941 VDD.n2131 VDD.n2110 228
R942 VDD.n4415 VDD.n2131 228
R943 VDD.n4415 VDD.n2138 228
R944 VDD.n4411 VDD.n2138 228
R945 VDD.n4411 VDD.n2141 228
R946 VDD.n2163 VDD.n2141 228
R947 VDD.n4396 VDD.n2163 228
R948 VDD.n4396 VDD.n2169 228
R949 VDD.n4392 VDD.n2169 228
R950 VDD.n4392 VDD.n2172 228
R951 VDD.n2185 VDD.n2172 228
R952 VDD.n2210 VDD.n2185 228
R953 VDD.n2210 VDD.n2202 228
R954 VDD.n4371 VDD.n2202 228
R955 VDD.n4371 VDD.n2208 228
R956 VDD.n4367 VDD.n2208 228
R957 VDD.n4367 VDD.n2214 228
R958 VDD.n2460 VDD.n2459 220.383
R959 VDD.n8715 VDD.n8714 218.173
R960 VDD.n8291 VDD.n8261 218.173
R961 VDD.n8794 VDD.n8748 218.173
R962 VDD.n8391 VDD.n8257 218.173
R963 VDD.n7860 VDD.n7859 218.173
R964 VDD.n7436 VDD.n7406 218.173
R965 VDD.n7939 VDD.n7893 218.173
R966 VDD.n7536 VDD.n7402 218.173
R967 VDD.n7006 VDD.n7005 218.173
R968 VDD.n6582 VDD.n6552 218.173
R969 VDD.n7085 VDD.n7039 218.173
R970 VDD.n6682 VDD.n6548 218.173
R971 VDD.n6151 VDD.n6150 218.173
R972 VDD.n5727 VDD.n5697 218.173
R973 VDD.n6230 VDD.n6184 218.173
R974 VDD.n5827 VDD.n5693 218.173
R975 VDD.n5666 VDD.t134 217.947
R976 VDD.n6517 VDD.t22 217.947
R977 VDD.n7375 VDD.t56 217.947
R978 VDD.n8226 VDD.t30 217.947
R979 VDD.n2460 VDD.n2340 213.983
R980 VDD.n8570 VDD.n8540 205.079
R981 VDD.n8570 VDD.n8569 205.079
R982 VDD.n8569 VDD.n8568 205.079
R983 VDD.n8568 VDD.n8541 205.079
R984 VDD.n8562 VDD.n8541 205.079
R985 VDD.n8562 VDD.n8561 205.079
R986 VDD.n8561 VDD.n8560 205.079
R987 VDD.n8560 VDD.n8545 205.079
R988 VDD.n8554 VDD.n8545 205.079
R989 VDD.n8554 VDD.n8553 205.079
R990 VDD.n8553 VDD.n8552 205.079
R991 VDD.n8552 VDD.n8277 205.079
R992 VDD.n8995 VDD.n8277 205.079
R993 VDD.n8649 VDD.n8498 205.079
R994 VDD.n8655 VDD.n8498 205.079
R995 VDD.n8656 VDD.n8655 205.079
R996 VDD.n8657 VDD.n8656 205.079
R997 VDD.n8657 VDD.n8494 205.079
R998 VDD.n8663 VDD.n8494 205.079
R999 VDD.n8664 VDD.n8663 205.079
R1000 VDD.n8665 VDD.n8664 205.079
R1001 VDD.n8665 VDD.n8490 205.079
R1002 VDD.n8671 VDD.n8490 205.079
R1003 VDD.n8672 VDD.n8671 205.079
R1004 VDD.n8674 VDD.n8672 205.079
R1005 VDD.n8674 VDD.n8673 205.079
R1006 VDD.n8993 VDD.n8279 205.079
R1007 VDD.n8987 VDD.n8279 205.079
R1008 VDD.n8987 VDD.n8986 205.079
R1009 VDD.n8986 VDD.n8985 205.079
R1010 VDD.n8985 VDD.n8407 205.079
R1011 VDD.n8979 VDD.n8407 205.079
R1012 VDD.n8979 VDD.n8978 205.079
R1013 VDD.n8978 VDD.n8977 205.079
R1014 VDD.n8977 VDD.n8411 205.079
R1015 VDD.n8971 VDD.n8411 205.079
R1016 VDD.n8971 VDD.n8970 205.079
R1017 VDD.n8970 VDD.n8969 205.079
R1018 VDD.n8969 VDD.n8415 205.079
R1019 VDD.n8871 VDD.n8464 205.079
R1020 VDD.n8872 VDD.n8871 205.079
R1021 VDD.n8873 VDD.n8872 205.079
R1022 VDD.n8873 VDD.n8460 205.079
R1023 VDD.n8879 VDD.n8460 205.079
R1024 VDD.n8880 VDD.n8879 205.079
R1025 VDD.n8881 VDD.n8880 205.079
R1026 VDD.n8881 VDD.n8456 205.079
R1027 VDD.n8887 VDD.n8456 205.079
R1028 VDD.n8888 VDD.n8887 205.079
R1029 VDD.n8889 VDD.n8888 205.079
R1030 VDD.n8889 VDD.n8451 205.079
R1031 VDD.n8896 VDD.n8451 205.079
R1032 VDD.n7715 VDD.n7685 205.079
R1033 VDD.n7715 VDD.n7714 205.079
R1034 VDD.n7714 VDD.n7713 205.079
R1035 VDD.n7713 VDD.n7686 205.079
R1036 VDD.n7707 VDD.n7686 205.079
R1037 VDD.n7707 VDD.n7706 205.079
R1038 VDD.n7706 VDD.n7705 205.079
R1039 VDD.n7705 VDD.n7690 205.079
R1040 VDD.n7699 VDD.n7690 205.079
R1041 VDD.n7699 VDD.n7698 205.079
R1042 VDD.n7698 VDD.n7697 205.079
R1043 VDD.n7697 VDD.n7422 205.079
R1044 VDD.n8140 VDD.n7422 205.079
R1045 VDD.n7794 VDD.n7643 205.079
R1046 VDD.n7800 VDD.n7643 205.079
R1047 VDD.n7801 VDD.n7800 205.079
R1048 VDD.n7802 VDD.n7801 205.079
R1049 VDD.n7802 VDD.n7639 205.079
R1050 VDD.n7808 VDD.n7639 205.079
R1051 VDD.n7809 VDD.n7808 205.079
R1052 VDD.n7810 VDD.n7809 205.079
R1053 VDD.n7810 VDD.n7635 205.079
R1054 VDD.n7816 VDD.n7635 205.079
R1055 VDD.n7817 VDD.n7816 205.079
R1056 VDD.n7819 VDD.n7817 205.079
R1057 VDD.n7819 VDD.n7818 205.079
R1058 VDD.n8138 VDD.n7424 205.079
R1059 VDD.n8132 VDD.n7424 205.079
R1060 VDD.n8132 VDD.n8131 205.079
R1061 VDD.n8131 VDD.n8130 205.079
R1062 VDD.n8130 VDD.n7552 205.079
R1063 VDD.n8124 VDD.n7552 205.079
R1064 VDD.n8124 VDD.n8123 205.079
R1065 VDD.n8123 VDD.n8122 205.079
R1066 VDD.n8122 VDD.n7556 205.079
R1067 VDD.n8116 VDD.n7556 205.079
R1068 VDD.n8116 VDD.n8115 205.079
R1069 VDD.n8115 VDD.n8114 205.079
R1070 VDD.n8114 VDD.n7560 205.079
R1071 VDD.n8016 VDD.n7609 205.079
R1072 VDD.n8017 VDD.n8016 205.079
R1073 VDD.n8018 VDD.n8017 205.079
R1074 VDD.n8018 VDD.n7605 205.079
R1075 VDD.n8024 VDD.n7605 205.079
R1076 VDD.n8025 VDD.n8024 205.079
R1077 VDD.n8026 VDD.n8025 205.079
R1078 VDD.n8026 VDD.n7601 205.079
R1079 VDD.n8032 VDD.n7601 205.079
R1080 VDD.n8033 VDD.n8032 205.079
R1081 VDD.n8034 VDD.n8033 205.079
R1082 VDD.n8034 VDD.n7596 205.079
R1083 VDD.n8041 VDD.n7596 205.079
R1084 VDD.n6861 VDD.n6831 205.079
R1085 VDD.n6861 VDD.n6860 205.079
R1086 VDD.n6860 VDD.n6859 205.079
R1087 VDD.n6859 VDD.n6832 205.079
R1088 VDD.n6853 VDD.n6832 205.079
R1089 VDD.n6853 VDD.n6852 205.079
R1090 VDD.n6852 VDD.n6851 205.079
R1091 VDD.n6851 VDD.n6836 205.079
R1092 VDD.n6845 VDD.n6836 205.079
R1093 VDD.n6845 VDD.n6844 205.079
R1094 VDD.n6844 VDD.n6843 205.079
R1095 VDD.n6843 VDD.n6568 205.079
R1096 VDD.n7286 VDD.n6568 205.079
R1097 VDD.n6940 VDD.n6789 205.079
R1098 VDD.n6946 VDD.n6789 205.079
R1099 VDD.n6947 VDD.n6946 205.079
R1100 VDD.n6948 VDD.n6947 205.079
R1101 VDD.n6948 VDD.n6785 205.079
R1102 VDD.n6954 VDD.n6785 205.079
R1103 VDD.n6955 VDD.n6954 205.079
R1104 VDD.n6956 VDD.n6955 205.079
R1105 VDD.n6956 VDD.n6781 205.079
R1106 VDD.n6962 VDD.n6781 205.079
R1107 VDD.n6963 VDD.n6962 205.079
R1108 VDD.n6965 VDD.n6963 205.079
R1109 VDD.n6965 VDD.n6964 205.079
R1110 VDD.n7284 VDD.n6570 205.079
R1111 VDD.n7278 VDD.n6570 205.079
R1112 VDD.n7278 VDD.n7277 205.079
R1113 VDD.n7277 VDD.n7276 205.079
R1114 VDD.n7276 VDD.n6698 205.079
R1115 VDD.n7270 VDD.n6698 205.079
R1116 VDD.n7270 VDD.n7269 205.079
R1117 VDD.n7269 VDD.n7268 205.079
R1118 VDD.n7268 VDD.n6702 205.079
R1119 VDD.n7262 VDD.n6702 205.079
R1120 VDD.n7262 VDD.n7261 205.079
R1121 VDD.n7261 VDD.n7260 205.079
R1122 VDD.n7260 VDD.n6706 205.079
R1123 VDD.n7162 VDD.n6755 205.079
R1124 VDD.n7163 VDD.n7162 205.079
R1125 VDD.n7164 VDD.n7163 205.079
R1126 VDD.n7164 VDD.n6751 205.079
R1127 VDD.n7170 VDD.n6751 205.079
R1128 VDD.n7171 VDD.n7170 205.079
R1129 VDD.n7172 VDD.n7171 205.079
R1130 VDD.n7172 VDD.n6747 205.079
R1131 VDD.n7178 VDD.n6747 205.079
R1132 VDD.n7179 VDD.n7178 205.079
R1133 VDD.n7180 VDD.n7179 205.079
R1134 VDD.n7180 VDD.n6742 205.079
R1135 VDD.n7187 VDD.n6742 205.079
R1136 VDD.n6006 VDD.n5976 205.079
R1137 VDD.n6006 VDD.n6005 205.079
R1138 VDD.n6005 VDD.n6004 205.079
R1139 VDD.n6004 VDD.n5977 205.079
R1140 VDD.n5998 VDD.n5977 205.079
R1141 VDD.n5998 VDD.n5997 205.079
R1142 VDD.n5997 VDD.n5996 205.079
R1143 VDD.n5996 VDD.n5981 205.079
R1144 VDD.n5990 VDD.n5981 205.079
R1145 VDD.n5990 VDD.n5989 205.079
R1146 VDD.n5989 VDD.n5988 205.079
R1147 VDD.n5988 VDD.n5713 205.079
R1148 VDD.n6431 VDD.n5713 205.079
R1149 VDD.n6085 VDD.n5934 205.079
R1150 VDD.n6091 VDD.n5934 205.079
R1151 VDD.n6092 VDD.n6091 205.079
R1152 VDD.n6093 VDD.n6092 205.079
R1153 VDD.n6093 VDD.n5930 205.079
R1154 VDD.n6099 VDD.n5930 205.079
R1155 VDD.n6100 VDD.n6099 205.079
R1156 VDD.n6101 VDD.n6100 205.079
R1157 VDD.n6101 VDD.n5926 205.079
R1158 VDD.n6107 VDD.n5926 205.079
R1159 VDD.n6108 VDD.n6107 205.079
R1160 VDD.n6110 VDD.n6108 205.079
R1161 VDD.n6110 VDD.n6109 205.079
R1162 VDD.n6429 VDD.n5715 205.079
R1163 VDD.n6423 VDD.n5715 205.079
R1164 VDD.n6423 VDD.n6422 205.079
R1165 VDD.n6422 VDD.n6421 205.079
R1166 VDD.n6421 VDD.n5843 205.079
R1167 VDD.n6415 VDD.n5843 205.079
R1168 VDD.n6415 VDD.n6414 205.079
R1169 VDD.n6414 VDD.n6413 205.079
R1170 VDD.n6413 VDD.n5847 205.079
R1171 VDD.n6407 VDD.n5847 205.079
R1172 VDD.n6407 VDD.n6406 205.079
R1173 VDD.n6406 VDD.n6405 205.079
R1174 VDD.n6405 VDD.n5851 205.079
R1175 VDD.n6307 VDD.n5900 205.079
R1176 VDD.n6308 VDD.n6307 205.079
R1177 VDD.n6309 VDD.n6308 205.079
R1178 VDD.n6309 VDD.n5896 205.079
R1179 VDD.n6315 VDD.n5896 205.079
R1180 VDD.n6316 VDD.n6315 205.079
R1181 VDD.n6317 VDD.n6316 205.079
R1182 VDD.n6317 VDD.n5892 205.079
R1183 VDD.n6323 VDD.n5892 205.079
R1184 VDD.n6324 VDD.n6323 205.079
R1185 VDD.n6325 VDD.n6324 205.079
R1186 VDD.n6325 VDD.n5887 205.079
R1187 VDD.n6332 VDD.n5887 205.079
R1188 VDD.n5363 VDD.n5362 205.079
R1189 VDD.n5362 VDD.n5361 205.079
R1190 VDD.n5361 VDD.n330 205.079
R1191 VDD.n5352 VDD.n330 205.079
R1192 VDD.n5352 VDD.n5351 205.079
R1193 VDD.n5351 VDD.n5350 205.079
R1194 VDD.n5350 VDD.n339 205.079
R1195 VDD.n5341 VDD.n339 205.079
R1196 VDD.n5341 VDD.n5340 205.079
R1197 VDD.n5340 VDD.n5339 205.079
R1198 VDD.n5339 VDD.n346 205.079
R1199 VDD.n5330 VDD.n346 205.079
R1200 VDD.n5330 VDD.n5329 205.079
R1201 VDD.n5329 VDD.n5328 205.079
R1202 VDD.n5328 VDD.n355 205.079
R1203 VDD.n5319 VDD.n355 205.079
R1204 VDD.n5319 VDD.n5318 205.079
R1205 VDD.n5318 VDD.n5317 205.079
R1206 VDD.n5317 VDD.n364 205.079
R1207 VDD.n5308 VDD.n364 205.079
R1208 VDD.n5308 VDD.n5307 205.079
R1209 VDD.n5307 VDD.n5306 205.079
R1210 VDD.n5306 VDD.n373 205.079
R1211 VDD.n384 VDD.n373 205.079
R1212 VDD.n5297 VDD.n384 205.079
R1213 VDD.n5297 VDD.n5296 205.079
R1214 VDD.n5296 VDD.n5295 205.079
R1215 VDD.n5295 VDD.n385 205.079
R1216 VDD.n5286 VDD.n385 205.079
R1217 VDD.n5284 VDD.n396 205.079
R1218 VDD.n5275 VDD.n396 205.079
R1219 VDD.n5275 VDD.n5274 205.079
R1220 VDD.n5274 VDD.n5273 205.079
R1221 VDD.n5273 VDD.n586 205.079
R1222 VDD.n597 VDD.n586 205.079
R1223 VDD.n5264 VDD.n597 205.079
R1224 VDD.n5264 VDD.n5263 205.079
R1225 VDD.n5263 VDD.n5262 205.079
R1226 VDD.n5262 VDD.n598 205.079
R1227 VDD.n5253 VDD.n598 205.079
R1228 VDD.n5253 VDD.n5252 205.079
R1229 VDD.n5252 VDD.n5251 205.079
R1230 VDD.n5251 VDD.n607 205.079
R1231 VDD.n5242 VDD.n607 205.079
R1232 VDD.n5242 VDD.n5241 205.079
R1233 VDD.n5241 VDD.n5240 205.079
R1234 VDD.n5240 VDD.n616 205.079
R1235 VDD.n5231 VDD.n616 205.079
R1236 VDD.n5231 VDD.n5230 205.079
R1237 VDD.n5230 VDD.n5229 205.079
R1238 VDD.n5229 VDD.n625 205.079
R1239 VDD.n5220 VDD.n625 205.079
R1240 VDD.n5220 VDD.n5219 205.079
R1241 VDD.n5219 VDD.n5218 205.079
R1242 VDD.n5218 VDD.n634 205.079
R1243 VDD.n5209 VDD.n634 205.079
R1244 VDD.n5209 VDD.n5208 205.079
R1245 VDD.n5208 VDD.n5207 205.079
R1246 VDD.n5207 VDD.n641 205.079
R1247 VDD.n5198 VDD.n641 205.079
R1248 VDD.n5198 VDD.n5197 205.079
R1249 VDD.n5197 VDD.n5196 205.079
R1250 VDD.n5196 VDD.n650 205.079
R1251 VDD.n5187 VDD.n650 205.079
R1252 VDD.n5187 VDD.n5186 205.079
R1253 VDD.n5186 VDD.n5185 205.079
R1254 VDD.n5185 VDD.n659 205.079
R1255 VDD.n5176 VDD.n659 205.079
R1256 VDD.n5176 VDD.n5175 205.079
R1257 VDD.n5175 VDD.n5174 205.079
R1258 VDD.n5174 VDD.n668 205.079
R1259 VDD.n678 VDD.n668 205.079
R1260 VDD.n5164 VDD.n678 205.079
R1261 VDD.n4718 VDD.n4717 205.079
R1262 VDD.n4717 VDD.n913 205.079
R1263 VDD.n4731 VDD.n913 205.079
R1264 VDD.n4732 VDD.n4731 205.079
R1265 VDD.n4733 VDD.n4732 205.079
R1266 VDD.n4733 VDD.n906 205.079
R1267 VDD.n4744 VDD.n906 205.079
R1268 VDD.n4745 VDD.n4744 205.079
R1269 VDD.n4746 VDD.n4745 205.079
R1270 VDD.n4746 VDD.n899 205.079
R1271 VDD.n4755 VDD.n899 205.079
R1272 VDD.n4756 VDD.n4755 205.079
R1273 VDD.n4757 VDD.n4756 205.079
R1274 VDD.n4757 VDD.n892 205.079
R1275 VDD.n4768 VDD.n892 205.079
R1276 VDD.n4769 VDD.n4768 205.079
R1277 VDD.n4770 VDD.n4769 205.079
R1278 VDD.n4770 VDD.n885 205.079
R1279 VDD.n4781 VDD.n885 205.079
R1280 VDD.n4782 VDD.n4781 205.079
R1281 VDD.n4783 VDD.n4782 205.079
R1282 VDD.n4783 VDD.n878 205.079
R1283 VDD.n4794 VDD.n878 205.079
R1284 VDD.n4795 VDD.n4794 205.079
R1285 VDD.n4796 VDD.n4795 205.079
R1286 VDD.n4796 VDD.n872 205.079
R1287 VDD.n4806 VDD.n872 205.079
R1288 VDD.n4807 VDD.n4806 205.079
R1289 VDD.n4808 VDD.n4807 205.079
R1290 VDD.n4808 VDD.n865 205.079
R1291 VDD.n4819 VDD.n865 205.079
R1292 VDD.n4820 VDD.n4819 205.079
R1293 VDD.n4821 VDD.n4820 205.079
R1294 VDD.n4821 VDD.n858 205.079
R1295 VDD.n4832 VDD.n858 205.079
R1296 VDD.n4833 VDD.n4832 205.079
R1297 VDD.n4834 VDD.n4833 205.079
R1298 VDD.n4834 VDD.n851 205.079
R1299 VDD.n4845 VDD.n851 205.079
R1300 VDD.n4846 VDD.n4845 205.079
R1301 VDD.n4847 VDD.n4846 205.079
R1302 VDD.n4847 VDD.n844 205.079
R1303 VDD.n4858 VDD.n844 205.079
R1304 VDD.n4859 VDD.n4858 205.079
R1305 VDD.n4860 VDD.n4859 205.079
R1306 VDD.n4860 VDD.n837 205.079
R1307 VDD.n4869 VDD.n837 205.079
R1308 VDD.n4870 VDD.n4869 205.079
R1309 VDD.n4871 VDD.n4870 205.079
R1310 VDD.n4871 VDD.n830 205.079
R1311 VDD.n4882 VDD.n830 205.079
R1312 VDD.n4883 VDD.n4882 205.079
R1313 VDD.n4884 VDD.n4883 205.079
R1314 VDD.n4884 VDD.n823 205.079
R1315 VDD.n4895 VDD.n823 205.079
R1316 VDD.n4896 VDD.n4895 205.079
R1317 VDD.n4897 VDD.n4896 205.079
R1318 VDD.n4897 VDD.n816 205.079
R1319 VDD.n4908 VDD.n816 205.079
R1320 VDD.n4909 VDD.n4908 205.079
R1321 VDD.n4910 VDD.n4909 205.079
R1322 VDD.n4910 VDD.n810 205.079
R1323 VDD.n4920 VDD.n810 205.079
R1324 VDD.n4921 VDD.n4920 205.079
R1325 VDD.n4922 VDD.n4921 205.079
R1326 VDD.n4922 VDD.n803 205.079
R1327 VDD.n4933 VDD.n803 205.079
R1328 VDD.n4934 VDD.n4933 205.079
R1329 VDD.n4935 VDD.n4934 205.079
R1330 VDD.n4935 VDD.n796 205.079
R1331 VDD.n4946 VDD.n796 205.079
R1332 VDD.n4947 VDD.n4946 205.079
R1333 VDD.n4948 VDD.n4947 205.079
R1334 VDD.n4948 VDD.n789 205.079
R1335 VDD.n4959 VDD.n789 205.079
R1336 VDD.n4960 VDD.n4959 205.079
R1337 VDD.n4961 VDD.n4960 205.079
R1338 VDD.n4961 VDD.n782 205.079
R1339 VDD.n4972 VDD.n782 205.079
R1340 VDD.n4973 VDD.n4972 205.079
R1341 VDD.n4974 VDD.n4973 205.079
R1342 VDD.n4974 VDD.n775 205.079
R1343 VDD.n4983 VDD.n775 205.079
R1344 VDD.n4984 VDD.n4983 205.079
R1345 VDD.n4985 VDD.n4984 205.079
R1346 VDD.n4985 VDD.n768 205.079
R1347 VDD.n4996 VDD.n768 205.079
R1348 VDD.n4997 VDD.n4996 205.079
R1349 VDD.n4998 VDD.n4997 205.079
R1350 VDD.n4998 VDD.n761 205.079
R1351 VDD.n5009 VDD.n761 205.079
R1352 VDD.n5010 VDD.n5009 205.079
R1353 VDD.n5011 VDD.n5010 205.079
R1354 VDD.n5011 VDD.n754 205.079
R1355 VDD.n5022 VDD.n754 205.079
R1356 VDD.n5023 VDD.n5022 205.079
R1357 VDD.n5024 VDD.n5023 205.079
R1358 VDD.n5024 VDD.n748 205.079
R1359 VDD.n5034 VDD.n748 205.079
R1360 VDD.n5035 VDD.n5034 205.079
R1361 VDD.n5036 VDD.n5035 205.079
R1362 VDD.n5036 VDD.n741 205.079
R1363 VDD.n5047 VDD.n741 205.079
R1364 VDD.n5048 VDD.n5047 205.079
R1365 VDD.n5049 VDD.n5048 205.079
R1366 VDD.n5049 VDD.n734 205.079
R1367 VDD.n5060 VDD.n734 205.079
R1368 VDD.n5061 VDD.n5060 205.079
R1369 VDD.n5062 VDD.n5061 205.079
R1370 VDD.n5062 VDD.n727 205.079
R1371 VDD.n5073 VDD.n727 205.079
R1372 VDD.n5074 VDD.n5073 205.079
R1373 VDD.n5075 VDD.n5074 205.079
R1374 VDD.n5075 VDD.n720 205.079
R1375 VDD.n5086 VDD.n720 205.079
R1376 VDD.n5087 VDD.n5086 205.079
R1377 VDD.n5088 VDD.n5087 205.079
R1378 VDD.n5088 VDD.n713 205.079
R1379 VDD.n5097 VDD.n713 205.079
R1380 VDD.n5098 VDD.n5097 205.079
R1381 VDD.n5099 VDD.n5098 205.079
R1382 VDD.n5099 VDD.n706 205.079
R1383 VDD.n5110 VDD.n706 205.079
R1384 VDD.n5111 VDD.n5110 205.079
R1385 VDD.n5112 VDD.n5111 205.079
R1386 VDD.n5112 VDD.n699 205.079
R1387 VDD.n5123 VDD.n699 205.079
R1388 VDD.n5124 VDD.n5123 205.079
R1389 VDD.n5125 VDD.n5124 205.079
R1390 VDD.n5125 VDD.n692 205.079
R1391 VDD.n5136 VDD.n692 205.079
R1392 VDD.n5137 VDD.n5136 205.079
R1393 VDD.n5138 VDD.n5137 205.079
R1394 VDD.n5138 VDD.n686 205.079
R1395 VDD.n5148 VDD.n686 205.079
R1396 VDD.n5149 VDD.n5148 205.079
R1397 VDD.n5151 VDD.n5149 205.079
R1398 VDD.n5151 VDD.n5150 205.079
R1399 VDD.n5150 VDD.n679 205.079
R1400 VDD.n4579 VDD.n4578 205.079
R1401 VDD.n4579 VDD.n994 205.079
R1402 VDD.n4590 VDD.n994 205.079
R1403 VDD.n4591 VDD.n4590 205.079
R1404 VDD.n4592 VDD.n4591 205.079
R1405 VDD.n4592 VDD.n988 205.079
R1406 VDD.n4602 VDD.n988 205.079
R1407 VDD.n4603 VDD.n4602 205.079
R1408 VDD.n4604 VDD.n4603 205.079
R1409 VDD.n4604 VDD.n980 205.079
R1410 VDD.n4613 VDD.n980 205.079
R1411 VDD.n4614 VDD.n4613 205.079
R1412 VDD.n4615 VDD.n4614 205.079
R1413 VDD.n4615 VDD.n973 205.079
R1414 VDD.n4626 VDD.n973 205.079
R1415 VDD.n4627 VDD.n4626 205.079
R1416 VDD.n4628 VDD.n4627 205.079
R1417 VDD.n4628 VDD.n966 205.079
R1418 VDD.n4639 VDD.n966 205.079
R1419 VDD.n4640 VDD.n4639 205.079
R1420 VDD.n4641 VDD.n4640 205.079
R1421 VDD.n4641 VDD.n959 205.079
R1422 VDD.n4652 VDD.n959 205.079
R1423 VDD.n4653 VDD.n4652 205.079
R1424 VDD.n4654 VDD.n4653 205.079
R1425 VDD.n4654 VDD.n952 205.079
R1426 VDD.n4662 VDD.n952 205.079
R1427 VDD.n4663 VDD.n4662 205.079
R1428 VDD.n4664 VDD.n4663 205.079
R1429 VDD.n4664 VDD.n945 205.079
R1430 VDD.n4675 VDD.n945 205.079
R1431 VDD.n4676 VDD.n4675 205.079
R1432 VDD.n4677 VDD.n4676 205.079
R1433 VDD.n4677 VDD.n938 205.079
R1434 VDD.n4688 VDD.n938 205.079
R1435 VDD.n4689 VDD.n4688 205.079
R1436 VDD.n4690 VDD.n4689 205.079
R1437 VDD.n4690 VDD.n931 205.079
R1438 VDD.n4701 VDD.n931 205.079
R1439 VDD.n4702 VDD.n4701 205.079
R1440 VDD.n4703 VDD.n4702 205.079
R1441 VDD.n4703 VDD.n922 205.079
R1442 VDD.n4714 VDD.n922 205.079
R1443 VDD.n8904 VDD.n8446 203.786
R1444 VDD.n8905 VDD.n8904 203.786
R1445 VDD.n8906 VDD.n8905 203.786
R1446 VDD.n8906 VDD.n8442 203.786
R1447 VDD.n8912 VDD.n8442 203.786
R1448 VDD.n8913 VDD.n8912 203.786
R1449 VDD.n8914 VDD.n8913 203.786
R1450 VDD.n8914 VDD.n8438 203.786
R1451 VDD.n8920 VDD.n8438 203.786
R1452 VDD.n8921 VDD.n8920 203.786
R1453 VDD.n8922 VDD.n8921 203.786
R1454 VDD.n8922 VDD.n8434 203.786
R1455 VDD.n8928 VDD.n8434 203.786
R1456 VDD.n8929 VDD.n8928 203.786
R1457 VDD.n8930 VDD.n8929 203.786
R1458 VDD.n8930 VDD.n8430 203.786
R1459 VDD.n8936 VDD.n8430 203.786
R1460 VDD.n8937 VDD.n8936 203.786
R1461 VDD.n8938 VDD.n8937 203.786
R1462 VDD.n8938 VDD.n8426 203.786
R1463 VDD.n8944 VDD.n8426 203.786
R1464 VDD.n8945 VDD.n8944 203.786
R1465 VDD.n8946 VDD.n8945 203.786
R1466 VDD.n8946 VDD.n8422 203.786
R1467 VDD.n8952 VDD.n8422 203.786
R1468 VDD.n8953 VDD.n8952 203.786
R1469 VDD.n8956 VDD.n8953 203.786
R1470 VDD.n8956 VDD.n8955 203.786
R1471 VDD.n8049 VDD.n7591 203.786
R1472 VDD.n8050 VDD.n8049 203.786
R1473 VDD.n8051 VDD.n8050 203.786
R1474 VDD.n8051 VDD.n7587 203.786
R1475 VDD.n8057 VDD.n7587 203.786
R1476 VDD.n8058 VDD.n8057 203.786
R1477 VDD.n8059 VDD.n8058 203.786
R1478 VDD.n8059 VDD.n7583 203.786
R1479 VDD.n8065 VDD.n7583 203.786
R1480 VDD.n8066 VDD.n8065 203.786
R1481 VDD.n8067 VDD.n8066 203.786
R1482 VDD.n8067 VDD.n7579 203.786
R1483 VDD.n8073 VDD.n7579 203.786
R1484 VDD.n8074 VDD.n8073 203.786
R1485 VDD.n8075 VDD.n8074 203.786
R1486 VDD.n8075 VDD.n7575 203.786
R1487 VDD.n8081 VDD.n7575 203.786
R1488 VDD.n8082 VDD.n8081 203.786
R1489 VDD.n8083 VDD.n8082 203.786
R1490 VDD.n8083 VDD.n7571 203.786
R1491 VDD.n8089 VDD.n7571 203.786
R1492 VDD.n8090 VDD.n8089 203.786
R1493 VDD.n8091 VDD.n8090 203.786
R1494 VDD.n8091 VDD.n7567 203.786
R1495 VDD.n8097 VDD.n7567 203.786
R1496 VDD.n8098 VDD.n8097 203.786
R1497 VDD.n8101 VDD.n8098 203.786
R1498 VDD.n8101 VDD.n8100 203.786
R1499 VDD.n7195 VDD.n6737 203.786
R1500 VDD.n7196 VDD.n7195 203.786
R1501 VDD.n7197 VDD.n7196 203.786
R1502 VDD.n7197 VDD.n6733 203.786
R1503 VDD.n7203 VDD.n6733 203.786
R1504 VDD.n7204 VDD.n7203 203.786
R1505 VDD.n7205 VDD.n7204 203.786
R1506 VDD.n7205 VDD.n6729 203.786
R1507 VDD.n7211 VDD.n6729 203.786
R1508 VDD.n7212 VDD.n7211 203.786
R1509 VDD.n7213 VDD.n7212 203.786
R1510 VDD.n7213 VDD.n6725 203.786
R1511 VDD.n7219 VDD.n6725 203.786
R1512 VDD.n7220 VDD.n7219 203.786
R1513 VDD.n7221 VDD.n7220 203.786
R1514 VDD.n7221 VDD.n6721 203.786
R1515 VDD.n7227 VDD.n6721 203.786
R1516 VDD.n7228 VDD.n7227 203.786
R1517 VDD.n7229 VDD.n7228 203.786
R1518 VDD.n7229 VDD.n6717 203.786
R1519 VDD.n7235 VDD.n6717 203.786
R1520 VDD.n7236 VDD.n7235 203.786
R1521 VDD.n7237 VDD.n7236 203.786
R1522 VDD.n7237 VDD.n6713 203.786
R1523 VDD.n7243 VDD.n6713 203.786
R1524 VDD.n7244 VDD.n7243 203.786
R1525 VDD.n7247 VDD.n7244 203.786
R1526 VDD.n7247 VDD.n7246 203.786
R1527 VDD.n6340 VDD.n5882 203.786
R1528 VDD.n6341 VDD.n6340 203.786
R1529 VDD.n6342 VDD.n6341 203.786
R1530 VDD.n6342 VDD.n5878 203.786
R1531 VDD.n6348 VDD.n5878 203.786
R1532 VDD.n6349 VDD.n6348 203.786
R1533 VDD.n6350 VDD.n6349 203.786
R1534 VDD.n6350 VDD.n5874 203.786
R1535 VDD.n6356 VDD.n5874 203.786
R1536 VDD.n6357 VDD.n6356 203.786
R1537 VDD.n6358 VDD.n6357 203.786
R1538 VDD.n6358 VDD.n5870 203.786
R1539 VDD.n6364 VDD.n5870 203.786
R1540 VDD.n6365 VDD.n6364 203.786
R1541 VDD.n6366 VDD.n6365 203.786
R1542 VDD.n6366 VDD.n5866 203.786
R1543 VDD.n6372 VDD.n5866 203.786
R1544 VDD.n6373 VDD.n6372 203.786
R1545 VDD.n6374 VDD.n6373 203.786
R1546 VDD.n6374 VDD.n5862 203.786
R1547 VDD.n6380 VDD.n5862 203.786
R1548 VDD.n6381 VDD.n6380 203.786
R1549 VDD.n6382 VDD.n6381 203.786
R1550 VDD.n6382 VDD.n5858 203.786
R1551 VDD.n6388 VDD.n5858 203.786
R1552 VDD.n6389 VDD.n6388 203.786
R1553 VDD.n6392 VDD.n6389 203.786
R1554 VDD.n6392 VDD.n6391 203.786
R1555 VDD.n4720 VDD.n4719 198.731
R1556 VDD.n5161 VDD.n680 195.649
R1557 VDD.n4715 VDD.n4714 193.017
R1558 VDD.n5444 VDD.n282 186.405
R1559 VDD.n2350 VDD.n2349 185
R1560 VDD.n2348 VDD.n2347 185
R1561 VDD.n267 VDD.n265 185
R1562 VDD.n5474 VDD.n5459 185
R1563 VDD.n5472 VDD.n5459 185
R1564 VDD.n5459 VDD.n250 185
R1565 VDD.n5500 VDD.n247 185
R1566 VDD.n5503 VDD.n247 185
R1567 VDD.n2446 VDD.n247 185
R1568 VDD.n2455 VDD.n245 185
R1569 VDD.n2446 VDD.n245 185
R1570 VDD.n5503 VDD.n245 185
R1571 VDD.n5500 VDD.n245 185
R1572 VDD.n2455 VDD.n247 185
R1573 VDD.n2622 VDD.n2621 185
R1574 VDD.n2622 VDD.n2600 185
R1575 VDD.n2621 VDD.n2597 185
R1576 VDD.n2600 VDD.n2597 185
R1577 VDD.n2621 VDD.n2620 185
R1578 VDD.n4001 VDD.n2482 185
R1579 VDD.n4001 VDD.n2488 185
R1580 VDD.n3993 VDD.n2488 185
R1581 VDD.n3993 VDD.n2482 185
R1582 VDD.n2489 VDD.n2482 185
R1583 VDD.n2489 VDD.n2488 185
R1584 VDD.n4009 VDD.n394 185
R1585 VDD.n4007 VDD.n394 185
R1586 VDD.n2481 VDD.n394 185
R1587 VDD.n3951 VDD.n2496 185
R1588 VDD.n2496 VDD.n2014 185
R1589 VDD.n3950 VDD.n2014 185
R1590 VDD.n3952 VDD.n2014 185
R1591 VDD.n3947 VDD.n2014 185
R1592 VDD.n3952 VDD.n3951 185
R1593 VDD.n2503 VDD.n2014 185
R1594 VDD.n2502 VDD.n2014 185
R1595 VDD.n3991 VDD.n2492 179.883
R1596 VDD.n5641 VDD.n5618 175.386
R1597 VDD.n5668 VDD.n5642 175.386
R1598 VDD.n6489 VDD.n6488 175.386
R1599 VDD.n6504 VDD.n6470 175.386
R1600 VDD.n7350 VDD.n7327 175.386
R1601 VDD.n7377 VDD.n7351 175.386
R1602 VDD.n8198 VDD.n8197 175.386
R1603 VDD.n8213 VDD.n8179 175.386
R1604 VDD.n3609 VDD.n3608 174.535
R1605 VDD.n2650 VDD.n2649 174.535
R1606 VDD.n3597 VDD.n2657 174.535
R1607 VDD.n3595 VDD.n2658 174.535
R1608 VDD.n3586 VDD.n3585 174.535
R1609 VDD.n3168 VDD.n3167 174.535
R1610 VDD.n3123 VDD.n3122 174.535
R1611 VDD.n3153 VDD.n3126 174.535
R1612 VDD.n3151 VDD.n3127 174.535
R1613 VDD.n3142 VDD.n3141 174.535
R1614 VDD.n3788 VDD.n3787 174.535
R1615 VDD.n3782 VDD.n3781 174.535
R1616 VDD.n2939 VDD.n2928 174.535
R1617 VDD.n2931 VDD.n2930 174.535
R1618 VDD.n2999 VDD.n2998 174.535
R1619 VDD.n2992 VDD.n2991 174.535
R1620 VDD.n2987 VDD.n2986 174.535
R1621 VDD.n89 VDD.n47 174.535
R1622 VDD.n85 VDD.n84 174.535
R1623 VDD.n76 VDD.n75 174.535
R1624 VDD.n68 VDD.n63 174.535
R1625 VDD.n5548 VDD.n5530 174.535
R1626 VDD.n5592 VDD.n5591 174.535
R1627 VDD.n5582 VDD.n5566 174.535
R1628 VDD.n5580 VDD.n5567 174.535
R1629 VDD.n192 VDD.n178 174.535
R1630 VDD.n233 VDD.n232 174.535
R1631 VDD.n222 VDD.n221 174.535
R1632 VDD.n214 VDD.n209 174.535
R1633 VDD.n5627 VDD.t68 171.452
R1634 VDD.t144 VDD.n6487 171.452
R1635 VDD.n7336 VDD.t14 171.452
R1636 VDD.t65 VDD.n8196 171.452
R1637 VDD.n1860 VDD.n1859 171
R1638 VDD.n8994 VDD.n8993 168.889
R1639 VDD.n8468 VDD.n8464 168.889
R1640 VDD.n8139 VDD.n8138 168.889
R1641 VDD.n7613 VDD.n7609 168.889
R1642 VDD.n7285 VDD.n7284 168.889
R1643 VDD.n6759 VDD.n6755 168.889
R1644 VDD.n6430 VDD.n6429 168.889
R1645 VDD.n5904 VDD.n5900 168.889
R1646 VDD.n1470 VDD.n1398 167.919
R1647 VDD.n4715 VDD.n921 165.874
R1648 VDD.n8898 VDD.n8897 164.827
R1649 VDD.n8043 VDD.n8042 164.827
R1650 VDD.n7189 VDD.n7188 164.827
R1651 VDD.n6334 VDD.n6333 164.827
R1652 VDD.n8954 VDD.n8415 162.857
R1653 VDD.n8897 VDD.n8896 162.857
R1654 VDD.n8099 VDD.n7560 162.857
R1655 VDD.n8042 VDD.n8041 162.857
R1656 VDD.n7245 VDD.n6706 162.857
R1657 VDD.n7188 VDD.n7187 162.857
R1658 VDD.n6390 VDD.n5851 162.857
R1659 VDD.n6333 VDD.n6332 162.857
R1660 VDD.n5163 VDD.n5162 162.857
R1661 VDD.n8954 VDD.n8418 161.831
R1662 VDD.n8099 VDD.n7563 161.831
R1663 VDD.n7245 VDD.n6709 161.831
R1664 VDD.n6390 VDD.n5854 161.831
R1665 VDD.n5630 VDD.t69 160.743
R1666 VDD.n6479 VDD.t145 160.743
R1667 VDD.n7339 VDD.t15 160.743
R1668 VDD.n8188 VDD.t66 160.743
R1669 VDD.n8853 VDD.n8468 160.256
R1670 VDD.n7998 VDD.n7613 160.256
R1671 VDD.n7144 VDD.n6759 160.256
R1672 VDD.n6289 VDD.n5904 160.256
R1673 VDD.n3985 VDD.n2496 159.156
R1674 VDD.n8647 VDD.n8503 159.113
R1675 VDD.n8633 VDD.n8503 159.113
R1676 VDD.n8633 VDD.n8632 159.113
R1677 VDD.n8632 VDD.n8631 159.113
R1678 VDD.n8631 VDD.n8508 159.113
R1679 VDD.n8625 VDD.n8508 159.113
R1680 VDD.n8625 VDD.n8624 159.113
R1681 VDD.n8624 VDD.n8623 159.113
R1682 VDD.n8623 VDD.n8512 159.113
R1683 VDD.n8617 VDD.n8512 159.113
R1684 VDD.n8617 VDD.n8616 159.113
R1685 VDD.n8616 VDD.n8615 159.113
R1686 VDD.n8615 VDD.n8516 159.113
R1687 VDD.n8609 VDD.n8516 159.113
R1688 VDD.n8609 VDD.n8608 159.113
R1689 VDD.n8608 VDD.n8607 159.113
R1690 VDD.n8607 VDD.n8520 159.113
R1691 VDD.n8601 VDD.n8520 159.113
R1692 VDD.n8601 VDD.n8600 159.113
R1693 VDD.n8600 VDD.n8599 159.113
R1694 VDD.n8599 VDD.n8524 159.113
R1695 VDD.n8593 VDD.n8524 159.113
R1696 VDD.n8593 VDD.n8592 159.113
R1697 VDD.n8592 VDD.n8591 159.113
R1698 VDD.n8591 VDD.n8528 159.113
R1699 VDD.n8585 VDD.n8528 159.113
R1700 VDD.n8585 VDD.n8584 159.113
R1701 VDD.n8584 VDD.n8583 159.113
R1702 VDD.n7792 VDD.n7648 159.113
R1703 VDD.n7778 VDD.n7648 159.113
R1704 VDD.n7778 VDD.n7777 159.113
R1705 VDD.n7777 VDD.n7776 159.113
R1706 VDD.n7776 VDD.n7653 159.113
R1707 VDD.n7770 VDD.n7653 159.113
R1708 VDD.n7770 VDD.n7769 159.113
R1709 VDD.n7769 VDD.n7768 159.113
R1710 VDD.n7768 VDD.n7657 159.113
R1711 VDD.n7762 VDD.n7657 159.113
R1712 VDD.n7762 VDD.n7761 159.113
R1713 VDD.n7761 VDD.n7760 159.113
R1714 VDD.n7760 VDD.n7661 159.113
R1715 VDD.n7754 VDD.n7661 159.113
R1716 VDD.n7754 VDD.n7753 159.113
R1717 VDD.n7753 VDD.n7752 159.113
R1718 VDD.n7752 VDD.n7665 159.113
R1719 VDD.n7746 VDD.n7665 159.113
R1720 VDD.n7746 VDD.n7745 159.113
R1721 VDD.n7745 VDD.n7744 159.113
R1722 VDD.n7744 VDD.n7669 159.113
R1723 VDD.n7738 VDD.n7669 159.113
R1724 VDD.n7738 VDD.n7737 159.113
R1725 VDD.n7737 VDD.n7736 159.113
R1726 VDD.n7736 VDD.n7673 159.113
R1727 VDD.n7730 VDD.n7673 159.113
R1728 VDD.n7730 VDD.n7729 159.113
R1729 VDD.n7729 VDD.n7728 159.113
R1730 VDD.n6938 VDD.n6794 159.113
R1731 VDD.n6924 VDD.n6794 159.113
R1732 VDD.n6924 VDD.n6923 159.113
R1733 VDD.n6923 VDD.n6922 159.113
R1734 VDD.n6922 VDD.n6799 159.113
R1735 VDD.n6916 VDD.n6799 159.113
R1736 VDD.n6916 VDD.n6915 159.113
R1737 VDD.n6915 VDD.n6914 159.113
R1738 VDD.n6914 VDD.n6803 159.113
R1739 VDD.n6908 VDD.n6803 159.113
R1740 VDD.n6908 VDD.n6907 159.113
R1741 VDD.n6907 VDD.n6906 159.113
R1742 VDD.n6906 VDD.n6807 159.113
R1743 VDD.n6900 VDD.n6807 159.113
R1744 VDD.n6900 VDD.n6899 159.113
R1745 VDD.n6899 VDD.n6898 159.113
R1746 VDD.n6898 VDD.n6811 159.113
R1747 VDD.n6892 VDD.n6811 159.113
R1748 VDD.n6892 VDD.n6891 159.113
R1749 VDD.n6891 VDD.n6890 159.113
R1750 VDD.n6890 VDD.n6815 159.113
R1751 VDD.n6884 VDD.n6815 159.113
R1752 VDD.n6884 VDD.n6883 159.113
R1753 VDD.n6883 VDD.n6882 159.113
R1754 VDD.n6882 VDD.n6819 159.113
R1755 VDD.n6876 VDD.n6819 159.113
R1756 VDD.n6876 VDD.n6875 159.113
R1757 VDD.n6875 VDD.n6874 159.113
R1758 VDD.n6083 VDD.n5939 159.113
R1759 VDD.n6069 VDD.n5939 159.113
R1760 VDD.n6069 VDD.n6068 159.113
R1761 VDD.n6068 VDD.n6067 159.113
R1762 VDD.n6067 VDD.n5944 159.113
R1763 VDD.n6061 VDD.n5944 159.113
R1764 VDD.n6061 VDD.n6060 159.113
R1765 VDD.n6060 VDD.n6059 159.113
R1766 VDD.n6059 VDD.n5948 159.113
R1767 VDD.n6053 VDD.n5948 159.113
R1768 VDD.n6053 VDD.n6052 159.113
R1769 VDD.n6052 VDD.n6051 159.113
R1770 VDD.n6051 VDD.n5952 159.113
R1771 VDD.n6045 VDD.n5952 159.113
R1772 VDD.n6045 VDD.n6044 159.113
R1773 VDD.n6044 VDD.n6043 159.113
R1774 VDD.n6043 VDD.n5956 159.113
R1775 VDD.n6037 VDD.n5956 159.113
R1776 VDD.n6037 VDD.n6036 159.113
R1777 VDD.n6036 VDD.n6035 159.113
R1778 VDD.n6035 VDD.n5960 159.113
R1779 VDD.n6029 VDD.n5960 159.113
R1780 VDD.n6029 VDD.n6028 159.113
R1781 VDD.n6028 VDD.n6027 159.113
R1782 VDD.n6027 VDD.n5964 159.113
R1783 VDD.n6021 VDD.n5964 159.113
R1784 VDD.n6021 VDD.n6020 159.113
R1785 VDD.n6020 VDD.n6019 159.113
R1786 VDD.n5622 VDD.t71 158.225
R1787 VDD.n6500 VDD.t147 158.225
R1788 VDD.n7331 VDD.t17 158.225
R1789 VDD.n8209 VDD.t64 158.225
R1790 VDD.n8994 VDD.n8278 154.488
R1791 VDD.n8139 VDD.n7423 154.488
R1792 VDD.n7285 VDD.n6569 154.488
R1793 VDD.n6430 VDD.n5714 154.488
R1794 VDD.n5498 VDD.n250 153.975
R1795 VDD.n3496 VDD.n3493 152
R1796 VDD.n3495 VDD.n3494 152
R1797 VDD.n3513 VDD.n3507 152
R1798 VDD.n3512 VDD.n3511 152
R1799 VDD.n3198 VDD.n3195 152
R1800 VDD.n3197 VDD.n3196 152
R1801 VDD.n3215 VDD.n3209 152
R1802 VDD.n3214 VDD.n3213 152
R1803 VDD.n3746 VDD.n3743 152
R1804 VDD.n3745 VDD.n3744 152
R1805 VDD.n3844 VDD.n3843 152
R1806 VDD.n3839 VDD.n3737 152
R1807 VDD.n3838 VDD.n3837 152
R1808 VDD.n3842 VDD.n3841 152
R1809 VDD.n3882 VDD.n3881 152
R1810 VDD.n3883 VDD.n3877 152
R1811 VDD.n3864 VDD.n3863 152
R1812 VDD.n3861 VDD.n3860 152
R1813 VDD.n3862 VDD.n3709 152
R1814 VDD.n3865 VDD.n3710 152
R1815 VDD.n2825 VDD.n2824 152
R1816 VDD.n2827 VDD.n2826 152
R1817 VDD.n2967 VDD.n2966 152
R1818 VDD.n2969 VDD.n2968 152
R1819 VDD.t142 VDD.t141 151.181
R1820 VDD.t141 VDD.t140 151.181
R1821 VDD.t98 VDD.t83 151.181
R1822 VDD.t44 VDD.t98 151.181
R1823 VDD.t99 VDD.t44 151.181
R1824 VDD.t126 VDD.t99 151.181
R1825 VDD.t4 VDD.t126 151.181
R1826 VDD.t8 VDD.t4 151.181
R1827 VDD.t115 VDD.t8 151.181
R1828 VDD.n8646 VDD.n8504 141.731
R1829 VDD.n8582 VDD.n8533 141.731
R1830 VDD.n7791 VDD.n7649 141.731
R1831 VDD.n7727 VDD.n7678 141.731
R1832 VDD.n6937 VDD.n6795 141.731
R1833 VDD.n6873 VDD.n6824 141.731
R1834 VDD.n6082 VDD.n5940 141.731
R1835 VDD.n6018 VDD.n5969 141.731
R1836 VDD.n8899 VDD.n8447 140.19
R1837 VDD.n8961 VDD.n8419 140.19
R1838 VDD.n8044 VDD.n7592 140.19
R1839 VDD.n8106 VDD.n7564 140.19
R1840 VDD.n7190 VDD.n6738 140.19
R1841 VDD.n7252 VDD.n6710 140.19
R1842 VDD.n6335 VDD.n5883 140.19
R1843 VDD.n6397 VDD.n5855 140.19
R1844 VDD.n8799 VDD.n8715 133.655
R1845 VDD.n8810 VDD.n8748 133.655
R1846 VDD.n8745 VDD.n8724 133.655
R1847 VDD.n8741 VDD.n8723 133.655
R1848 VDD.n8739 VDD.n8738 133.655
R1849 VDD.n8735 VDD.n8734 133.655
R1850 VDD.n8300 VDD.n8292 133.655
R1851 VDD.n8838 VDD.n8693 133.655
R1852 VDD.n8830 VDD.n8693 133.655
R1853 VDD.n8830 VDD.n8700 133.655
R1854 VDD.n8822 VDD.n8700 133.655
R1855 VDD.n8822 VDD.n8710 133.655
R1856 VDD.n8733 VDD.n8732 133.655
R1857 VDD.n8732 VDD.n8265 133.655
R1858 VDD.n9007 VDD.n8265 133.655
R1859 VDD.n9007 VDD.n9006 133.655
R1860 VDD.n9006 VDD.n8266 133.655
R1861 VDD.n8851 VDD.n8682 133.655
R1862 VDD.n8843 VDD.n8688 133.655
R1863 VDD.n8703 VDD.n8681 133.655
R1864 VDD.n8828 VDD.n8703 133.655
R1865 VDD.n8828 VDD.n8704 133.655
R1866 VDD.n8824 VDD.n8704 133.655
R1867 VDD.n8824 VDD.n8707 133.655
R1868 VDD.n8729 VDD.n8728 133.655
R1869 VDD.n8728 VDD.n8727 133.655
R1870 VDD.n8727 VDD.n8268 133.655
R1871 VDD.n9004 VDD.n8268 133.655
R1872 VDD.n9004 VDD.n8269 133.655
R1873 VDD.n8774 VDD.n8773 133.655
R1874 VDD.n8780 VDD.n8779 133.655
R1875 VDD.n8835 VDD.n8697 133.655
R1876 VDD.n8835 VDD.n8698 133.655
R1877 VDD.n8714 VDD.n8698 133.655
R1878 VDD.n8817 VDD.n8719 133.655
R1879 VDD.n8719 VDD.n8249 133.655
R1880 VDD.n9018 VDD.n8249 133.655
R1881 VDD.n9018 VDD.n8250 133.655
R1882 VDD.n9010 VDD.n8250 133.655
R1883 VDD.n8396 VDD.n8291 133.655
R1884 VDD.n8399 VDD.n8287 133.655
R1885 VDD.n8331 VDD.n8330 133.655
R1886 VDD.n8322 VDD.n8320 133.655
R1887 VDD.n8789 VDD.n8696 133.655
R1888 VDD.n8793 VDD.n8696 133.655
R1889 VDD.n8794 VDD.n8793 133.655
R1890 VDD.n8815 VDD.n8751 133.655
R1891 VDD.n8751 VDD.n8253 133.655
R1892 VDD.n9016 VDD.n8253 133.655
R1893 VDD.n9016 VDD.n8254 133.655
R1894 VDD.n9012 VDD.n8254 133.655
R1895 VDD.n8394 VDD.n8391 133.655
R1896 VDD.n8394 VDD.n8284 133.655
R1897 VDD.n8401 VDD.n8284 133.655
R1898 VDD.n8357 VDD.n8261 133.655
R1899 VDD.n8346 VDD.n8257 133.655
R1900 VDD.n7944 VDD.n7860 133.655
R1901 VDD.n7955 VDD.n7893 133.655
R1902 VDD.n7890 VDD.n7869 133.655
R1903 VDD.n7886 VDD.n7868 133.655
R1904 VDD.n7884 VDD.n7883 133.655
R1905 VDD.n7880 VDD.n7879 133.655
R1906 VDD.n7445 VDD.n7437 133.655
R1907 VDD.n7983 VDD.n7838 133.655
R1908 VDD.n7975 VDD.n7838 133.655
R1909 VDD.n7975 VDD.n7845 133.655
R1910 VDD.n7967 VDD.n7845 133.655
R1911 VDD.n7967 VDD.n7855 133.655
R1912 VDD.n7878 VDD.n7877 133.655
R1913 VDD.n7877 VDD.n7410 133.655
R1914 VDD.n8152 VDD.n7410 133.655
R1915 VDD.n8152 VDD.n8151 133.655
R1916 VDD.n8151 VDD.n7411 133.655
R1917 VDD.n7996 VDD.n7827 133.655
R1918 VDD.n7988 VDD.n7833 133.655
R1919 VDD.n7848 VDD.n7826 133.655
R1920 VDD.n7973 VDD.n7848 133.655
R1921 VDD.n7973 VDD.n7849 133.655
R1922 VDD.n7969 VDD.n7849 133.655
R1923 VDD.n7969 VDD.n7852 133.655
R1924 VDD.n7874 VDD.n7873 133.655
R1925 VDD.n7873 VDD.n7872 133.655
R1926 VDD.n7872 VDD.n7413 133.655
R1927 VDD.n8149 VDD.n7413 133.655
R1928 VDD.n8149 VDD.n7414 133.655
R1929 VDD.n7919 VDD.n7918 133.655
R1930 VDD.n7925 VDD.n7924 133.655
R1931 VDD.n7980 VDD.n7842 133.655
R1932 VDD.n7980 VDD.n7843 133.655
R1933 VDD.n7859 VDD.n7843 133.655
R1934 VDD.n7962 VDD.n7864 133.655
R1935 VDD.n7864 VDD.n7394 133.655
R1936 VDD.n8163 VDD.n7394 133.655
R1937 VDD.n8163 VDD.n7395 133.655
R1938 VDD.n8155 VDD.n7395 133.655
R1939 VDD.n7541 VDD.n7436 133.655
R1940 VDD.n7544 VDD.n7432 133.655
R1941 VDD.n7476 VDD.n7475 133.655
R1942 VDD.n7467 VDD.n7465 133.655
R1943 VDD.n7934 VDD.n7841 133.655
R1944 VDD.n7938 VDD.n7841 133.655
R1945 VDD.n7939 VDD.n7938 133.655
R1946 VDD.n7960 VDD.n7896 133.655
R1947 VDD.n7896 VDD.n7398 133.655
R1948 VDD.n8161 VDD.n7398 133.655
R1949 VDD.n8161 VDD.n7399 133.655
R1950 VDD.n8157 VDD.n7399 133.655
R1951 VDD.n7539 VDD.n7536 133.655
R1952 VDD.n7539 VDD.n7429 133.655
R1953 VDD.n7546 VDD.n7429 133.655
R1954 VDD.n7502 VDD.n7406 133.655
R1955 VDD.n7491 VDD.n7402 133.655
R1956 VDD.n7090 VDD.n7006 133.655
R1957 VDD.n7101 VDD.n7039 133.655
R1958 VDD.n7036 VDD.n7015 133.655
R1959 VDD.n7032 VDD.n7014 133.655
R1960 VDD.n7030 VDD.n7029 133.655
R1961 VDD.n7026 VDD.n7025 133.655
R1962 VDD.n6591 VDD.n6583 133.655
R1963 VDD.n7129 VDD.n6984 133.655
R1964 VDD.n7121 VDD.n6984 133.655
R1965 VDD.n7121 VDD.n6991 133.655
R1966 VDD.n7113 VDD.n6991 133.655
R1967 VDD.n7113 VDD.n7001 133.655
R1968 VDD.n7024 VDD.n7023 133.655
R1969 VDD.n7023 VDD.n6556 133.655
R1970 VDD.n7298 VDD.n6556 133.655
R1971 VDD.n7298 VDD.n7297 133.655
R1972 VDD.n7297 VDD.n6557 133.655
R1973 VDD.n7142 VDD.n6973 133.655
R1974 VDD.n7134 VDD.n6979 133.655
R1975 VDD.n6994 VDD.n6972 133.655
R1976 VDD.n7119 VDD.n6994 133.655
R1977 VDD.n7119 VDD.n6995 133.655
R1978 VDD.n7115 VDD.n6995 133.655
R1979 VDD.n7115 VDD.n6998 133.655
R1980 VDD.n7020 VDD.n7019 133.655
R1981 VDD.n7019 VDD.n7018 133.655
R1982 VDD.n7018 VDD.n6559 133.655
R1983 VDD.n7295 VDD.n6559 133.655
R1984 VDD.n7295 VDD.n6560 133.655
R1985 VDD.n7065 VDD.n7064 133.655
R1986 VDD.n7071 VDD.n7070 133.655
R1987 VDD.n7126 VDD.n6988 133.655
R1988 VDD.n7126 VDD.n6989 133.655
R1989 VDD.n7005 VDD.n6989 133.655
R1990 VDD.n7108 VDD.n7010 133.655
R1991 VDD.n7010 VDD.n6540 133.655
R1992 VDD.n7309 VDD.n6540 133.655
R1993 VDD.n7309 VDD.n6541 133.655
R1994 VDD.n7301 VDD.n6541 133.655
R1995 VDD.n6687 VDD.n6582 133.655
R1996 VDD.n6690 VDD.n6578 133.655
R1997 VDD.n6622 VDD.n6621 133.655
R1998 VDD.n6613 VDD.n6611 133.655
R1999 VDD.n7080 VDD.n6987 133.655
R2000 VDD.n7084 VDD.n6987 133.655
R2001 VDD.n7085 VDD.n7084 133.655
R2002 VDD.n7106 VDD.n7042 133.655
R2003 VDD.n7042 VDD.n6544 133.655
R2004 VDD.n7307 VDD.n6544 133.655
R2005 VDD.n7307 VDD.n6545 133.655
R2006 VDD.n7303 VDD.n6545 133.655
R2007 VDD.n6685 VDD.n6682 133.655
R2008 VDD.n6685 VDD.n6575 133.655
R2009 VDD.n6692 VDD.n6575 133.655
R2010 VDD.n6648 VDD.n6552 133.655
R2011 VDD.n6637 VDD.n6548 133.655
R2012 VDD.n6235 VDD.n6151 133.655
R2013 VDD.n6246 VDD.n6184 133.655
R2014 VDD.n6181 VDD.n6160 133.655
R2015 VDD.n6177 VDD.n6159 133.655
R2016 VDD.n6175 VDD.n6174 133.655
R2017 VDD.n6171 VDD.n6170 133.655
R2018 VDD.n5736 VDD.n5728 133.655
R2019 VDD.n6274 VDD.n6129 133.655
R2020 VDD.n6266 VDD.n6129 133.655
R2021 VDD.n6266 VDD.n6136 133.655
R2022 VDD.n6258 VDD.n6136 133.655
R2023 VDD.n6258 VDD.n6146 133.655
R2024 VDD.n6169 VDD.n6168 133.655
R2025 VDD.n6168 VDD.n5701 133.655
R2026 VDD.n6443 VDD.n5701 133.655
R2027 VDD.n6443 VDD.n6442 133.655
R2028 VDD.n6442 VDD.n5702 133.655
R2029 VDD.n6287 VDD.n6118 133.655
R2030 VDD.n6279 VDD.n6124 133.655
R2031 VDD.n6139 VDD.n6117 133.655
R2032 VDD.n6264 VDD.n6139 133.655
R2033 VDD.n6264 VDD.n6140 133.655
R2034 VDD.n6260 VDD.n6140 133.655
R2035 VDD.n6260 VDD.n6143 133.655
R2036 VDD.n6165 VDD.n6164 133.655
R2037 VDD.n6164 VDD.n6163 133.655
R2038 VDD.n6163 VDD.n5704 133.655
R2039 VDD.n6440 VDD.n5704 133.655
R2040 VDD.n6440 VDD.n5705 133.655
R2041 VDD.n6210 VDD.n6209 133.655
R2042 VDD.n6216 VDD.n6215 133.655
R2043 VDD.n6271 VDD.n6133 133.655
R2044 VDD.n6271 VDD.n6134 133.655
R2045 VDD.n6150 VDD.n6134 133.655
R2046 VDD.n6253 VDD.n6155 133.655
R2047 VDD.n6155 VDD.n5685 133.655
R2048 VDD.n6454 VDD.n5685 133.655
R2049 VDD.n6454 VDD.n5686 133.655
R2050 VDD.n6446 VDD.n5686 133.655
R2051 VDD.n5832 VDD.n5727 133.655
R2052 VDD.n5835 VDD.n5723 133.655
R2053 VDD.n5767 VDD.n5766 133.655
R2054 VDD.n5758 VDD.n5756 133.655
R2055 VDD.n6225 VDD.n6132 133.655
R2056 VDD.n6229 VDD.n6132 133.655
R2057 VDD.n6230 VDD.n6229 133.655
R2058 VDD.n6251 VDD.n6187 133.655
R2059 VDD.n6187 VDD.n5689 133.655
R2060 VDD.n6452 VDD.n5689 133.655
R2061 VDD.n6452 VDD.n5690 133.655
R2062 VDD.n6448 VDD.n5690 133.655
R2063 VDD.n5830 VDD.n5827 133.655
R2064 VDD.n5830 VDD.n5720 133.655
R2065 VDD.n5837 VDD.n5720 133.655
R2066 VDD.n5793 VDD.n5697 133.655
R2067 VDD.n5782 VDD.n5693 133.655
R2068 VDD.n8648 VDD.n8502 128.696
R2069 VDD.n7793 VDD.n7647 128.696
R2070 VDD.n6939 VDD.n6793 128.696
R2071 VDD.n6084 VDD.n5938 128.696
R2072 VDD.n2488 VDD.t115 126.425
R2073 VDD.n8536 VDD.n8532 126.356
R2074 VDD.n7681 VDD.n7677 126.356
R2075 VDD.n6827 VDD.n6823 126.356
R2076 VDD.n5972 VDD.n5968 126.356
R2077 VDD.n5286 VDD.n5285 123.651
R2078 VDD.t89 VDD.n5666 117.838
R2079 VDD.n6517 VDD.t36 117.838
R2080 VDD.t18 VDD.n7375 117.838
R2081 VDD.n8226 VDD.t73 117.838
R2082 VDD.n4718 VDD.n4715 117.62
R2083 VDD.n2925 VDD.t120 116.841
R2084 VDD.n64 VDD.t55 116.841
R2085 VDD.t51 VDD.n5569 116.841
R2086 VDD.n3582 VDD.t107 116.841
R2087 VDD.n3138 VDD.t117 116.841
R2088 VDD.t109 VDD.n3764 116.841
R2089 VDD.n210 VDD.t7 116.841
R2090 VDD.n8634 VDD.n8505 104.757
R2091 VDD.n8634 VDD.n8507 104.757
R2092 VDD.n8630 VDD.n8507 104.757
R2093 VDD.n8630 VDD.n8509 104.757
R2094 VDD.n8626 VDD.n8509 104.757
R2095 VDD.n8626 VDD.n8511 104.757
R2096 VDD.n8622 VDD.n8511 104.757
R2097 VDD.n8622 VDD.n8513 104.757
R2098 VDD.n8618 VDD.n8513 104.757
R2099 VDD.n8618 VDD.n8515 104.757
R2100 VDD.n8614 VDD.n8515 104.757
R2101 VDD.n8614 VDD.n8517 104.757
R2102 VDD.n8610 VDD.n8517 104.757
R2103 VDD.n8610 VDD.n8519 104.757
R2104 VDD.n8606 VDD.n8519 104.757
R2105 VDD.n8606 VDD.n8521 104.757
R2106 VDD.n8602 VDD.n8521 104.757
R2107 VDD.n8602 VDD.n8523 104.757
R2108 VDD.n8598 VDD.n8523 104.757
R2109 VDD.n8598 VDD.n8525 104.757
R2110 VDD.n8594 VDD.n8525 104.757
R2111 VDD.n8594 VDD.n8527 104.757
R2112 VDD.n8590 VDD.n8527 104.757
R2113 VDD.n8590 VDD.n8529 104.757
R2114 VDD.n8586 VDD.n8529 104.757
R2115 VDD.n8586 VDD.n8531 104.757
R2116 VDD.n8582 VDD.n8531 104.757
R2117 VDD.n8650 VDD.n8501 104.757
R2118 VDD.n8650 VDD.n8499 104.757
R2119 VDD.n8654 VDD.n8499 104.757
R2120 VDD.n8654 VDD.n8497 104.757
R2121 VDD.n8658 VDD.n8497 104.757
R2122 VDD.n8658 VDD.n8495 104.757
R2123 VDD.n8662 VDD.n8495 104.757
R2124 VDD.n8662 VDD.n8493 104.757
R2125 VDD.n8666 VDD.n8493 104.757
R2126 VDD.n8666 VDD.n8491 104.757
R2127 VDD.n8670 VDD.n8491 104.757
R2128 VDD.n8670 VDD.n8489 104.757
R2129 VDD.n8675 VDD.n8489 104.757
R2130 VDD.n8675 VDD.n8487 104.757
R2131 VDD.n8862 VDD.n8487 104.757
R2132 VDD.n8841 VDD.n8479 104.757
R2133 VDD.n8758 VDD.n8479 104.757
R2134 VDD.n8762 VDD.n8761 104.757
R2135 VDD.n8866 VDD.n8465 104.757
R2136 VDD.n8870 VDD.n8465 104.757
R2137 VDD.n8870 VDD.n8463 104.757
R2138 VDD.n8874 VDD.n8463 104.757
R2139 VDD.n8874 VDD.n8461 104.757
R2140 VDD.n8878 VDD.n8461 104.757
R2141 VDD.n8878 VDD.n8459 104.757
R2142 VDD.n8882 VDD.n8459 104.757
R2143 VDD.n8882 VDD.n8457 104.757
R2144 VDD.n8886 VDD.n8457 104.757
R2145 VDD.n8886 VDD.n8455 104.757
R2146 VDD.n8890 VDD.n8455 104.757
R2147 VDD.n8890 VDD.n8452 104.757
R2148 VDD.n8895 VDD.n8452 104.757
R2149 VDD.n8895 VDD.n8453 104.757
R2150 VDD.n8899 VDD.n8449 104.757
R2151 VDD.n8903 VDD.n8447 104.757
R2152 VDD.n8903 VDD.n8445 104.757
R2153 VDD.n8907 VDD.n8445 104.757
R2154 VDD.n8907 VDD.n8443 104.757
R2155 VDD.n8911 VDD.n8443 104.757
R2156 VDD.n8911 VDD.n8441 104.757
R2157 VDD.n8915 VDD.n8441 104.757
R2158 VDD.n8915 VDD.n8439 104.757
R2159 VDD.n8919 VDD.n8439 104.757
R2160 VDD.n8919 VDD.n8437 104.757
R2161 VDD.n8923 VDD.n8437 104.757
R2162 VDD.n8923 VDD.n8435 104.757
R2163 VDD.n8927 VDD.n8435 104.757
R2164 VDD.n8927 VDD.n8433 104.757
R2165 VDD.n8931 VDD.n8433 104.757
R2166 VDD.n8931 VDD.n8431 104.757
R2167 VDD.n8935 VDD.n8431 104.757
R2168 VDD.n8935 VDD.n8429 104.757
R2169 VDD.n8939 VDD.n8429 104.757
R2170 VDD.n8939 VDD.n8427 104.757
R2171 VDD.n8943 VDD.n8427 104.757
R2172 VDD.n8943 VDD.n8425 104.757
R2173 VDD.n8947 VDD.n8425 104.757
R2174 VDD.n8947 VDD.n8423 104.757
R2175 VDD.n8951 VDD.n8423 104.757
R2176 VDD.n8951 VDD.n8421 104.757
R2177 VDD.n8957 VDD.n8421 104.757
R2178 VDD.n8957 VDD.n8419 104.757
R2179 VDD.n8578 VDD.n8577 104.757
R2180 VDD.n8575 VDD.n8537 104.757
R2181 VDD.n8571 VDD.n8537 104.757
R2182 VDD.n8571 VDD.n8539 104.757
R2183 VDD.n8567 VDD.n8539 104.757
R2184 VDD.n8567 VDD.n8542 104.757
R2185 VDD.n8563 VDD.n8542 104.757
R2186 VDD.n8563 VDD.n8544 104.757
R2187 VDD.n8559 VDD.n8544 104.757
R2188 VDD.n8559 VDD.n8546 104.757
R2189 VDD.n8555 VDD.n8546 104.757
R2190 VDD.n8555 VDD.n8548 104.757
R2191 VDD.n8551 VDD.n8548 104.757
R2192 VDD.n8551 VDD.n8275 104.757
R2193 VDD.n8996 VDD.n8275 104.757
R2194 VDD.n8997 VDD.n8996 104.757
R2195 VDD.n8383 VDD.n8298 104.757
R2196 VDD.n8381 VDD.n8299 104.757
R2197 VDD.n8373 VDD.n8372 104.757
R2198 VDD.n8368 VDD.n8367 104.757
R2199 VDD.n8336 VDD.n8305 104.757
R2200 VDD.n8327 VDD.n8311 104.757
R2201 VDD.n8325 VDD.n8312 104.757
R2202 VDD.n8316 VDD.n8315 104.757
R2203 VDD.n8992 VDD.n8280 104.757
R2204 VDD.n8992 VDD.n8281 104.757
R2205 VDD.n8988 VDD.n8281 104.757
R2206 VDD.n8988 VDD.n8406 104.757
R2207 VDD.n8984 VDD.n8406 104.757
R2208 VDD.n8984 VDD.n8408 104.757
R2209 VDD.n8980 VDD.n8408 104.757
R2210 VDD.n8980 VDD.n8410 104.757
R2211 VDD.n8976 VDD.n8410 104.757
R2212 VDD.n8976 VDD.n8412 104.757
R2213 VDD.n8972 VDD.n8412 104.757
R2214 VDD.n8972 VDD.n8414 104.757
R2215 VDD.n8968 VDD.n8414 104.757
R2216 VDD.n8968 VDD.n8416 104.757
R2217 VDD.n8964 VDD.n8416 104.757
R2218 VDD.n8962 VDD.n8961 104.757
R2219 VDD.n7779 VDD.n7650 104.757
R2220 VDD.n7779 VDD.n7652 104.757
R2221 VDD.n7775 VDD.n7652 104.757
R2222 VDD.n7775 VDD.n7654 104.757
R2223 VDD.n7771 VDD.n7654 104.757
R2224 VDD.n7771 VDD.n7656 104.757
R2225 VDD.n7767 VDD.n7656 104.757
R2226 VDD.n7767 VDD.n7658 104.757
R2227 VDD.n7763 VDD.n7658 104.757
R2228 VDD.n7763 VDD.n7660 104.757
R2229 VDD.n7759 VDD.n7660 104.757
R2230 VDD.n7759 VDD.n7662 104.757
R2231 VDD.n7755 VDD.n7662 104.757
R2232 VDD.n7755 VDD.n7664 104.757
R2233 VDD.n7751 VDD.n7664 104.757
R2234 VDD.n7751 VDD.n7666 104.757
R2235 VDD.n7747 VDD.n7666 104.757
R2236 VDD.n7747 VDD.n7668 104.757
R2237 VDD.n7743 VDD.n7668 104.757
R2238 VDD.n7743 VDD.n7670 104.757
R2239 VDD.n7739 VDD.n7670 104.757
R2240 VDD.n7739 VDD.n7672 104.757
R2241 VDD.n7735 VDD.n7672 104.757
R2242 VDD.n7735 VDD.n7674 104.757
R2243 VDD.n7731 VDD.n7674 104.757
R2244 VDD.n7731 VDD.n7676 104.757
R2245 VDD.n7727 VDD.n7676 104.757
R2246 VDD.n7795 VDD.n7646 104.757
R2247 VDD.n7795 VDD.n7644 104.757
R2248 VDD.n7799 VDD.n7644 104.757
R2249 VDD.n7799 VDD.n7642 104.757
R2250 VDD.n7803 VDD.n7642 104.757
R2251 VDD.n7803 VDD.n7640 104.757
R2252 VDD.n7807 VDD.n7640 104.757
R2253 VDD.n7807 VDD.n7638 104.757
R2254 VDD.n7811 VDD.n7638 104.757
R2255 VDD.n7811 VDD.n7636 104.757
R2256 VDD.n7815 VDD.n7636 104.757
R2257 VDD.n7815 VDD.n7634 104.757
R2258 VDD.n7820 VDD.n7634 104.757
R2259 VDD.n7820 VDD.n7632 104.757
R2260 VDD.n8007 VDD.n7632 104.757
R2261 VDD.n7986 VDD.n7624 104.757
R2262 VDD.n7903 VDD.n7624 104.757
R2263 VDD.n7907 VDD.n7906 104.757
R2264 VDD.n8011 VDD.n7610 104.757
R2265 VDD.n8015 VDD.n7610 104.757
R2266 VDD.n8015 VDD.n7608 104.757
R2267 VDD.n8019 VDD.n7608 104.757
R2268 VDD.n8019 VDD.n7606 104.757
R2269 VDD.n8023 VDD.n7606 104.757
R2270 VDD.n8023 VDD.n7604 104.757
R2271 VDD.n8027 VDD.n7604 104.757
R2272 VDD.n8027 VDD.n7602 104.757
R2273 VDD.n8031 VDD.n7602 104.757
R2274 VDD.n8031 VDD.n7600 104.757
R2275 VDD.n8035 VDD.n7600 104.757
R2276 VDD.n8035 VDD.n7597 104.757
R2277 VDD.n8040 VDD.n7597 104.757
R2278 VDD.n8040 VDD.n7598 104.757
R2279 VDD.n8044 VDD.n7594 104.757
R2280 VDD.n8048 VDD.n7592 104.757
R2281 VDD.n8048 VDD.n7590 104.757
R2282 VDD.n8052 VDD.n7590 104.757
R2283 VDD.n8052 VDD.n7588 104.757
R2284 VDD.n8056 VDD.n7588 104.757
R2285 VDD.n8056 VDD.n7586 104.757
R2286 VDD.n8060 VDD.n7586 104.757
R2287 VDD.n8060 VDD.n7584 104.757
R2288 VDD.n8064 VDD.n7584 104.757
R2289 VDD.n8064 VDD.n7582 104.757
R2290 VDD.n8068 VDD.n7582 104.757
R2291 VDD.n8068 VDD.n7580 104.757
R2292 VDD.n8072 VDD.n7580 104.757
R2293 VDD.n8072 VDD.n7578 104.757
R2294 VDD.n8076 VDD.n7578 104.757
R2295 VDD.n8076 VDD.n7576 104.757
R2296 VDD.n8080 VDD.n7576 104.757
R2297 VDD.n8080 VDD.n7574 104.757
R2298 VDD.n8084 VDD.n7574 104.757
R2299 VDD.n8084 VDD.n7572 104.757
R2300 VDD.n8088 VDD.n7572 104.757
R2301 VDD.n8088 VDD.n7570 104.757
R2302 VDD.n8092 VDD.n7570 104.757
R2303 VDD.n8092 VDD.n7568 104.757
R2304 VDD.n8096 VDD.n7568 104.757
R2305 VDD.n8096 VDD.n7566 104.757
R2306 VDD.n8102 VDD.n7566 104.757
R2307 VDD.n8102 VDD.n7564 104.757
R2308 VDD.n7723 VDD.n7722 104.757
R2309 VDD.n7720 VDD.n7682 104.757
R2310 VDD.n7716 VDD.n7682 104.757
R2311 VDD.n7716 VDD.n7684 104.757
R2312 VDD.n7712 VDD.n7684 104.757
R2313 VDD.n7712 VDD.n7687 104.757
R2314 VDD.n7708 VDD.n7687 104.757
R2315 VDD.n7708 VDD.n7689 104.757
R2316 VDD.n7704 VDD.n7689 104.757
R2317 VDD.n7704 VDD.n7691 104.757
R2318 VDD.n7700 VDD.n7691 104.757
R2319 VDD.n7700 VDD.n7693 104.757
R2320 VDD.n7696 VDD.n7693 104.757
R2321 VDD.n7696 VDD.n7420 104.757
R2322 VDD.n8141 VDD.n7420 104.757
R2323 VDD.n8142 VDD.n8141 104.757
R2324 VDD.n7528 VDD.n7443 104.757
R2325 VDD.n7526 VDD.n7444 104.757
R2326 VDD.n7518 VDD.n7517 104.757
R2327 VDD.n7513 VDD.n7512 104.757
R2328 VDD.n7481 VDD.n7450 104.757
R2329 VDD.n7472 VDD.n7456 104.757
R2330 VDD.n7470 VDD.n7457 104.757
R2331 VDD.n7461 VDD.n7460 104.757
R2332 VDD.n8137 VDD.n7425 104.757
R2333 VDD.n8137 VDD.n7426 104.757
R2334 VDD.n8133 VDD.n7426 104.757
R2335 VDD.n8133 VDD.n7551 104.757
R2336 VDD.n8129 VDD.n7551 104.757
R2337 VDD.n8129 VDD.n7553 104.757
R2338 VDD.n8125 VDD.n7553 104.757
R2339 VDD.n8125 VDD.n7555 104.757
R2340 VDD.n8121 VDD.n7555 104.757
R2341 VDD.n8121 VDD.n7557 104.757
R2342 VDD.n8117 VDD.n7557 104.757
R2343 VDD.n8117 VDD.n7559 104.757
R2344 VDD.n8113 VDD.n7559 104.757
R2345 VDD.n8113 VDD.n7561 104.757
R2346 VDD.n8109 VDD.n7561 104.757
R2347 VDD.n8107 VDD.n8106 104.757
R2348 VDD.n6925 VDD.n6796 104.757
R2349 VDD.n6925 VDD.n6798 104.757
R2350 VDD.n6921 VDD.n6798 104.757
R2351 VDD.n6921 VDD.n6800 104.757
R2352 VDD.n6917 VDD.n6800 104.757
R2353 VDD.n6917 VDD.n6802 104.757
R2354 VDD.n6913 VDD.n6802 104.757
R2355 VDD.n6913 VDD.n6804 104.757
R2356 VDD.n6909 VDD.n6804 104.757
R2357 VDD.n6909 VDD.n6806 104.757
R2358 VDD.n6905 VDD.n6806 104.757
R2359 VDD.n6905 VDD.n6808 104.757
R2360 VDD.n6901 VDD.n6808 104.757
R2361 VDD.n6901 VDD.n6810 104.757
R2362 VDD.n6897 VDD.n6810 104.757
R2363 VDD.n6897 VDD.n6812 104.757
R2364 VDD.n6893 VDD.n6812 104.757
R2365 VDD.n6893 VDD.n6814 104.757
R2366 VDD.n6889 VDD.n6814 104.757
R2367 VDD.n6889 VDD.n6816 104.757
R2368 VDD.n6885 VDD.n6816 104.757
R2369 VDD.n6885 VDD.n6818 104.757
R2370 VDD.n6881 VDD.n6818 104.757
R2371 VDD.n6881 VDD.n6820 104.757
R2372 VDD.n6877 VDD.n6820 104.757
R2373 VDD.n6877 VDD.n6822 104.757
R2374 VDD.n6873 VDD.n6822 104.757
R2375 VDD.n6941 VDD.n6792 104.757
R2376 VDD.n6941 VDD.n6790 104.757
R2377 VDD.n6945 VDD.n6790 104.757
R2378 VDD.n6945 VDD.n6788 104.757
R2379 VDD.n6949 VDD.n6788 104.757
R2380 VDD.n6949 VDD.n6786 104.757
R2381 VDD.n6953 VDD.n6786 104.757
R2382 VDD.n6953 VDD.n6784 104.757
R2383 VDD.n6957 VDD.n6784 104.757
R2384 VDD.n6957 VDD.n6782 104.757
R2385 VDD.n6961 VDD.n6782 104.757
R2386 VDD.n6961 VDD.n6780 104.757
R2387 VDD.n6966 VDD.n6780 104.757
R2388 VDD.n6966 VDD.n6778 104.757
R2389 VDD.n7153 VDD.n6778 104.757
R2390 VDD.n7132 VDD.n6770 104.757
R2391 VDD.n7049 VDD.n6770 104.757
R2392 VDD.n7053 VDD.n7052 104.757
R2393 VDD.n7157 VDD.n6756 104.757
R2394 VDD.n7161 VDD.n6756 104.757
R2395 VDD.n7161 VDD.n6754 104.757
R2396 VDD.n7165 VDD.n6754 104.757
R2397 VDD.n7165 VDD.n6752 104.757
R2398 VDD.n7169 VDD.n6752 104.757
R2399 VDD.n7169 VDD.n6750 104.757
R2400 VDD.n7173 VDD.n6750 104.757
R2401 VDD.n7173 VDD.n6748 104.757
R2402 VDD.n7177 VDD.n6748 104.757
R2403 VDD.n7177 VDD.n6746 104.757
R2404 VDD.n7181 VDD.n6746 104.757
R2405 VDD.n7181 VDD.n6743 104.757
R2406 VDD.n7186 VDD.n6743 104.757
R2407 VDD.n7186 VDD.n6744 104.757
R2408 VDD.n7190 VDD.n6740 104.757
R2409 VDD.n7194 VDD.n6738 104.757
R2410 VDD.n7194 VDD.n6736 104.757
R2411 VDD.n7198 VDD.n6736 104.757
R2412 VDD.n7198 VDD.n6734 104.757
R2413 VDD.n7202 VDD.n6734 104.757
R2414 VDD.n7202 VDD.n6732 104.757
R2415 VDD.n7206 VDD.n6732 104.757
R2416 VDD.n7206 VDD.n6730 104.757
R2417 VDD.n7210 VDD.n6730 104.757
R2418 VDD.n7210 VDD.n6728 104.757
R2419 VDD.n7214 VDD.n6728 104.757
R2420 VDD.n7214 VDD.n6726 104.757
R2421 VDD.n7218 VDD.n6726 104.757
R2422 VDD.n7218 VDD.n6724 104.757
R2423 VDD.n7222 VDD.n6724 104.757
R2424 VDD.n7222 VDD.n6722 104.757
R2425 VDD.n7226 VDD.n6722 104.757
R2426 VDD.n7226 VDD.n6720 104.757
R2427 VDD.n7230 VDD.n6720 104.757
R2428 VDD.n7230 VDD.n6718 104.757
R2429 VDD.n7234 VDD.n6718 104.757
R2430 VDD.n7234 VDD.n6716 104.757
R2431 VDD.n7238 VDD.n6716 104.757
R2432 VDD.n7238 VDD.n6714 104.757
R2433 VDD.n7242 VDD.n6714 104.757
R2434 VDD.n7242 VDD.n6712 104.757
R2435 VDD.n7248 VDD.n6712 104.757
R2436 VDD.n7248 VDD.n6710 104.757
R2437 VDD.n6869 VDD.n6868 104.757
R2438 VDD.n6866 VDD.n6828 104.757
R2439 VDD.n6862 VDD.n6828 104.757
R2440 VDD.n6862 VDD.n6830 104.757
R2441 VDD.n6858 VDD.n6830 104.757
R2442 VDD.n6858 VDD.n6833 104.757
R2443 VDD.n6854 VDD.n6833 104.757
R2444 VDD.n6854 VDD.n6835 104.757
R2445 VDD.n6850 VDD.n6835 104.757
R2446 VDD.n6850 VDD.n6837 104.757
R2447 VDD.n6846 VDD.n6837 104.757
R2448 VDD.n6846 VDD.n6839 104.757
R2449 VDD.n6842 VDD.n6839 104.757
R2450 VDD.n6842 VDD.n6566 104.757
R2451 VDD.n7287 VDD.n6566 104.757
R2452 VDD.n7288 VDD.n7287 104.757
R2453 VDD.n6674 VDD.n6589 104.757
R2454 VDD.n6672 VDD.n6590 104.757
R2455 VDD.n6664 VDD.n6663 104.757
R2456 VDD.n6659 VDD.n6658 104.757
R2457 VDD.n6627 VDD.n6596 104.757
R2458 VDD.n6618 VDD.n6602 104.757
R2459 VDD.n6616 VDD.n6603 104.757
R2460 VDD.n6607 VDD.n6606 104.757
R2461 VDD.n7283 VDD.n6571 104.757
R2462 VDD.n7283 VDD.n6572 104.757
R2463 VDD.n7279 VDD.n6572 104.757
R2464 VDD.n7279 VDD.n6697 104.757
R2465 VDD.n7275 VDD.n6697 104.757
R2466 VDD.n7275 VDD.n6699 104.757
R2467 VDD.n7271 VDD.n6699 104.757
R2468 VDD.n7271 VDD.n6701 104.757
R2469 VDD.n7267 VDD.n6701 104.757
R2470 VDD.n7267 VDD.n6703 104.757
R2471 VDD.n7263 VDD.n6703 104.757
R2472 VDD.n7263 VDD.n6705 104.757
R2473 VDD.n7259 VDD.n6705 104.757
R2474 VDD.n7259 VDD.n6707 104.757
R2475 VDD.n7255 VDD.n6707 104.757
R2476 VDD.n7253 VDD.n7252 104.757
R2477 VDD.n6070 VDD.n5941 104.757
R2478 VDD.n6070 VDD.n5943 104.757
R2479 VDD.n6066 VDD.n5943 104.757
R2480 VDD.n6066 VDD.n5945 104.757
R2481 VDD.n6062 VDD.n5945 104.757
R2482 VDD.n6062 VDD.n5947 104.757
R2483 VDD.n6058 VDD.n5947 104.757
R2484 VDD.n6058 VDD.n5949 104.757
R2485 VDD.n6054 VDD.n5949 104.757
R2486 VDD.n6054 VDD.n5951 104.757
R2487 VDD.n6050 VDD.n5951 104.757
R2488 VDD.n6050 VDD.n5953 104.757
R2489 VDD.n6046 VDD.n5953 104.757
R2490 VDD.n6046 VDD.n5955 104.757
R2491 VDD.n6042 VDD.n5955 104.757
R2492 VDD.n6042 VDD.n5957 104.757
R2493 VDD.n6038 VDD.n5957 104.757
R2494 VDD.n6038 VDD.n5959 104.757
R2495 VDD.n6034 VDD.n5959 104.757
R2496 VDD.n6034 VDD.n5961 104.757
R2497 VDD.n6030 VDD.n5961 104.757
R2498 VDD.n6030 VDD.n5963 104.757
R2499 VDD.n6026 VDD.n5963 104.757
R2500 VDD.n6026 VDD.n5965 104.757
R2501 VDD.n6022 VDD.n5965 104.757
R2502 VDD.n6022 VDD.n5967 104.757
R2503 VDD.n6018 VDD.n5967 104.757
R2504 VDD.n6086 VDD.n5937 104.757
R2505 VDD.n6086 VDD.n5935 104.757
R2506 VDD.n6090 VDD.n5935 104.757
R2507 VDD.n6090 VDD.n5933 104.757
R2508 VDD.n6094 VDD.n5933 104.757
R2509 VDD.n6094 VDD.n5931 104.757
R2510 VDD.n6098 VDD.n5931 104.757
R2511 VDD.n6098 VDD.n5929 104.757
R2512 VDD.n6102 VDD.n5929 104.757
R2513 VDD.n6102 VDD.n5927 104.757
R2514 VDD.n6106 VDD.n5927 104.757
R2515 VDD.n6106 VDD.n5925 104.757
R2516 VDD.n6111 VDD.n5925 104.757
R2517 VDD.n6111 VDD.n5923 104.757
R2518 VDD.n6298 VDD.n5923 104.757
R2519 VDD.n6277 VDD.n5915 104.757
R2520 VDD.n6194 VDD.n5915 104.757
R2521 VDD.n6198 VDD.n6197 104.757
R2522 VDD.n6302 VDD.n5901 104.757
R2523 VDD.n6306 VDD.n5901 104.757
R2524 VDD.n6306 VDD.n5899 104.757
R2525 VDD.n6310 VDD.n5899 104.757
R2526 VDD.n6310 VDD.n5897 104.757
R2527 VDD.n6314 VDD.n5897 104.757
R2528 VDD.n6314 VDD.n5895 104.757
R2529 VDD.n6318 VDD.n5895 104.757
R2530 VDD.n6318 VDD.n5893 104.757
R2531 VDD.n6322 VDD.n5893 104.757
R2532 VDD.n6322 VDD.n5891 104.757
R2533 VDD.n6326 VDD.n5891 104.757
R2534 VDD.n6326 VDD.n5888 104.757
R2535 VDD.n6331 VDD.n5888 104.757
R2536 VDD.n6331 VDD.n5889 104.757
R2537 VDD.n6335 VDD.n5885 104.757
R2538 VDD.n6339 VDD.n5883 104.757
R2539 VDD.n6339 VDD.n5881 104.757
R2540 VDD.n6343 VDD.n5881 104.757
R2541 VDD.n6343 VDD.n5879 104.757
R2542 VDD.n6347 VDD.n5879 104.757
R2543 VDD.n6347 VDD.n5877 104.757
R2544 VDD.n6351 VDD.n5877 104.757
R2545 VDD.n6351 VDD.n5875 104.757
R2546 VDD.n6355 VDD.n5875 104.757
R2547 VDD.n6355 VDD.n5873 104.757
R2548 VDD.n6359 VDD.n5873 104.757
R2549 VDD.n6359 VDD.n5871 104.757
R2550 VDD.n6363 VDD.n5871 104.757
R2551 VDD.n6363 VDD.n5869 104.757
R2552 VDD.n6367 VDD.n5869 104.757
R2553 VDD.n6367 VDD.n5867 104.757
R2554 VDD.n6371 VDD.n5867 104.757
R2555 VDD.n6371 VDD.n5865 104.757
R2556 VDD.n6375 VDD.n5865 104.757
R2557 VDD.n6375 VDD.n5863 104.757
R2558 VDD.n6379 VDD.n5863 104.757
R2559 VDD.n6379 VDD.n5861 104.757
R2560 VDD.n6383 VDD.n5861 104.757
R2561 VDD.n6383 VDD.n5859 104.757
R2562 VDD.n6387 VDD.n5859 104.757
R2563 VDD.n6387 VDD.n5857 104.757
R2564 VDD.n6393 VDD.n5857 104.757
R2565 VDD.n6393 VDD.n5855 104.757
R2566 VDD.n6014 VDD.n6013 104.757
R2567 VDD.n6011 VDD.n5973 104.757
R2568 VDD.n6007 VDD.n5973 104.757
R2569 VDD.n6007 VDD.n5975 104.757
R2570 VDD.n6003 VDD.n5975 104.757
R2571 VDD.n6003 VDD.n5978 104.757
R2572 VDD.n5999 VDD.n5978 104.757
R2573 VDD.n5999 VDD.n5980 104.757
R2574 VDD.n5995 VDD.n5980 104.757
R2575 VDD.n5995 VDD.n5982 104.757
R2576 VDD.n5991 VDD.n5982 104.757
R2577 VDD.n5991 VDD.n5984 104.757
R2578 VDD.n5987 VDD.n5984 104.757
R2579 VDD.n5987 VDD.n5711 104.757
R2580 VDD.n6432 VDD.n5711 104.757
R2581 VDD.n6433 VDD.n6432 104.757
R2582 VDD.n5819 VDD.n5734 104.757
R2583 VDD.n5817 VDD.n5735 104.757
R2584 VDD.n5809 VDD.n5808 104.757
R2585 VDD.n5804 VDD.n5803 104.757
R2586 VDD.n5772 VDD.n5741 104.757
R2587 VDD.n5763 VDD.n5747 104.757
R2588 VDD.n5761 VDD.n5748 104.757
R2589 VDD.n5752 VDD.n5751 104.757
R2590 VDD.n6428 VDD.n5716 104.757
R2591 VDD.n6428 VDD.n5717 104.757
R2592 VDD.n6424 VDD.n5717 104.757
R2593 VDD.n6424 VDD.n5842 104.757
R2594 VDD.n6420 VDD.n5842 104.757
R2595 VDD.n6420 VDD.n5844 104.757
R2596 VDD.n6416 VDD.n5844 104.757
R2597 VDD.n6416 VDD.n5846 104.757
R2598 VDD.n6412 VDD.n5846 104.757
R2599 VDD.n6412 VDD.n5848 104.757
R2600 VDD.n6408 VDD.n5848 104.757
R2601 VDD.n6408 VDD.n5850 104.757
R2602 VDD.n6404 VDD.n5850 104.757
R2603 VDD.n6404 VDD.n5852 104.757
R2604 VDD.n6400 VDD.n5852 104.757
R2605 VDD.n6398 VDD.n6397 104.757
R2606 VDD.n1400 VDD.n1399 104.757
R2607 VDD.n1461 VDD.n1460 104.757
R2608 VDD.n1450 VDD.n1449 104.757
R2609 VDD.n1443 VDD.n1442 104.757
R2610 VDD.n1432 VDD.n1431 104.757
R2611 VDD.n1425 VDD.n1424 104.757
R2612 VDD.n1475 VDD.n1389 104.757
R2613 VDD.n1475 VDD.n1390 104.757
R2614 VDD.n1390 VDD.n1003 104.757
R2615 VDD.n4575 VDD.n1003 104.757
R2616 VDD.n4575 VDD.n1004 104.757
R2617 VDD.n1906 VDD.n1004 104.757
R2618 VDD.n1907 VDD.n1906 104.757
R2619 VDD.n1908 VDD.n1907 104.757
R2620 VDD.n4556 VDD.n1908 104.757
R2621 VDD.n4556 VDD.n1909 104.757
R2622 VDD.n1937 VDD.n1909 104.757
R2623 VDD.n1938 VDD.n1937 104.757
R2624 VDD.n1939 VDD.n1938 104.757
R2625 VDD.n4537 VDD.n1939 104.757
R2626 VDD.n4537 VDD.n1940 104.757
R2627 VDD.n1969 VDD.n1940 104.757
R2628 VDD.n1969 VDD.n1958 104.757
R2629 VDD.n4522 VDD.n1958 104.757
R2630 VDD.n4522 VDD.n4521 104.757
R2631 VDD.n4521 VDD.n1959 104.757
R2632 VDD.n4512 VDD.n1959 104.757
R2633 VDD.n4512 VDD.n1978 104.757
R2634 VDD.n2009 VDD.n1978 104.757
R2635 VDD.n2010 VDD.n2009 104.757
R2636 VDD.n2011 VDD.n2010 104.757
R2637 VDD.n4493 VDD.n2011 104.757
R2638 VDD.n4493 VDD.n2012 104.757
R2639 VDD.n2042 VDD.n2012 104.757
R2640 VDD.n2043 VDD.n2042 104.757
R2641 VDD.n2044 VDD.n2043 104.757
R2642 VDD.n4474 VDD.n2044 104.757
R2643 VDD.n4474 VDD.n2045 104.757
R2644 VDD.n2091 VDD.n2045 104.757
R2645 VDD.n2092 VDD.n2091 104.757
R2646 VDD.n2093 VDD.n2092 104.757
R2647 VDD.n2094 VDD.n2093 104.757
R2648 VDD.n2095 VDD.n2094 104.757
R2649 VDD.n2096 VDD.n2095 104.757
R2650 VDD.n2097 VDD.n2096 104.757
R2651 VDD.n4440 VDD.n2097 104.757
R2652 VDD.n4440 VDD.n2098 104.757
R2653 VDD.n2126 VDD.n2098 104.757
R2654 VDD.n2127 VDD.n2126 104.757
R2655 VDD.n2128 VDD.n2127 104.757
R2656 VDD.n4421 VDD.n2128 104.757
R2657 VDD.n4421 VDD.n2129 104.757
R2658 VDD.n2157 VDD.n2129 104.757
R2659 VDD.n2158 VDD.n2157 104.757
R2660 VDD.n2159 VDD.n2158 104.757
R2661 VDD.n4402 VDD.n2159 104.757
R2662 VDD.n4402 VDD.n2160 104.757
R2663 VDD.n2190 VDD.n2160 104.757
R2664 VDD.n2190 VDD.n2179 104.757
R2665 VDD.n4387 VDD.n2179 104.757
R2666 VDD.n4387 VDD.n4386 104.757
R2667 VDD.n4386 VDD.n2180 104.757
R2668 VDD.n4377 VDD.n2180 104.757
R2669 VDD.n4377 VDD.n2199 104.757
R2670 VDD.n2230 VDD.n2199 104.757
R2671 VDD.n2231 VDD.n2230 104.757
R2672 VDD.n2232 VDD.n2231 104.757
R2673 VDD.n4358 VDD.n2232 104.757
R2674 VDD.n4358 VDD.n2233 104.757
R2675 VDD.n2470 VDD.n2469 104.757
R2676 VDD.n2466 VDD.n2463 104.757
R2677 VDD.n4022 VDD.n2365 104.757
R2678 VDD.n4288 VDD.n2365 104.757
R2679 VDD.n4288 VDD.n2366 104.757
R2680 VDD.n4284 VDD.n2366 104.757
R2681 VDD.n4284 VDD.n2369 104.757
R2682 VDD.n4277 VDD.n2369 104.757
R2683 VDD.n4277 VDD.n2374 104.757
R2684 VDD.n4273 VDD.n2374 104.757
R2685 VDD.n4273 VDD.n2376 104.757
R2686 VDD.n4266 VDD.n2376 104.757
R2687 VDD.n4266 VDD.n2383 104.757
R2688 VDD.n4262 VDD.n2383 104.757
R2689 VDD.n4262 VDD.n2385 104.757
R2690 VDD.n4255 VDD.n2385 104.757
R2691 VDD.n4255 VDD.n2392 104.757
R2692 VDD.n4251 VDD.n2392 104.757
R2693 VDD.n4251 VDD.n2394 104.757
R2694 VDD.n4244 VDD.n2394 104.757
R2695 VDD.n4244 VDD.n2401 104.757
R2696 VDD.n4240 VDD.n2401 104.757
R2697 VDD.n4240 VDD.n2402 104.757
R2698 VDD.n2409 VDD.n2402 104.757
R2699 VDD.n4232 VDD.n2409 104.757
R2700 VDD.n4232 VDD.n2410 104.757
R2701 VDD.n4228 VDD.n2410 104.757
R2702 VDD.n4228 VDD.n2414 104.757
R2703 VDD.n4221 VDD.n2414 104.757
R2704 VDD.n4221 VDD.n2421 104.757
R2705 VDD.n4217 VDD.n2421 104.757
R2706 VDD.n4217 VDD.n2423 104.757
R2707 VDD.n4210 VDD.n2423 104.757
R2708 VDD.n4210 VDD.n2430 104.757
R2709 VDD.n4206 VDD.n2430 104.757
R2710 VDD.n4206 VDD.n2432 104.757
R2711 VDD.n4199 VDD.n2432 104.757
R2712 VDD.n4199 VDD.n2439 104.757
R2713 VDD.n4083 VDD.n2439 104.757
R2714 VDD.n4093 VDD.n4083 104.757
R2715 VDD.n4093 VDD.n4081 104.757
R2716 VDD.n4097 VDD.n4081 104.757
R2717 VDD.n4097 VDD.n4076 104.757
R2718 VDD.n4106 VDD.n4076 104.757
R2719 VDD.n4106 VDD.n4074 104.757
R2720 VDD.n4110 VDD.n4074 104.757
R2721 VDD.n4110 VDD.n4069 104.757
R2722 VDD.n4119 VDD.n4069 104.757
R2723 VDD.n4119 VDD.n4067 104.757
R2724 VDD.n4124 VDD.n4067 104.757
R2725 VDD.n4124 VDD.n4062 104.757
R2726 VDD.n4133 VDD.n4062 104.757
R2727 VDD.n4133 VDD.n4061 104.757
R2728 VDD.n4137 VDD.n4061 104.757
R2729 VDD.n4137 VDD.n4057 104.757
R2730 VDD.n4145 VDD.n4057 104.757
R2731 VDD.n4145 VDD.n4055 104.757
R2732 VDD.n4149 VDD.n4055 104.757
R2733 VDD.n4149 VDD.n4049 104.757
R2734 VDD.n4157 VDD.n4049 104.757
R2735 VDD.n4157 VDD.n4047 104.757
R2736 VDD.n4161 VDD.n4047 104.757
R2737 VDD.n4161 VDD.n4042 104.757
R2738 VDD.n4170 VDD.n4042 104.757
R2739 VDD.n4170 VDD.n4040 104.757
R2740 VDD.n4174 VDD.n4040 104.757
R2741 VDD.n4174 VDD.n4035 104.757
R2742 VDD.n4183 VDD.n4035 104.757
R2743 VDD.n4183 VDD.n4032 104.757
R2744 VDD.n4188 VDD.n4032 104.757
R2745 VDD.n4188 VDD.n4033 104.757
R2746 VDD.n4033 VDD.n271 104.757
R2747 VDD.n5458 VDD.n271 104.757
R2748 VDD.n5458 VDD.n272 104.757
R2749 VDD.n5441 VDD.n272 104.757
R2750 VDD.n5444 VDD.n5441 104.757
R2751 VDD.n1470 VDD.n1376 104.757
R2752 VDD.n1482 VDD.n1376 104.757
R2753 VDD.n1483 VDD.n1482 104.757
R2754 VDD.n1483 VDD.n1370 104.757
R2755 VDD.n1495 VDD.n1370 104.757
R2756 VDD.n1495 VDD.n1363 104.757
R2757 VDD.n1503 VDD.n1363 104.757
R2758 VDD.n1503 VDD.n1354 104.757
R2759 VDD.n1514 VDD.n1354 104.757
R2760 VDD.n1515 VDD.n1514 104.757
R2761 VDD.n1515 VDD.n1348 104.757
R2762 VDD.n1527 VDD.n1348 104.757
R2763 VDD.n1527 VDD.n1342 104.757
R2764 VDD.n1539 VDD.n1342 104.757
R2765 VDD.n1539 VDD.n1335 104.757
R2766 VDD.n1547 VDD.n1335 104.757
R2767 VDD.n1547 VDD.n1326 104.757
R2768 VDD.n1558 VDD.n1326 104.757
R2769 VDD.n1559 VDD.n1558 104.757
R2770 VDD.n1559 VDD.n1319 104.757
R2771 VDD.n1570 VDD.n1319 104.757
R2772 VDD.n1570 VDD.n1312 104.757
R2773 VDD.n1578 VDD.n1312 104.757
R2774 VDD.n1578 VDD.n1303 104.757
R2775 VDD.n1589 VDD.n1303 104.757
R2776 VDD.n1590 VDD.n1589 104.757
R2777 VDD.n1590 VDD.n1297 104.757
R2778 VDD.n1602 VDD.n1297 104.757
R2779 VDD.n1602 VDD.n1291 104.757
R2780 VDD.n1614 VDD.n1291 104.757
R2781 VDD.n1614 VDD.n1278 104.757
R2782 VDD.n1813 VDD.n1278 104.757
R2783 VDD.n1813 VDD.n1279 104.757
R2784 VDD.n1803 VDD.n1279 104.757
R2785 VDD.n1803 VDD.n1802 104.757
R2786 VDD.n1802 VDD.n1624 104.757
R2787 VDD.n1640 VDD.n1624 104.757
R2788 VDD.n1788 VDD.n1640 104.757
R2789 VDD.n1788 VDD.n1787 104.757
R2790 VDD.n1787 VDD.n1641 104.757
R2791 VDD.n1656 VDD.n1641 104.757
R2792 VDD.n1774 VDD.n1656 104.757
R2793 VDD.n1774 VDD.n1773 104.757
R2794 VDD.n1773 VDD.n1657 104.757
R2795 VDD.n1673 VDD.n1657 104.757
R2796 VDD.n1759 VDD.n1673 104.757
R2797 VDD.n1759 VDD.n1758 104.757
R2798 VDD.n1758 VDD.n1674 104.757
R2799 VDD.n1690 VDD.n1674 104.757
R2800 VDD.n1744 VDD.n1690 104.757
R2801 VDD.n1744 VDD.n1743 104.757
R2802 VDD.n1743 VDD.n1691 104.757
R2803 VDD.n1728 VDD.n1691 104.757
R2804 VDD.n1729 VDD.n1728 104.757
R2805 VDD.n1729 VDD.n1044 104.757
R2806 VDD.n1882 VDD.n1044 104.757
R2807 VDD.n1882 VDD.n1045 104.757
R2808 VDD.n1875 VDD.n1045 104.757
R2809 VDD.n1875 VDD.n1051 104.757
R2810 VDD.n1871 VDD.n1051 104.757
R2811 VDD.n1871 VDD.n1053 104.757
R2812 VDD.n1864 VDD.n1053 104.757
R2813 VDD.n1864 VDD.n1058 104.757
R2814 VDD.n1818 VDD.n1817 104.757
R2815 VDD.n1165 VDD.n1000 104.757
R2816 VDD.n4580 VDD.n1000 104.757
R2817 VDD.n4580 VDD.n995 104.757
R2818 VDD.n4589 VDD.n995 104.757
R2819 VDD.n4589 VDD.n993 104.757
R2820 VDD.n4593 VDD.n993 104.757
R2821 VDD.n4593 VDD.n989 104.757
R2822 VDD.n4601 VDD.n989 104.757
R2823 VDD.n4601 VDD.n987 104.757
R2824 VDD.n4605 VDD.n987 104.757
R2825 VDD.n4605 VDD.n981 104.757
R2826 VDD.n4612 VDD.n981 104.757
R2827 VDD.n4612 VDD.n979 104.757
R2828 VDD.n4616 VDD.n979 104.757
R2829 VDD.n4616 VDD.n974 104.757
R2830 VDD.n4625 VDD.n974 104.757
R2831 VDD.n4625 VDD.n972 104.757
R2832 VDD.n4629 VDD.n972 104.757
R2833 VDD.n4629 VDD.n967 104.757
R2834 VDD.n4638 VDD.n967 104.757
R2835 VDD.n4638 VDD.n965 104.757
R2836 VDD.n4642 VDD.n965 104.757
R2837 VDD.n4642 VDD.n960 104.757
R2838 VDD.n4651 VDD.n960 104.757
R2839 VDD.n4651 VDD.n958 104.757
R2840 VDD.n4655 VDD.n958 104.757
R2841 VDD.n4655 VDD.n953 104.757
R2842 VDD.n4661 VDD.n953 104.757
R2843 VDD.n4661 VDD.n951 104.757
R2844 VDD.n4665 VDD.n951 104.757
R2845 VDD.n4665 VDD.n946 104.757
R2846 VDD.n4674 VDD.n946 104.757
R2847 VDD.n4674 VDD.n944 104.757
R2848 VDD.n4678 VDD.n944 104.757
R2849 VDD.n4678 VDD.n939 104.757
R2850 VDD.n4687 VDD.n939 104.757
R2851 VDD.n4687 VDD.n937 104.757
R2852 VDD.n4691 VDD.n937 104.757
R2853 VDD.n4691 VDD.n932 104.757
R2854 VDD.n4700 VDD.n932 104.757
R2855 VDD.n4700 VDD.n930 104.757
R2856 VDD.n4704 VDD.n930 104.757
R2857 VDD.n4704 VDD.n923 104.757
R2858 VDD.n4713 VDD.n923 104.757
R2859 VDD.n4713 VDD.n926 104.757
R2860 VDD.n4716 VDD.n914 104.757
R2861 VDD.n4730 VDD.n914 104.757
R2862 VDD.n4730 VDD.n912 104.757
R2863 VDD.n4734 VDD.n912 104.757
R2864 VDD.n4734 VDD.n907 104.757
R2865 VDD.n4743 VDD.n907 104.757
R2866 VDD.n4743 VDD.n905 104.757
R2867 VDD.n4747 VDD.n905 104.757
R2868 VDD.n4747 VDD.n900 104.757
R2869 VDD.n4754 VDD.n900 104.757
R2870 VDD.n4754 VDD.n898 104.757
R2871 VDD.n4758 VDD.n898 104.757
R2872 VDD.n4758 VDD.n893 104.757
R2873 VDD.n4767 VDD.n893 104.757
R2874 VDD.n4767 VDD.n891 104.757
R2875 VDD.n4771 VDD.n891 104.757
R2876 VDD.n4771 VDD.n886 104.757
R2877 VDD.n4780 VDD.n886 104.757
R2878 VDD.n4780 VDD.n884 104.757
R2879 VDD.n4784 VDD.n884 104.757
R2880 VDD.n4784 VDD.n879 104.757
R2881 VDD.n4793 VDD.n879 104.757
R2882 VDD.n4793 VDD.n877 104.757
R2883 VDD.n4797 VDD.n877 104.757
R2884 VDD.n4797 VDD.n873 104.757
R2885 VDD.n4805 VDD.n873 104.757
R2886 VDD.n4805 VDD.n871 104.757
R2887 VDD.n4809 VDD.n871 104.757
R2888 VDD.n4809 VDD.n866 104.757
R2889 VDD.n4818 VDD.n866 104.757
R2890 VDD.n4818 VDD.n864 104.757
R2891 VDD.n4822 VDD.n864 104.757
R2892 VDD.n4822 VDD.n859 104.757
R2893 VDD.n4831 VDD.n859 104.757
R2894 VDD.n4831 VDD.n857 104.757
R2895 VDD.n4835 VDD.n857 104.757
R2896 VDD.n4835 VDD.n852 104.757
R2897 VDD.n4844 VDD.n852 104.757
R2898 VDD.n4844 VDD.n850 104.757
R2899 VDD.n4848 VDD.n850 104.757
R2900 VDD.n4848 VDD.n845 104.757
R2901 VDD.n4857 VDD.n845 104.757
R2902 VDD.n4857 VDD.n843 104.757
R2903 VDD.n4861 VDD.n843 104.757
R2904 VDD.n4861 VDD.n838 104.757
R2905 VDD.n4868 VDD.n838 104.757
R2906 VDD.n4868 VDD.n836 104.757
R2907 VDD.n4872 VDD.n836 104.757
R2908 VDD.n4872 VDD.n831 104.757
R2909 VDD.n4881 VDD.n831 104.757
R2910 VDD.n4881 VDD.n829 104.757
R2911 VDD.n4885 VDD.n829 104.757
R2912 VDD.n4885 VDD.n824 104.757
R2913 VDD.n4894 VDD.n824 104.757
R2914 VDD.n4894 VDD.n822 104.757
R2915 VDD.n4898 VDD.n822 104.757
R2916 VDD.n4898 VDD.n817 104.757
R2917 VDD.n4907 VDD.n817 104.757
R2918 VDD.n4907 VDD.n815 104.757
R2919 VDD.n4911 VDD.n815 104.757
R2920 VDD.n4911 VDD.n811 104.757
R2921 VDD.n4919 VDD.n811 104.757
R2922 VDD.n4919 VDD.n809 104.757
R2923 VDD.n4923 VDD.n809 104.757
R2924 VDD.n4923 VDD.n804 104.757
R2925 VDD.n4932 VDD.n804 104.757
R2926 VDD.n4932 VDD.n802 104.757
R2927 VDD.n4936 VDD.n802 104.757
R2928 VDD.n4936 VDD.n797 104.757
R2929 VDD.n4945 VDD.n797 104.757
R2930 VDD.n4945 VDD.n795 104.757
R2931 VDD.n4949 VDD.n795 104.757
R2932 VDD.n4949 VDD.n790 104.757
R2933 VDD.n4958 VDD.n790 104.757
R2934 VDD.n4958 VDD.n788 104.757
R2935 VDD.n4962 VDD.n788 104.757
R2936 VDD.n4962 VDD.n783 104.757
R2937 VDD.n4971 VDD.n783 104.757
R2938 VDD.n4971 VDD.n781 104.757
R2939 VDD.n4975 VDD.n781 104.757
R2940 VDD.n4975 VDD.n776 104.757
R2941 VDD.n4982 VDD.n776 104.757
R2942 VDD.n4982 VDD.n774 104.757
R2943 VDD.n4986 VDD.n774 104.757
R2944 VDD.n4986 VDD.n769 104.757
R2945 VDD.n4995 VDD.n769 104.757
R2946 VDD.n4995 VDD.n767 104.757
R2947 VDD.n4999 VDD.n767 104.757
R2948 VDD.n4999 VDD.n762 104.757
R2949 VDD.n5008 VDD.n762 104.757
R2950 VDD.n5008 VDD.n760 104.757
R2951 VDD.n5012 VDD.n760 104.757
R2952 VDD.n5012 VDD.n755 104.757
R2953 VDD.n5021 VDD.n755 104.757
R2954 VDD.n5021 VDD.n753 104.757
R2955 VDD.n5025 VDD.n753 104.757
R2956 VDD.n5025 VDD.n749 104.757
R2957 VDD.n5033 VDD.n749 104.757
R2958 VDD.n5033 VDD.n747 104.757
R2959 VDD.n5037 VDD.n747 104.757
R2960 VDD.n5037 VDD.n742 104.757
R2961 VDD.n5046 VDD.n742 104.757
R2962 VDD.n5046 VDD.n740 104.757
R2963 VDD.n5050 VDD.n740 104.757
R2964 VDD.n5050 VDD.n735 104.757
R2965 VDD.n5059 VDD.n735 104.757
R2966 VDD.n5059 VDD.n733 104.757
R2967 VDD.n5063 VDD.n733 104.757
R2968 VDD.n5063 VDD.n728 104.757
R2969 VDD.n5072 VDD.n728 104.757
R2970 VDD.n5072 VDD.n726 104.757
R2971 VDD.n5076 VDD.n726 104.757
R2972 VDD.n5076 VDD.n721 104.757
R2973 VDD.n5085 VDD.n721 104.757
R2974 VDD.n5085 VDD.n719 104.757
R2975 VDD.n5089 VDD.n719 104.757
R2976 VDD.n5089 VDD.n714 104.757
R2977 VDD.n5096 VDD.n714 104.757
R2978 VDD.n5096 VDD.n712 104.757
R2979 VDD.n5100 VDD.n712 104.757
R2980 VDD.n5100 VDD.n707 104.757
R2981 VDD.n5109 VDD.n707 104.757
R2982 VDD.n5109 VDD.n705 104.757
R2983 VDD.n5113 VDD.n705 104.757
R2984 VDD.n5113 VDD.n700 104.757
R2985 VDD.n5122 VDD.n700 104.757
R2986 VDD.n5122 VDD.n698 104.757
R2987 VDD.n5126 VDD.n698 104.757
R2988 VDD.n5126 VDD.n693 104.757
R2989 VDD.n5135 VDD.n693 104.757
R2990 VDD.n5135 VDD.n691 104.757
R2991 VDD.n5139 VDD.n691 104.757
R2992 VDD.n5139 VDD.n687 104.757
R2993 VDD.n5147 VDD.n687 104.757
R2994 VDD.n5147 VDD.n684 104.757
R2995 VDD.n5152 VDD.n684 104.757
R2996 VDD.n5152 VDD.n685 104.757
R2997 VDD.n685 VDD.n680 104.757
R2998 VDD.n5451 VDD.n279 104.757
R2999 VDD.n5438 VDD.n280 104.757
R3000 VDD.n5431 VDD.n295 104.757
R3001 VDD.n5428 VDD.n5427 104.757
R3002 VDD.n5420 VDD.n5419 104.757
R3003 VDD.n5416 VDD.n5415 104.757
R3004 VDD.n5408 VDD.n5407 104.757
R3005 VDD.n5404 VDD.n5403 104.757
R3006 VDD.n314 VDD.n313 104.757
R3007 VDD.n5396 VDD.n5395 104.757
R3008 VDD.n5388 VDD.n5387 104.757
R3009 VDD.n5384 VDD.n5383 104.757
R3010 VDD.n5376 VDD.n5375 104.757
R3011 VDD.n5372 VDD.n5371 104.757
R3012 VDD.n5364 VDD.n328 104.757
R3013 VDD.n5364 VDD.n329 104.757
R3014 VDD.n5360 VDD.n329 104.757
R3015 VDD.n5360 VDD.n331 104.757
R3016 VDD.n5353 VDD.n331 104.757
R3017 VDD.n5353 VDD.n338 104.757
R3018 VDD.n5349 VDD.n338 104.757
R3019 VDD.n5349 VDD.n340 104.757
R3020 VDD.n5342 VDD.n340 104.757
R3021 VDD.n5342 VDD.n345 104.757
R3022 VDD.n5338 VDD.n345 104.757
R3023 VDD.n5338 VDD.n347 104.757
R3024 VDD.n5331 VDD.n347 104.757
R3025 VDD.n5331 VDD.n354 104.757
R3026 VDD.n5327 VDD.n354 104.757
R3027 VDD.n5327 VDD.n356 104.757
R3028 VDD.n5320 VDD.n356 104.757
R3029 VDD.n5320 VDD.n363 104.757
R3030 VDD.n5316 VDD.n363 104.757
R3031 VDD.n5316 VDD.n365 104.757
R3032 VDD.n5309 VDD.n365 104.757
R3033 VDD.n5309 VDD.n372 104.757
R3034 VDD.n5305 VDD.n372 104.757
R3035 VDD.n5305 VDD.n374 104.757
R3036 VDD.n382 VDD.n374 104.757
R3037 VDD.n5298 VDD.n382 104.757
R3038 VDD.n5298 VDD.n383 104.757
R3039 VDD.n5294 VDD.n383 104.757
R3040 VDD.n5294 VDD.n386 104.757
R3041 VDD.n5287 VDD.n386 104.757
R3042 VDD.n5287 VDD.n393 104.757
R3043 VDD.n458 VDD.n456 104.757
R3044 VDD.n465 VDD.n447 104.757
R3045 VDD.n468 VDD.n467 104.757
R3046 VDD.n477 VDD.n475 104.757
R3047 VDD.n485 VDD.n439 104.757
R3048 VDD.n489 VDD.n487 104.757
R3049 VDD.n496 VDD.n435 104.757
R3050 VDD.n499 VDD.n498 104.757
R3051 VDD.n508 VDD.n506 104.757
R3052 VDD.n515 VDD.n427 104.757
R3053 VDD.n518 VDD.n517 104.757
R3054 VDD.n527 VDD.n525 104.757
R3055 VDD.n534 VDD.n419 104.757
R3056 VDD.n538 VDD.n537 104.757
R3057 VDD.n546 VDD.n415 104.757
R3058 VDD.n549 VDD.n548 104.757
R3059 VDD.n558 VDD.n556 104.757
R3060 VDD.n565 VDD.n407 104.757
R3061 VDD.n568 VDD.n567 104.757
R3062 VDD.n577 VDD.n575 104.757
R3063 VDD.n5283 VDD.n397 104.757
R3064 VDD.n5283 VDD.n398 104.757
R3065 VDD.n5276 VDD.n398 104.757
R3066 VDD.n5276 VDD.n585 104.757
R3067 VDD.n5272 VDD.n585 104.757
R3068 VDD.n5272 VDD.n587 104.757
R3069 VDD.n595 VDD.n587 104.757
R3070 VDD.n5265 VDD.n595 104.757
R3071 VDD.n5265 VDD.n596 104.757
R3072 VDD.n5261 VDD.n596 104.757
R3073 VDD.n5261 VDD.n599 104.757
R3074 VDD.n5254 VDD.n599 104.757
R3075 VDD.n5254 VDD.n606 104.757
R3076 VDD.n5250 VDD.n606 104.757
R3077 VDD.n5250 VDD.n608 104.757
R3078 VDD.n5243 VDD.n608 104.757
R3079 VDD.n5243 VDD.n615 104.757
R3080 VDD.n5239 VDD.n615 104.757
R3081 VDD.n5239 VDD.n617 104.757
R3082 VDD.n5232 VDD.n617 104.757
R3083 VDD.n5232 VDD.n624 104.757
R3084 VDD.n5228 VDD.n624 104.757
R3085 VDD.n5228 VDD.n626 104.757
R3086 VDD.n5221 VDD.n626 104.757
R3087 VDD.n5221 VDD.n633 104.757
R3088 VDD.n5217 VDD.n633 104.757
R3089 VDD.n5217 VDD.n635 104.757
R3090 VDD.n5210 VDD.n635 104.757
R3091 VDD.n5210 VDD.n640 104.757
R3092 VDD.n5206 VDD.n640 104.757
R3093 VDD.n5206 VDD.n642 104.757
R3094 VDD.n5199 VDD.n642 104.757
R3095 VDD.n5199 VDD.n649 104.757
R3096 VDD.n5195 VDD.n649 104.757
R3097 VDD.n5195 VDD.n651 104.757
R3098 VDD.n5188 VDD.n651 104.757
R3099 VDD.n5188 VDD.n658 104.757
R3100 VDD.n5184 VDD.n658 104.757
R3101 VDD.n5184 VDD.n660 104.757
R3102 VDD.n5177 VDD.n660 104.757
R3103 VDD.n5177 VDD.n667 104.757
R3104 VDD.n5173 VDD.n667 104.757
R3105 VDD.n5173 VDD.n669 104.757
R3106 VDD.n676 VDD.n669 104.757
R3107 VDD.n5165 VDD.n676 104.757
R3108 VDD.n5165 VDD.n677 104.757
R3109 VDD.n5363 VDD.n281 99.5243
R3110 VDD.n2612 VDD.n2611 98.9686
R3111 VDD.n8582 VDD.n8581 96.8641
R3112 VDD.n7727 VDD.n7726 96.8641
R3113 VDD.n6873 VDD.n6872 96.8641
R3114 VDD.n6018 VDD.n6017 96.8641
R3115 VDD.t70 VDD.n5641 96.8274
R3116 VDD.n6489 VDD.t146 96.8274
R3117 VDD.t16 VDD.n7350 96.8274
R3118 VDD.n8198 VDD.t63 96.8274
R3119 VDD.n8540 VDD.n8532 96.5084
R3120 VDD.n8649 VDD.n8648 96.5084
R3121 VDD.n7685 VDD.n7677 96.5084
R3122 VDD.n7794 VDD.n7793 96.5084
R3123 VDD.n6831 VDD.n6823 96.5084
R3124 VDD.n6940 VDD.n6939 96.5084
R3125 VDD.n5976 VDD.n5968 96.5084
R3126 VDD.n6085 VDD.n6084 96.5084
R3127 VDD.n8681 VDD.n8678 92.5005
R3128 VDD.n8837 VDD.n8681 92.5005
R3129 VDD.n9002 VDD.n8269 92.5005
R3130 VDD.n8389 VDD.n8269 92.5005
R3131 VDD.n9004 VDD.n9003 92.5005
R3132 VDD.n9005 VDD.n9004 92.5005
R3133 VDD.n8270 VDD.n8268 92.5005
R3134 VDD.n8268 VDD.n8260 92.5005
R3135 VDD.n8727 VDD.n8726 92.5005
R3136 VDD.n8727 VDD.n8259 92.5005
R3137 VDD.n8728 VDD.n8725 92.5005
R3138 VDD.n8728 VDD.n8252 92.5005
R3139 VDD.n8730 VDD.n8729 92.5005
R3140 VDD.n8729 VDD.n8251 92.5005
R3141 VDD.n8743 VDD.n8723 92.5005
R3142 VDD.n8742 VDD.n8741 92.5005
R3143 VDD.n8740 VDD.n8739 92.5005
R3144 VDD.n8738 VDD.n8737 92.5005
R3145 VDD.n8736 VDD.n8735 92.5005
R3146 VDD.n8745 VDD.n8744 92.5005
R3147 VDD.n8707 VDD.n8706 92.5005
R3148 VDD.n8720 VDD.n8707 92.5005
R3149 VDD.n8825 VDD.n8824 92.5005
R3150 VDD.n8824 VDD.n8823 92.5005
R3151 VDD.n8826 VDD.n8704 92.5005
R3152 VDD.n8708 VDD.n8704 92.5005
R3153 VDD.n8828 VDD.n8827 92.5005
R3154 VDD.n8829 VDD.n8828 92.5005
R3155 VDD.n8705 VDD.n8703 92.5005
R3156 VDD.n8703 VDD.n8695 92.5005
R3157 VDD.n8868 VDD.n8465 92.5005
R3158 VDD.n8465 VDD.n8464 92.5005
R3159 VDD.n8891 VDD.n8890 92.5005
R3160 VDD.n8890 VDD.n8889 92.5005
R3161 VDD.n8455 VDD.n8454 92.5005
R3162 VDD.n8888 VDD.n8455 92.5005
R3163 VDD.n8886 VDD.n8885 92.5005
R3164 VDD.n8887 VDD.n8886 92.5005
R3165 VDD.n8884 VDD.n8457 92.5005
R3166 VDD.n8457 VDD.n8456 92.5005
R3167 VDD.n8883 VDD.n8882 92.5005
R3168 VDD.n8882 VDD.n8881 92.5005
R3169 VDD.n8459 VDD.n8458 92.5005
R3170 VDD.n8880 VDD.n8459 92.5005
R3171 VDD.n8878 VDD.n8877 92.5005
R3172 VDD.n8879 VDD.n8878 92.5005
R3173 VDD.n8876 VDD.n8461 92.5005
R3174 VDD.n8461 VDD.n8460 92.5005
R3175 VDD.n8875 VDD.n8874 92.5005
R3176 VDD.n8874 VDD.n8873 92.5005
R3177 VDD.n8463 VDD.n8462 92.5005
R3178 VDD.n8872 VDD.n8463 92.5005
R3179 VDD.n8870 VDD.n8869 92.5005
R3180 VDD.n8871 VDD.n8870 92.5005
R3181 VDD.n8892 VDD.n8452 92.5005
R3182 VDD.n8452 VDD.n8451 92.5005
R3183 VDD.n8895 VDD.n8894 92.5005
R3184 VDD.n8896 VDD.n8895 92.5005
R3185 VDD.n8893 VDD.n8453 92.5005
R3186 VDD.n8449 VDD.n8448 92.5005
R3187 VDD.n8900 VDD.n8899 92.5005
R3188 VDD.n8899 VDD.n8898 92.5005
R3189 VDD.n8903 VDD.n8902 92.5005
R3190 VDD.n8904 VDD.n8903 92.5005
R3191 VDD.n8445 VDD.n8444 92.5005
R3192 VDD.n8905 VDD.n8445 92.5005
R3193 VDD.n8908 VDD.n8907 92.5005
R3194 VDD.n8907 VDD.n8906 92.5005
R3195 VDD.n8909 VDD.n8443 92.5005
R3196 VDD.n8443 VDD.n8442 92.5005
R3197 VDD.n8911 VDD.n8910 92.5005
R3198 VDD.n8912 VDD.n8911 92.5005
R3199 VDD.n8441 VDD.n8440 92.5005
R3200 VDD.n8913 VDD.n8441 92.5005
R3201 VDD.n8916 VDD.n8915 92.5005
R3202 VDD.n8915 VDD.n8914 92.5005
R3203 VDD.n8917 VDD.n8439 92.5005
R3204 VDD.n8439 VDD.n8438 92.5005
R3205 VDD.n8919 VDD.n8918 92.5005
R3206 VDD.n8920 VDD.n8919 92.5005
R3207 VDD.n8437 VDD.n8436 92.5005
R3208 VDD.n8921 VDD.n8437 92.5005
R3209 VDD.n8924 VDD.n8923 92.5005
R3210 VDD.n8923 VDD.n8922 92.5005
R3211 VDD.n8925 VDD.n8435 92.5005
R3212 VDD.n8435 VDD.n8434 92.5005
R3213 VDD.n8927 VDD.n8926 92.5005
R3214 VDD.n8928 VDD.n8927 92.5005
R3215 VDD.n8433 VDD.n8432 92.5005
R3216 VDD.n8929 VDD.n8433 92.5005
R3217 VDD.n8932 VDD.n8931 92.5005
R3218 VDD.n8931 VDD.n8930 92.5005
R3219 VDD.n8933 VDD.n8431 92.5005
R3220 VDD.n8431 VDD.n8430 92.5005
R3221 VDD.n8935 VDD.n8934 92.5005
R3222 VDD.n8936 VDD.n8935 92.5005
R3223 VDD.n8429 VDD.n8428 92.5005
R3224 VDD.n8937 VDD.n8429 92.5005
R3225 VDD.n8940 VDD.n8939 92.5005
R3226 VDD.n8939 VDD.n8938 92.5005
R3227 VDD.n8941 VDD.n8427 92.5005
R3228 VDD.n8427 VDD.n8426 92.5005
R3229 VDD.n8943 VDD.n8942 92.5005
R3230 VDD.n8944 VDD.n8943 92.5005
R3231 VDD.n8425 VDD.n8424 92.5005
R3232 VDD.n8945 VDD.n8425 92.5005
R3233 VDD.n8948 VDD.n8947 92.5005
R3234 VDD.n8947 VDD.n8946 92.5005
R3235 VDD.n8949 VDD.n8423 92.5005
R3236 VDD.n8423 VDD.n8422 92.5005
R3237 VDD.n8951 VDD.n8950 92.5005
R3238 VDD.n8952 VDD.n8951 92.5005
R3239 VDD.n8421 VDD.n8420 92.5005
R3240 VDD.n8953 VDD.n8421 92.5005
R3241 VDD.n8958 VDD.n8957 92.5005
R3242 VDD.n8957 VDD.n8956 92.5005
R3243 VDD.n8959 VDD.n8419 92.5005
R3244 VDD.n8955 VDD.n8419 92.5005
R3245 VDD.n8901 VDD.n8447 92.5005
R3246 VDD.n8447 VDD.n8446 92.5005
R3247 VDD.n8973 VDD.n8972 92.5005
R3248 VDD.n8972 VDD.n8971 92.5005
R3249 VDD.n8974 VDD.n8412 92.5005
R3250 VDD.n8412 VDD.n8411 92.5005
R3251 VDD.n8976 VDD.n8975 92.5005
R3252 VDD.n8977 VDD.n8976 92.5005
R3253 VDD.n8410 VDD.n8409 92.5005
R3254 VDD.n8978 VDD.n8410 92.5005
R3255 VDD.n8981 VDD.n8980 92.5005
R3256 VDD.n8980 VDD.n8979 92.5005
R3257 VDD.n8982 VDD.n8408 92.5005
R3258 VDD.n8408 VDD.n8407 92.5005
R3259 VDD.n8984 VDD.n8983 92.5005
R3260 VDD.n8985 VDD.n8984 92.5005
R3261 VDD.n8406 VDD.n8405 92.5005
R3262 VDD.n8986 VDD.n8406 92.5005
R3263 VDD.n8989 VDD.n8988 92.5005
R3264 VDD.n8988 VDD.n8987 92.5005
R3265 VDD.n8990 VDD.n8281 92.5005
R3266 VDD.n8281 VDD.n8279 92.5005
R3267 VDD.n8992 VDD.n8991 92.5005
R3268 VDD.n8993 VDD.n8992 92.5005
R3269 VDD.n8968 VDD.n8967 92.5005
R3270 VDD.n8969 VDD.n8968 92.5005
R3271 VDD.n8966 VDD.n8416 92.5005
R3272 VDD.n8416 VDD.n8415 92.5005
R3273 VDD.n8965 VDD.n8964 92.5005
R3274 VDD.n8962 VDD.n8417 92.5005
R3275 VDD.n8961 VDD.n8960 92.5005
R3276 VDD.n8961 VDD.n8418 92.5005
R3277 VDD.n8414 VDD.n8413 92.5005
R3278 VDD.n8970 VDD.n8414 92.5005
R3279 VDD.n8404 VDD.n8280 92.5005
R3280 VDD.n8336 VDD.n8335 92.5005
R3281 VDD.n8333 VDD.n8305 92.5005
R3282 VDD.n8311 VDD.n8306 92.5005
R3283 VDD.n8328 VDD.n8327 92.5005
R3284 VDD.n8325 VDD.n8324 92.5005
R3285 VDD.n8319 VDD.n8312 92.5005
R3286 VDD.n8317 VDD.n8316 92.5005
R3287 VDD.n8315 VDD.n8282 92.5005
R3288 VDD.n8338 VDD.n8290 92.5005
R3289 VDD.n8340 VDD.n8289 92.5005
R3290 VDD.n8365 VDD.n8364 92.5005
R3291 VDD.n8298 VDD.n8272 92.5005
R3292 VDD.n8384 VDD.n8383 92.5005
R3293 VDD.n8381 VDD.n8380 92.5005
R3294 VDD.n8377 VDD.n8299 92.5005
R3295 VDD.n8374 VDD.n8373 92.5005
R3296 VDD.n8372 VDD.n8371 92.5005
R3297 VDD.n8301 VDD.n8300 92.5005
R3298 VDD.n8376 VDD.n8375 92.5005
R3299 VDD.n8379 VDD.n8378 92.5005
R3300 VDD.n8297 VDD.n8296 92.5005
R3301 VDD.n8386 VDD.n8385 92.5005
R3302 VDD.n8997 VDD.n8271 92.5005
R3303 VDD.n9000 VDD.n8999 92.5005
R3304 VDD.n8370 VDD.n8292 92.5005
R3305 VDD.n8388 VDD.n8292 92.5005
R3306 VDD.n8369 VDD.n8368 92.5005
R3307 VDD.n8367 VDD.n8304 92.5005
R3308 VDD.n8583 VDD.n8582 92.5005
R3309 VDD.n8580 VDD.n8533 92.5005
R3310 VDD.n8579 VDD.n8578 92.5005
R3311 VDD.n8577 VDD.n8534 92.5005
R3312 VDD.n8575 VDD.n8574 92.5005
R3313 VDD.n8573 VDD.n8537 92.5005
R3314 VDD.n8540 VDD.n8537 92.5005
R3315 VDD.n8572 VDD.n8571 92.5005
R3316 VDD.n8571 VDD.n8570 92.5005
R3317 VDD.n8539 VDD.n8538 92.5005
R3318 VDD.n8569 VDD.n8539 92.5005
R3319 VDD.n8567 VDD.n8566 92.5005
R3320 VDD.n8568 VDD.n8567 92.5005
R3321 VDD.n8565 VDD.n8542 92.5005
R3322 VDD.n8542 VDD.n8541 92.5005
R3323 VDD.n8564 VDD.n8563 92.5005
R3324 VDD.n8563 VDD.n8562 92.5005
R3325 VDD.n8544 VDD.n8543 92.5005
R3326 VDD.n8561 VDD.n8544 92.5005
R3327 VDD.n8559 VDD.n8558 92.5005
R3328 VDD.n8560 VDD.n8559 92.5005
R3329 VDD.n8557 VDD.n8546 92.5005
R3330 VDD.n8546 VDD.n8545 92.5005
R3331 VDD.n8556 VDD.n8555 92.5005
R3332 VDD.n8555 VDD.n8554 92.5005
R3333 VDD.n8548 VDD.n8547 92.5005
R3334 VDD.n8553 VDD.n8548 92.5005
R3335 VDD.n8551 VDD.n8550 92.5005
R3336 VDD.n8552 VDD.n8551 92.5005
R3337 VDD.n8549 VDD.n8275 92.5005
R3338 VDD.n8277 VDD.n8275 92.5005
R3339 VDD.n8996 VDD.n8276 92.5005
R3340 VDD.n8996 VDD.n8995 92.5005
R3341 VDD.n8635 VDD.n8634 92.5005
R3342 VDD.n8634 VDD.n8633 92.5005
R3343 VDD.n8507 VDD.n8506 92.5005
R3344 VDD.n8632 VDD.n8507 92.5005
R3345 VDD.n8630 VDD.n8629 92.5005
R3346 VDD.n8631 VDD.n8630 92.5005
R3347 VDD.n8628 VDD.n8509 92.5005
R3348 VDD.n8509 VDD.n8508 92.5005
R3349 VDD.n8627 VDD.n8626 92.5005
R3350 VDD.n8626 VDD.n8625 92.5005
R3351 VDD.n8511 VDD.n8510 92.5005
R3352 VDD.n8624 VDD.n8511 92.5005
R3353 VDD.n8622 VDD.n8621 92.5005
R3354 VDD.n8623 VDD.n8622 92.5005
R3355 VDD.n8620 VDD.n8513 92.5005
R3356 VDD.n8513 VDD.n8512 92.5005
R3357 VDD.n8619 VDD.n8618 92.5005
R3358 VDD.n8618 VDD.n8617 92.5005
R3359 VDD.n8515 VDD.n8514 92.5005
R3360 VDD.n8616 VDD.n8515 92.5005
R3361 VDD.n8614 VDD.n8613 92.5005
R3362 VDD.n8615 VDD.n8614 92.5005
R3363 VDD.n8612 VDD.n8517 92.5005
R3364 VDD.n8517 VDD.n8516 92.5005
R3365 VDD.n8611 VDD.n8610 92.5005
R3366 VDD.n8610 VDD.n8609 92.5005
R3367 VDD.n8519 VDD.n8518 92.5005
R3368 VDD.n8608 VDD.n8519 92.5005
R3369 VDD.n8606 VDD.n8605 92.5005
R3370 VDD.n8607 VDD.n8606 92.5005
R3371 VDD.n8604 VDD.n8521 92.5005
R3372 VDD.n8521 VDD.n8520 92.5005
R3373 VDD.n8603 VDD.n8602 92.5005
R3374 VDD.n8602 VDD.n8601 92.5005
R3375 VDD.n8523 VDD.n8522 92.5005
R3376 VDD.n8600 VDD.n8523 92.5005
R3377 VDD.n8598 VDD.n8597 92.5005
R3378 VDD.n8599 VDD.n8598 92.5005
R3379 VDD.n8596 VDD.n8525 92.5005
R3380 VDD.n8525 VDD.n8524 92.5005
R3381 VDD.n8595 VDD.n8594 92.5005
R3382 VDD.n8594 VDD.n8593 92.5005
R3383 VDD.n8527 VDD.n8526 92.5005
R3384 VDD.n8592 VDD.n8527 92.5005
R3385 VDD.n8590 VDD.n8589 92.5005
R3386 VDD.n8591 VDD.n8590 92.5005
R3387 VDD.n8588 VDD.n8529 92.5005
R3388 VDD.n8529 VDD.n8528 92.5005
R3389 VDD.n8587 VDD.n8586 92.5005
R3390 VDD.n8586 VDD.n8585 92.5005
R3391 VDD.n8531 VDD.n8530 92.5005
R3392 VDD.n8584 VDD.n8531 92.5005
R3393 VDD.n8643 VDD.n8504 92.5005
R3394 VDD.n8647 VDD.n8646 92.5005
R3395 VDD.n8505 VDD.n8503 92.5005
R3396 VDD.n8677 VDD.n8487 92.5005
R3397 VDD.n8673 VDD.n8487 92.5005
R3398 VDD.n8676 VDD.n8675 92.5005
R3399 VDD.n8675 VDD.n8674 92.5005
R3400 VDD.n8489 VDD.n8488 92.5005
R3401 VDD.n8672 VDD.n8489 92.5005
R3402 VDD.n8670 VDD.n8669 92.5005
R3403 VDD.n8671 VDD.n8670 92.5005
R3404 VDD.n8668 VDD.n8491 92.5005
R3405 VDD.n8491 VDD.n8490 92.5005
R3406 VDD.n8667 VDD.n8666 92.5005
R3407 VDD.n8666 VDD.n8665 92.5005
R3408 VDD.n8493 VDD.n8492 92.5005
R3409 VDD.n8664 VDD.n8493 92.5005
R3410 VDD.n8662 VDD.n8661 92.5005
R3411 VDD.n8663 VDD.n8662 92.5005
R3412 VDD.n8660 VDD.n8495 92.5005
R3413 VDD.n8495 VDD.n8494 92.5005
R3414 VDD.n8659 VDD.n8658 92.5005
R3415 VDD.n8658 VDD.n8657 92.5005
R3416 VDD.n8497 VDD.n8496 92.5005
R3417 VDD.n8656 VDD.n8497 92.5005
R3418 VDD.n8654 VDD.n8653 92.5005
R3419 VDD.n8655 VDD.n8654 92.5005
R3420 VDD.n8652 VDD.n8499 92.5005
R3421 VDD.n8499 VDD.n8498 92.5005
R3422 VDD.n8651 VDD.n8650 92.5005
R3423 VDD.n8650 VDD.n8649 92.5005
R3424 VDD.n8501 VDD.n8500 92.5005
R3425 VDD.n8639 VDD.n8636 92.5005
R3426 VDD.n8642 VDD.n8641 92.5005
R3427 VDD.n8867 VDD.n8866 92.5005
R3428 VDD.n8784 VDD.n8467 92.5005
R3429 VDD.n8786 VDD.n8785 92.5005
R3430 VDD.n8783 VDD.n8782 92.5005
R3431 VDD.n8753 VDD.n8752 92.5005
R3432 VDD.n8777 VDD.n8776 92.5005
R3433 VDD.n8755 VDD.n8754 92.5005
R3434 VDD.n8771 VDD.n8770 92.5005
R3435 VDD.n8767 VDD.n8766 92.5005
R3436 VDD.n8765 VDD.n8764 92.5005
R3437 VDD.n8842 VDD.n8841 92.5005
R3438 VDD.n8846 VDD.n8845 92.5005
R3439 VDD.n8849 VDD.n8848 92.5005
R3440 VDD.n8691 VDD.n8690 92.5005
R3441 VDD.n8680 VDD.n8679 92.5005
R3442 VDD.n8858 VDD.n8857 92.5005
R3443 VDD.n8859 VDD.n8486 92.5005
R3444 VDD.n8862 VDD.n8861 92.5005
R3445 VDD.n8856 VDD.n8855 92.5005
R3446 VDD.n8689 VDD.n8682 92.5005
R3447 VDD.n8851 VDD.n8850 92.5005
R3448 VDD.n8847 VDD.n8688 92.5005
R3449 VDD.n8844 VDD.n8843 92.5005
R3450 VDD.n8692 VDD.n8479 92.5005
R3451 VDD.n8864 VDD.n8479 92.5005
R3452 VDD.n8840 VDD.n8839 92.5005
R3453 VDD.n8759 VDD.n8758 92.5005
R3454 VDD.n8761 VDD.n8760 92.5005
R3455 VDD.n8763 VDD.n8762 92.5005
R3456 VDD.n8769 VDD.n8768 92.5005
R3457 VDD.n8788 VDD.n8787 92.5005
R3458 VDD.n8781 VDD.n8780 92.5005
R3459 VDD.n8779 VDD.n8778 92.5005
R3460 VDD.n8775 VDD.n8774 92.5005
R3461 VDD.n8773 VDD.n8772 92.5005
R3462 VDD.n8396 VDD.n8395 92.5005
R3463 VDD.n8287 VDD.n8286 92.5005
R3464 VDD.n8399 VDD.n8398 92.5005
R3465 VDD.n8400 VDD.n8399 92.5005
R3466 VDD.n8332 VDD.n8331 92.5005
R3467 VDD.n8330 VDD.n8329 92.5005
R3468 VDD.n8320 VDD.n8309 92.5005
R3469 VDD.n8323 VDD.n8322 92.5005
R3470 VDD.n8318 VDD.n8285 92.5005
R3471 VDD.n8334 VDD.n8288 92.5005
R3472 VDD.n8346 VDD.n8345 92.5005
R3473 VDD.n8348 VDD.n8344 92.5005
R3474 VDD.n8351 VDD.n8350 92.5005
R3475 VDD.n8353 VDD.n8352 92.5005
R3476 VDD.n8355 VDD.n8342 92.5005
R3477 VDD.n8358 VDD.n8357 92.5005
R3478 VDD.n8402 VDD.n8401 92.5005
R3479 VDD.n8401 VDD.n8400 92.5005
R3480 VDD.n8284 VDD.n8283 92.5005
R3481 VDD.n8286 VDD.n8284 92.5005
R3482 VDD.n8394 VDD.n8393 92.5005
R3483 VDD.n8395 VDD.n8394 92.5005
R3484 VDD.n8392 VDD.n8391 92.5005
R3485 VDD.n8391 VDD.n8390 92.5005
R3486 VDD.n9013 VDD.n9012 92.5005
R3487 VDD.n9012 VDD.n9011 92.5005
R3488 VDD.n9014 VDD.n8254 92.5005
R3489 VDD.n8258 VDD.n8254 92.5005
R3490 VDD.n9016 VDD.n9015 92.5005
R3491 VDD.n9017 VDD.n9016 92.5005
R3492 VDD.n8255 VDD.n8253 92.5005
R3493 VDD.n8749 VDD.n8253 92.5005
R3494 VDD.n8813 VDD.n8751 92.5005
R3495 VDD.n8751 VDD.n8750 92.5005
R3496 VDD.n8815 VDD.n8814 92.5005
R3497 VDD.n8816 VDD.n8815 92.5005
R3498 VDD.n8795 VDD.n8794 92.5005
R3499 VDD.n8794 VDD.n8702 92.5005
R3500 VDD.n8793 VDD.n8792 92.5005
R3501 VDD.n8793 VDD.n8701 92.5005
R3502 VDD.n8791 VDD.n8696 92.5005
R3503 VDD.n8836 VDD.n8696 92.5005
R3504 VDD.n8790 VDD.n8789 92.5005
R3505 VDD.n8789 VDD.n8683 92.5005
R3506 VDD.n8811 VDD.n8810 92.5005
R3507 VDD.n8808 VDD.n8796 92.5005
R3508 VDD.n8806 VDD.n8805 92.5005
R3509 VDD.n8804 VDD.n8803 92.5005
R3510 VDD.n8801 VDD.n8798 92.5005
R3511 VDD.n8799 VDD.n8712 92.5005
R3512 VDD.n8756 VDD.n8697 92.5005
R3513 VDD.n8697 VDD.n8683 92.5005
R3514 VDD.n8835 VDD.n8834 92.5005
R3515 VDD.n8836 VDD.n8835 92.5005
R3516 VDD.n8832 VDD.n8698 92.5005
R3517 VDD.n8701 VDD.n8698 92.5005
R3518 VDD.n8714 VDD.n8699 92.5005
R3519 VDD.n8714 VDD.n8702 92.5005
R3520 VDD.n8818 VDD.n8817 92.5005
R3521 VDD.n8817 VDD.n8816 92.5005
R3522 VDD.n8719 VDD.n8718 92.5005
R3523 VDD.n8750 VDD.n8719 92.5005
R3524 VDD.n8717 VDD.n8249 92.5005
R3525 VDD.n8749 VDD.n8249 92.5005
R3526 VDD.n9019 VDD.n9018 92.5005
R3527 VDD.n9018 VDD.n9017 92.5005
R3528 VDD.n8262 VDD.n8250 92.5005
R3529 VDD.n8258 VDD.n8250 92.5005
R3530 VDD.n9010 VDD.n9009 92.5005
R3531 VDD.n9011 VDD.n9010 92.5005
R3532 VDD.n8361 VDD.n8291 92.5005
R3533 VDD.n8390 VDD.n8291 92.5005
R3534 VDD.n8833 VDD.n8693 92.5005
R3535 VDD.n8695 VDD.n8693 92.5005
R3536 VDD.n8831 VDD.n8830 92.5005
R3537 VDD.n8830 VDD.n8829 92.5005
R3538 VDD.n8711 VDD.n8700 92.5005
R3539 VDD.n8708 VDD.n8700 92.5005
R3540 VDD.n8822 VDD.n8821 92.5005
R3541 VDD.n8823 VDD.n8822 92.5005
R3542 VDD.n8819 VDD.n8710 92.5005
R3543 VDD.n8720 VDD.n8710 92.5005
R3544 VDD.n8733 VDD.n8247 92.5005
R3545 VDD.n8733 VDD.n8251 92.5005
R3546 VDD.n8732 VDD.n8248 92.5005
R3547 VDD.n8732 VDD.n8252 92.5005
R3548 VDD.n8265 VDD.n8263 92.5005
R3549 VDD.n8265 VDD.n8259 92.5005
R3550 VDD.n9008 VDD.n9007 92.5005
R3551 VDD.n9007 VDD.n8260 92.5005
R3552 VDD.n9006 VDD.n8264 92.5005
R3553 VDD.n9006 VDD.n9005 92.5005
R3554 VDD.n8360 VDD.n8266 92.5005
R3555 VDD.n8389 VDD.n8266 92.5005
R3556 VDD.n8838 VDD.n8694 92.5005
R3557 VDD.n8838 VDD.n8837 92.5005
R3558 VDD.n7826 VDD.n7823 92.5005
R3559 VDD.n7982 VDD.n7826 92.5005
R3560 VDD.n8147 VDD.n7414 92.5005
R3561 VDD.n7534 VDD.n7414 92.5005
R3562 VDD.n8149 VDD.n8148 92.5005
R3563 VDD.n8150 VDD.n8149 92.5005
R3564 VDD.n7415 VDD.n7413 92.5005
R3565 VDD.n7413 VDD.n7405 92.5005
R3566 VDD.n7872 VDD.n7871 92.5005
R3567 VDD.n7872 VDD.n7404 92.5005
R3568 VDD.n7873 VDD.n7870 92.5005
R3569 VDD.n7873 VDD.n7397 92.5005
R3570 VDD.n7875 VDD.n7874 92.5005
R3571 VDD.n7874 VDD.n7396 92.5005
R3572 VDD.n7888 VDD.n7868 92.5005
R3573 VDD.n7887 VDD.n7886 92.5005
R3574 VDD.n7885 VDD.n7884 92.5005
R3575 VDD.n7883 VDD.n7882 92.5005
R3576 VDD.n7881 VDD.n7880 92.5005
R3577 VDD.n7890 VDD.n7889 92.5005
R3578 VDD.n7852 VDD.n7851 92.5005
R3579 VDD.n7865 VDD.n7852 92.5005
R3580 VDD.n7970 VDD.n7969 92.5005
R3581 VDD.n7969 VDD.n7968 92.5005
R3582 VDD.n7971 VDD.n7849 92.5005
R3583 VDD.n7853 VDD.n7849 92.5005
R3584 VDD.n7973 VDD.n7972 92.5005
R3585 VDD.n7974 VDD.n7973 92.5005
R3586 VDD.n7850 VDD.n7848 92.5005
R3587 VDD.n7848 VDD.n7840 92.5005
R3588 VDD.n8013 VDD.n7610 92.5005
R3589 VDD.n7610 VDD.n7609 92.5005
R3590 VDD.n8036 VDD.n8035 92.5005
R3591 VDD.n8035 VDD.n8034 92.5005
R3592 VDD.n7600 VDD.n7599 92.5005
R3593 VDD.n8033 VDD.n7600 92.5005
R3594 VDD.n8031 VDD.n8030 92.5005
R3595 VDD.n8032 VDD.n8031 92.5005
R3596 VDD.n8029 VDD.n7602 92.5005
R3597 VDD.n7602 VDD.n7601 92.5005
R3598 VDD.n8028 VDD.n8027 92.5005
R3599 VDD.n8027 VDD.n8026 92.5005
R3600 VDD.n7604 VDD.n7603 92.5005
R3601 VDD.n8025 VDD.n7604 92.5005
R3602 VDD.n8023 VDD.n8022 92.5005
R3603 VDD.n8024 VDD.n8023 92.5005
R3604 VDD.n8021 VDD.n7606 92.5005
R3605 VDD.n7606 VDD.n7605 92.5005
R3606 VDD.n8020 VDD.n8019 92.5005
R3607 VDD.n8019 VDD.n8018 92.5005
R3608 VDD.n7608 VDD.n7607 92.5005
R3609 VDD.n8017 VDD.n7608 92.5005
R3610 VDD.n8015 VDD.n8014 92.5005
R3611 VDD.n8016 VDD.n8015 92.5005
R3612 VDD.n8037 VDD.n7597 92.5005
R3613 VDD.n7597 VDD.n7596 92.5005
R3614 VDD.n8040 VDD.n8039 92.5005
R3615 VDD.n8041 VDD.n8040 92.5005
R3616 VDD.n8038 VDD.n7598 92.5005
R3617 VDD.n7594 VDD.n7593 92.5005
R3618 VDD.n8045 VDD.n8044 92.5005
R3619 VDD.n8044 VDD.n8043 92.5005
R3620 VDD.n8048 VDD.n8047 92.5005
R3621 VDD.n8049 VDD.n8048 92.5005
R3622 VDD.n7590 VDD.n7589 92.5005
R3623 VDD.n8050 VDD.n7590 92.5005
R3624 VDD.n8053 VDD.n8052 92.5005
R3625 VDD.n8052 VDD.n8051 92.5005
R3626 VDD.n8054 VDD.n7588 92.5005
R3627 VDD.n7588 VDD.n7587 92.5005
R3628 VDD.n8056 VDD.n8055 92.5005
R3629 VDD.n8057 VDD.n8056 92.5005
R3630 VDD.n7586 VDD.n7585 92.5005
R3631 VDD.n8058 VDD.n7586 92.5005
R3632 VDD.n8061 VDD.n8060 92.5005
R3633 VDD.n8060 VDD.n8059 92.5005
R3634 VDD.n8062 VDD.n7584 92.5005
R3635 VDD.n7584 VDD.n7583 92.5005
R3636 VDD.n8064 VDD.n8063 92.5005
R3637 VDD.n8065 VDD.n8064 92.5005
R3638 VDD.n7582 VDD.n7581 92.5005
R3639 VDD.n8066 VDD.n7582 92.5005
R3640 VDD.n8069 VDD.n8068 92.5005
R3641 VDD.n8068 VDD.n8067 92.5005
R3642 VDD.n8070 VDD.n7580 92.5005
R3643 VDD.n7580 VDD.n7579 92.5005
R3644 VDD.n8072 VDD.n8071 92.5005
R3645 VDD.n8073 VDD.n8072 92.5005
R3646 VDD.n7578 VDD.n7577 92.5005
R3647 VDD.n8074 VDD.n7578 92.5005
R3648 VDD.n8077 VDD.n8076 92.5005
R3649 VDD.n8076 VDD.n8075 92.5005
R3650 VDD.n8078 VDD.n7576 92.5005
R3651 VDD.n7576 VDD.n7575 92.5005
R3652 VDD.n8080 VDD.n8079 92.5005
R3653 VDD.n8081 VDD.n8080 92.5005
R3654 VDD.n7574 VDD.n7573 92.5005
R3655 VDD.n8082 VDD.n7574 92.5005
R3656 VDD.n8085 VDD.n8084 92.5005
R3657 VDD.n8084 VDD.n8083 92.5005
R3658 VDD.n8086 VDD.n7572 92.5005
R3659 VDD.n7572 VDD.n7571 92.5005
R3660 VDD.n8088 VDD.n8087 92.5005
R3661 VDD.n8089 VDD.n8088 92.5005
R3662 VDD.n7570 VDD.n7569 92.5005
R3663 VDD.n8090 VDD.n7570 92.5005
R3664 VDD.n8093 VDD.n8092 92.5005
R3665 VDD.n8092 VDD.n8091 92.5005
R3666 VDD.n8094 VDD.n7568 92.5005
R3667 VDD.n7568 VDD.n7567 92.5005
R3668 VDD.n8096 VDD.n8095 92.5005
R3669 VDD.n8097 VDD.n8096 92.5005
R3670 VDD.n7566 VDD.n7565 92.5005
R3671 VDD.n8098 VDD.n7566 92.5005
R3672 VDD.n8103 VDD.n8102 92.5005
R3673 VDD.n8102 VDD.n8101 92.5005
R3674 VDD.n8104 VDD.n7564 92.5005
R3675 VDD.n8100 VDD.n7564 92.5005
R3676 VDD.n8046 VDD.n7592 92.5005
R3677 VDD.n7592 VDD.n7591 92.5005
R3678 VDD.n8118 VDD.n8117 92.5005
R3679 VDD.n8117 VDD.n8116 92.5005
R3680 VDD.n8119 VDD.n7557 92.5005
R3681 VDD.n7557 VDD.n7556 92.5005
R3682 VDD.n8121 VDD.n8120 92.5005
R3683 VDD.n8122 VDD.n8121 92.5005
R3684 VDD.n7555 VDD.n7554 92.5005
R3685 VDD.n8123 VDD.n7555 92.5005
R3686 VDD.n8126 VDD.n8125 92.5005
R3687 VDD.n8125 VDD.n8124 92.5005
R3688 VDD.n8127 VDD.n7553 92.5005
R3689 VDD.n7553 VDD.n7552 92.5005
R3690 VDD.n8129 VDD.n8128 92.5005
R3691 VDD.n8130 VDD.n8129 92.5005
R3692 VDD.n7551 VDD.n7550 92.5005
R3693 VDD.n8131 VDD.n7551 92.5005
R3694 VDD.n8134 VDD.n8133 92.5005
R3695 VDD.n8133 VDD.n8132 92.5005
R3696 VDD.n8135 VDD.n7426 92.5005
R3697 VDD.n7426 VDD.n7424 92.5005
R3698 VDD.n8137 VDD.n8136 92.5005
R3699 VDD.n8138 VDD.n8137 92.5005
R3700 VDD.n8113 VDD.n8112 92.5005
R3701 VDD.n8114 VDD.n8113 92.5005
R3702 VDD.n8111 VDD.n7561 92.5005
R3703 VDD.n7561 VDD.n7560 92.5005
R3704 VDD.n8110 VDD.n8109 92.5005
R3705 VDD.n8107 VDD.n7562 92.5005
R3706 VDD.n8106 VDD.n8105 92.5005
R3707 VDD.n8106 VDD.n7563 92.5005
R3708 VDD.n7559 VDD.n7558 92.5005
R3709 VDD.n8115 VDD.n7559 92.5005
R3710 VDD.n7549 VDD.n7425 92.5005
R3711 VDD.n7481 VDD.n7480 92.5005
R3712 VDD.n7478 VDD.n7450 92.5005
R3713 VDD.n7456 VDD.n7451 92.5005
R3714 VDD.n7473 VDD.n7472 92.5005
R3715 VDD.n7470 VDD.n7469 92.5005
R3716 VDD.n7464 VDD.n7457 92.5005
R3717 VDD.n7462 VDD.n7461 92.5005
R3718 VDD.n7460 VDD.n7427 92.5005
R3719 VDD.n7483 VDD.n7435 92.5005
R3720 VDD.n7485 VDD.n7434 92.5005
R3721 VDD.n7510 VDD.n7509 92.5005
R3722 VDD.n7443 VDD.n7417 92.5005
R3723 VDD.n7529 VDD.n7528 92.5005
R3724 VDD.n7526 VDD.n7525 92.5005
R3725 VDD.n7522 VDD.n7444 92.5005
R3726 VDD.n7519 VDD.n7518 92.5005
R3727 VDD.n7517 VDD.n7516 92.5005
R3728 VDD.n7446 VDD.n7445 92.5005
R3729 VDD.n7521 VDD.n7520 92.5005
R3730 VDD.n7524 VDD.n7523 92.5005
R3731 VDD.n7442 VDD.n7441 92.5005
R3732 VDD.n7531 VDD.n7530 92.5005
R3733 VDD.n8142 VDD.n7416 92.5005
R3734 VDD.n8145 VDD.n8144 92.5005
R3735 VDD.n7515 VDD.n7437 92.5005
R3736 VDD.n7533 VDD.n7437 92.5005
R3737 VDD.n7514 VDD.n7513 92.5005
R3738 VDD.n7512 VDD.n7449 92.5005
R3739 VDD.n7728 VDD.n7727 92.5005
R3740 VDD.n7725 VDD.n7678 92.5005
R3741 VDD.n7724 VDD.n7723 92.5005
R3742 VDD.n7722 VDD.n7679 92.5005
R3743 VDD.n7720 VDD.n7719 92.5005
R3744 VDD.n7718 VDD.n7682 92.5005
R3745 VDD.n7685 VDD.n7682 92.5005
R3746 VDD.n7717 VDD.n7716 92.5005
R3747 VDD.n7716 VDD.n7715 92.5005
R3748 VDD.n7684 VDD.n7683 92.5005
R3749 VDD.n7714 VDD.n7684 92.5005
R3750 VDD.n7712 VDD.n7711 92.5005
R3751 VDD.n7713 VDD.n7712 92.5005
R3752 VDD.n7710 VDD.n7687 92.5005
R3753 VDD.n7687 VDD.n7686 92.5005
R3754 VDD.n7709 VDD.n7708 92.5005
R3755 VDD.n7708 VDD.n7707 92.5005
R3756 VDD.n7689 VDD.n7688 92.5005
R3757 VDD.n7706 VDD.n7689 92.5005
R3758 VDD.n7704 VDD.n7703 92.5005
R3759 VDD.n7705 VDD.n7704 92.5005
R3760 VDD.n7702 VDD.n7691 92.5005
R3761 VDD.n7691 VDD.n7690 92.5005
R3762 VDD.n7701 VDD.n7700 92.5005
R3763 VDD.n7700 VDD.n7699 92.5005
R3764 VDD.n7693 VDD.n7692 92.5005
R3765 VDD.n7698 VDD.n7693 92.5005
R3766 VDD.n7696 VDD.n7695 92.5005
R3767 VDD.n7697 VDD.n7696 92.5005
R3768 VDD.n7694 VDD.n7420 92.5005
R3769 VDD.n7422 VDD.n7420 92.5005
R3770 VDD.n8141 VDD.n7421 92.5005
R3771 VDD.n8141 VDD.n8140 92.5005
R3772 VDD.n7780 VDD.n7779 92.5005
R3773 VDD.n7779 VDD.n7778 92.5005
R3774 VDD.n7652 VDD.n7651 92.5005
R3775 VDD.n7777 VDD.n7652 92.5005
R3776 VDD.n7775 VDD.n7774 92.5005
R3777 VDD.n7776 VDD.n7775 92.5005
R3778 VDD.n7773 VDD.n7654 92.5005
R3779 VDD.n7654 VDD.n7653 92.5005
R3780 VDD.n7772 VDD.n7771 92.5005
R3781 VDD.n7771 VDD.n7770 92.5005
R3782 VDD.n7656 VDD.n7655 92.5005
R3783 VDD.n7769 VDD.n7656 92.5005
R3784 VDD.n7767 VDD.n7766 92.5005
R3785 VDD.n7768 VDD.n7767 92.5005
R3786 VDD.n7765 VDD.n7658 92.5005
R3787 VDD.n7658 VDD.n7657 92.5005
R3788 VDD.n7764 VDD.n7763 92.5005
R3789 VDD.n7763 VDD.n7762 92.5005
R3790 VDD.n7660 VDD.n7659 92.5005
R3791 VDD.n7761 VDD.n7660 92.5005
R3792 VDD.n7759 VDD.n7758 92.5005
R3793 VDD.n7760 VDD.n7759 92.5005
R3794 VDD.n7757 VDD.n7662 92.5005
R3795 VDD.n7662 VDD.n7661 92.5005
R3796 VDD.n7756 VDD.n7755 92.5005
R3797 VDD.n7755 VDD.n7754 92.5005
R3798 VDD.n7664 VDD.n7663 92.5005
R3799 VDD.n7753 VDD.n7664 92.5005
R3800 VDD.n7751 VDD.n7750 92.5005
R3801 VDD.n7752 VDD.n7751 92.5005
R3802 VDD.n7749 VDD.n7666 92.5005
R3803 VDD.n7666 VDD.n7665 92.5005
R3804 VDD.n7748 VDD.n7747 92.5005
R3805 VDD.n7747 VDD.n7746 92.5005
R3806 VDD.n7668 VDD.n7667 92.5005
R3807 VDD.n7745 VDD.n7668 92.5005
R3808 VDD.n7743 VDD.n7742 92.5005
R3809 VDD.n7744 VDD.n7743 92.5005
R3810 VDD.n7741 VDD.n7670 92.5005
R3811 VDD.n7670 VDD.n7669 92.5005
R3812 VDD.n7740 VDD.n7739 92.5005
R3813 VDD.n7739 VDD.n7738 92.5005
R3814 VDD.n7672 VDD.n7671 92.5005
R3815 VDD.n7737 VDD.n7672 92.5005
R3816 VDD.n7735 VDD.n7734 92.5005
R3817 VDD.n7736 VDD.n7735 92.5005
R3818 VDD.n7733 VDD.n7674 92.5005
R3819 VDD.n7674 VDD.n7673 92.5005
R3820 VDD.n7732 VDD.n7731 92.5005
R3821 VDD.n7731 VDD.n7730 92.5005
R3822 VDD.n7676 VDD.n7675 92.5005
R3823 VDD.n7729 VDD.n7676 92.5005
R3824 VDD.n7788 VDD.n7649 92.5005
R3825 VDD.n7792 VDD.n7791 92.5005
R3826 VDD.n7650 VDD.n7648 92.5005
R3827 VDD.n7822 VDD.n7632 92.5005
R3828 VDD.n7818 VDD.n7632 92.5005
R3829 VDD.n7821 VDD.n7820 92.5005
R3830 VDD.n7820 VDD.n7819 92.5005
R3831 VDD.n7634 VDD.n7633 92.5005
R3832 VDD.n7817 VDD.n7634 92.5005
R3833 VDD.n7815 VDD.n7814 92.5005
R3834 VDD.n7816 VDD.n7815 92.5005
R3835 VDD.n7813 VDD.n7636 92.5005
R3836 VDD.n7636 VDD.n7635 92.5005
R3837 VDD.n7812 VDD.n7811 92.5005
R3838 VDD.n7811 VDD.n7810 92.5005
R3839 VDD.n7638 VDD.n7637 92.5005
R3840 VDD.n7809 VDD.n7638 92.5005
R3841 VDD.n7807 VDD.n7806 92.5005
R3842 VDD.n7808 VDD.n7807 92.5005
R3843 VDD.n7805 VDD.n7640 92.5005
R3844 VDD.n7640 VDD.n7639 92.5005
R3845 VDD.n7804 VDD.n7803 92.5005
R3846 VDD.n7803 VDD.n7802 92.5005
R3847 VDD.n7642 VDD.n7641 92.5005
R3848 VDD.n7801 VDD.n7642 92.5005
R3849 VDD.n7799 VDD.n7798 92.5005
R3850 VDD.n7800 VDD.n7799 92.5005
R3851 VDD.n7797 VDD.n7644 92.5005
R3852 VDD.n7644 VDD.n7643 92.5005
R3853 VDD.n7796 VDD.n7795 92.5005
R3854 VDD.n7795 VDD.n7794 92.5005
R3855 VDD.n7646 VDD.n7645 92.5005
R3856 VDD.n7784 VDD.n7781 92.5005
R3857 VDD.n7787 VDD.n7786 92.5005
R3858 VDD.n8012 VDD.n8011 92.5005
R3859 VDD.n7929 VDD.n7612 92.5005
R3860 VDD.n7931 VDD.n7930 92.5005
R3861 VDD.n7928 VDD.n7927 92.5005
R3862 VDD.n7898 VDD.n7897 92.5005
R3863 VDD.n7922 VDD.n7921 92.5005
R3864 VDD.n7900 VDD.n7899 92.5005
R3865 VDD.n7916 VDD.n7915 92.5005
R3866 VDD.n7912 VDD.n7911 92.5005
R3867 VDD.n7910 VDD.n7909 92.5005
R3868 VDD.n7987 VDD.n7986 92.5005
R3869 VDD.n7991 VDD.n7990 92.5005
R3870 VDD.n7994 VDD.n7993 92.5005
R3871 VDD.n7836 VDD.n7835 92.5005
R3872 VDD.n7825 VDD.n7824 92.5005
R3873 VDD.n8003 VDD.n8002 92.5005
R3874 VDD.n8004 VDD.n7631 92.5005
R3875 VDD.n8007 VDD.n8006 92.5005
R3876 VDD.n8001 VDD.n8000 92.5005
R3877 VDD.n7834 VDD.n7827 92.5005
R3878 VDD.n7996 VDD.n7995 92.5005
R3879 VDD.n7992 VDD.n7833 92.5005
R3880 VDD.n7989 VDD.n7988 92.5005
R3881 VDD.n7837 VDD.n7624 92.5005
R3882 VDD.n8009 VDD.n7624 92.5005
R3883 VDD.n7985 VDD.n7984 92.5005
R3884 VDD.n7904 VDD.n7903 92.5005
R3885 VDD.n7906 VDD.n7905 92.5005
R3886 VDD.n7908 VDD.n7907 92.5005
R3887 VDD.n7914 VDD.n7913 92.5005
R3888 VDD.n7933 VDD.n7932 92.5005
R3889 VDD.n7926 VDD.n7925 92.5005
R3890 VDD.n7924 VDD.n7923 92.5005
R3891 VDD.n7920 VDD.n7919 92.5005
R3892 VDD.n7918 VDD.n7917 92.5005
R3893 VDD.n7541 VDD.n7540 92.5005
R3894 VDD.n7432 VDD.n7431 92.5005
R3895 VDD.n7544 VDD.n7543 92.5005
R3896 VDD.n7545 VDD.n7544 92.5005
R3897 VDD.n7477 VDD.n7476 92.5005
R3898 VDD.n7475 VDD.n7474 92.5005
R3899 VDD.n7465 VDD.n7454 92.5005
R3900 VDD.n7468 VDD.n7467 92.5005
R3901 VDD.n7463 VDD.n7430 92.5005
R3902 VDD.n7479 VDD.n7433 92.5005
R3903 VDD.n7491 VDD.n7490 92.5005
R3904 VDD.n7493 VDD.n7489 92.5005
R3905 VDD.n7496 VDD.n7495 92.5005
R3906 VDD.n7498 VDD.n7497 92.5005
R3907 VDD.n7500 VDD.n7487 92.5005
R3908 VDD.n7503 VDD.n7502 92.5005
R3909 VDD.n7547 VDD.n7546 92.5005
R3910 VDD.n7546 VDD.n7545 92.5005
R3911 VDD.n7429 VDD.n7428 92.5005
R3912 VDD.n7431 VDD.n7429 92.5005
R3913 VDD.n7539 VDD.n7538 92.5005
R3914 VDD.n7540 VDD.n7539 92.5005
R3915 VDD.n7537 VDD.n7536 92.5005
R3916 VDD.n7536 VDD.n7535 92.5005
R3917 VDD.n8158 VDD.n8157 92.5005
R3918 VDD.n8157 VDD.n8156 92.5005
R3919 VDD.n8159 VDD.n7399 92.5005
R3920 VDD.n7403 VDD.n7399 92.5005
R3921 VDD.n8161 VDD.n8160 92.5005
R3922 VDD.n8162 VDD.n8161 92.5005
R3923 VDD.n7400 VDD.n7398 92.5005
R3924 VDD.n7894 VDD.n7398 92.5005
R3925 VDD.n7958 VDD.n7896 92.5005
R3926 VDD.n7896 VDD.n7895 92.5005
R3927 VDD.n7960 VDD.n7959 92.5005
R3928 VDD.n7961 VDD.n7960 92.5005
R3929 VDD.n7940 VDD.n7939 92.5005
R3930 VDD.n7939 VDD.n7847 92.5005
R3931 VDD.n7938 VDD.n7937 92.5005
R3932 VDD.n7938 VDD.n7846 92.5005
R3933 VDD.n7936 VDD.n7841 92.5005
R3934 VDD.n7981 VDD.n7841 92.5005
R3935 VDD.n7935 VDD.n7934 92.5005
R3936 VDD.n7934 VDD.n7828 92.5005
R3937 VDD.n7956 VDD.n7955 92.5005
R3938 VDD.n7953 VDD.n7941 92.5005
R3939 VDD.n7951 VDD.n7950 92.5005
R3940 VDD.n7949 VDD.n7948 92.5005
R3941 VDD.n7946 VDD.n7943 92.5005
R3942 VDD.n7944 VDD.n7857 92.5005
R3943 VDD.n7901 VDD.n7842 92.5005
R3944 VDD.n7842 VDD.n7828 92.5005
R3945 VDD.n7980 VDD.n7979 92.5005
R3946 VDD.n7981 VDD.n7980 92.5005
R3947 VDD.n7977 VDD.n7843 92.5005
R3948 VDD.n7846 VDD.n7843 92.5005
R3949 VDD.n7859 VDD.n7844 92.5005
R3950 VDD.n7859 VDD.n7847 92.5005
R3951 VDD.n7963 VDD.n7962 92.5005
R3952 VDD.n7962 VDD.n7961 92.5005
R3953 VDD.n7864 VDD.n7863 92.5005
R3954 VDD.n7895 VDD.n7864 92.5005
R3955 VDD.n7862 VDD.n7394 92.5005
R3956 VDD.n7894 VDD.n7394 92.5005
R3957 VDD.n8164 VDD.n8163 92.5005
R3958 VDD.n8163 VDD.n8162 92.5005
R3959 VDD.n7407 VDD.n7395 92.5005
R3960 VDD.n7403 VDD.n7395 92.5005
R3961 VDD.n8155 VDD.n8154 92.5005
R3962 VDD.n8156 VDD.n8155 92.5005
R3963 VDD.n7506 VDD.n7436 92.5005
R3964 VDD.n7535 VDD.n7436 92.5005
R3965 VDD.n7978 VDD.n7838 92.5005
R3966 VDD.n7840 VDD.n7838 92.5005
R3967 VDD.n7976 VDD.n7975 92.5005
R3968 VDD.n7975 VDD.n7974 92.5005
R3969 VDD.n7856 VDD.n7845 92.5005
R3970 VDD.n7853 VDD.n7845 92.5005
R3971 VDD.n7967 VDD.n7966 92.5005
R3972 VDD.n7968 VDD.n7967 92.5005
R3973 VDD.n7964 VDD.n7855 92.5005
R3974 VDD.n7865 VDD.n7855 92.5005
R3975 VDD.n7878 VDD.n7392 92.5005
R3976 VDD.n7878 VDD.n7396 92.5005
R3977 VDD.n7877 VDD.n7393 92.5005
R3978 VDD.n7877 VDD.n7397 92.5005
R3979 VDD.n7410 VDD.n7408 92.5005
R3980 VDD.n7410 VDD.n7404 92.5005
R3981 VDD.n8153 VDD.n8152 92.5005
R3982 VDD.n8152 VDD.n7405 92.5005
R3983 VDD.n8151 VDD.n7409 92.5005
R3984 VDD.n8151 VDD.n8150 92.5005
R3985 VDD.n7505 VDD.n7411 92.5005
R3986 VDD.n7534 VDD.n7411 92.5005
R3987 VDD.n7983 VDD.n7839 92.5005
R3988 VDD.n7983 VDD.n7982 92.5005
R3989 VDD.n6972 VDD.n6969 92.5005
R3990 VDD.n7128 VDD.n6972 92.5005
R3991 VDD.n7293 VDD.n6560 92.5005
R3992 VDD.n6680 VDD.n6560 92.5005
R3993 VDD.n7295 VDD.n7294 92.5005
R3994 VDD.n7296 VDD.n7295 92.5005
R3995 VDD.n6561 VDD.n6559 92.5005
R3996 VDD.n6559 VDD.n6551 92.5005
R3997 VDD.n7018 VDD.n7017 92.5005
R3998 VDD.n7018 VDD.n6550 92.5005
R3999 VDD.n7019 VDD.n7016 92.5005
R4000 VDD.n7019 VDD.n6543 92.5005
R4001 VDD.n7021 VDD.n7020 92.5005
R4002 VDD.n7020 VDD.n6542 92.5005
R4003 VDD.n7034 VDD.n7014 92.5005
R4004 VDD.n7033 VDD.n7032 92.5005
R4005 VDD.n7031 VDD.n7030 92.5005
R4006 VDD.n7029 VDD.n7028 92.5005
R4007 VDD.n7027 VDD.n7026 92.5005
R4008 VDD.n7036 VDD.n7035 92.5005
R4009 VDD.n6998 VDD.n6997 92.5005
R4010 VDD.n7011 VDD.n6998 92.5005
R4011 VDD.n7116 VDD.n7115 92.5005
R4012 VDD.n7115 VDD.n7114 92.5005
R4013 VDD.n7117 VDD.n6995 92.5005
R4014 VDD.n6999 VDD.n6995 92.5005
R4015 VDD.n7119 VDD.n7118 92.5005
R4016 VDD.n7120 VDD.n7119 92.5005
R4017 VDD.n6996 VDD.n6994 92.5005
R4018 VDD.n6994 VDD.n6986 92.5005
R4019 VDD.n7159 VDD.n6756 92.5005
R4020 VDD.n6756 VDD.n6755 92.5005
R4021 VDD.n7182 VDD.n7181 92.5005
R4022 VDD.n7181 VDD.n7180 92.5005
R4023 VDD.n6746 VDD.n6745 92.5005
R4024 VDD.n7179 VDD.n6746 92.5005
R4025 VDD.n7177 VDD.n7176 92.5005
R4026 VDD.n7178 VDD.n7177 92.5005
R4027 VDD.n7175 VDD.n6748 92.5005
R4028 VDD.n6748 VDD.n6747 92.5005
R4029 VDD.n7174 VDD.n7173 92.5005
R4030 VDD.n7173 VDD.n7172 92.5005
R4031 VDD.n6750 VDD.n6749 92.5005
R4032 VDD.n7171 VDD.n6750 92.5005
R4033 VDD.n7169 VDD.n7168 92.5005
R4034 VDD.n7170 VDD.n7169 92.5005
R4035 VDD.n7167 VDD.n6752 92.5005
R4036 VDD.n6752 VDD.n6751 92.5005
R4037 VDD.n7166 VDD.n7165 92.5005
R4038 VDD.n7165 VDD.n7164 92.5005
R4039 VDD.n6754 VDD.n6753 92.5005
R4040 VDD.n7163 VDD.n6754 92.5005
R4041 VDD.n7161 VDD.n7160 92.5005
R4042 VDD.n7162 VDD.n7161 92.5005
R4043 VDD.n7183 VDD.n6743 92.5005
R4044 VDD.n6743 VDD.n6742 92.5005
R4045 VDD.n7186 VDD.n7185 92.5005
R4046 VDD.n7187 VDD.n7186 92.5005
R4047 VDD.n7184 VDD.n6744 92.5005
R4048 VDD.n6740 VDD.n6739 92.5005
R4049 VDD.n7191 VDD.n7190 92.5005
R4050 VDD.n7190 VDD.n7189 92.5005
R4051 VDD.n7194 VDD.n7193 92.5005
R4052 VDD.n7195 VDD.n7194 92.5005
R4053 VDD.n6736 VDD.n6735 92.5005
R4054 VDD.n7196 VDD.n6736 92.5005
R4055 VDD.n7199 VDD.n7198 92.5005
R4056 VDD.n7198 VDD.n7197 92.5005
R4057 VDD.n7200 VDD.n6734 92.5005
R4058 VDD.n6734 VDD.n6733 92.5005
R4059 VDD.n7202 VDD.n7201 92.5005
R4060 VDD.n7203 VDD.n7202 92.5005
R4061 VDD.n6732 VDD.n6731 92.5005
R4062 VDD.n7204 VDD.n6732 92.5005
R4063 VDD.n7207 VDD.n7206 92.5005
R4064 VDD.n7206 VDD.n7205 92.5005
R4065 VDD.n7208 VDD.n6730 92.5005
R4066 VDD.n6730 VDD.n6729 92.5005
R4067 VDD.n7210 VDD.n7209 92.5005
R4068 VDD.n7211 VDD.n7210 92.5005
R4069 VDD.n6728 VDD.n6727 92.5005
R4070 VDD.n7212 VDD.n6728 92.5005
R4071 VDD.n7215 VDD.n7214 92.5005
R4072 VDD.n7214 VDD.n7213 92.5005
R4073 VDD.n7216 VDD.n6726 92.5005
R4074 VDD.n6726 VDD.n6725 92.5005
R4075 VDD.n7218 VDD.n7217 92.5005
R4076 VDD.n7219 VDD.n7218 92.5005
R4077 VDD.n6724 VDD.n6723 92.5005
R4078 VDD.n7220 VDD.n6724 92.5005
R4079 VDD.n7223 VDD.n7222 92.5005
R4080 VDD.n7222 VDD.n7221 92.5005
R4081 VDD.n7224 VDD.n6722 92.5005
R4082 VDD.n6722 VDD.n6721 92.5005
R4083 VDD.n7226 VDD.n7225 92.5005
R4084 VDD.n7227 VDD.n7226 92.5005
R4085 VDD.n6720 VDD.n6719 92.5005
R4086 VDD.n7228 VDD.n6720 92.5005
R4087 VDD.n7231 VDD.n7230 92.5005
R4088 VDD.n7230 VDD.n7229 92.5005
R4089 VDD.n7232 VDD.n6718 92.5005
R4090 VDD.n6718 VDD.n6717 92.5005
R4091 VDD.n7234 VDD.n7233 92.5005
R4092 VDD.n7235 VDD.n7234 92.5005
R4093 VDD.n6716 VDD.n6715 92.5005
R4094 VDD.n7236 VDD.n6716 92.5005
R4095 VDD.n7239 VDD.n7238 92.5005
R4096 VDD.n7238 VDD.n7237 92.5005
R4097 VDD.n7240 VDD.n6714 92.5005
R4098 VDD.n6714 VDD.n6713 92.5005
R4099 VDD.n7242 VDD.n7241 92.5005
R4100 VDD.n7243 VDD.n7242 92.5005
R4101 VDD.n6712 VDD.n6711 92.5005
R4102 VDD.n7244 VDD.n6712 92.5005
R4103 VDD.n7249 VDD.n7248 92.5005
R4104 VDD.n7248 VDD.n7247 92.5005
R4105 VDD.n7250 VDD.n6710 92.5005
R4106 VDD.n7246 VDD.n6710 92.5005
R4107 VDD.n7192 VDD.n6738 92.5005
R4108 VDD.n6738 VDD.n6737 92.5005
R4109 VDD.n7264 VDD.n7263 92.5005
R4110 VDD.n7263 VDD.n7262 92.5005
R4111 VDD.n7265 VDD.n6703 92.5005
R4112 VDD.n6703 VDD.n6702 92.5005
R4113 VDD.n7267 VDD.n7266 92.5005
R4114 VDD.n7268 VDD.n7267 92.5005
R4115 VDD.n6701 VDD.n6700 92.5005
R4116 VDD.n7269 VDD.n6701 92.5005
R4117 VDD.n7272 VDD.n7271 92.5005
R4118 VDD.n7271 VDD.n7270 92.5005
R4119 VDD.n7273 VDD.n6699 92.5005
R4120 VDD.n6699 VDD.n6698 92.5005
R4121 VDD.n7275 VDD.n7274 92.5005
R4122 VDD.n7276 VDD.n7275 92.5005
R4123 VDD.n6697 VDD.n6696 92.5005
R4124 VDD.n7277 VDD.n6697 92.5005
R4125 VDD.n7280 VDD.n7279 92.5005
R4126 VDD.n7279 VDD.n7278 92.5005
R4127 VDD.n7281 VDD.n6572 92.5005
R4128 VDD.n6572 VDD.n6570 92.5005
R4129 VDD.n7283 VDD.n7282 92.5005
R4130 VDD.n7284 VDD.n7283 92.5005
R4131 VDD.n7259 VDD.n7258 92.5005
R4132 VDD.n7260 VDD.n7259 92.5005
R4133 VDD.n7257 VDD.n6707 92.5005
R4134 VDD.n6707 VDD.n6706 92.5005
R4135 VDD.n7256 VDD.n7255 92.5005
R4136 VDD.n7253 VDD.n6708 92.5005
R4137 VDD.n7252 VDD.n7251 92.5005
R4138 VDD.n7252 VDD.n6709 92.5005
R4139 VDD.n6705 VDD.n6704 92.5005
R4140 VDD.n7261 VDD.n6705 92.5005
R4141 VDD.n6695 VDD.n6571 92.5005
R4142 VDD.n6627 VDD.n6626 92.5005
R4143 VDD.n6624 VDD.n6596 92.5005
R4144 VDD.n6602 VDD.n6597 92.5005
R4145 VDD.n6619 VDD.n6618 92.5005
R4146 VDD.n6616 VDD.n6615 92.5005
R4147 VDD.n6610 VDD.n6603 92.5005
R4148 VDD.n6608 VDD.n6607 92.5005
R4149 VDD.n6606 VDD.n6573 92.5005
R4150 VDD.n6629 VDD.n6581 92.5005
R4151 VDD.n6631 VDD.n6580 92.5005
R4152 VDD.n6656 VDD.n6655 92.5005
R4153 VDD.n6589 VDD.n6563 92.5005
R4154 VDD.n6675 VDD.n6674 92.5005
R4155 VDD.n6672 VDD.n6671 92.5005
R4156 VDD.n6668 VDD.n6590 92.5005
R4157 VDD.n6665 VDD.n6664 92.5005
R4158 VDD.n6663 VDD.n6662 92.5005
R4159 VDD.n6592 VDD.n6591 92.5005
R4160 VDD.n6667 VDD.n6666 92.5005
R4161 VDD.n6670 VDD.n6669 92.5005
R4162 VDD.n6588 VDD.n6587 92.5005
R4163 VDD.n6677 VDD.n6676 92.5005
R4164 VDD.n7288 VDD.n6562 92.5005
R4165 VDD.n7291 VDD.n7290 92.5005
R4166 VDD.n6661 VDD.n6583 92.5005
R4167 VDD.n6679 VDD.n6583 92.5005
R4168 VDD.n6660 VDD.n6659 92.5005
R4169 VDD.n6658 VDD.n6595 92.5005
R4170 VDD.n6874 VDD.n6873 92.5005
R4171 VDD.n6871 VDD.n6824 92.5005
R4172 VDD.n6870 VDD.n6869 92.5005
R4173 VDD.n6868 VDD.n6825 92.5005
R4174 VDD.n6866 VDD.n6865 92.5005
R4175 VDD.n6864 VDD.n6828 92.5005
R4176 VDD.n6831 VDD.n6828 92.5005
R4177 VDD.n6863 VDD.n6862 92.5005
R4178 VDD.n6862 VDD.n6861 92.5005
R4179 VDD.n6830 VDD.n6829 92.5005
R4180 VDD.n6860 VDD.n6830 92.5005
R4181 VDD.n6858 VDD.n6857 92.5005
R4182 VDD.n6859 VDD.n6858 92.5005
R4183 VDD.n6856 VDD.n6833 92.5005
R4184 VDD.n6833 VDD.n6832 92.5005
R4185 VDD.n6855 VDD.n6854 92.5005
R4186 VDD.n6854 VDD.n6853 92.5005
R4187 VDD.n6835 VDD.n6834 92.5005
R4188 VDD.n6852 VDD.n6835 92.5005
R4189 VDD.n6850 VDD.n6849 92.5005
R4190 VDD.n6851 VDD.n6850 92.5005
R4191 VDD.n6848 VDD.n6837 92.5005
R4192 VDD.n6837 VDD.n6836 92.5005
R4193 VDD.n6847 VDD.n6846 92.5005
R4194 VDD.n6846 VDD.n6845 92.5005
R4195 VDD.n6839 VDD.n6838 92.5005
R4196 VDD.n6844 VDD.n6839 92.5005
R4197 VDD.n6842 VDD.n6841 92.5005
R4198 VDD.n6843 VDD.n6842 92.5005
R4199 VDD.n6840 VDD.n6566 92.5005
R4200 VDD.n6568 VDD.n6566 92.5005
R4201 VDD.n7287 VDD.n6567 92.5005
R4202 VDD.n7287 VDD.n7286 92.5005
R4203 VDD.n6926 VDD.n6925 92.5005
R4204 VDD.n6925 VDD.n6924 92.5005
R4205 VDD.n6798 VDD.n6797 92.5005
R4206 VDD.n6923 VDD.n6798 92.5005
R4207 VDD.n6921 VDD.n6920 92.5005
R4208 VDD.n6922 VDD.n6921 92.5005
R4209 VDD.n6919 VDD.n6800 92.5005
R4210 VDD.n6800 VDD.n6799 92.5005
R4211 VDD.n6918 VDD.n6917 92.5005
R4212 VDD.n6917 VDD.n6916 92.5005
R4213 VDD.n6802 VDD.n6801 92.5005
R4214 VDD.n6915 VDD.n6802 92.5005
R4215 VDD.n6913 VDD.n6912 92.5005
R4216 VDD.n6914 VDD.n6913 92.5005
R4217 VDD.n6911 VDD.n6804 92.5005
R4218 VDD.n6804 VDD.n6803 92.5005
R4219 VDD.n6910 VDD.n6909 92.5005
R4220 VDD.n6909 VDD.n6908 92.5005
R4221 VDD.n6806 VDD.n6805 92.5005
R4222 VDD.n6907 VDD.n6806 92.5005
R4223 VDD.n6905 VDD.n6904 92.5005
R4224 VDD.n6906 VDD.n6905 92.5005
R4225 VDD.n6903 VDD.n6808 92.5005
R4226 VDD.n6808 VDD.n6807 92.5005
R4227 VDD.n6902 VDD.n6901 92.5005
R4228 VDD.n6901 VDD.n6900 92.5005
R4229 VDD.n6810 VDD.n6809 92.5005
R4230 VDD.n6899 VDD.n6810 92.5005
R4231 VDD.n6897 VDD.n6896 92.5005
R4232 VDD.n6898 VDD.n6897 92.5005
R4233 VDD.n6895 VDD.n6812 92.5005
R4234 VDD.n6812 VDD.n6811 92.5005
R4235 VDD.n6894 VDD.n6893 92.5005
R4236 VDD.n6893 VDD.n6892 92.5005
R4237 VDD.n6814 VDD.n6813 92.5005
R4238 VDD.n6891 VDD.n6814 92.5005
R4239 VDD.n6889 VDD.n6888 92.5005
R4240 VDD.n6890 VDD.n6889 92.5005
R4241 VDD.n6887 VDD.n6816 92.5005
R4242 VDD.n6816 VDD.n6815 92.5005
R4243 VDD.n6886 VDD.n6885 92.5005
R4244 VDD.n6885 VDD.n6884 92.5005
R4245 VDD.n6818 VDD.n6817 92.5005
R4246 VDD.n6883 VDD.n6818 92.5005
R4247 VDD.n6881 VDD.n6880 92.5005
R4248 VDD.n6882 VDD.n6881 92.5005
R4249 VDD.n6879 VDD.n6820 92.5005
R4250 VDD.n6820 VDD.n6819 92.5005
R4251 VDD.n6878 VDD.n6877 92.5005
R4252 VDD.n6877 VDD.n6876 92.5005
R4253 VDD.n6822 VDD.n6821 92.5005
R4254 VDD.n6875 VDD.n6822 92.5005
R4255 VDD.n6934 VDD.n6795 92.5005
R4256 VDD.n6938 VDD.n6937 92.5005
R4257 VDD.n6796 VDD.n6794 92.5005
R4258 VDD.n6968 VDD.n6778 92.5005
R4259 VDD.n6964 VDD.n6778 92.5005
R4260 VDD.n6967 VDD.n6966 92.5005
R4261 VDD.n6966 VDD.n6965 92.5005
R4262 VDD.n6780 VDD.n6779 92.5005
R4263 VDD.n6963 VDD.n6780 92.5005
R4264 VDD.n6961 VDD.n6960 92.5005
R4265 VDD.n6962 VDD.n6961 92.5005
R4266 VDD.n6959 VDD.n6782 92.5005
R4267 VDD.n6782 VDD.n6781 92.5005
R4268 VDD.n6958 VDD.n6957 92.5005
R4269 VDD.n6957 VDD.n6956 92.5005
R4270 VDD.n6784 VDD.n6783 92.5005
R4271 VDD.n6955 VDD.n6784 92.5005
R4272 VDD.n6953 VDD.n6952 92.5005
R4273 VDD.n6954 VDD.n6953 92.5005
R4274 VDD.n6951 VDD.n6786 92.5005
R4275 VDD.n6786 VDD.n6785 92.5005
R4276 VDD.n6950 VDD.n6949 92.5005
R4277 VDD.n6949 VDD.n6948 92.5005
R4278 VDD.n6788 VDD.n6787 92.5005
R4279 VDD.n6947 VDD.n6788 92.5005
R4280 VDD.n6945 VDD.n6944 92.5005
R4281 VDD.n6946 VDD.n6945 92.5005
R4282 VDD.n6943 VDD.n6790 92.5005
R4283 VDD.n6790 VDD.n6789 92.5005
R4284 VDD.n6942 VDD.n6941 92.5005
R4285 VDD.n6941 VDD.n6940 92.5005
R4286 VDD.n6792 VDD.n6791 92.5005
R4287 VDD.n6930 VDD.n6927 92.5005
R4288 VDD.n6933 VDD.n6932 92.5005
R4289 VDD.n7158 VDD.n7157 92.5005
R4290 VDD.n7075 VDD.n6758 92.5005
R4291 VDD.n7077 VDD.n7076 92.5005
R4292 VDD.n7074 VDD.n7073 92.5005
R4293 VDD.n7044 VDD.n7043 92.5005
R4294 VDD.n7068 VDD.n7067 92.5005
R4295 VDD.n7046 VDD.n7045 92.5005
R4296 VDD.n7062 VDD.n7061 92.5005
R4297 VDD.n7058 VDD.n7057 92.5005
R4298 VDD.n7056 VDD.n7055 92.5005
R4299 VDD.n7133 VDD.n7132 92.5005
R4300 VDD.n7137 VDD.n7136 92.5005
R4301 VDD.n7140 VDD.n7139 92.5005
R4302 VDD.n6982 VDD.n6981 92.5005
R4303 VDD.n6971 VDD.n6970 92.5005
R4304 VDD.n7149 VDD.n7148 92.5005
R4305 VDD.n7150 VDD.n6777 92.5005
R4306 VDD.n7153 VDD.n7152 92.5005
R4307 VDD.n7147 VDD.n7146 92.5005
R4308 VDD.n6980 VDD.n6973 92.5005
R4309 VDD.n7142 VDD.n7141 92.5005
R4310 VDD.n7138 VDD.n6979 92.5005
R4311 VDD.n7135 VDD.n7134 92.5005
R4312 VDD.n6983 VDD.n6770 92.5005
R4313 VDD.n7155 VDD.n6770 92.5005
R4314 VDD.n7131 VDD.n7130 92.5005
R4315 VDD.n7050 VDD.n7049 92.5005
R4316 VDD.n7052 VDD.n7051 92.5005
R4317 VDD.n7054 VDD.n7053 92.5005
R4318 VDD.n7060 VDD.n7059 92.5005
R4319 VDD.n7079 VDD.n7078 92.5005
R4320 VDD.n7072 VDD.n7071 92.5005
R4321 VDD.n7070 VDD.n7069 92.5005
R4322 VDD.n7066 VDD.n7065 92.5005
R4323 VDD.n7064 VDD.n7063 92.5005
R4324 VDD.n6687 VDD.n6686 92.5005
R4325 VDD.n6578 VDD.n6577 92.5005
R4326 VDD.n6690 VDD.n6689 92.5005
R4327 VDD.n6691 VDD.n6690 92.5005
R4328 VDD.n6623 VDD.n6622 92.5005
R4329 VDD.n6621 VDD.n6620 92.5005
R4330 VDD.n6611 VDD.n6600 92.5005
R4331 VDD.n6614 VDD.n6613 92.5005
R4332 VDD.n6609 VDD.n6576 92.5005
R4333 VDD.n6625 VDD.n6579 92.5005
R4334 VDD.n6637 VDD.n6636 92.5005
R4335 VDD.n6639 VDD.n6635 92.5005
R4336 VDD.n6642 VDD.n6641 92.5005
R4337 VDD.n6644 VDD.n6643 92.5005
R4338 VDD.n6646 VDD.n6633 92.5005
R4339 VDD.n6649 VDD.n6648 92.5005
R4340 VDD.n6693 VDD.n6692 92.5005
R4341 VDD.n6692 VDD.n6691 92.5005
R4342 VDD.n6575 VDD.n6574 92.5005
R4343 VDD.n6577 VDD.n6575 92.5005
R4344 VDD.n6685 VDD.n6684 92.5005
R4345 VDD.n6686 VDD.n6685 92.5005
R4346 VDD.n6683 VDD.n6682 92.5005
R4347 VDD.n6682 VDD.n6681 92.5005
R4348 VDD.n7304 VDD.n7303 92.5005
R4349 VDD.n7303 VDD.n7302 92.5005
R4350 VDD.n7305 VDD.n6545 92.5005
R4351 VDD.n6549 VDD.n6545 92.5005
R4352 VDD.n7307 VDD.n7306 92.5005
R4353 VDD.n7308 VDD.n7307 92.5005
R4354 VDD.n6546 VDD.n6544 92.5005
R4355 VDD.n7040 VDD.n6544 92.5005
R4356 VDD.n7104 VDD.n7042 92.5005
R4357 VDD.n7042 VDD.n7041 92.5005
R4358 VDD.n7106 VDD.n7105 92.5005
R4359 VDD.n7107 VDD.n7106 92.5005
R4360 VDD.n7086 VDD.n7085 92.5005
R4361 VDD.n7085 VDD.n6993 92.5005
R4362 VDD.n7084 VDD.n7083 92.5005
R4363 VDD.n7084 VDD.n6992 92.5005
R4364 VDD.n7082 VDD.n6987 92.5005
R4365 VDD.n7127 VDD.n6987 92.5005
R4366 VDD.n7081 VDD.n7080 92.5005
R4367 VDD.n7080 VDD.n6974 92.5005
R4368 VDD.n7102 VDD.n7101 92.5005
R4369 VDD.n7099 VDD.n7087 92.5005
R4370 VDD.n7097 VDD.n7096 92.5005
R4371 VDD.n7095 VDD.n7094 92.5005
R4372 VDD.n7092 VDD.n7089 92.5005
R4373 VDD.n7090 VDD.n7003 92.5005
R4374 VDD.n7047 VDD.n6988 92.5005
R4375 VDD.n6988 VDD.n6974 92.5005
R4376 VDD.n7126 VDD.n7125 92.5005
R4377 VDD.n7127 VDD.n7126 92.5005
R4378 VDD.n7123 VDD.n6989 92.5005
R4379 VDD.n6992 VDD.n6989 92.5005
R4380 VDD.n7005 VDD.n6990 92.5005
R4381 VDD.n7005 VDD.n6993 92.5005
R4382 VDD.n7109 VDD.n7108 92.5005
R4383 VDD.n7108 VDD.n7107 92.5005
R4384 VDD.n7010 VDD.n7009 92.5005
R4385 VDD.n7041 VDD.n7010 92.5005
R4386 VDD.n7008 VDD.n6540 92.5005
R4387 VDD.n7040 VDD.n6540 92.5005
R4388 VDD.n7310 VDD.n7309 92.5005
R4389 VDD.n7309 VDD.n7308 92.5005
R4390 VDD.n6553 VDD.n6541 92.5005
R4391 VDD.n6549 VDD.n6541 92.5005
R4392 VDD.n7301 VDD.n7300 92.5005
R4393 VDD.n7302 VDD.n7301 92.5005
R4394 VDD.n6652 VDD.n6582 92.5005
R4395 VDD.n6681 VDD.n6582 92.5005
R4396 VDD.n7124 VDD.n6984 92.5005
R4397 VDD.n6986 VDD.n6984 92.5005
R4398 VDD.n7122 VDD.n7121 92.5005
R4399 VDD.n7121 VDD.n7120 92.5005
R4400 VDD.n7002 VDD.n6991 92.5005
R4401 VDD.n6999 VDD.n6991 92.5005
R4402 VDD.n7113 VDD.n7112 92.5005
R4403 VDD.n7114 VDD.n7113 92.5005
R4404 VDD.n7110 VDD.n7001 92.5005
R4405 VDD.n7011 VDD.n7001 92.5005
R4406 VDD.n7024 VDD.n6538 92.5005
R4407 VDD.n7024 VDD.n6542 92.5005
R4408 VDD.n7023 VDD.n6539 92.5005
R4409 VDD.n7023 VDD.n6543 92.5005
R4410 VDD.n6556 VDD.n6554 92.5005
R4411 VDD.n6556 VDD.n6550 92.5005
R4412 VDD.n7299 VDD.n7298 92.5005
R4413 VDD.n7298 VDD.n6551 92.5005
R4414 VDD.n7297 VDD.n6555 92.5005
R4415 VDD.n7297 VDD.n7296 92.5005
R4416 VDD.n6651 VDD.n6557 92.5005
R4417 VDD.n6680 VDD.n6557 92.5005
R4418 VDD.n7129 VDD.n6985 92.5005
R4419 VDD.n7129 VDD.n7128 92.5005
R4420 VDD.n6117 VDD.n6114 92.5005
R4421 VDD.n6273 VDD.n6117 92.5005
R4422 VDD.n6438 VDD.n5705 92.5005
R4423 VDD.n5825 VDD.n5705 92.5005
R4424 VDD.n6440 VDD.n6439 92.5005
R4425 VDD.n6441 VDD.n6440 92.5005
R4426 VDD.n5706 VDD.n5704 92.5005
R4427 VDD.n5704 VDD.n5696 92.5005
R4428 VDD.n6163 VDD.n6162 92.5005
R4429 VDD.n6163 VDD.n5695 92.5005
R4430 VDD.n6164 VDD.n6161 92.5005
R4431 VDD.n6164 VDD.n5688 92.5005
R4432 VDD.n6166 VDD.n6165 92.5005
R4433 VDD.n6165 VDD.n5687 92.5005
R4434 VDD.n6179 VDD.n6159 92.5005
R4435 VDD.n6178 VDD.n6177 92.5005
R4436 VDD.n6176 VDD.n6175 92.5005
R4437 VDD.n6174 VDD.n6173 92.5005
R4438 VDD.n6172 VDD.n6171 92.5005
R4439 VDD.n6181 VDD.n6180 92.5005
R4440 VDD.n6143 VDD.n6142 92.5005
R4441 VDD.n6156 VDD.n6143 92.5005
R4442 VDD.n6261 VDD.n6260 92.5005
R4443 VDD.n6260 VDD.n6259 92.5005
R4444 VDD.n6262 VDD.n6140 92.5005
R4445 VDD.n6144 VDD.n6140 92.5005
R4446 VDD.n6264 VDD.n6263 92.5005
R4447 VDD.n6265 VDD.n6264 92.5005
R4448 VDD.n6141 VDD.n6139 92.5005
R4449 VDD.n6139 VDD.n6131 92.5005
R4450 VDD.n6304 VDD.n5901 92.5005
R4451 VDD.n5901 VDD.n5900 92.5005
R4452 VDD.n6327 VDD.n6326 92.5005
R4453 VDD.n6326 VDD.n6325 92.5005
R4454 VDD.n5891 VDD.n5890 92.5005
R4455 VDD.n6324 VDD.n5891 92.5005
R4456 VDD.n6322 VDD.n6321 92.5005
R4457 VDD.n6323 VDD.n6322 92.5005
R4458 VDD.n6320 VDD.n5893 92.5005
R4459 VDD.n5893 VDD.n5892 92.5005
R4460 VDD.n6319 VDD.n6318 92.5005
R4461 VDD.n6318 VDD.n6317 92.5005
R4462 VDD.n5895 VDD.n5894 92.5005
R4463 VDD.n6316 VDD.n5895 92.5005
R4464 VDD.n6314 VDD.n6313 92.5005
R4465 VDD.n6315 VDD.n6314 92.5005
R4466 VDD.n6312 VDD.n5897 92.5005
R4467 VDD.n5897 VDD.n5896 92.5005
R4468 VDD.n6311 VDD.n6310 92.5005
R4469 VDD.n6310 VDD.n6309 92.5005
R4470 VDD.n5899 VDD.n5898 92.5005
R4471 VDD.n6308 VDD.n5899 92.5005
R4472 VDD.n6306 VDD.n6305 92.5005
R4473 VDD.n6307 VDD.n6306 92.5005
R4474 VDD.n6328 VDD.n5888 92.5005
R4475 VDD.n5888 VDD.n5887 92.5005
R4476 VDD.n6331 VDD.n6330 92.5005
R4477 VDD.n6332 VDD.n6331 92.5005
R4478 VDD.n6329 VDD.n5889 92.5005
R4479 VDD.n5885 VDD.n5884 92.5005
R4480 VDD.n6336 VDD.n6335 92.5005
R4481 VDD.n6335 VDD.n6334 92.5005
R4482 VDD.n6339 VDD.n6338 92.5005
R4483 VDD.n6340 VDD.n6339 92.5005
R4484 VDD.n5881 VDD.n5880 92.5005
R4485 VDD.n6341 VDD.n5881 92.5005
R4486 VDD.n6344 VDD.n6343 92.5005
R4487 VDD.n6343 VDD.n6342 92.5005
R4488 VDD.n6345 VDD.n5879 92.5005
R4489 VDD.n5879 VDD.n5878 92.5005
R4490 VDD.n6347 VDD.n6346 92.5005
R4491 VDD.n6348 VDD.n6347 92.5005
R4492 VDD.n5877 VDD.n5876 92.5005
R4493 VDD.n6349 VDD.n5877 92.5005
R4494 VDD.n6352 VDD.n6351 92.5005
R4495 VDD.n6351 VDD.n6350 92.5005
R4496 VDD.n6353 VDD.n5875 92.5005
R4497 VDD.n5875 VDD.n5874 92.5005
R4498 VDD.n6355 VDD.n6354 92.5005
R4499 VDD.n6356 VDD.n6355 92.5005
R4500 VDD.n5873 VDD.n5872 92.5005
R4501 VDD.n6357 VDD.n5873 92.5005
R4502 VDD.n6360 VDD.n6359 92.5005
R4503 VDD.n6359 VDD.n6358 92.5005
R4504 VDD.n6361 VDD.n5871 92.5005
R4505 VDD.n5871 VDD.n5870 92.5005
R4506 VDD.n6363 VDD.n6362 92.5005
R4507 VDD.n6364 VDD.n6363 92.5005
R4508 VDD.n5869 VDD.n5868 92.5005
R4509 VDD.n6365 VDD.n5869 92.5005
R4510 VDD.n6368 VDD.n6367 92.5005
R4511 VDD.n6367 VDD.n6366 92.5005
R4512 VDD.n6369 VDD.n5867 92.5005
R4513 VDD.n5867 VDD.n5866 92.5005
R4514 VDD.n6371 VDD.n6370 92.5005
R4515 VDD.n6372 VDD.n6371 92.5005
R4516 VDD.n5865 VDD.n5864 92.5005
R4517 VDD.n6373 VDD.n5865 92.5005
R4518 VDD.n6376 VDD.n6375 92.5005
R4519 VDD.n6375 VDD.n6374 92.5005
R4520 VDD.n6377 VDD.n5863 92.5005
R4521 VDD.n5863 VDD.n5862 92.5005
R4522 VDD.n6379 VDD.n6378 92.5005
R4523 VDD.n6380 VDD.n6379 92.5005
R4524 VDD.n5861 VDD.n5860 92.5005
R4525 VDD.n6381 VDD.n5861 92.5005
R4526 VDD.n6384 VDD.n6383 92.5005
R4527 VDD.n6383 VDD.n6382 92.5005
R4528 VDD.n6385 VDD.n5859 92.5005
R4529 VDD.n5859 VDD.n5858 92.5005
R4530 VDD.n6387 VDD.n6386 92.5005
R4531 VDD.n6388 VDD.n6387 92.5005
R4532 VDD.n5857 VDD.n5856 92.5005
R4533 VDD.n6389 VDD.n5857 92.5005
R4534 VDD.n6394 VDD.n6393 92.5005
R4535 VDD.n6393 VDD.n6392 92.5005
R4536 VDD.n6395 VDD.n5855 92.5005
R4537 VDD.n6391 VDD.n5855 92.5005
R4538 VDD.n6337 VDD.n5883 92.5005
R4539 VDD.n5883 VDD.n5882 92.5005
R4540 VDD.n6409 VDD.n6408 92.5005
R4541 VDD.n6408 VDD.n6407 92.5005
R4542 VDD.n6410 VDD.n5848 92.5005
R4543 VDD.n5848 VDD.n5847 92.5005
R4544 VDD.n6412 VDD.n6411 92.5005
R4545 VDD.n6413 VDD.n6412 92.5005
R4546 VDD.n5846 VDD.n5845 92.5005
R4547 VDD.n6414 VDD.n5846 92.5005
R4548 VDD.n6417 VDD.n6416 92.5005
R4549 VDD.n6416 VDD.n6415 92.5005
R4550 VDD.n6418 VDD.n5844 92.5005
R4551 VDD.n5844 VDD.n5843 92.5005
R4552 VDD.n6420 VDD.n6419 92.5005
R4553 VDD.n6421 VDD.n6420 92.5005
R4554 VDD.n5842 VDD.n5841 92.5005
R4555 VDD.n6422 VDD.n5842 92.5005
R4556 VDD.n6425 VDD.n6424 92.5005
R4557 VDD.n6424 VDD.n6423 92.5005
R4558 VDD.n6426 VDD.n5717 92.5005
R4559 VDD.n5717 VDD.n5715 92.5005
R4560 VDD.n6428 VDD.n6427 92.5005
R4561 VDD.n6429 VDD.n6428 92.5005
R4562 VDD.n6404 VDD.n6403 92.5005
R4563 VDD.n6405 VDD.n6404 92.5005
R4564 VDD.n6402 VDD.n5852 92.5005
R4565 VDD.n5852 VDD.n5851 92.5005
R4566 VDD.n6401 VDD.n6400 92.5005
R4567 VDD.n6398 VDD.n5853 92.5005
R4568 VDD.n6397 VDD.n6396 92.5005
R4569 VDD.n6397 VDD.n5854 92.5005
R4570 VDD.n5850 VDD.n5849 92.5005
R4571 VDD.n6406 VDD.n5850 92.5005
R4572 VDD.n5840 VDD.n5716 92.5005
R4573 VDD.n5772 VDD.n5771 92.5005
R4574 VDD.n5769 VDD.n5741 92.5005
R4575 VDD.n5747 VDD.n5742 92.5005
R4576 VDD.n5764 VDD.n5763 92.5005
R4577 VDD.n5761 VDD.n5760 92.5005
R4578 VDD.n5755 VDD.n5748 92.5005
R4579 VDD.n5753 VDD.n5752 92.5005
R4580 VDD.n5751 VDD.n5718 92.5005
R4581 VDD.n5774 VDD.n5726 92.5005
R4582 VDD.n5776 VDD.n5725 92.5005
R4583 VDD.n5801 VDD.n5800 92.5005
R4584 VDD.n5734 VDD.n5708 92.5005
R4585 VDD.n5820 VDD.n5819 92.5005
R4586 VDD.n5817 VDD.n5816 92.5005
R4587 VDD.n5813 VDD.n5735 92.5005
R4588 VDD.n5810 VDD.n5809 92.5005
R4589 VDD.n5808 VDD.n5807 92.5005
R4590 VDD.n5737 VDD.n5736 92.5005
R4591 VDD.n5812 VDD.n5811 92.5005
R4592 VDD.n5815 VDD.n5814 92.5005
R4593 VDD.n5733 VDD.n5732 92.5005
R4594 VDD.n5822 VDD.n5821 92.5005
R4595 VDD.n6433 VDD.n5707 92.5005
R4596 VDD.n6436 VDD.n6435 92.5005
R4597 VDD.n5806 VDD.n5728 92.5005
R4598 VDD.n5824 VDD.n5728 92.5005
R4599 VDD.n5805 VDD.n5804 92.5005
R4600 VDD.n5803 VDD.n5740 92.5005
R4601 VDD.n6019 VDD.n6018 92.5005
R4602 VDD.n6016 VDD.n5969 92.5005
R4603 VDD.n6015 VDD.n6014 92.5005
R4604 VDD.n6013 VDD.n5970 92.5005
R4605 VDD.n6011 VDD.n6010 92.5005
R4606 VDD.n6009 VDD.n5973 92.5005
R4607 VDD.n5976 VDD.n5973 92.5005
R4608 VDD.n6008 VDD.n6007 92.5005
R4609 VDD.n6007 VDD.n6006 92.5005
R4610 VDD.n5975 VDD.n5974 92.5005
R4611 VDD.n6005 VDD.n5975 92.5005
R4612 VDD.n6003 VDD.n6002 92.5005
R4613 VDD.n6004 VDD.n6003 92.5005
R4614 VDD.n6001 VDD.n5978 92.5005
R4615 VDD.n5978 VDD.n5977 92.5005
R4616 VDD.n6000 VDD.n5999 92.5005
R4617 VDD.n5999 VDD.n5998 92.5005
R4618 VDD.n5980 VDD.n5979 92.5005
R4619 VDD.n5997 VDD.n5980 92.5005
R4620 VDD.n5995 VDD.n5994 92.5005
R4621 VDD.n5996 VDD.n5995 92.5005
R4622 VDD.n5993 VDD.n5982 92.5005
R4623 VDD.n5982 VDD.n5981 92.5005
R4624 VDD.n5992 VDD.n5991 92.5005
R4625 VDD.n5991 VDD.n5990 92.5005
R4626 VDD.n5984 VDD.n5983 92.5005
R4627 VDD.n5989 VDD.n5984 92.5005
R4628 VDD.n5987 VDD.n5986 92.5005
R4629 VDD.n5988 VDD.n5987 92.5005
R4630 VDD.n5985 VDD.n5711 92.5005
R4631 VDD.n5713 VDD.n5711 92.5005
R4632 VDD.n6432 VDD.n5712 92.5005
R4633 VDD.n6432 VDD.n6431 92.5005
R4634 VDD.n6071 VDD.n6070 92.5005
R4635 VDD.n6070 VDD.n6069 92.5005
R4636 VDD.n5943 VDD.n5942 92.5005
R4637 VDD.n6068 VDD.n5943 92.5005
R4638 VDD.n6066 VDD.n6065 92.5005
R4639 VDD.n6067 VDD.n6066 92.5005
R4640 VDD.n6064 VDD.n5945 92.5005
R4641 VDD.n5945 VDD.n5944 92.5005
R4642 VDD.n6063 VDD.n6062 92.5005
R4643 VDD.n6062 VDD.n6061 92.5005
R4644 VDD.n5947 VDD.n5946 92.5005
R4645 VDD.n6060 VDD.n5947 92.5005
R4646 VDD.n6058 VDD.n6057 92.5005
R4647 VDD.n6059 VDD.n6058 92.5005
R4648 VDD.n6056 VDD.n5949 92.5005
R4649 VDD.n5949 VDD.n5948 92.5005
R4650 VDD.n6055 VDD.n6054 92.5005
R4651 VDD.n6054 VDD.n6053 92.5005
R4652 VDD.n5951 VDD.n5950 92.5005
R4653 VDD.n6052 VDD.n5951 92.5005
R4654 VDD.n6050 VDD.n6049 92.5005
R4655 VDD.n6051 VDD.n6050 92.5005
R4656 VDD.n6048 VDD.n5953 92.5005
R4657 VDD.n5953 VDD.n5952 92.5005
R4658 VDD.n6047 VDD.n6046 92.5005
R4659 VDD.n6046 VDD.n6045 92.5005
R4660 VDD.n5955 VDD.n5954 92.5005
R4661 VDD.n6044 VDD.n5955 92.5005
R4662 VDD.n6042 VDD.n6041 92.5005
R4663 VDD.n6043 VDD.n6042 92.5005
R4664 VDD.n6040 VDD.n5957 92.5005
R4665 VDD.n5957 VDD.n5956 92.5005
R4666 VDD.n6039 VDD.n6038 92.5005
R4667 VDD.n6038 VDD.n6037 92.5005
R4668 VDD.n5959 VDD.n5958 92.5005
R4669 VDD.n6036 VDD.n5959 92.5005
R4670 VDD.n6034 VDD.n6033 92.5005
R4671 VDD.n6035 VDD.n6034 92.5005
R4672 VDD.n6032 VDD.n5961 92.5005
R4673 VDD.n5961 VDD.n5960 92.5005
R4674 VDD.n6031 VDD.n6030 92.5005
R4675 VDD.n6030 VDD.n6029 92.5005
R4676 VDD.n5963 VDD.n5962 92.5005
R4677 VDD.n6028 VDD.n5963 92.5005
R4678 VDD.n6026 VDD.n6025 92.5005
R4679 VDD.n6027 VDD.n6026 92.5005
R4680 VDD.n6024 VDD.n5965 92.5005
R4681 VDD.n5965 VDD.n5964 92.5005
R4682 VDD.n6023 VDD.n6022 92.5005
R4683 VDD.n6022 VDD.n6021 92.5005
R4684 VDD.n5967 VDD.n5966 92.5005
R4685 VDD.n6020 VDD.n5967 92.5005
R4686 VDD.n6079 VDD.n5940 92.5005
R4687 VDD.n6083 VDD.n6082 92.5005
R4688 VDD.n5941 VDD.n5939 92.5005
R4689 VDD.n6113 VDD.n5923 92.5005
R4690 VDD.n6109 VDD.n5923 92.5005
R4691 VDD.n6112 VDD.n6111 92.5005
R4692 VDD.n6111 VDD.n6110 92.5005
R4693 VDD.n5925 VDD.n5924 92.5005
R4694 VDD.n6108 VDD.n5925 92.5005
R4695 VDD.n6106 VDD.n6105 92.5005
R4696 VDD.n6107 VDD.n6106 92.5005
R4697 VDD.n6104 VDD.n5927 92.5005
R4698 VDD.n5927 VDD.n5926 92.5005
R4699 VDD.n6103 VDD.n6102 92.5005
R4700 VDD.n6102 VDD.n6101 92.5005
R4701 VDD.n5929 VDD.n5928 92.5005
R4702 VDD.n6100 VDD.n5929 92.5005
R4703 VDD.n6098 VDD.n6097 92.5005
R4704 VDD.n6099 VDD.n6098 92.5005
R4705 VDD.n6096 VDD.n5931 92.5005
R4706 VDD.n5931 VDD.n5930 92.5005
R4707 VDD.n6095 VDD.n6094 92.5005
R4708 VDD.n6094 VDD.n6093 92.5005
R4709 VDD.n5933 VDD.n5932 92.5005
R4710 VDD.n6092 VDD.n5933 92.5005
R4711 VDD.n6090 VDD.n6089 92.5005
R4712 VDD.n6091 VDD.n6090 92.5005
R4713 VDD.n6088 VDD.n5935 92.5005
R4714 VDD.n5935 VDD.n5934 92.5005
R4715 VDD.n6087 VDD.n6086 92.5005
R4716 VDD.n6086 VDD.n6085 92.5005
R4717 VDD.n5937 VDD.n5936 92.5005
R4718 VDD.n6075 VDD.n6072 92.5005
R4719 VDD.n6078 VDD.n6077 92.5005
R4720 VDD.n6303 VDD.n6302 92.5005
R4721 VDD.n6220 VDD.n5903 92.5005
R4722 VDD.n6222 VDD.n6221 92.5005
R4723 VDD.n6219 VDD.n6218 92.5005
R4724 VDD.n6189 VDD.n6188 92.5005
R4725 VDD.n6213 VDD.n6212 92.5005
R4726 VDD.n6191 VDD.n6190 92.5005
R4727 VDD.n6207 VDD.n6206 92.5005
R4728 VDD.n6203 VDD.n6202 92.5005
R4729 VDD.n6201 VDD.n6200 92.5005
R4730 VDD.n6278 VDD.n6277 92.5005
R4731 VDD.n6282 VDD.n6281 92.5005
R4732 VDD.n6285 VDD.n6284 92.5005
R4733 VDD.n6127 VDD.n6126 92.5005
R4734 VDD.n6116 VDD.n6115 92.5005
R4735 VDD.n6294 VDD.n6293 92.5005
R4736 VDD.n6295 VDD.n5922 92.5005
R4737 VDD.n6298 VDD.n6297 92.5005
R4738 VDD.n6292 VDD.n6291 92.5005
R4739 VDD.n6125 VDD.n6118 92.5005
R4740 VDD.n6287 VDD.n6286 92.5005
R4741 VDD.n6283 VDD.n6124 92.5005
R4742 VDD.n6280 VDD.n6279 92.5005
R4743 VDD.n6128 VDD.n5915 92.5005
R4744 VDD.n6300 VDD.n5915 92.5005
R4745 VDD.n6276 VDD.n6275 92.5005
R4746 VDD.n6195 VDD.n6194 92.5005
R4747 VDD.n6197 VDD.n6196 92.5005
R4748 VDD.n6199 VDD.n6198 92.5005
R4749 VDD.n6205 VDD.n6204 92.5005
R4750 VDD.n6224 VDD.n6223 92.5005
R4751 VDD.n6217 VDD.n6216 92.5005
R4752 VDD.n6215 VDD.n6214 92.5005
R4753 VDD.n6211 VDD.n6210 92.5005
R4754 VDD.n6209 VDD.n6208 92.5005
R4755 VDD.n5832 VDD.n5831 92.5005
R4756 VDD.n5723 VDD.n5722 92.5005
R4757 VDD.n5835 VDD.n5834 92.5005
R4758 VDD.n5836 VDD.n5835 92.5005
R4759 VDD.n5768 VDD.n5767 92.5005
R4760 VDD.n5766 VDD.n5765 92.5005
R4761 VDD.n5756 VDD.n5745 92.5005
R4762 VDD.n5759 VDD.n5758 92.5005
R4763 VDD.n5754 VDD.n5721 92.5005
R4764 VDD.n5770 VDD.n5724 92.5005
R4765 VDD.n5782 VDD.n5781 92.5005
R4766 VDD.n5784 VDD.n5780 92.5005
R4767 VDD.n5787 VDD.n5786 92.5005
R4768 VDD.n5789 VDD.n5788 92.5005
R4769 VDD.n5791 VDD.n5778 92.5005
R4770 VDD.n5794 VDD.n5793 92.5005
R4771 VDD.n5838 VDD.n5837 92.5005
R4772 VDD.n5837 VDD.n5836 92.5005
R4773 VDD.n5720 VDD.n5719 92.5005
R4774 VDD.n5722 VDD.n5720 92.5005
R4775 VDD.n5830 VDD.n5829 92.5005
R4776 VDD.n5831 VDD.n5830 92.5005
R4777 VDD.n5828 VDD.n5827 92.5005
R4778 VDD.n5827 VDD.n5826 92.5005
R4779 VDD.n6449 VDD.n6448 92.5005
R4780 VDD.n6448 VDD.n6447 92.5005
R4781 VDD.n6450 VDD.n5690 92.5005
R4782 VDD.n5694 VDD.n5690 92.5005
R4783 VDD.n6452 VDD.n6451 92.5005
R4784 VDD.n6453 VDD.n6452 92.5005
R4785 VDD.n5691 VDD.n5689 92.5005
R4786 VDD.n6185 VDD.n5689 92.5005
R4787 VDD.n6249 VDD.n6187 92.5005
R4788 VDD.n6187 VDD.n6186 92.5005
R4789 VDD.n6251 VDD.n6250 92.5005
R4790 VDD.n6252 VDD.n6251 92.5005
R4791 VDD.n6231 VDD.n6230 92.5005
R4792 VDD.n6230 VDD.n6138 92.5005
R4793 VDD.n6229 VDD.n6228 92.5005
R4794 VDD.n6229 VDD.n6137 92.5005
R4795 VDD.n6227 VDD.n6132 92.5005
R4796 VDD.n6272 VDD.n6132 92.5005
R4797 VDD.n6226 VDD.n6225 92.5005
R4798 VDD.n6225 VDD.n6119 92.5005
R4799 VDD.n6247 VDD.n6246 92.5005
R4800 VDD.n6244 VDD.n6232 92.5005
R4801 VDD.n6242 VDD.n6241 92.5005
R4802 VDD.n6240 VDD.n6239 92.5005
R4803 VDD.n6237 VDD.n6234 92.5005
R4804 VDD.n6235 VDD.n6148 92.5005
R4805 VDD.n6192 VDD.n6133 92.5005
R4806 VDD.n6133 VDD.n6119 92.5005
R4807 VDD.n6271 VDD.n6270 92.5005
R4808 VDD.n6272 VDD.n6271 92.5005
R4809 VDD.n6268 VDD.n6134 92.5005
R4810 VDD.n6137 VDD.n6134 92.5005
R4811 VDD.n6150 VDD.n6135 92.5005
R4812 VDD.n6150 VDD.n6138 92.5005
R4813 VDD.n6254 VDD.n6253 92.5005
R4814 VDD.n6253 VDD.n6252 92.5005
R4815 VDD.n6155 VDD.n6154 92.5005
R4816 VDD.n6186 VDD.n6155 92.5005
R4817 VDD.n6153 VDD.n5685 92.5005
R4818 VDD.n6185 VDD.n5685 92.5005
R4819 VDD.n6455 VDD.n6454 92.5005
R4820 VDD.n6454 VDD.n6453 92.5005
R4821 VDD.n5698 VDD.n5686 92.5005
R4822 VDD.n5694 VDD.n5686 92.5005
R4823 VDD.n6446 VDD.n6445 92.5005
R4824 VDD.n6447 VDD.n6446 92.5005
R4825 VDD.n5797 VDD.n5727 92.5005
R4826 VDD.n5826 VDD.n5727 92.5005
R4827 VDD.n6269 VDD.n6129 92.5005
R4828 VDD.n6131 VDD.n6129 92.5005
R4829 VDD.n6267 VDD.n6266 92.5005
R4830 VDD.n6266 VDD.n6265 92.5005
R4831 VDD.n6147 VDD.n6136 92.5005
R4832 VDD.n6144 VDD.n6136 92.5005
R4833 VDD.n6258 VDD.n6257 92.5005
R4834 VDD.n6259 VDD.n6258 92.5005
R4835 VDD.n6255 VDD.n6146 92.5005
R4836 VDD.n6156 VDD.n6146 92.5005
R4837 VDD.n6169 VDD.n5683 92.5005
R4838 VDD.n6169 VDD.n5687 92.5005
R4839 VDD.n6168 VDD.n5684 92.5005
R4840 VDD.n6168 VDD.n5688 92.5005
R4841 VDD.n5701 VDD.n5699 92.5005
R4842 VDD.n5701 VDD.n5695 92.5005
R4843 VDD.n6444 VDD.n6443 92.5005
R4844 VDD.n6443 VDD.n5696 92.5005
R4845 VDD.n6442 VDD.n5700 92.5005
R4846 VDD.n6442 VDD.n6441 92.5005
R4847 VDD.n5796 VDD.n5702 92.5005
R4848 VDD.n5825 VDD.n5702 92.5005
R4849 VDD.n6274 VDD.n6130 92.5005
R4850 VDD.n6274 VDD.n6273 92.5005
R4851 VDD.n5449 VDD.n282 92.5005
R4852 VDD.n274 VDD.n272 92.5005
R4853 VDD.n272 VDD.n270 92.5005
R4854 VDD.n5441 VDD.n5440 92.5005
R4855 VDD.n5442 VDD.n5441 92.5005
R4856 VDD.n5445 VDD.n5444 92.5005
R4857 VDD.n5444 VDD.n5443 92.5005
R4858 VDD.n4289 VDD.n4288 92.5005
R4859 VDD.n4288 VDD.n4287 92.5005
R4860 VDD.n2366 VDD.n2364 92.5005
R4861 VDD.n4286 VDD.n2366 92.5005
R4862 VDD.n4284 VDD.n4283 92.5005
R4863 VDD.n4285 VDD.n4284 92.5005
R4864 VDD.n2371 VDD.n2369 92.5005
R4865 VDD.n2369 VDD.n2368 92.5005
R4866 VDD.n4278 VDD.n4277 92.5005
R4867 VDD.n4277 VDD.n4276 92.5005
R4868 VDD.n2377 VDD.n2374 92.5005
R4869 VDD.n4275 VDD.n2374 92.5005
R4870 VDD.n4273 VDD.n4272 92.5005
R4871 VDD.n4274 VDD.n4273 92.5005
R4872 VDD.n2379 VDD.n2376 92.5005
R4873 VDD.n2376 VDD.n2375 92.5005
R4874 VDD.n4267 VDD.n4266 92.5005
R4875 VDD.n4266 VDD.n4265 92.5005
R4876 VDD.n2386 VDD.n2383 92.5005
R4877 VDD.n4264 VDD.n2383 92.5005
R4878 VDD.n4262 VDD.n4261 92.5005
R4879 VDD.n4263 VDD.n4262 92.5005
R4880 VDD.n2388 VDD.n2385 92.5005
R4881 VDD.n2385 VDD.n2384 92.5005
R4882 VDD.n4256 VDD.n4255 92.5005
R4883 VDD.n4255 VDD.n4254 92.5005
R4884 VDD.n2395 VDD.n2392 92.5005
R4885 VDD.n4253 VDD.n2392 92.5005
R4886 VDD.n4251 VDD.n4250 92.5005
R4887 VDD.n4252 VDD.n4251 92.5005
R4888 VDD.n2397 VDD.n2394 92.5005
R4889 VDD.n2394 VDD.n2393 92.5005
R4890 VDD.n4245 VDD.n4244 92.5005
R4891 VDD.n4244 VDD.n4243 92.5005
R4892 VDD.n2403 VDD.n2401 92.5005
R4893 VDD.n4242 VDD.n2401 92.5005
R4894 VDD.n4240 VDD.n4239 92.5005
R4895 VDD.n4241 VDD.n4240 92.5005
R4896 VDD.n4238 VDD.n2402 92.5005
R4897 VDD.n2411 VDD.n2402 92.5005
R4898 VDD.n2409 VDD.n2405 92.5005
R4899 VDD.n2412 VDD.n2409 92.5005
R4900 VDD.n4233 VDD.n4232 92.5005
R4901 VDD.n4232 VDD.n4231 92.5005
R4902 VDD.n2415 VDD.n2410 92.5005
R4903 VDD.n4230 VDD.n2410 92.5005
R4904 VDD.n4228 VDD.n4227 92.5005
R4905 VDD.n4229 VDD.n4228 92.5005
R4906 VDD.n2417 VDD.n2414 92.5005
R4907 VDD.n2414 VDD.n2413 92.5005
R4908 VDD.n4222 VDD.n4221 92.5005
R4909 VDD.n4221 VDD.n4220 92.5005
R4910 VDD.n2424 VDD.n2421 92.5005
R4911 VDD.n4219 VDD.n2421 92.5005
R4912 VDD.n4217 VDD.n4216 92.5005
R4913 VDD.n4218 VDD.n4217 92.5005
R4914 VDD.n2426 VDD.n2423 92.5005
R4915 VDD.n2423 VDD.n2422 92.5005
R4916 VDD.n4211 VDD.n4210 92.5005
R4917 VDD.n4210 VDD.n4209 92.5005
R4918 VDD.n2433 VDD.n2430 92.5005
R4919 VDD.n4208 VDD.n2430 92.5005
R4920 VDD.n4206 VDD.n4205 92.5005
R4921 VDD.n4207 VDD.n4206 92.5005
R4922 VDD.n2435 VDD.n2432 92.5005
R4923 VDD.n2432 VDD.n2431 92.5005
R4924 VDD.n4200 VDD.n4199 92.5005
R4925 VDD.n4199 VDD.n4198 92.5005
R4926 VDD.n4086 VDD.n2439 92.5005
R4927 VDD.n2440 VDD.n2439 92.5005
R4928 VDD.n4084 VDD.n4083 92.5005
R4929 VDD.n4083 VDD.n4082 92.5005
R4930 VDD.n4093 VDD.n4092 92.5005
R4931 VDD.n4094 VDD.n4093 92.5005
R4932 VDD.n4091 VDD.n4081 92.5005
R4933 VDD.n4095 VDD.n4081 92.5005
R4934 VDD.n4098 VDD.n4097 92.5005
R4935 VDD.n4097 VDD.n4096 92.5005
R4936 VDD.n4099 VDD.n4076 92.5005
R4937 VDD.n4076 VDD.n4075 92.5005
R4938 VDD.n4106 VDD.n4105 92.5005
R4939 VDD.n4107 VDD.n4106 92.5005
R4940 VDD.n4078 VDD.n4074 92.5005
R4941 VDD.n4108 VDD.n4074 92.5005
R4942 VDD.n4111 VDD.n4110 92.5005
R4943 VDD.n4110 VDD.n4109 92.5005
R4944 VDD.n4112 VDD.n4069 92.5005
R4945 VDD.n4069 VDD.n4068 92.5005
R4946 VDD.n4119 VDD.n4118 92.5005
R4947 VDD.n4120 VDD.n4119 92.5005
R4948 VDD.n4071 VDD.n4067 92.5005
R4949 VDD.n4121 VDD.n4067 92.5005
R4950 VDD.n4125 VDD.n4124 92.5005
R4951 VDD.n4124 VDD.n4123 92.5005
R4952 VDD.n4126 VDD.n4062 92.5005
R4953 VDD.n4122 VDD.n4062 92.5005
R4954 VDD.n4133 VDD.n4132 92.5005
R4955 VDD.n4134 VDD.n4133 92.5005
R4956 VDD.n4064 VDD.n4061 92.5005
R4957 VDD.n4135 VDD.n4061 92.5005
R4958 VDD.n4138 VDD.n4137 92.5005
R4959 VDD.n4137 VDD.n4136 92.5005
R4960 VDD.n4058 VDD.n4057 92.5005
R4961 VDD.n4057 VDD.n4056 92.5005
R4962 VDD.n4145 VDD.n4144 92.5005
R4963 VDD.n4146 VDD.n4145 92.5005
R4964 VDD.n4055 VDD.n4053 92.5005
R4965 VDD.n4147 VDD.n4055 92.5005
R4966 VDD.n4150 VDD.n4149 92.5005
R4967 VDD.n4149 VDD.n4148 92.5005
R4968 VDD.n4054 VDD.n4049 92.5005
R4969 VDD.n4049 VDD.n4048 92.5005
R4970 VDD.n4157 VDD.n4156 92.5005
R4971 VDD.n4158 VDD.n4157 92.5005
R4972 VDD.n4051 VDD.n4047 92.5005
R4973 VDD.n4159 VDD.n4047 92.5005
R4974 VDD.n4162 VDD.n4161 92.5005
R4975 VDD.n4161 VDD.n4160 92.5005
R4976 VDD.n4163 VDD.n4042 92.5005
R4977 VDD.n4042 VDD.n4041 92.5005
R4978 VDD.n4170 VDD.n4169 92.5005
R4979 VDD.n4171 VDD.n4170 92.5005
R4980 VDD.n4044 VDD.n4040 92.5005
R4981 VDD.n4172 VDD.n4040 92.5005
R4982 VDD.n4175 VDD.n4174 92.5005
R4983 VDD.n4174 VDD.n4173 92.5005
R4984 VDD.n4176 VDD.n4035 92.5005
R4985 VDD.n4035 VDD.n4034 92.5005
R4986 VDD.n4183 VDD.n4182 92.5005
R4987 VDD.n4184 VDD.n4183 92.5005
R4988 VDD.n4037 VDD.n4032 92.5005
R4989 VDD.n4185 VDD.n4032 92.5005
R4990 VDD.n4189 VDD.n4188 92.5005
R4991 VDD.n4188 VDD.n4187 92.5005
R4992 VDD.n4033 VDD.n4029 92.5005
R4993 VDD.n4186 VDD.n4033 92.5005
R4994 VDD.n4194 VDD.n271 92.5005
R4995 VDD.n271 VDD.n268 92.5005
R4996 VDD.n5458 VDD.n5457 92.5005
R4997 VDD.n5459 VDD.n5458 92.5005
R4998 VDD.n1887 VDD.n1886 92.5005
R4999 VDD.n1036 VDD.n1035 92.5005
R5000 VDD.n1707 VDD.n1706 92.5005
R5001 VDD.n1709 VDD.n1708 92.5005
R5002 VDD.n1711 VDD.n1710 92.5005
R5003 VDD.n1713 VDD.n1712 92.5005
R5004 VDD.n1715 VDD.n1714 92.5005
R5005 VDD.n1717 VDD.n1716 92.5005
R5006 VDD.n1719 VDD.n1718 92.5005
R5007 VDD.n1721 VDD.n1720 92.5005
R5008 VDD.n1723 VDD.n1722 92.5005
R5009 VDD.n1725 VDD.n1724 92.5005
R5010 VDD.n2471 VDD.n2470 92.5005
R5011 VDD.n2469 VDD.n2468 92.5005
R5012 VDD.n2467 VDD.n2466 92.5005
R5013 VDD.n2463 VDD.n2462 92.5005
R5014 VDD.n4023 VDD.n4022 92.5005
R5015 VDD.n4020 VDD.n2365 92.5005
R5016 VDD.n2367 VDD.n2365 92.5005
R5017 VDD.n1404 VDD.n1403 92.5005
R5018 VDD.n1456 VDD.n1405 92.5005
R5019 VDD.n1458 VDD.n1457 92.5005
R5020 VDD.n1446 VDD.n1409 92.5005
R5021 VDD.n1448 VDD.n1447 92.5005
R5022 VDD.n1438 VDD.n1410 92.5005
R5023 VDD.n1440 VDD.n1439 92.5005
R5024 VDD.n1428 VDD.n1415 92.5005
R5025 VDD.n1430 VDD.n1429 92.5005
R5026 VDD.n1417 VDD.n1416 92.5005
R5027 VDD.n1422 VDD.n1386 92.5005
R5028 VDD.n1478 VDD.n1477 92.5005
R5029 VDD.n1467 VDD.n1399 92.5005
R5030 VDD.n1401 VDD.n1400 92.5005
R5031 VDD.n1462 VDD.n1461 92.5005
R5032 VDD.n1460 VDD.n1459 92.5005
R5033 VDD.n1449 VDD.n1407 92.5005
R5034 VDD.n1451 VDD.n1450 92.5005
R5035 VDD.n1444 VDD.n1443 92.5005
R5036 VDD.n1442 VDD.n1441 92.5005
R5037 VDD.n1431 VDD.n1412 92.5005
R5038 VDD.n1433 VDD.n1432 92.5005
R5039 VDD.n1426 VDD.n1425 92.5005
R5040 VDD.n1424 VDD.n1423 92.5005
R5041 VDD.n1421 VDD.n1389 92.5005
R5042 VDD.n1476 VDD.n1475 92.5005
R5043 VDD.n1475 VDD.n1474 92.5005
R5044 VDD.n1468 VDD.n1376 92.5005
R5045 VDD.n1380 VDD.n1376 92.5005
R5046 VDD.n1482 VDD.n1379 92.5005
R5047 VDD.n1482 VDD.n1481 92.5005
R5048 VDD.n1488 VDD.n1487 92.5005
R5049 VDD.n1487 VDD.n1486 92.5005
R5050 VDD.n1371 VDD.n1365 92.5005
R5051 VDD.n1369 VDD.n1365 92.5005
R5052 VDD.n1498 VDD.n1368 92.5005
R5053 VDD.n1498 VDD.n1497 92.5005
R5054 VDD.n1499 VDD.n1362 92.5005
R5055 VDD.n1500 VDD.n1499 92.5005
R5056 VDD.n1505 VDD.n1359 92.5005
R5057 VDD.n1501 VDD.n1359 92.5005
R5058 VDD.n1511 VDD.n1510 92.5005
R5059 VDD.n1512 VDD.n1511 92.5005
R5060 VDD.n1355 VDD.n1352 92.5005
R5061 VDD.n1353 VDD.n1352 92.5005
R5062 VDD.n1520 VDD.n1519 92.5005
R5063 VDD.n1519 VDD.n1518 92.5005
R5064 VDD.n1525 VDD.n1346 92.5005
R5065 VDD.n1347 VDD.n1346 92.5005
R5066 VDD.n1532 VDD.n1531 92.5005
R5067 VDD.n1531 VDD.n1530 92.5005
R5068 VDD.n1343 VDD.n1337 92.5005
R5069 VDD.n1341 VDD.n1337 92.5005
R5070 VDD.n1542 VDD.n1340 92.5005
R5071 VDD.n1542 VDD.n1541 92.5005
R5072 VDD.n1543 VDD.n1334 92.5005
R5073 VDD.n1544 VDD.n1543 92.5005
R5074 VDD.n1549 VDD.n1331 92.5005
R5075 VDD.n1545 VDD.n1331 92.5005
R5076 VDD.n1555 VDD.n1554 92.5005
R5077 VDD.n1556 VDD.n1555 92.5005
R5078 VDD.n1327 VDD.n1324 92.5005
R5079 VDD.n1325 VDD.n1324 92.5005
R5080 VDD.n1564 VDD.n1563 92.5005
R5081 VDD.n1563 VDD.n1562 92.5005
R5082 VDD.n1320 VDD.n1314 92.5005
R5083 VDD.n1318 VDD.n1314 92.5005
R5084 VDD.n1573 VDD.n1317 92.5005
R5085 VDD.n1573 VDD.n1572 92.5005
R5086 VDD.n1574 VDD.n1311 92.5005
R5087 VDD.n1575 VDD.n1574 92.5005
R5088 VDD.n1580 VDD.n1308 92.5005
R5089 VDD.n1576 VDD.n1308 92.5005
R5090 VDD.n1586 VDD.n1585 92.5005
R5091 VDD.n1587 VDD.n1586 92.5005
R5092 VDD.n1304 VDD.n1301 92.5005
R5093 VDD.n1302 VDD.n1301 92.5005
R5094 VDD.n1595 VDD.n1594 92.5005
R5095 VDD.n1594 VDD.n1593 92.5005
R5096 VDD.n1600 VDD.n1295 92.5005
R5097 VDD.n1296 VDD.n1295 92.5005
R5098 VDD.n1607 VDD.n1606 92.5005
R5099 VDD.n1606 VDD.n1605 92.5005
R5100 VDD.n1292 VDD.n1286 92.5005
R5101 VDD.n1290 VDD.n1286 92.5005
R5102 VDD.n1618 VDD.n1289 92.5005
R5103 VDD.n1618 VDD.n1617 92.5005
R5104 VDD.n1619 VDD.n1280 92.5005
R5105 VDD.n1619 VDD.n1276 92.5005
R5106 VDD.n1620 VDD.n1281 92.5005
R5107 VDD.n1620 VDD.n1277 92.5005
R5108 VDD.n1807 VDD.n1806 92.5005
R5109 VDD.n1806 VDD.n1805 92.5005
R5110 VDD.n1626 VDD.n1621 92.5005
R5111 VDD.n1623 VDD.n1621 92.5005
R5112 VDD.n1799 VDD.n1798 92.5005
R5113 VDD.n1800 VDD.n1799 92.5005
R5114 VDD.n1631 VDD.n1629 92.5005
R5115 VDD.n1637 VDD.n1629 92.5005
R5116 VDD.n1792 VDD.n1791 92.5005
R5117 VDD.n1791 VDD.n1790 92.5005
R5118 VDD.n1642 VDD.n1636 92.5005
R5119 VDD.n1639 VDD.n1636 92.5005
R5120 VDD.n1784 VDD.n1783 92.5005
R5121 VDD.n1785 VDD.n1784 92.5005
R5122 VDD.n1649 VDD.n1646 92.5005
R5123 VDD.n1653 VDD.n1646 92.5005
R5124 VDD.n1778 VDD.n1777 92.5005
R5125 VDD.n1777 VDD.n1776 92.5005
R5126 VDD.n1659 VDD.n1652 92.5005
R5127 VDD.n1655 VDD.n1652 92.5005
R5128 VDD.n1770 VDD.n1769 92.5005
R5129 VDD.n1771 VDD.n1770 92.5005
R5130 VDD.n1664 VDD.n1662 92.5005
R5131 VDD.n1670 VDD.n1662 92.5005
R5132 VDD.n1763 VDD.n1762 92.5005
R5133 VDD.n1762 VDD.n1761 92.5005
R5134 VDD.n1676 VDD.n1669 92.5005
R5135 VDD.n1672 VDD.n1669 92.5005
R5136 VDD.n1755 VDD.n1754 92.5005
R5137 VDD.n1756 VDD.n1755 92.5005
R5138 VDD.n1681 VDD.n1679 92.5005
R5139 VDD.n1687 VDD.n1679 92.5005
R5140 VDD.n1748 VDD.n1747 92.5005
R5141 VDD.n1747 VDD.n1746 92.5005
R5142 VDD.n1693 VDD.n1686 92.5005
R5143 VDD.n1689 VDD.n1686 92.5005
R5144 VDD.n1740 VDD.n1739 92.5005
R5145 VDD.n1741 VDD.n1740 92.5005
R5146 VDD.n1698 VDD.n1696 92.5005
R5147 VDD.n1726 VDD.n1696 92.5005
R5148 VDD.n1733 VDD.n1732 92.5005
R5149 VDD.n1732 VDD.n1731 92.5005
R5150 VDD.n1882 VDD.n1881 92.5005
R5151 VDD.n1883 VDD.n1882 92.5005
R5152 VDD.n1704 VDD.n1044 92.5005
R5153 VDD.n1044 VDD.n1037 92.5005
R5154 VDD.n1729 VDD.n1702 92.5005
R5155 VDD.n1730 VDD.n1729 92.5005
R5156 VDD.n1728 VDD.n1701 92.5005
R5157 VDD.n1728 VDD.n1727 92.5005
R5158 VDD.n1738 VDD.n1691 92.5005
R5159 VDD.n1695 VDD.n1691 92.5005
R5160 VDD.n1743 VDD.n1694 92.5005
R5161 VDD.n1743 VDD.n1742 92.5005
R5162 VDD.n1744 VDD.n1685 92.5005
R5163 VDD.n1745 VDD.n1744 92.5005
R5164 VDD.n1690 VDD.n1684 92.5005
R5165 VDD.n1690 VDD.n1688 92.5005
R5166 VDD.n1753 VDD.n1674 92.5005
R5167 VDD.n1678 VDD.n1674 92.5005
R5168 VDD.n1758 VDD.n1677 92.5005
R5169 VDD.n1758 VDD.n1757 92.5005
R5170 VDD.n1759 VDD.n1668 92.5005
R5171 VDD.n1760 VDD.n1759 92.5005
R5172 VDD.n1673 VDD.n1667 92.5005
R5173 VDD.n1673 VDD.n1671 92.5005
R5174 VDD.n1768 VDD.n1657 92.5005
R5175 VDD.n1661 VDD.n1657 92.5005
R5176 VDD.n1773 VDD.n1660 92.5005
R5177 VDD.n1773 VDD.n1772 92.5005
R5178 VDD.n1774 VDD.n1651 92.5005
R5179 VDD.n1775 VDD.n1774 92.5005
R5180 VDD.n1656 VDD.n1650 92.5005
R5181 VDD.n1656 VDD.n1654 92.5005
R5182 VDD.n1647 VDD.n1641 92.5005
R5183 VDD.n1645 VDD.n1641 92.5005
R5184 VDD.n1787 VDD.n1644 92.5005
R5185 VDD.n1787 VDD.n1786 92.5005
R5186 VDD.n1788 VDD.n1635 92.5005
R5187 VDD.n1789 VDD.n1788 92.5005
R5188 VDD.n1640 VDD.n1634 92.5005
R5189 VDD.n1640 VDD.n1638 92.5005
R5190 VDD.n1797 VDD.n1624 92.5005
R5191 VDD.n1628 VDD.n1624 92.5005
R5192 VDD.n1802 VDD.n1627 92.5005
R5193 VDD.n1802 VDD.n1801 92.5005
R5194 VDD.n1803 VDD.n1285 92.5005
R5195 VDD.n1804 VDD.n1803 92.5005
R5196 VDD.n1284 VDD.n1279 92.5005
R5197 VDD.n1622 VDD.n1279 92.5005
R5198 VDD.n1813 VDD.n1812 92.5005
R5199 VDD.n1814 VDD.n1813 92.5005
R5200 VDD.n1288 VDD.n1278 92.5005
R5201 VDD.n1616 VDD.n1278 92.5005
R5202 VDD.n1614 VDD.n1613 92.5005
R5203 VDD.n1615 VDD.n1614 92.5005
R5204 VDD.n1608 VDD.n1291 92.5005
R5205 VDD.n1604 VDD.n1291 92.5005
R5206 VDD.n1602 VDD.n1601 92.5005
R5207 VDD.n1603 VDD.n1602 92.5005
R5208 VDD.n1298 VDD.n1297 92.5005
R5209 VDD.n1592 VDD.n1297 92.5005
R5210 VDD.n1590 VDD.n1300 92.5005
R5211 VDD.n1591 VDD.n1590 92.5005
R5212 VDD.n1589 VDD.n1306 92.5005
R5213 VDD.n1589 VDD.n1588 92.5005
R5214 VDD.n1309 VDD.n1303 92.5005
R5215 VDD.n1307 VDD.n1303 92.5005
R5216 VDD.n1579 VDD.n1578 92.5005
R5217 VDD.n1578 VDD.n1577 92.5005
R5218 VDD.n1315 VDD.n1312 92.5005
R5219 VDD.n1313 VDD.n1312 92.5005
R5220 VDD.n1570 VDD.n1569 92.5005
R5221 VDD.n1571 VDD.n1570 92.5005
R5222 VDD.n1323 VDD.n1319 92.5005
R5223 VDD.n1561 VDD.n1319 92.5005
R5224 VDD.n1559 VDD.n1322 92.5005
R5225 VDD.n1560 VDD.n1559 92.5005
R5226 VDD.n1558 VDD.n1329 92.5005
R5227 VDD.n1558 VDD.n1557 92.5005
R5228 VDD.n1332 VDD.n1326 92.5005
R5229 VDD.n1330 VDD.n1326 92.5005
R5230 VDD.n1548 VDD.n1547 92.5005
R5231 VDD.n1547 VDD.n1546 92.5005
R5232 VDD.n1339 VDD.n1335 92.5005
R5233 VDD.n1336 VDD.n1335 92.5005
R5234 VDD.n1539 VDD.n1538 92.5005
R5235 VDD.n1540 VDD.n1539 92.5005
R5236 VDD.n1533 VDD.n1342 92.5005
R5237 VDD.n1529 VDD.n1342 92.5005
R5238 VDD.n1527 VDD.n1526 92.5005
R5239 VDD.n1528 VDD.n1527 92.5005
R5240 VDD.n1349 VDD.n1348 92.5005
R5241 VDD.n1517 VDD.n1348 92.5005
R5242 VDD.n1515 VDD.n1351 92.5005
R5243 VDD.n1516 VDD.n1515 92.5005
R5244 VDD.n1514 VDD.n1357 92.5005
R5245 VDD.n1514 VDD.n1513 92.5005
R5246 VDD.n1360 VDD.n1354 92.5005
R5247 VDD.n1358 VDD.n1354 92.5005
R5248 VDD.n1504 VDD.n1503 92.5005
R5249 VDD.n1503 VDD.n1502 92.5005
R5250 VDD.n1367 VDD.n1363 92.5005
R5251 VDD.n1364 VDD.n1363 92.5005
R5252 VDD.n1495 VDD.n1494 92.5005
R5253 VDD.n1496 VDD.n1495 92.5005
R5254 VDD.n1489 VDD.n1370 92.5005
R5255 VDD.n1485 VDD.n1370 92.5005
R5256 VDD.n1483 VDD.n1373 92.5005
R5257 VDD.n1484 VDD.n1483 92.5005
R5258 VDD.n1378 VDD.n1374 92.5005
R5259 VDD.n1375 VDD.n1374 92.5005
R5260 VDD.n1471 VDD.n1470 92.5005
R5261 VDD.n1470 VDD.n1391 92.5005
R5262 VDD.n1474 VDD.n1398 92.5005
R5263 VDD.n1865 VDD.n1864 92.5005
R5264 VDD.n1864 VDD.n1863 92.5005
R5265 VDD.n1055 VDD.n1053 92.5005
R5266 VDD.n1053 VDD.n1052 92.5005
R5267 VDD.n1871 VDD.n1870 92.5005
R5268 VDD.n1872 VDD.n1871 92.5005
R5269 VDD.n1051 VDD.n1050 92.5005
R5270 VDD.n1873 VDD.n1051 92.5005
R5271 VDD.n1876 VDD.n1875 92.5005
R5272 VDD.n1875 VDD.n1874 92.5005
R5273 VDD.n1047 VDD.n1045 92.5005
R5274 VDD.n1045 VDD.n1043 92.5005
R5275 VDD.n1819 VDD.n1818 92.5005
R5276 VDD.n1086 VDD.n1083 92.5005
R5277 VDD.n1825 VDD.n1824 92.5005
R5278 VDD.n1828 VDD.n1827 92.5005
R5279 VDD.n1080 VDD.n1077 92.5005
R5280 VDD.n1834 VDD.n1833 92.5005
R5281 VDD.n1836 VDD.n1072 92.5005
R5282 VDD.n1839 VDD.n1838 92.5005
R5283 VDD.n1073 VDD.n1070 92.5005
R5284 VDD.n1845 VDD.n1844 92.5005
R5285 VDD.n1848 VDD.n1847 92.5005
R5286 VDD.n1067 VDD.n1064 92.5005
R5287 VDD.n1854 VDD.n1853 92.5005
R5288 VDD.n1857 VDD.n1856 92.5005
R5289 VDD.n1859 VDD.n1858 92.5005
R5290 VDD.n1861 VDD.n1860 92.5005
R5291 VDD.n1862 VDD.n1058 92.5005
R5292 VDD.n279 VDD.n277 92.5005
R5293 VDD.n5452 VDD.n5451 92.5005
R5294 VDD.n296 VDD.n280 92.5005
R5295 VDD.n5438 VDD.n5437 92.5005
R5296 VDD.n298 VDD.n295 92.5005
R5297 VDD.n5432 VDD.n5431 92.5005
R5298 VDD.n5429 VDD.n5428 92.5005
R5299 VDD.n5427 VDD.n5426 92.5005
R5300 VDD.n5419 VDD.n302 92.5005
R5301 VDD.n5421 VDD.n5420 92.5005
R5302 VDD.n5417 VDD.n5416 92.5005
R5303 VDD.n5415 VDD.n5414 92.5005
R5304 VDD.n5407 VDD.n306 92.5005
R5305 VDD.n5409 VDD.n5408 92.5005
R5306 VDD.n5405 VDD.n5404 92.5005
R5307 VDD.n5403 VDD.n5402 92.5005
R5308 VDD.n313 VDD.n310 92.5005
R5309 VDD.n315 VDD.n314 92.5005
R5310 VDD.n5397 VDD.n5396 92.5005
R5311 VDD.n5395 VDD.n5394 92.5005
R5312 VDD.n5387 VDD.n317 92.5005
R5313 VDD.n5389 VDD.n5388 92.5005
R5314 VDD.n5385 VDD.n5384 92.5005
R5315 VDD.n5383 VDD.n5382 92.5005
R5316 VDD.n5375 VDD.n320 92.5005
R5317 VDD.n5377 VDD.n5376 92.5005
R5318 VDD.n5373 VDD.n5372 92.5005
R5319 VDD.n5371 VDD.n5370 92.5005
R5320 VDD.n328 VDD.n324 92.5005
R5321 VDD.n5365 VDD.n5364 92.5005
R5322 VDD.n5364 VDD.n5363 92.5005
R5323 VDD.n332 VDD.n329 92.5005
R5324 VDD.n5362 VDD.n329 92.5005
R5325 VDD.n5360 VDD.n5359 92.5005
R5326 VDD.n5361 VDD.n5360 92.5005
R5327 VDD.n334 VDD.n331 92.5005
R5328 VDD.n331 VDD.n330 92.5005
R5329 VDD.n5354 VDD.n5353 92.5005
R5330 VDD.n5353 VDD.n5352 92.5005
R5331 VDD.n341 VDD.n338 92.5005
R5332 VDD.n5351 VDD.n338 92.5005
R5333 VDD.n5349 VDD.n5348 92.5005
R5334 VDD.n5350 VDD.n5349 92.5005
R5335 VDD.n342 VDD.n340 92.5005
R5336 VDD.n340 VDD.n339 92.5005
R5337 VDD.n5343 VDD.n5342 92.5005
R5338 VDD.n5342 VDD.n5341 92.5005
R5339 VDD.n348 VDD.n345 92.5005
R5340 VDD.n5340 VDD.n345 92.5005
R5341 VDD.n5338 VDD.n5337 92.5005
R5342 VDD.n5339 VDD.n5338 92.5005
R5343 VDD.n350 VDD.n347 92.5005
R5344 VDD.n347 VDD.n346 92.5005
R5345 VDD.n5332 VDD.n5331 92.5005
R5346 VDD.n5331 VDD.n5330 92.5005
R5347 VDD.n357 VDD.n354 92.5005
R5348 VDD.n5329 VDD.n354 92.5005
R5349 VDD.n5327 VDD.n5326 92.5005
R5350 VDD.n5328 VDD.n5327 92.5005
R5351 VDD.n359 VDD.n356 92.5005
R5352 VDD.n356 VDD.n355 92.5005
R5353 VDD.n5321 VDD.n5320 92.5005
R5354 VDD.n5320 VDD.n5319 92.5005
R5355 VDD.n366 VDD.n363 92.5005
R5356 VDD.n5318 VDD.n363 92.5005
R5357 VDD.n5316 VDD.n5315 92.5005
R5358 VDD.n5317 VDD.n5316 92.5005
R5359 VDD.n368 VDD.n365 92.5005
R5360 VDD.n365 VDD.n364 92.5005
R5361 VDD.n5310 VDD.n5309 92.5005
R5362 VDD.n5309 VDD.n5308 92.5005
R5363 VDD.n375 VDD.n372 92.5005
R5364 VDD.n5307 VDD.n372 92.5005
R5365 VDD.n5305 VDD.n5304 92.5005
R5366 VDD.n5306 VDD.n5305 92.5005
R5367 VDD.n377 VDD.n374 92.5005
R5368 VDD.n374 VDD.n373 92.5005
R5369 VDD.n382 VDD.n380 92.5005
R5370 VDD.n384 VDD.n382 92.5005
R5371 VDD.n5299 VDD.n5298 92.5005
R5372 VDD.n5298 VDD.n5297 92.5005
R5373 VDD.n387 VDD.n383 92.5005
R5374 VDD.n5296 VDD.n383 92.5005
R5375 VDD.n5294 VDD.n5293 92.5005
R5376 VDD.n5295 VDD.n5294 92.5005
R5377 VDD.n389 VDD.n386 92.5005
R5378 VDD.n386 VDD.n385 92.5005
R5379 VDD.n5288 VDD.n5287 92.5005
R5380 VDD.n5287 VDD.n5286 92.5005
R5381 VDD.n579 VDD.n397 92.5005
R5382 VDD.n452 VDD.n393 92.5005
R5383 VDD.n456 VDD.n455 92.5005
R5384 VDD.n459 VDD.n458 92.5005
R5385 VDD.n448 VDD.n447 92.5005
R5386 VDD.n465 VDD.n464 92.5005
R5387 VDD.n469 VDD.n468 92.5005
R5388 VDD.n467 VDD.n444 92.5005
R5389 VDD.n475 VDD.n474 92.5005
R5390 VDD.n478 VDD.n477 92.5005
R5391 VDD.n440 VDD.n439 92.5005
R5392 VDD.n485 VDD.n484 92.5005
R5393 VDD.n487 VDD.n438 92.5005
R5394 VDD.n490 VDD.n489 92.5005
R5395 VDD.n436 VDD.n435 92.5005
R5396 VDD.n496 VDD.n495 92.5005
R5397 VDD.n500 VDD.n499 92.5005
R5398 VDD.n498 VDD.n432 92.5005
R5399 VDD.n506 VDD.n505 92.5005
R5400 VDD.n509 VDD.n508 92.5005
R5401 VDD.n428 VDD.n427 92.5005
R5402 VDD.n515 VDD.n514 92.5005
R5403 VDD.n519 VDD.n518 92.5005
R5404 VDD.n517 VDD.n424 92.5005
R5405 VDD.n525 VDD.n524 92.5005
R5406 VDD.n528 VDD.n527 92.5005
R5407 VDD.n420 VDD.n419 92.5005
R5408 VDD.n534 VDD.n533 92.5005
R5409 VDD.n539 VDD.n538 92.5005
R5410 VDD.n537 VDD.n416 92.5005
R5411 VDD.n544 VDD.n415 92.5005
R5412 VDD.n546 VDD.n545 92.5005
R5413 VDD.n550 VDD.n549 92.5005
R5414 VDD.n548 VDD.n412 92.5005
R5415 VDD.n556 VDD.n555 92.5005
R5416 VDD.n559 VDD.n558 92.5005
R5417 VDD.n408 VDD.n407 92.5005
R5418 VDD.n565 VDD.n564 92.5005
R5419 VDD.n569 VDD.n568 92.5005
R5420 VDD.n567 VDD.n404 92.5005
R5421 VDD.n575 VDD.n574 92.5005
R5422 VDD.n578 VDD.n577 92.5005
R5423 VDD.n5283 VDD.n5282 92.5005
R5424 VDD.n5284 VDD.n5283 92.5005
R5425 VDD.n400 VDD.n398 92.5005
R5426 VDD.n398 VDD.n396 92.5005
R5427 VDD.n5277 VDD.n5276 92.5005
R5428 VDD.n5276 VDD.n5275 92.5005
R5429 VDD.n588 VDD.n585 92.5005
R5430 VDD.n5274 VDD.n585 92.5005
R5431 VDD.n5272 VDD.n5271 92.5005
R5432 VDD.n5273 VDD.n5272 92.5005
R5433 VDD.n590 VDD.n587 92.5005
R5434 VDD.n587 VDD.n586 92.5005
R5435 VDD.n595 VDD.n593 92.5005
R5436 VDD.n597 VDD.n595 92.5005
R5437 VDD.n5266 VDD.n5265 92.5005
R5438 VDD.n5265 VDD.n5264 92.5005
R5439 VDD.n600 VDD.n596 92.5005
R5440 VDD.n5263 VDD.n596 92.5005
R5441 VDD.n5261 VDD.n5260 92.5005
R5442 VDD.n5262 VDD.n5261 92.5005
R5443 VDD.n602 VDD.n599 92.5005
R5444 VDD.n599 VDD.n598 92.5005
R5445 VDD.n5255 VDD.n5254 92.5005
R5446 VDD.n5254 VDD.n5253 92.5005
R5447 VDD.n609 VDD.n606 92.5005
R5448 VDD.n5252 VDD.n606 92.5005
R5449 VDD.n5250 VDD.n5249 92.5005
R5450 VDD.n5251 VDD.n5250 92.5005
R5451 VDD.n611 VDD.n608 92.5005
R5452 VDD.n608 VDD.n607 92.5005
R5453 VDD.n5244 VDD.n5243 92.5005
R5454 VDD.n5243 VDD.n5242 92.5005
R5455 VDD.n618 VDD.n615 92.5005
R5456 VDD.n5241 VDD.n615 92.5005
R5457 VDD.n5239 VDD.n5238 92.5005
R5458 VDD.n5240 VDD.n5239 92.5005
R5459 VDD.n620 VDD.n617 92.5005
R5460 VDD.n617 VDD.n616 92.5005
R5461 VDD.n5233 VDD.n5232 92.5005
R5462 VDD.n5232 VDD.n5231 92.5005
R5463 VDD.n627 VDD.n624 92.5005
R5464 VDD.n5230 VDD.n624 92.5005
R5465 VDD.n5228 VDD.n5227 92.5005
R5466 VDD.n5229 VDD.n5228 92.5005
R5467 VDD.n629 VDD.n626 92.5005
R5468 VDD.n626 VDD.n625 92.5005
R5469 VDD.n5222 VDD.n5221 92.5005
R5470 VDD.n5221 VDD.n5220 92.5005
R5471 VDD.n633 VDD.n632 92.5005
R5472 VDD.n5219 VDD.n633 92.5005
R5473 VDD.n5217 VDD.n5216 92.5005
R5474 VDD.n5218 VDD.n5217 92.5005
R5475 VDD.n637 VDD.n635 92.5005
R5476 VDD.n635 VDD.n634 92.5005
R5477 VDD.n5211 VDD.n5210 92.5005
R5478 VDD.n5210 VDD.n5209 92.5005
R5479 VDD.n643 VDD.n640 92.5005
R5480 VDD.n5208 VDD.n640 92.5005
R5481 VDD.n5206 VDD.n5205 92.5005
R5482 VDD.n5207 VDD.n5206 92.5005
R5483 VDD.n645 VDD.n642 92.5005
R5484 VDD.n642 VDD.n641 92.5005
R5485 VDD.n5200 VDD.n5199 92.5005
R5486 VDD.n5199 VDD.n5198 92.5005
R5487 VDD.n652 VDD.n649 92.5005
R5488 VDD.n5197 VDD.n649 92.5005
R5489 VDD.n5195 VDD.n5194 92.5005
R5490 VDD.n5196 VDD.n5195 92.5005
R5491 VDD.n654 VDD.n651 92.5005
R5492 VDD.n651 VDD.n650 92.5005
R5493 VDD.n5189 VDD.n5188 92.5005
R5494 VDD.n5188 VDD.n5187 92.5005
R5495 VDD.n661 VDD.n658 92.5005
R5496 VDD.n5186 VDD.n658 92.5005
R5497 VDD.n5184 VDD.n5183 92.5005
R5498 VDD.n5185 VDD.n5184 92.5005
R5499 VDD.n663 VDD.n660 92.5005
R5500 VDD.n660 VDD.n659 92.5005
R5501 VDD.n5178 VDD.n5177 92.5005
R5502 VDD.n5177 VDD.n5176 92.5005
R5503 VDD.n670 VDD.n667 92.5005
R5504 VDD.n5175 VDD.n667 92.5005
R5505 VDD.n5173 VDD.n5172 92.5005
R5506 VDD.n5174 VDD.n5173 92.5005
R5507 VDD.n5171 VDD.n669 92.5005
R5508 VDD.n669 VDD.n668 92.5005
R5509 VDD.n676 VDD.n672 92.5005
R5510 VDD.n678 VDD.n676 92.5005
R5511 VDD.n5166 VDD.n5165 92.5005
R5512 VDD.n5165 VDD.n5164 92.5005
R5513 VDD.n4721 VDD.n4720 92.5005
R5514 VDD.n924 VDD.n918 92.5005
R5515 VDD.n4710 VDD.n926 92.5005
R5516 VDD.n5162 VDD.n677 92.5005
R5517 VDD.n5162 VDD.n5161 92.5005
R5518 VDD.n5158 VDD.n680 92.5005
R5519 VDD.n680 VDD.n679 92.5005
R5520 VDD.n685 VDD.n681 92.5005
R5521 VDD.n5150 VDD.n685 92.5005
R5522 VDD.n5153 VDD.n5152 92.5005
R5523 VDD.n5152 VDD.n5151 92.5005
R5524 VDD.n684 VDD.n683 92.5005
R5525 VDD.n5149 VDD.n684 92.5005
R5526 VDD.n5147 VDD.n5146 92.5005
R5527 VDD.n5148 VDD.n5147 92.5005
R5528 VDD.n688 VDD.n687 92.5005
R5529 VDD.n687 VDD.n686 92.5005
R5530 VDD.n5140 VDD.n5139 92.5005
R5531 VDD.n5139 VDD.n5138 92.5005
R5532 VDD.n695 VDD.n691 92.5005
R5533 VDD.n5137 VDD.n691 92.5005
R5534 VDD.n5135 VDD.n5134 92.5005
R5535 VDD.n5136 VDD.n5135 92.5005
R5536 VDD.n5128 VDD.n693 92.5005
R5537 VDD.n693 VDD.n692 92.5005
R5538 VDD.n5127 VDD.n5126 92.5005
R5539 VDD.n5126 VDD.n5125 92.5005
R5540 VDD.n702 VDD.n698 92.5005
R5541 VDD.n5124 VDD.n698 92.5005
R5542 VDD.n5122 VDD.n5121 92.5005
R5543 VDD.n5123 VDD.n5122 92.5005
R5544 VDD.n5115 VDD.n700 92.5005
R5545 VDD.n700 VDD.n699 92.5005
R5546 VDD.n5114 VDD.n5113 92.5005
R5547 VDD.n5113 VDD.n5112 92.5005
R5548 VDD.n709 VDD.n705 92.5005
R5549 VDD.n5111 VDD.n705 92.5005
R5550 VDD.n5109 VDD.n5108 92.5005
R5551 VDD.n5110 VDD.n5109 92.5005
R5552 VDD.n5102 VDD.n707 92.5005
R5553 VDD.n707 VDD.n706 92.5005
R5554 VDD.n5101 VDD.n5100 92.5005
R5555 VDD.n5100 VDD.n5099 92.5005
R5556 VDD.n716 VDD.n712 92.5005
R5557 VDD.n5098 VDD.n712 92.5005
R5558 VDD.n5096 VDD.n5095 92.5005
R5559 VDD.n5097 VDD.n5096 92.5005
R5560 VDD.n715 VDD.n714 92.5005
R5561 VDD.n714 VDD.n713 92.5005
R5562 VDD.n5090 VDD.n5089 92.5005
R5563 VDD.n5089 VDD.n5088 92.5005
R5564 VDD.n723 VDD.n719 92.5005
R5565 VDD.n5087 VDD.n719 92.5005
R5566 VDD.n5085 VDD.n5084 92.5005
R5567 VDD.n5086 VDD.n5085 92.5005
R5568 VDD.n5078 VDD.n721 92.5005
R5569 VDD.n721 VDD.n720 92.5005
R5570 VDD.n5077 VDD.n5076 92.5005
R5571 VDD.n5076 VDD.n5075 92.5005
R5572 VDD.n730 VDD.n726 92.5005
R5573 VDD.n5074 VDD.n726 92.5005
R5574 VDD.n5072 VDD.n5071 92.5005
R5575 VDD.n5073 VDD.n5072 92.5005
R5576 VDD.n5065 VDD.n728 92.5005
R5577 VDD.n728 VDD.n727 92.5005
R5578 VDD.n5064 VDD.n5063 92.5005
R5579 VDD.n5063 VDD.n5062 92.5005
R5580 VDD.n737 VDD.n733 92.5005
R5581 VDD.n5061 VDD.n733 92.5005
R5582 VDD.n5059 VDD.n5058 92.5005
R5583 VDD.n5060 VDD.n5059 92.5005
R5584 VDD.n5052 VDD.n735 92.5005
R5585 VDD.n735 VDD.n734 92.5005
R5586 VDD.n5051 VDD.n5050 92.5005
R5587 VDD.n5050 VDD.n5049 92.5005
R5588 VDD.n744 VDD.n740 92.5005
R5589 VDD.n5048 VDD.n740 92.5005
R5590 VDD.n5046 VDD.n5045 92.5005
R5591 VDD.n5047 VDD.n5046 92.5005
R5592 VDD.n5039 VDD.n742 92.5005
R5593 VDD.n742 VDD.n741 92.5005
R5594 VDD.n5038 VDD.n5037 92.5005
R5595 VDD.n5037 VDD.n5036 92.5005
R5596 VDD.n747 VDD.n746 92.5005
R5597 VDD.n5035 VDD.n747 92.5005
R5598 VDD.n5033 VDD.n5032 92.5005
R5599 VDD.n5034 VDD.n5033 92.5005
R5600 VDD.n750 VDD.n749 92.5005
R5601 VDD.n749 VDD.n748 92.5005
R5602 VDD.n5026 VDD.n5025 92.5005
R5603 VDD.n5025 VDD.n5024 92.5005
R5604 VDD.n757 VDD.n753 92.5005
R5605 VDD.n5023 VDD.n753 92.5005
R5606 VDD.n5021 VDD.n5020 92.5005
R5607 VDD.n5022 VDD.n5021 92.5005
R5608 VDD.n5014 VDD.n755 92.5005
R5609 VDD.n755 VDD.n754 92.5005
R5610 VDD.n5013 VDD.n5012 92.5005
R5611 VDD.n5012 VDD.n5011 92.5005
R5612 VDD.n764 VDD.n760 92.5005
R5613 VDD.n5010 VDD.n760 92.5005
R5614 VDD.n5008 VDD.n5007 92.5005
R5615 VDD.n5009 VDD.n5008 92.5005
R5616 VDD.n5001 VDD.n762 92.5005
R5617 VDD.n762 VDD.n761 92.5005
R5618 VDD.n5000 VDD.n4999 92.5005
R5619 VDD.n4999 VDD.n4998 92.5005
R5620 VDD.n771 VDD.n767 92.5005
R5621 VDD.n4997 VDD.n767 92.5005
R5622 VDD.n4995 VDD.n4994 92.5005
R5623 VDD.n4996 VDD.n4995 92.5005
R5624 VDD.n4988 VDD.n769 92.5005
R5625 VDD.n769 VDD.n768 92.5005
R5626 VDD.n4987 VDD.n4986 92.5005
R5627 VDD.n4986 VDD.n4985 92.5005
R5628 VDD.n778 VDD.n774 92.5005
R5629 VDD.n4984 VDD.n774 92.5005
R5630 VDD.n4982 VDD.n4981 92.5005
R5631 VDD.n4983 VDD.n4982 92.5005
R5632 VDD.n777 VDD.n776 92.5005
R5633 VDD.n776 VDD.n775 92.5005
R5634 VDD.n4976 VDD.n4975 92.5005
R5635 VDD.n4975 VDD.n4974 92.5005
R5636 VDD.n785 VDD.n781 92.5005
R5637 VDD.n4973 VDD.n781 92.5005
R5638 VDD.n4971 VDD.n4970 92.5005
R5639 VDD.n4972 VDD.n4971 92.5005
R5640 VDD.n4964 VDD.n783 92.5005
R5641 VDD.n783 VDD.n782 92.5005
R5642 VDD.n4963 VDD.n4962 92.5005
R5643 VDD.n4962 VDD.n4961 92.5005
R5644 VDD.n792 VDD.n788 92.5005
R5645 VDD.n4960 VDD.n788 92.5005
R5646 VDD.n4958 VDD.n4957 92.5005
R5647 VDD.n4959 VDD.n4958 92.5005
R5648 VDD.n4951 VDD.n790 92.5005
R5649 VDD.n790 VDD.n789 92.5005
R5650 VDD.n4950 VDD.n4949 92.5005
R5651 VDD.n4949 VDD.n4948 92.5005
R5652 VDD.n799 VDD.n795 92.5005
R5653 VDD.n4947 VDD.n795 92.5005
R5654 VDD.n4945 VDD.n4944 92.5005
R5655 VDD.n4946 VDD.n4945 92.5005
R5656 VDD.n4938 VDD.n797 92.5005
R5657 VDD.n797 VDD.n796 92.5005
R5658 VDD.n4937 VDD.n4936 92.5005
R5659 VDD.n4936 VDD.n4935 92.5005
R5660 VDD.n806 VDD.n802 92.5005
R5661 VDD.n4934 VDD.n802 92.5005
R5662 VDD.n4932 VDD.n4931 92.5005
R5663 VDD.n4933 VDD.n4932 92.5005
R5664 VDD.n4925 VDD.n804 92.5005
R5665 VDD.n804 VDD.n803 92.5005
R5666 VDD.n4924 VDD.n4923 92.5005
R5667 VDD.n4923 VDD.n4922 92.5005
R5668 VDD.n809 VDD.n808 92.5005
R5669 VDD.n4921 VDD.n809 92.5005
R5670 VDD.n4919 VDD.n4918 92.5005
R5671 VDD.n4920 VDD.n4919 92.5005
R5672 VDD.n812 VDD.n811 92.5005
R5673 VDD.n811 VDD.n810 92.5005
R5674 VDD.n4912 VDD.n4911 92.5005
R5675 VDD.n4911 VDD.n4910 92.5005
R5676 VDD.n819 VDD.n815 92.5005
R5677 VDD.n4909 VDD.n815 92.5005
R5678 VDD.n4907 VDD.n4906 92.5005
R5679 VDD.n4908 VDD.n4907 92.5005
R5680 VDD.n4900 VDD.n817 92.5005
R5681 VDD.n817 VDD.n816 92.5005
R5682 VDD.n4899 VDD.n4898 92.5005
R5683 VDD.n4898 VDD.n4897 92.5005
R5684 VDD.n826 VDD.n822 92.5005
R5685 VDD.n4896 VDD.n822 92.5005
R5686 VDD.n4894 VDD.n4893 92.5005
R5687 VDD.n4895 VDD.n4894 92.5005
R5688 VDD.n4887 VDD.n824 92.5005
R5689 VDD.n824 VDD.n823 92.5005
R5690 VDD.n4886 VDD.n4885 92.5005
R5691 VDD.n4885 VDD.n4884 92.5005
R5692 VDD.n833 VDD.n829 92.5005
R5693 VDD.n4883 VDD.n829 92.5005
R5694 VDD.n4881 VDD.n4880 92.5005
R5695 VDD.n4882 VDD.n4881 92.5005
R5696 VDD.n4874 VDD.n831 92.5005
R5697 VDD.n831 VDD.n830 92.5005
R5698 VDD.n4873 VDD.n4872 92.5005
R5699 VDD.n4872 VDD.n4871 92.5005
R5700 VDD.n840 VDD.n836 92.5005
R5701 VDD.n4870 VDD.n836 92.5005
R5702 VDD.n4868 VDD.n4867 92.5005
R5703 VDD.n4869 VDD.n4868 92.5005
R5704 VDD.n839 VDD.n838 92.5005
R5705 VDD.n838 VDD.n837 92.5005
R5706 VDD.n4862 VDD.n4861 92.5005
R5707 VDD.n4861 VDD.n4860 92.5005
R5708 VDD.n847 VDD.n843 92.5005
R5709 VDD.n4859 VDD.n843 92.5005
R5710 VDD.n4857 VDD.n4856 92.5005
R5711 VDD.n4858 VDD.n4857 92.5005
R5712 VDD.n4850 VDD.n845 92.5005
R5713 VDD.n845 VDD.n844 92.5005
R5714 VDD.n4849 VDD.n4848 92.5005
R5715 VDD.n4848 VDD.n4847 92.5005
R5716 VDD.n854 VDD.n850 92.5005
R5717 VDD.n4846 VDD.n850 92.5005
R5718 VDD.n4844 VDD.n4843 92.5005
R5719 VDD.n4845 VDD.n4844 92.5005
R5720 VDD.n4837 VDD.n852 92.5005
R5721 VDD.n852 VDD.n851 92.5005
R5722 VDD.n4836 VDD.n4835 92.5005
R5723 VDD.n4835 VDD.n4834 92.5005
R5724 VDD.n861 VDD.n857 92.5005
R5725 VDD.n4833 VDD.n857 92.5005
R5726 VDD.n4831 VDD.n4830 92.5005
R5727 VDD.n4832 VDD.n4831 92.5005
R5728 VDD.n4824 VDD.n859 92.5005
R5729 VDD.n859 VDD.n858 92.5005
R5730 VDD.n4823 VDD.n4822 92.5005
R5731 VDD.n4822 VDD.n4821 92.5005
R5732 VDD.n868 VDD.n864 92.5005
R5733 VDD.n4820 VDD.n864 92.5005
R5734 VDD.n4818 VDD.n4817 92.5005
R5735 VDD.n4819 VDD.n4818 92.5005
R5736 VDD.n4811 VDD.n866 92.5005
R5737 VDD.n866 VDD.n865 92.5005
R5738 VDD.n4810 VDD.n4809 92.5005
R5739 VDD.n4809 VDD.n4808 92.5005
R5740 VDD.n871 VDD.n870 92.5005
R5741 VDD.n4807 VDD.n871 92.5005
R5742 VDD.n4805 VDD.n4804 92.5005
R5743 VDD.n4806 VDD.n4805 92.5005
R5744 VDD.n874 VDD.n873 92.5005
R5745 VDD.n873 VDD.n872 92.5005
R5746 VDD.n4798 VDD.n4797 92.5005
R5747 VDD.n4797 VDD.n4796 92.5005
R5748 VDD.n881 VDD.n877 92.5005
R5749 VDD.n4795 VDD.n877 92.5005
R5750 VDD.n4793 VDD.n4792 92.5005
R5751 VDD.n4794 VDD.n4793 92.5005
R5752 VDD.n4786 VDD.n879 92.5005
R5753 VDD.n879 VDD.n878 92.5005
R5754 VDD.n4785 VDD.n4784 92.5005
R5755 VDD.n4784 VDD.n4783 92.5005
R5756 VDD.n888 VDD.n884 92.5005
R5757 VDD.n4782 VDD.n884 92.5005
R5758 VDD.n4780 VDD.n4779 92.5005
R5759 VDD.n4781 VDD.n4780 92.5005
R5760 VDD.n4773 VDD.n886 92.5005
R5761 VDD.n886 VDD.n885 92.5005
R5762 VDD.n4772 VDD.n4771 92.5005
R5763 VDD.n4771 VDD.n4770 92.5005
R5764 VDD.n895 VDD.n891 92.5005
R5765 VDD.n4769 VDD.n891 92.5005
R5766 VDD.n4767 VDD.n4766 92.5005
R5767 VDD.n4768 VDD.n4767 92.5005
R5768 VDD.n4760 VDD.n893 92.5005
R5769 VDD.n893 VDD.n892 92.5005
R5770 VDD.n4759 VDD.n4758 92.5005
R5771 VDD.n4758 VDD.n4757 92.5005
R5772 VDD.n902 VDD.n898 92.5005
R5773 VDD.n4756 VDD.n898 92.5005
R5774 VDD.n4754 VDD.n4753 92.5005
R5775 VDD.n4755 VDD.n4754 92.5005
R5776 VDD.n901 VDD.n900 92.5005
R5777 VDD.n900 VDD.n899 92.5005
R5778 VDD.n4748 VDD.n4747 92.5005
R5779 VDD.n4747 VDD.n4746 92.5005
R5780 VDD.n909 VDD.n905 92.5005
R5781 VDD.n4745 VDD.n905 92.5005
R5782 VDD.n4743 VDD.n4742 92.5005
R5783 VDD.n4744 VDD.n4743 92.5005
R5784 VDD.n4736 VDD.n907 92.5005
R5785 VDD.n907 VDD.n906 92.5005
R5786 VDD.n4735 VDD.n4734 92.5005
R5787 VDD.n4734 VDD.n4733 92.5005
R5788 VDD.n916 VDD.n912 92.5005
R5789 VDD.n4732 VDD.n912 92.5005
R5790 VDD.n4730 VDD.n4729 92.5005
R5791 VDD.n4731 VDD.n4730 92.5005
R5792 VDD.n4723 VDD.n914 92.5005
R5793 VDD.n914 VDD.n913 92.5005
R5794 VDD.n4717 VDD.n4716 92.5005
R5795 VDD.n4719 VDD.n4718 92.5005
R5796 VDD.n4713 VDD.n4712 92.5005
R5797 VDD.n4714 VDD.n4713 92.5005
R5798 VDD.n927 VDD.n923 92.5005
R5799 VDD.n923 VDD.n922 92.5005
R5800 VDD.n4705 VDD.n4704 92.5005
R5801 VDD.n4704 VDD.n4703 92.5005
R5802 VDD.n934 VDD.n930 92.5005
R5803 VDD.n4702 VDD.n930 92.5005
R5804 VDD.n4700 VDD.n4699 92.5005
R5805 VDD.n4701 VDD.n4700 92.5005
R5806 VDD.n4693 VDD.n932 92.5005
R5807 VDD.n932 VDD.n931 92.5005
R5808 VDD.n4692 VDD.n4691 92.5005
R5809 VDD.n4691 VDD.n4690 92.5005
R5810 VDD.n941 VDD.n937 92.5005
R5811 VDD.n4689 VDD.n937 92.5005
R5812 VDD.n4687 VDD.n4686 92.5005
R5813 VDD.n4688 VDD.n4687 92.5005
R5814 VDD.n4680 VDD.n939 92.5005
R5815 VDD.n939 VDD.n938 92.5005
R5816 VDD.n4679 VDD.n4678 92.5005
R5817 VDD.n4678 VDD.n4677 92.5005
R5818 VDD.n948 VDD.n944 92.5005
R5819 VDD.n4676 VDD.n944 92.5005
R5820 VDD.n4674 VDD.n4673 92.5005
R5821 VDD.n4675 VDD.n4674 92.5005
R5822 VDD.n4667 VDD.n946 92.5005
R5823 VDD.n946 VDD.n945 92.5005
R5824 VDD.n4666 VDD.n4665 92.5005
R5825 VDD.n4665 VDD.n4664 92.5005
R5826 VDD.n955 VDD.n951 92.5005
R5827 VDD.n4663 VDD.n951 92.5005
R5828 VDD.n4661 VDD.n4660 92.5005
R5829 VDD.n4662 VDD.n4661 92.5005
R5830 VDD.n954 VDD.n953 92.5005
R5831 VDD.n953 VDD.n952 92.5005
R5832 VDD.n4656 VDD.n4655 92.5005
R5833 VDD.n4655 VDD.n4654 92.5005
R5834 VDD.n962 VDD.n958 92.5005
R5835 VDD.n4653 VDD.n958 92.5005
R5836 VDD.n4651 VDD.n4650 92.5005
R5837 VDD.n4652 VDD.n4651 92.5005
R5838 VDD.n4644 VDD.n960 92.5005
R5839 VDD.n960 VDD.n959 92.5005
R5840 VDD.n4643 VDD.n4642 92.5005
R5841 VDD.n4642 VDD.n4641 92.5005
R5842 VDD.n969 VDD.n965 92.5005
R5843 VDD.n4640 VDD.n965 92.5005
R5844 VDD.n4638 VDD.n4637 92.5005
R5845 VDD.n4639 VDD.n4638 92.5005
R5846 VDD.n4631 VDD.n967 92.5005
R5847 VDD.n967 VDD.n966 92.5005
R5848 VDD.n4630 VDD.n4629 92.5005
R5849 VDD.n4629 VDD.n4628 92.5005
R5850 VDD.n976 VDD.n972 92.5005
R5851 VDD.n4627 VDD.n972 92.5005
R5852 VDD.n4625 VDD.n4624 92.5005
R5853 VDD.n4626 VDD.n4625 92.5005
R5854 VDD.n4618 VDD.n974 92.5005
R5855 VDD.n974 VDD.n973 92.5005
R5856 VDD.n4617 VDD.n4616 92.5005
R5857 VDD.n4616 VDD.n4615 92.5005
R5858 VDD.n983 VDD.n979 92.5005
R5859 VDD.n4614 VDD.n979 92.5005
R5860 VDD.n4612 VDD.n4611 92.5005
R5861 VDD.n4613 VDD.n4612 92.5005
R5862 VDD.n986 VDD.n981 92.5005
R5863 VDD.n981 VDD.n980 92.5005
R5864 VDD.n4606 VDD.n4605 92.5005
R5865 VDD.n4605 VDD.n4604 92.5005
R5866 VDD.n987 VDD.n985 92.5005
R5867 VDD.n4603 VDD.n987 92.5005
R5868 VDD.n4601 VDD.n4600 92.5005
R5869 VDD.n4602 VDD.n4601 92.5005
R5870 VDD.n990 VDD.n989 92.5005
R5871 VDD.n989 VDD.n988 92.5005
R5872 VDD.n4594 VDD.n4593 92.5005
R5873 VDD.n4593 VDD.n4592 92.5005
R5874 VDD.n997 VDD.n993 92.5005
R5875 VDD.n4591 VDD.n993 92.5005
R5876 VDD.n4589 VDD.n4588 92.5005
R5877 VDD.n4590 VDD.n4589 92.5005
R5878 VDD.n4582 VDD.n995 92.5005
R5879 VDD.n995 VDD.n994 92.5005
R5880 VDD.n4581 VDD.n4580 92.5005
R5881 VDD.n4580 VDD.n4579 92.5005
R5882 VDD.n1161 VDD.n1000 92.5005
R5883 VDD.n4578 VDD.n1000 92.5005
R5884 VDD.n2291 VDD.n2290 92.5005
R5885 VDD.n2293 VDD.n2292 92.5005
R5886 VDD.n2295 VDD.n2294 92.5005
R5887 VDD.n2297 VDD.n2296 92.5005
R5888 VDD.n2299 VDD.n2298 92.5005
R5889 VDD.n2301 VDD.n2300 92.5005
R5890 VDD.n2303 VDD.n2302 92.5005
R5891 VDD.n2305 VDD.n2304 92.5005
R5892 VDD.n2307 VDD.n2306 92.5005
R5893 VDD.n2309 VDD.n2308 92.5005
R5894 VDD.n2311 VDD.n2310 92.5005
R5895 VDD.n2313 VDD.n2312 92.5005
R5896 VDD.n2315 VDD.n2314 92.5005
R5897 VDD.n2317 VDD.n2316 92.5005
R5898 VDD.n2319 VDD.n2318 92.5005
R5899 VDD.n2321 VDD.n2320 92.5005
R5900 VDD.n2323 VDD.n2322 92.5005
R5901 VDD.n2325 VDD.n2324 92.5005
R5902 VDD.n2327 VDD.n2326 92.5005
R5903 VDD.n2329 VDD.n2328 92.5005
R5904 VDD.n2331 VDD.n2330 92.5005
R5905 VDD.n2333 VDD.n2332 92.5005
R5906 VDD.n2335 VDD.n2334 92.5005
R5907 VDD.n2337 VDD.n2336 92.5005
R5908 VDD.n2339 VDD.n2338 92.5005
R5909 VDD.n4304 VDD.n4303 92.5005
R5910 VDD.n4306 VDD.n4305 92.5005
R5911 VDD.n4308 VDD.n4307 92.5005
R5912 VDD.n4310 VDD.n4309 92.5005
R5913 VDD.n4312 VDD.n4311 92.5005
R5914 VDD.n4314 VDD.n4313 92.5005
R5915 VDD.n4316 VDD.n4315 92.5005
R5916 VDD.n4318 VDD.n4317 92.5005
R5917 VDD.n4320 VDD.n4319 92.5005
R5918 VDD.n4322 VDD.n4321 92.5005
R5919 VDD.n4324 VDD.n4323 92.5005
R5920 VDD.n4326 VDD.n4325 92.5005
R5921 VDD.n4328 VDD.n4327 92.5005
R5922 VDD.n4331 VDD.n4330 92.5005
R5923 VDD.n4333 VDD.n4332 92.5005
R5924 VDD.n4335 VDD.n4334 92.5005
R5925 VDD.n4337 VDD.n4336 92.5005
R5926 VDD.n4339 VDD.n4338 92.5005
R5927 VDD.n4341 VDD.n4340 92.5005
R5928 VDD.n4343 VDD.n4342 92.5005
R5929 VDD.n4345 VDD.n4344 92.5005
R5930 VDD.n4347 VDD.n4346 92.5005
R5931 VDD.n4349 VDD.n4348 92.5005
R5932 VDD.n4351 VDD.n4350 92.5005
R5933 VDD.n4352 VDD.n2286 92.5005
R5934 VDD.n4354 VDD.n4353 92.5005
R5935 VDD.n2289 VDD.n2236 92.5005
R5936 VDD.n4356 VDD.n2236 92.5005
R5937 VDD.n2214 VDD.n2213 92.5005
R5938 VDD.n2234 VDD.n2214 92.5005
R5939 VDD.n4368 VDD.n4367 92.5005
R5940 VDD.n4367 VDD.n4366 92.5005
R5941 VDD.n4369 VDD.n2208 92.5005
R5942 VDD.n2215 VDD.n2208 92.5005
R5943 VDD.n4371 VDD.n4370 92.5005
R5944 VDD.n4372 VDD.n4371 92.5005
R5945 VDD.n2212 VDD.n2202 92.5005
R5946 VDD.n4375 VDD.n2202 92.5005
R5947 VDD.n2211 VDD.n2210 92.5005
R5948 VDD.n2210 VDD.n2200 92.5005
R5949 VDD.n2209 VDD.n2185 92.5005
R5950 VDD.n4384 VDD.n2185 92.5005
R5951 VDD.n2172 VDD.n2171 92.5005
R5952 VDD.n2183 VDD.n2172 92.5005
R5953 VDD.n4393 VDD.n4392 92.5005
R5954 VDD.n4392 VDD.n4391 92.5005
R5955 VDD.n4394 VDD.n2169 92.5005
R5956 VDD.n2173 VDD.n2169 92.5005
R5957 VDD.n4396 VDD.n4395 92.5005
R5958 VDD.n4397 VDD.n4396 92.5005
R5959 VDD.n2170 VDD.n2163 92.5005
R5960 VDD.n4400 VDD.n2163 92.5005
R5961 VDD.n2141 VDD.n2140 92.5005
R5962 VDD.n2161 VDD.n2141 92.5005
R5963 VDD.n4412 VDD.n4411 92.5005
R5964 VDD.n4411 VDD.n4410 92.5005
R5965 VDD.n4413 VDD.n2138 92.5005
R5966 VDD.n2142 VDD.n2138 92.5005
R5967 VDD.n4415 VDD.n4414 92.5005
R5968 VDD.n4416 VDD.n4415 92.5005
R5969 VDD.n2139 VDD.n2131 92.5005
R5970 VDD.n4419 VDD.n2131 92.5005
R5971 VDD.n2110 VDD.n2109 92.5005
R5972 VDD.n2130 VDD.n2110 92.5005
R5973 VDD.n4431 VDD.n4430 92.5005
R5974 VDD.n4430 VDD.n4429 92.5005
R5975 VDD.n4432 VDD.n2107 92.5005
R5976 VDD.n2111 VDD.n2107 92.5005
R5977 VDD.n4434 VDD.n4433 92.5005
R5978 VDD.n4435 VDD.n4434 92.5005
R5979 VDD.n2108 VDD.n2101 92.5005
R5980 VDD.n4438 VDD.n2101 92.5005
R5981 VDD.n2073 VDD.n2072 92.5005
R5982 VDD.n2099 VDD.n2073 92.5005
R5983 VDD.n4450 VDD.n4449 92.5005
R5984 VDD.n4449 VDD.n4448 92.5005
R5985 VDD.n4451 VDD.n2071 92.5005
R5986 VDD.n2074 VDD.n2071 92.5005
R5987 VDD.n4453 VDD.n4452 92.5005
R5988 VDD.n4454 VDD.n4453 92.5005
R5989 VDD.n2056 VDD.n2055 92.5005
R5990 VDD.n2068 VDD.n2056 92.5005
R5991 VDD.n4465 VDD.n4464 92.5005
R5992 VDD.n4464 VDD.n4463 92.5005
R5993 VDD.n4466 VDD.n2053 92.5005
R5994 VDD.n2089 VDD.n2053 92.5005
R5995 VDD.n4468 VDD.n4467 92.5005
R5996 VDD.n4469 VDD.n4468 92.5005
R5997 VDD.n2054 VDD.n2048 92.5005
R5998 VDD.n4472 VDD.n2048 92.5005
R5999 VDD.n2026 VDD.n2025 92.5005
R6000 VDD.n2046 VDD.n2026 92.5005
R6001 VDD.n4484 VDD.n4483 92.5005
R6002 VDD.n4483 VDD.n4482 92.5005
R6003 VDD.n4485 VDD.n2023 92.5005
R6004 VDD.n2027 VDD.n2023 92.5005
R6005 VDD.n4487 VDD.n4486 92.5005
R6006 VDD.n4488 VDD.n4487 92.5005
R6007 VDD.n2024 VDD.n2016 92.5005
R6008 VDD.n4491 VDD.n2016 92.5005
R6009 VDD.n1993 VDD.n1992 92.5005
R6010 VDD.n2013 VDD.n1993 92.5005
R6011 VDD.n4503 VDD.n4502 92.5005
R6012 VDD.n4502 VDD.n4501 92.5005
R6013 VDD.n4504 VDD.n1987 92.5005
R6014 VDD.n1994 VDD.n1987 92.5005
R6015 VDD.n4506 VDD.n4505 92.5005
R6016 VDD.n4507 VDD.n4506 92.5005
R6017 VDD.n1991 VDD.n1981 92.5005
R6018 VDD.n4510 VDD.n1981 92.5005
R6019 VDD.n1990 VDD.n1989 92.5005
R6020 VDD.n1989 VDD.n1979 92.5005
R6021 VDD.n1988 VDD.n1964 92.5005
R6022 VDD.n4519 VDD.n1964 92.5005
R6023 VDD.n1952 VDD.n1951 92.5005
R6024 VDD.n1962 VDD.n1952 92.5005
R6025 VDD.n4528 VDD.n4527 92.5005
R6026 VDD.n4527 VDD.n4526 92.5005
R6027 VDD.n4529 VDD.n1949 92.5005
R6028 VDD.n2607 VDD.n1949 92.5005
R6029 VDD.n4531 VDD.n4530 92.5005
R6030 VDD.n4532 VDD.n4531 92.5005
R6031 VDD.n1950 VDD.n1943 92.5005
R6032 VDD.n4535 VDD.n1943 92.5005
R6033 VDD.n1921 VDD.n1920 92.5005
R6034 VDD.n1941 VDD.n1921 92.5005
R6035 VDD.n4547 VDD.n4546 92.5005
R6036 VDD.n4546 VDD.n4545 92.5005
R6037 VDD.n4548 VDD.n1918 92.5005
R6038 VDD.n1922 VDD.n1918 92.5005
R6039 VDD.n4550 VDD.n4549 92.5005
R6040 VDD.n4551 VDD.n4550 92.5005
R6041 VDD.n1919 VDD.n1912 92.5005
R6042 VDD.n4554 VDD.n1912 92.5005
R6043 VDD.n1017 VDD.n1016 92.5005
R6044 VDD.n1910 VDD.n1017 92.5005
R6045 VDD.n4566 VDD.n4565 92.5005
R6046 VDD.n4565 VDD.n4564 92.5005
R6047 VDD.n4567 VDD.n1014 92.5005
R6048 VDD.n2602 VDD.n1014 92.5005
R6049 VDD.n4569 VDD.n4568 92.5005
R6050 VDD.n4570 VDD.n4569 92.5005
R6051 VDD.n1015 VDD.n1013 92.5005
R6052 VDD.n1013 VDD.n1002 92.5005
R6053 VDD.n1889 VDD.n1034 92.5005
R6054 VDD.n1034 VDD.n1001 92.5005
R6055 VDD.n1891 VDD.n1890 92.5005
R6056 VDD.n1892 VDD.n1891 92.5005
R6057 VDD.n1888 VDD.n1033 92.5005
R6058 VDD.n1816 VDD.n1033 92.5005
R6059 VDD.n1165 VDD.n1164 92.5005
R6060 VDD.n1168 VDD.n1167 92.5005
R6061 VDD.n1159 VDD.n1156 92.5005
R6062 VDD.n1174 VDD.n1173 92.5005
R6063 VDD.n1177 VDD.n1176 92.5005
R6064 VDD.n1153 VDD.n1149 92.5005
R6065 VDD.n1183 VDD.n1182 92.5005
R6066 VDD.n1185 VDD.n1145 92.5005
R6067 VDD.n1188 VDD.n1187 92.5005
R6068 VDD.n1190 VDD.n1189 92.5005
R6069 VDD.n1193 VDD.n1192 92.5005
R6070 VDD.n1142 VDD.n1139 92.5005
R6071 VDD.n1199 VDD.n1198 92.5005
R6072 VDD.n1202 VDD.n1201 92.5005
R6073 VDD.n1136 VDD.n1133 92.5005
R6074 VDD.n1208 VDD.n1207 92.5005
R6075 VDD.n1211 VDD.n1210 92.5005
R6076 VDD.n1130 VDD.n1127 92.5005
R6077 VDD.n1217 VDD.n1216 92.5005
R6078 VDD.n1220 VDD.n1219 92.5005
R6079 VDD.n1124 VDD.n1121 92.5005
R6080 VDD.n1226 VDD.n1225 92.5005
R6081 VDD.n1229 VDD.n1228 92.5005
R6082 VDD.n1118 VDD.n1114 92.5005
R6083 VDD.n1235 VDD.n1234 92.5005
R6084 VDD.n1237 VDD.n1110 92.5005
R6085 VDD.n1240 VDD.n1239 92.5005
R6086 VDD.n1242 VDD.n1241 92.5005
R6087 VDD.n1245 VDD.n1244 92.5005
R6088 VDD.n1107 VDD.n1104 92.5005
R6089 VDD.n1251 VDD.n1250 92.5005
R6090 VDD.n1254 VDD.n1253 92.5005
R6091 VDD.n1101 VDD.n1098 92.5005
R6092 VDD.n1260 VDD.n1259 92.5005
R6093 VDD.n1263 VDD.n1262 92.5005
R6094 VDD.n1095 VDD.n1091 92.5005
R6095 VDD.n1268 VDD.n1088 92.5005
R6096 VDD.n1817 VDD.n1275 92.5005
R6097 VDD.n1817 VDD.n1816 92.5005
R6098 VDD.n1388 VDD.n1029 92.5005
R6099 VDD.n1816 VDD.n1029 92.5005
R6100 VDD.n1894 VDD.n1893 92.5005
R6101 VDD.n1893 VDD.n1892 92.5005
R6102 VDD.n1895 VDD.n1007 92.5005
R6103 VDD.n1007 VDD.n1001 92.5005
R6104 VDD.n4573 VDD.n4572 92.5005
R6105 VDD.n4572 VDD.n1002 92.5005
R6106 VDD.n4571 VDD.n1010 92.5005
R6107 VDD.n4571 VDD.n4570 92.5005
R6108 VDD.n1904 VDD.n1008 92.5005
R6109 VDD.n2602 VDD.n1008 92.5005
R6110 VDD.n4563 VDD.n4562 92.5005
R6111 VDD.n4564 VDD.n4563 92.5005
R6112 VDD.n1025 VDD.n1020 92.5005
R6113 VDD.n1910 VDD.n1020 92.5005
R6114 VDD.n4553 VDD.n1026 92.5005
R6115 VDD.n4554 VDD.n4553 92.5005
R6116 VDD.n4552 VDD.n1916 92.5005
R6117 VDD.n4552 VDD.n4551 92.5005
R6118 VDD.n1935 VDD.n1913 92.5005
R6119 VDD.n1922 VDD.n1913 92.5005
R6120 VDD.n4544 VDD.n4543 92.5005
R6121 VDD.n4545 VDD.n4544 92.5005
R6122 VDD.n1930 VDD.n1925 92.5005
R6123 VDD.n1941 VDD.n1925 92.5005
R6124 VDD.n4534 VDD.n1931 92.5005
R6125 VDD.n4535 VDD.n4534 92.5005
R6126 VDD.n4533 VDD.n1947 92.5005
R6127 VDD.n4533 VDD.n4532 92.5005
R6128 VDD.n1971 VDD.n1944 92.5005
R6129 VDD.n2607 VDD.n1944 92.5005
R6130 VDD.n4525 VDD.n4524 92.5005
R6131 VDD.n4526 VDD.n4525 92.5005
R6132 VDD.n1960 VDD.n1955 92.5005
R6133 VDD.n1962 VDD.n1955 92.5005
R6134 VDD.n4518 VDD.n4517 92.5005
R6135 VDD.n4519 VDD.n4518 92.5005
R6136 VDD.n1976 VDD.n1965 92.5005
R6137 VDD.n1979 VDD.n1965 92.5005
R6138 VDD.n4509 VDD.n1977 92.5005
R6139 VDD.n4510 VDD.n4509 92.5005
R6140 VDD.n4508 VDD.n1985 92.5005
R6141 VDD.n4508 VDD.n4507 92.5005
R6142 VDD.n2007 VDD.n1982 92.5005
R6143 VDD.n1994 VDD.n1982 92.5005
R6144 VDD.n4500 VDD.n4499 92.5005
R6145 VDD.n4501 VDD.n4500 92.5005
R6146 VDD.n2002 VDD.n1997 92.5005
R6147 VDD.n2013 VDD.n1997 92.5005
R6148 VDD.n4490 VDD.n2003 92.5005
R6149 VDD.n4491 VDD.n4490 92.5005
R6150 VDD.n4489 VDD.n2020 92.5005
R6151 VDD.n4489 VDD.n4488 92.5005
R6152 VDD.n2040 VDD.n2017 92.5005
R6153 VDD.n2027 VDD.n2017 92.5005
R6154 VDD.n4481 VDD.n4480 92.5005
R6155 VDD.n4482 VDD.n4481 92.5005
R6156 VDD.n2035 VDD.n2030 92.5005
R6157 VDD.n2046 VDD.n2030 92.5005
R6158 VDD.n4471 VDD.n2036 92.5005
R6159 VDD.n4472 VDD.n4471 92.5005
R6160 VDD.n4470 VDD.n2052 92.5005
R6161 VDD.n4470 VDD.n4469 92.5005
R6162 VDD.n2087 VDD.n2049 92.5005
R6163 VDD.n2089 VDD.n2049 92.5005
R6164 VDD.n4462 VDD.n4461 92.5005
R6165 VDD.n4463 VDD.n4462 92.5005
R6166 VDD.n2064 VDD.n2059 92.5005
R6167 VDD.n2068 VDD.n2059 92.5005
R6168 VDD.n4456 VDD.n4455 92.5005
R6169 VDD.n4455 VDD.n4454 92.5005
R6170 VDD.n2078 VDD.n2067 92.5005
R6171 VDD.n2074 VDD.n2067 92.5005
R6172 VDD.n4447 VDD.n4446 92.5005
R6173 VDD.n4448 VDD.n4447 92.5005
R6174 VDD.n2082 VDD.n2077 92.5005
R6175 VDD.n2099 VDD.n2077 92.5005
R6176 VDD.n4437 VDD.n2083 92.5005
R6177 VDD.n4438 VDD.n4437 92.5005
R6178 VDD.n4436 VDD.n2105 92.5005
R6179 VDD.n4436 VDD.n4435 92.5005
R6180 VDD.n2124 VDD.n2102 92.5005
R6181 VDD.n2111 VDD.n2102 92.5005
R6182 VDD.n4428 VDD.n4427 92.5005
R6183 VDD.n4429 VDD.n4428 92.5005
R6184 VDD.n2119 VDD.n2114 92.5005
R6185 VDD.n2130 VDD.n2114 92.5005
R6186 VDD.n4418 VDD.n2120 92.5005
R6187 VDD.n4419 VDD.n4418 92.5005
R6188 VDD.n4417 VDD.n2135 92.5005
R6189 VDD.n4417 VDD.n4416 92.5005
R6190 VDD.n2155 VDD.n2132 92.5005
R6191 VDD.n2142 VDD.n2132 92.5005
R6192 VDD.n4409 VDD.n4408 92.5005
R6193 VDD.n4410 VDD.n4409 92.5005
R6194 VDD.n2150 VDD.n2145 92.5005
R6195 VDD.n2161 VDD.n2145 92.5005
R6196 VDD.n4399 VDD.n2151 92.5005
R6197 VDD.n4400 VDD.n4399 92.5005
R6198 VDD.n4398 VDD.n2167 92.5005
R6199 VDD.n4398 VDD.n4397 92.5005
R6200 VDD.n2192 VDD.n2164 92.5005
R6201 VDD.n2173 VDD.n2164 92.5005
R6202 VDD.n4390 VDD.n4389 92.5005
R6203 VDD.n4391 VDD.n4390 92.5005
R6204 VDD.n2181 VDD.n2176 92.5005
R6205 VDD.n2183 VDD.n2176 92.5005
R6206 VDD.n4383 VDD.n4382 92.5005
R6207 VDD.n4384 VDD.n4383 92.5005
R6208 VDD.n2197 VDD.n2186 92.5005
R6209 VDD.n2200 VDD.n2186 92.5005
R6210 VDD.n4374 VDD.n2198 92.5005
R6211 VDD.n4375 VDD.n4374 92.5005
R6212 VDD.n4373 VDD.n2206 92.5005
R6213 VDD.n4373 VDD.n4372 92.5005
R6214 VDD.n2228 VDD.n2203 92.5005
R6215 VDD.n2215 VDD.n2203 92.5005
R6216 VDD.n4365 VDD.n4364 92.5005
R6217 VDD.n4366 VDD.n4365 92.5005
R6218 VDD.n2223 VDD.n2218 92.5005
R6219 VDD.n2234 VDD.n2218 92.5005
R6220 VDD.n1390 VDD.n1028 92.5005
R6221 VDD.n1390 VDD.n1030 92.5005
R6222 VDD.n1896 VDD.n1003 92.5005
R6223 VDD.n1031 VDD.n1003 92.5005
R6224 VDD.n4575 VDD.n4574 92.5005
R6225 VDD.n4576 VDD.n4575 92.5005
R6226 VDD.n1009 VDD.n1004 92.5005
R6227 VDD.n1011 VDD.n1004 92.5005
R6228 VDD.n1906 VDD.n1905 92.5005
R6229 VDD.n1906 VDD.n1012 92.5005
R6230 VDD.n1907 VDD.n1021 92.5005
R6231 VDD.n1907 VDD.n1018 92.5005
R6232 VDD.n1908 VDD.n1022 92.5005
R6233 VDD.n2599 VDD.n1908 92.5005
R6234 VDD.n4557 VDD.n4556 92.5005
R6235 VDD.n4556 VDD.n4555 92.5005
R6236 VDD.n1915 VDD.n1909 92.5005
R6237 VDD.n1911 VDD.n1909 92.5005
R6238 VDD.n1937 VDD.n1936 92.5005
R6239 VDD.n1937 VDD.n1917 92.5005
R6240 VDD.n1938 VDD.n1926 92.5005
R6241 VDD.n1938 VDD.n1923 92.5005
R6242 VDD.n1939 VDD.n1927 92.5005
R6243 VDD.n1939 VDD.n1924 92.5005
R6244 VDD.n4538 VDD.n4537 92.5005
R6245 VDD.n4537 VDD.n4536 92.5005
R6246 VDD.n1946 VDD.n1940 92.5005
R6247 VDD.n1942 VDD.n1940 92.5005
R6248 VDD.n1970 VDD.n1969 92.5005
R6249 VDD.n1969 VDD.n1948 92.5005
R6250 VDD.n1958 VDD.n1956 92.5005
R6251 VDD.n1958 VDD.n1953 92.5005
R6252 VDD.n4523 VDD.n4522 92.5005
R6253 VDD.n4522 VDD.n1954 92.5005
R6254 VDD.n4521 VDD.n1961 92.5005
R6255 VDD.n4521 VDD.n4520 92.5005
R6256 VDD.n1966 VDD.n1959 92.5005
R6257 VDD.n1963 VDD.n1959 92.5005
R6258 VDD.n4513 VDD.n4512 92.5005
R6259 VDD.n4512 VDD.n4511 92.5005
R6260 VDD.n1984 VDD.n1978 92.5005
R6261 VDD.n1980 VDD.n1978 92.5005
R6262 VDD.n2009 VDD.n2008 92.5005
R6263 VDD.n2009 VDD.n1986 92.5005
R6264 VDD.n2010 VDD.n1998 92.5005
R6265 VDD.n2010 VDD.n1995 92.5005
R6266 VDD.n2011 VDD.n1999 92.5005
R6267 VDD.n2011 VDD.n1996 92.5005
R6268 VDD.n4494 VDD.n4493 92.5005
R6269 VDD.n4493 VDD.n4492 92.5005
R6270 VDD.n2019 VDD.n2012 92.5005
R6271 VDD.n2021 VDD.n2012 92.5005
R6272 VDD.n2042 VDD.n2041 92.5005
R6273 VDD.n2042 VDD.n2022 92.5005
R6274 VDD.n2043 VDD.n2031 92.5005
R6275 VDD.n2043 VDD.n2028 92.5005
R6276 VDD.n2044 VDD.n2032 92.5005
R6277 VDD.n2044 VDD.n2029 92.5005
R6278 VDD.n4475 VDD.n4474 92.5005
R6279 VDD.n4474 VDD.n4473 92.5005
R6280 VDD.n2051 VDD.n2045 92.5005
R6281 VDD.n2047 VDD.n2045 92.5005
R6282 VDD.n2091 VDD.n2088 92.5005
R6283 VDD.n2091 VDD.n2090 92.5005
R6284 VDD.n2092 VDD.n2060 92.5005
R6285 VDD.n2092 VDD.n2057 92.5005
R6286 VDD.n2093 VDD.n2061 92.5005
R6287 VDD.n2093 VDD.n2058 92.5005
R6288 VDD.n2094 VDD.n2065 92.5005
R6289 VDD.n2094 VDD.n2069 92.5005
R6290 VDD.n2095 VDD.n2066 92.5005
R6291 VDD.n2095 VDD.n2070 92.5005
R6292 VDD.n2096 VDD.n2079 92.5005
R6293 VDD.n2096 VDD.n2075 92.5005
R6294 VDD.n2097 VDD.n2080 92.5005
R6295 VDD.n2097 VDD.n2076 92.5005
R6296 VDD.n4441 VDD.n4440 92.5005
R6297 VDD.n4440 VDD.n4439 92.5005
R6298 VDD.n2104 VDD.n2098 92.5005
R6299 VDD.n2100 VDD.n2098 92.5005
R6300 VDD.n2126 VDD.n2125 92.5005
R6301 VDD.n2126 VDD.n2106 92.5005
R6302 VDD.n2127 VDD.n2115 92.5005
R6303 VDD.n2127 VDD.n2112 92.5005
R6304 VDD.n2128 VDD.n2116 92.5005
R6305 VDD.n2128 VDD.n2113 92.5005
R6306 VDD.n4422 VDD.n4421 92.5005
R6307 VDD.n4421 VDD.n4420 92.5005
R6308 VDD.n2134 VDD.n2129 92.5005
R6309 VDD.n2136 VDD.n2129 92.5005
R6310 VDD.n2157 VDD.n2156 92.5005
R6311 VDD.n2157 VDD.n2137 92.5005
R6312 VDD.n2158 VDD.n2146 92.5005
R6313 VDD.n2158 VDD.n2143 92.5005
R6314 VDD.n2159 VDD.n2147 92.5005
R6315 VDD.n2159 VDD.n2144 92.5005
R6316 VDD.n4403 VDD.n4402 92.5005
R6317 VDD.n4402 VDD.n4401 92.5005
R6318 VDD.n2166 VDD.n2160 92.5005
R6319 VDD.n2162 VDD.n2160 92.5005
R6320 VDD.n2191 VDD.n2190 92.5005
R6321 VDD.n2190 VDD.n2168 92.5005
R6322 VDD.n2179 VDD.n2177 92.5005
R6323 VDD.n2179 VDD.n2174 92.5005
R6324 VDD.n4388 VDD.n4387 92.5005
R6325 VDD.n4387 VDD.n2175 92.5005
R6326 VDD.n4386 VDD.n2182 92.5005
R6327 VDD.n4386 VDD.n4385 92.5005
R6328 VDD.n2187 VDD.n2180 92.5005
R6329 VDD.n2184 VDD.n2180 92.5005
R6330 VDD.n4378 VDD.n4377 92.5005
R6331 VDD.n4377 VDD.n4376 92.5005
R6332 VDD.n2205 VDD.n2199 92.5005
R6333 VDD.n2201 VDD.n2199 92.5005
R6334 VDD.n2230 VDD.n2229 92.5005
R6335 VDD.n2230 VDD.n2207 92.5005
R6336 VDD.n2231 VDD.n2219 92.5005
R6337 VDD.n2231 VDD.n2216 92.5005
R6338 VDD.n2232 VDD.n2220 92.5005
R6339 VDD.n2232 VDD.n2217 92.5005
R6340 VDD.n4359 VDD.n4358 92.5005
R6341 VDD.n4358 VDD.n4357 92.5005
R6342 VDD.n2235 VDD.n2233 92.5005
R6343 VDD.n4018 VDD.n4017 92.5005
R6344 VDD.n5653 VDD.t90 91.8719
R6345 VDD.n6522 VDD.t37 91.8719
R6346 VDD.n7362 VDD.t19 91.8719
R6347 VDD.n8231 VDD.t74 91.8719
R6348 VDD.n5163 VDD.n679 90.4767
R6349 VDD.n2351 VDD.n2350 86.0424
R6350 VDD.n5667 VDD.t91 84.4681
R6351 VDD.n6505 VDD.t38 84.4681
R6352 VDD.n7376 VDD.t20 84.4681
R6353 VDD.n8214 VDD.t75 84.4681
R6354 VDD.n4355 VDD.n2286 83.4438
R6355 VDD.n2292 VDD.n2237 83.4431
R6356 VDD.n5653 VDD.n5652 83.1021
R6357 VDD.n6522 VDD.n6521 83.1021
R6358 VDD.n7362 VDD.n7361 83.1021
R6359 VDD.n8231 VDD.n8230 83.1021
R6360 VDD.n2610 VDD.n2598 80.7889
R6361 VDD.n5642 VDD.t70 78.5582
R6362 VDD.t146 VDD.n6470 78.5582
R6363 VDD.n7351 VDD.t16 78.5582
R6364 VDD.t63 VDD.n8179 78.5582
R6365 VDD.n8995 VDD.n8994 78.4132
R6366 VDD.n8673 VDD.n8468 78.4132
R6367 VDD.n8140 VDD.n8139 78.4132
R6368 VDD.n7818 VDD.n7613 78.4132
R6369 VDD.n7286 VDD.n7285 78.4132
R6370 VDD.n6964 VDD.n6759 78.4132
R6371 VDD.n6431 VDD.n6430 78.4132
R6372 VDD.n6109 VDD.n5904 78.4132
R6373 VDD.t140 VDD.n4015 75.5912
R6374 VDD.n4015 VDD.t83 75.5912
R6375 VDD.n5285 VDD.n394 74.6009
R6376 VDD.n8339 VDD.n8274 72.0905
R6377 VDD.n8341 VDD.n8274 72.0905
R6378 VDD.n8640 VDD.n8502 72.0905
R6379 VDD.n8864 VDD.n8469 72.0905
R6380 VDD.n8864 VDD.n8470 72.0905
R6381 VDD.n8864 VDD.n8471 72.0905
R6382 VDD.n8864 VDD.n8472 72.0905
R6383 VDD.n8864 VDD.n8473 72.0905
R6384 VDD.n8864 VDD.n8474 72.0905
R6385 VDD.n8864 VDD.n8475 72.0905
R6386 VDD.n8864 VDD.n8476 72.0905
R6387 VDD.n8864 VDD.n8481 72.0905
R6388 VDD.n8864 VDD.n8482 72.0905
R6389 VDD.n8864 VDD.n8483 72.0905
R6390 VDD.n8864 VDD.n8484 72.0905
R6391 VDD.n8864 VDD.n8485 72.0905
R6392 VDD.n7484 VDD.n7419 72.0905
R6393 VDD.n7486 VDD.n7419 72.0905
R6394 VDD.n7785 VDD.n7647 72.0905
R6395 VDD.n8009 VDD.n7614 72.0905
R6396 VDD.n8009 VDD.n7615 72.0905
R6397 VDD.n8009 VDD.n7616 72.0905
R6398 VDD.n8009 VDD.n7617 72.0905
R6399 VDD.n8009 VDD.n7618 72.0905
R6400 VDD.n8009 VDD.n7619 72.0905
R6401 VDD.n8009 VDD.n7620 72.0905
R6402 VDD.n8009 VDD.n7621 72.0905
R6403 VDD.n8009 VDD.n7626 72.0905
R6404 VDD.n8009 VDD.n7627 72.0905
R6405 VDD.n8009 VDD.n7628 72.0905
R6406 VDD.n8009 VDD.n7629 72.0905
R6407 VDD.n8009 VDD.n7630 72.0905
R6408 VDD.n6630 VDD.n6565 72.0905
R6409 VDD.n6632 VDD.n6565 72.0905
R6410 VDD.n6931 VDD.n6793 72.0905
R6411 VDD.n7155 VDD.n6760 72.0905
R6412 VDD.n7155 VDD.n6761 72.0905
R6413 VDD.n7155 VDD.n6762 72.0905
R6414 VDD.n7155 VDD.n6763 72.0905
R6415 VDD.n7155 VDD.n6764 72.0905
R6416 VDD.n7155 VDD.n6765 72.0905
R6417 VDD.n7155 VDD.n6766 72.0905
R6418 VDD.n7155 VDD.n6767 72.0905
R6419 VDD.n7155 VDD.n6772 72.0905
R6420 VDD.n7155 VDD.n6773 72.0905
R6421 VDD.n7155 VDD.n6774 72.0905
R6422 VDD.n7155 VDD.n6775 72.0905
R6423 VDD.n7155 VDD.n6776 72.0905
R6424 VDD.n5775 VDD.n5710 72.0905
R6425 VDD.n5777 VDD.n5710 72.0905
R6426 VDD.n6076 VDD.n5938 72.0905
R6427 VDD.n6300 VDD.n5905 72.0905
R6428 VDD.n6300 VDD.n5906 72.0905
R6429 VDD.n6300 VDD.n5907 72.0905
R6430 VDD.n6300 VDD.n5908 72.0905
R6431 VDD.n6300 VDD.n5909 72.0905
R6432 VDD.n6300 VDD.n5910 72.0905
R6433 VDD.n6300 VDD.n5911 72.0905
R6434 VDD.n6300 VDD.n5912 72.0905
R6435 VDD.n6300 VDD.n5917 72.0905
R6436 VDD.n6300 VDD.n5918 72.0905
R6437 VDD.n6300 VDD.n5919 72.0905
R6438 VDD.n6300 VDD.n5920 72.0905
R6439 VDD.n6300 VDD.n5921 72.0905
R6440 VDD.n1082 VDD.n1059 72.0905
R6441 VDD.n1826 VDD.n1059 72.0905
R6442 VDD.n1081 VDD.n1059 72.0905
R6443 VDD.n1075 VDD.n1059 72.0905
R6444 VDD.n1835 VDD.n1059 72.0905
R6445 VDD.n1837 VDD.n1059 72.0905
R6446 VDD.n1074 VDD.n1059 72.0905
R6447 VDD.n1069 VDD.n1059 72.0905
R6448 VDD.n1846 VDD.n1059 72.0905
R6449 VDD.n1068 VDD.n1059 72.0905
R6450 VDD.n1063 VDD.n1059 72.0905
R6451 VDD.n1855 VDD.n1059 72.0905
R6452 VDD.n1160 VDD.n1032 72.0905
R6453 VDD.n1155 VDD.n1032 72.0905
R6454 VDD.n1175 VDD.n1032 72.0905
R6455 VDD.n1154 VDD.n1032 72.0905
R6456 VDD.n1147 VDD.n1032 72.0905
R6457 VDD.n1184 VDD.n1032 72.0905
R6458 VDD.n1186 VDD.n1032 72.0905
R6459 VDD.n1144 VDD.n1032 72.0905
R6460 VDD.n1191 VDD.n1032 72.0905
R6461 VDD.n1143 VDD.n1032 72.0905
R6462 VDD.n1138 VDD.n1032 72.0905
R6463 VDD.n1200 VDD.n1032 72.0905
R6464 VDD.n1137 VDD.n1032 72.0905
R6465 VDD.n1132 VDD.n1032 72.0905
R6466 VDD.n1209 VDD.n1032 72.0905
R6467 VDD.n1131 VDD.n1032 72.0905
R6468 VDD.n1126 VDD.n1032 72.0905
R6469 VDD.n1218 VDD.n1032 72.0905
R6470 VDD.n1125 VDD.n1032 72.0905
R6471 VDD.n1120 VDD.n1032 72.0905
R6472 VDD.n1227 VDD.n1032 72.0905
R6473 VDD.n1119 VDD.n1032 72.0905
R6474 VDD.n1112 VDD.n1032 72.0905
R6475 VDD.n1236 VDD.n1032 72.0905
R6476 VDD.n1238 VDD.n1032 72.0905
R6477 VDD.n1109 VDD.n1032 72.0905
R6478 VDD.n1243 VDD.n1032 72.0905
R6479 VDD.n1108 VDD.n1032 72.0905
R6480 VDD.n1103 VDD.n1032 72.0905
R6481 VDD.n1252 VDD.n1032 72.0905
R6482 VDD.n1102 VDD.n1032 72.0905
R6483 VDD.n1097 VDD.n1032 72.0905
R6484 VDD.n1261 VDD.n1032 72.0905
R6485 VDD.n1096 VDD.n1032 72.0905
R6486 VDD.n8853 VDD.n8683 71.1543
R6487 VDD.n8400 VDD.n8278 71.1543
R6488 VDD.n7998 VDD.n7828 71.1543
R6489 VDD.n7545 VDD.n7423 71.1543
R6490 VDD.n7144 VDD.n6974 71.1543
R6491 VDD.n6691 VDD.n6569 71.1543
R6492 VDD.n6289 VDD.n6119 71.1543
R6493 VDD.n5836 VDD.n5714 71.1543
R6494 VDD.n4350 VDD.n2285 70.5361
R6495 VDD.n4348 VDD.n2284 70.5361
R6496 VDD.n4346 VDD.n2283 70.5361
R6497 VDD.n4344 VDD.n2282 70.5361
R6498 VDD.n4342 VDD.n2281 70.5361
R6499 VDD.n4340 VDD.n2280 70.5361
R6500 VDD.n4338 VDD.n2279 70.5361
R6501 VDD.n4336 VDD.n2278 70.5361
R6502 VDD.n4334 VDD.n2277 70.5361
R6503 VDD.n4332 VDD.n2276 70.5361
R6504 VDD.n4330 VDD.n2275 70.5361
R6505 VDD.n4327 VDD.n2274 70.5361
R6506 VDD.n4325 VDD.n2273 70.5361
R6507 VDD.n4323 VDD.n2272 70.5361
R6508 VDD.n4321 VDD.n2271 70.5361
R6509 VDD.n4319 VDD.n2270 70.5361
R6510 VDD.n4317 VDD.n2269 70.5361
R6511 VDD.n4315 VDD.n2268 70.5361
R6512 VDD.n4313 VDD.n2267 70.5361
R6513 VDD.n4311 VDD.n2266 70.5361
R6514 VDD.n4309 VDD.n2265 70.5361
R6515 VDD.n4307 VDD.n2264 70.5361
R6516 VDD.n4305 VDD.n2263 70.5361
R6517 VDD.n4303 VDD.n2262 70.5361
R6518 VDD.n2338 VDD.n2261 70.5361
R6519 VDD.n2336 VDD.n2260 70.5361
R6520 VDD.n2334 VDD.n2259 70.5361
R6521 VDD.n2332 VDD.n2258 70.5361
R6522 VDD.n2330 VDD.n2257 70.5361
R6523 VDD.n2328 VDD.n2256 70.5361
R6524 VDD.n2326 VDD.n2255 70.5361
R6525 VDD.n2324 VDD.n2254 70.5361
R6526 VDD.n2322 VDD.n2253 70.5361
R6527 VDD.n2320 VDD.n2252 70.5361
R6528 VDD.n2318 VDD.n2251 70.5361
R6529 VDD.n2316 VDD.n2250 70.5361
R6530 VDD.n2314 VDD.n2249 70.5361
R6531 VDD.n2312 VDD.n2248 70.5361
R6532 VDD.n2310 VDD.n2247 70.5361
R6533 VDD.n2308 VDD.n2246 70.5361
R6534 VDD.n2306 VDD.n2245 70.5361
R6535 VDD.n2304 VDD.n2244 70.5361
R6536 VDD.n2302 VDD.n2243 70.5361
R6537 VDD.n2300 VDD.n2242 70.5361
R6538 VDD.n2298 VDD.n2241 70.5361
R6539 VDD.n2296 VDD.n2240 70.5361
R6540 VDD.n2294 VDD.n2239 70.5361
R6541 VDD.n2292 VDD.n2238 70.5361
R6542 VDD.n2294 VDD.n2238 70.5361
R6543 VDD.n2296 VDD.n2239 70.5361
R6544 VDD.n2298 VDD.n2240 70.5361
R6545 VDD.n2300 VDD.n2241 70.5361
R6546 VDD.n2302 VDD.n2242 70.5361
R6547 VDD.n2304 VDD.n2243 70.5361
R6548 VDD.n2306 VDD.n2244 70.5361
R6549 VDD.n2308 VDD.n2245 70.5361
R6550 VDD.n2310 VDD.n2246 70.5361
R6551 VDD.n2312 VDD.n2247 70.5361
R6552 VDD.n2314 VDD.n2248 70.5361
R6553 VDD.n2316 VDD.n2249 70.5361
R6554 VDD.n2318 VDD.n2250 70.5361
R6555 VDD.n2320 VDD.n2251 70.5361
R6556 VDD.n2322 VDD.n2252 70.5361
R6557 VDD.n2324 VDD.n2253 70.5361
R6558 VDD.n2326 VDD.n2254 70.5361
R6559 VDD.n2328 VDD.n2255 70.5361
R6560 VDD.n2330 VDD.n2256 70.5361
R6561 VDD.n2332 VDD.n2257 70.5361
R6562 VDD.n2334 VDD.n2258 70.5361
R6563 VDD.n2336 VDD.n2259 70.5361
R6564 VDD.n2338 VDD.n2260 70.5361
R6565 VDD.n4303 VDD.n2261 70.5361
R6566 VDD.n4305 VDD.n2262 70.5361
R6567 VDD.n4307 VDD.n2263 70.5361
R6568 VDD.n4309 VDD.n2264 70.5361
R6569 VDD.n4311 VDD.n2265 70.5361
R6570 VDD.n4313 VDD.n2266 70.5361
R6571 VDD.n4315 VDD.n2267 70.5361
R6572 VDD.n4317 VDD.n2268 70.5361
R6573 VDD.n4319 VDD.n2269 70.5361
R6574 VDD.n4321 VDD.n2270 70.5361
R6575 VDD.n4323 VDD.n2271 70.5361
R6576 VDD.n4325 VDD.n2272 70.5361
R6577 VDD.n4327 VDD.n2273 70.5361
R6578 VDD.n4330 VDD.n2274 70.5361
R6579 VDD.n4332 VDD.n2275 70.5361
R6580 VDD.n4334 VDD.n2276 70.5361
R6581 VDD.n4336 VDD.n2277 70.5361
R6582 VDD.n4338 VDD.n2278 70.5361
R6583 VDD.n4340 VDD.n2279 70.5361
R6584 VDD.n4342 VDD.n2280 70.5361
R6585 VDD.n4344 VDD.n2281 70.5361
R6586 VDD.n4346 VDD.n2282 70.5361
R6587 VDD.n4348 VDD.n2283 70.5361
R6588 VDD.n4350 VDD.n2284 70.5361
R6589 VDD.n2286 VDD.n2285 70.5361
R6590 VDD.n4006 VDD.n4005 69.0092
R6591 VDD.n3980 VDD.n2506 69.0092
R6592 VDD.n8388 VDD.n8294 67.9542
R6593 VDD.n8388 VDD.n8295 67.9542
R6594 VDD.n8349 VDD.n8267 67.9542
R6595 VDD.n8343 VDD.n8267 67.9542
R6596 VDD.n8354 VDD.n8267 67.9542
R6597 VDD.n8807 VDD.n8709 67.9542
R6598 VDD.n8797 VDD.n8709 67.9542
R6599 VDD.n8802 VDD.n8709 67.9542
R6600 VDD.n7533 VDD.n7439 67.9542
R6601 VDD.n7533 VDD.n7440 67.9542
R6602 VDD.n7494 VDD.n7412 67.9542
R6603 VDD.n7488 VDD.n7412 67.9542
R6604 VDD.n7499 VDD.n7412 67.9542
R6605 VDD.n7952 VDD.n7854 67.9542
R6606 VDD.n7942 VDD.n7854 67.9542
R6607 VDD.n7947 VDD.n7854 67.9542
R6608 VDD.n6679 VDD.n6585 67.9542
R6609 VDD.n6679 VDD.n6586 67.9542
R6610 VDD.n6640 VDD.n6558 67.9542
R6611 VDD.n6634 VDD.n6558 67.9542
R6612 VDD.n6645 VDD.n6558 67.9542
R6613 VDD.n7098 VDD.n7000 67.9542
R6614 VDD.n7088 VDD.n7000 67.9542
R6615 VDD.n7093 VDD.n7000 67.9542
R6616 VDD.n5824 VDD.n5730 67.9542
R6617 VDD.n5824 VDD.n5731 67.9542
R6618 VDD.n5785 VDD.n5703 67.9542
R6619 VDD.n5779 VDD.n5703 67.9542
R6620 VDD.n5790 VDD.n5703 67.9542
R6621 VDD.n6243 VDD.n6145 67.9542
R6622 VDD.n6233 VDD.n6145 67.9542
R6623 VDD.n6238 VDD.n6145 67.9542
R6624 VDD.n5448 VDD.n5447 66.8858
R6625 VDD.n1473 VDD.n1472 66.8856
R6626 VDD.n4010 VDD.n4009 64.4031
R6627 VDD.n3497 VDD.t105 60.2505
R6628 VDD.n3509 VDD.t123 60.2505
R6629 VDD.n3199 VDD.t121 60.2505
R6630 VDD.n3211 VDD.t114 60.2505
R6631 VDD.n3840 VDD.t102 60.2505
R6632 VDD.n3747 VDD.t108 60.2505
R6633 VDD.n3879 VDD.t110 60.2505
R6634 VDD.n3866 VDD.t112 60.2505
R6635 VDD.n2823 VDD.t125 60.2505
R6636 VDD.n2965 VDD.t118 60.2505
R6637 VDD.n8387 VDD.n8296 60.14
R6638 VDD.n8356 VDD.n8355 60.14
R6639 VDD.n8801 VDD.n8800 60.14
R6640 VDD.n7532 VDD.n7441 60.14
R6641 VDD.n7501 VDD.n7500 60.14
R6642 VDD.n7946 VDD.n7945 60.14
R6643 VDD.n6678 VDD.n6587 60.14
R6644 VDD.n6647 VDD.n6646 60.14
R6645 VDD.n7092 VDD.n7091 60.14
R6646 VDD.n5823 VDD.n5732 60.14
R6647 VDD.n5792 VDD.n5791 60.14
R6648 VDD.n6237 VDD.n6236 60.14
R6649 VDD.n8375 VDD.n8293 60.1394
R6650 VDD.n8348 VDD.n8347 60.1394
R6651 VDD.n8809 VDD.n8808 60.1394
R6652 VDD.n7520 VDD.n7438 60.1394
R6653 VDD.n7493 VDD.n7492 60.1394
R6654 VDD.n7954 VDD.n7953 60.1394
R6655 VDD.n6666 VDD.n6584 60.1394
R6656 VDD.n6639 VDD.n6638 60.1394
R6657 VDD.n7100 VDD.n7099 60.1394
R6658 VDD.n5811 VDD.n5729 60.1394
R6659 VDD.n5784 VDD.n5783 60.1394
R6660 VDD.n6245 VDD.n6244 60.1394
R6661 VDD.n2612 VDD.n2493 60.1048
R6662 VDD.n3987 VDD.n2493 60.1048
R6663 VDD.t107 VDD.n2668 59.2764
R6664 VDD.t117 VDD.n3137 59.2764
R6665 VDD.t109 VDD.n3792 59.2764
R6666 VDD.t120 VDD.n2924 59.2764
R6667 VDD.n66 VDD.t55 59.2764
R6668 VDD.n5571 VDD.t51 59.2764
R6669 VDD.n212 VDD.t7 59.2764
R6670 VDD.n4356 VDD.n2238 57.2334
R6671 VDD.n4356 VDD.n2239 57.2334
R6672 VDD.n4356 VDD.n2240 57.2334
R6673 VDD.n4356 VDD.n2241 57.2334
R6674 VDD.n4356 VDD.n2242 57.2334
R6675 VDD.n4356 VDD.n2243 57.2334
R6676 VDD.n4356 VDD.n2244 57.2334
R6677 VDD.n4356 VDD.n2245 57.2334
R6678 VDD.n4356 VDD.n2246 57.2334
R6679 VDD.n4356 VDD.n2247 57.2334
R6680 VDD.n4356 VDD.n2248 57.2334
R6681 VDD.n4356 VDD.n2249 57.2334
R6682 VDD.n4356 VDD.n2250 57.2334
R6683 VDD.n4356 VDD.n2251 57.2334
R6684 VDD.n4356 VDD.n2252 57.2334
R6685 VDD.n4356 VDD.n2253 57.2334
R6686 VDD.n4356 VDD.n2254 57.2334
R6687 VDD.n4356 VDD.n2255 57.2334
R6688 VDD.n4356 VDD.n2256 57.2334
R6689 VDD.n4356 VDD.n2257 57.2334
R6690 VDD.n4356 VDD.n2258 57.2334
R6691 VDD.n4356 VDD.n2259 57.2334
R6692 VDD.n4356 VDD.n2260 57.2334
R6693 VDD.n4356 VDD.n2261 57.2334
R6694 VDD.n4356 VDD.n2262 57.2334
R6695 VDD.n4356 VDD.n2263 57.2334
R6696 VDD.n4356 VDD.n2264 57.2334
R6697 VDD.n4356 VDD.n2265 57.2334
R6698 VDD.n4356 VDD.n2266 57.2334
R6699 VDD.n4356 VDD.n2267 57.2334
R6700 VDD.n4356 VDD.n2268 57.2334
R6701 VDD.n4356 VDD.n2269 57.2334
R6702 VDD.n4356 VDD.n2270 57.2334
R6703 VDD.n4356 VDD.n2271 57.2334
R6704 VDD.n4356 VDD.n2272 57.2334
R6705 VDD.n4356 VDD.n2273 57.2334
R6706 VDD.n4356 VDD.n2274 57.2334
R6707 VDD.n4356 VDD.n2275 57.2334
R6708 VDD.n4356 VDD.n2276 57.2334
R6709 VDD.n4356 VDD.n2277 57.2334
R6710 VDD.n4356 VDD.n2278 57.2334
R6711 VDD.n4356 VDD.n2279 57.2334
R6712 VDD.n4356 VDD.n2280 57.2334
R6713 VDD.n4356 VDD.n2281 57.2334
R6714 VDD.n4356 VDD.n2282 57.2334
R6715 VDD.n4356 VDD.n2283 57.2334
R6716 VDD.n4356 VDD.n2284 57.2334
R6717 VDD.n4356 VDD.n2285 57.2334
R6718 VDD.n4004 VDD.n2487 57.2295
R6719 VDD.n3948 VDD.n3945 57.2295
R6720 VDD.n8816 VDD.n8720 55.1287
R6721 VDD.n7961 VDD.n7865 55.1287
R6722 VDD.n7107 VDD.n7011 55.1287
R6723 VDD.n6252 VDD.n6156 55.1287
R6724 VDD.n1474 VDD.n1391 54.6255
R6725 VDD.n2352 VDD.n2351 54.3813
R6726 VDD.n1391 VDD.n1380 53.8338
R6727 VDD.n1730 VDD.n1037 53.8338
R6728 VDD.n1883 VDD.n1043 53.8338
R6729 VDD.n1874 VDD.n1043 53.8338
R6730 VDD.n1874 VDD.n1873 53.8338
R6731 VDD.n1873 VDD.n1872 53.8338
R6732 VDD.n1872 VDD.n1052 53.8338
R6733 VDD.n1863 VDD.n1052 53.8338
R6734 VDD.n1863 VDD.n1862 53.8338
R6735 VDD.n1862 VDD.n1861 53.8338
R6736 VDD.n2668 VDD.n2662 52.6902
R6737 VDD.n3137 VDD.n3131 52.6902
R6738 VDD.n3792 VDD.n3765 52.6902
R6739 VDD.n2924 VDD.n2921 52.6902
R6740 VDD.n67 VDD.n66 52.6902
R6741 VDD.n5572 VDD.n5571 52.6902
R6742 VDD.n213 VDD.n212 52.6902
R6743 VDD.n1403 VDD.n1381 51.067
R6744 VDD.n1457 VDD.n1382 51.067
R6745 VDD.n1447 VDD.n1383 51.067
R6746 VDD.n1439 VDD.n1384 51.067
R6747 VDD.n1429 VDD.n1385 51.067
R6748 VDD.n1479 VDD.n1386 51.067
R6749 VDD.n1456 VDD.n1381 51.0665
R6750 VDD.n1446 VDD.n1382 51.0665
R6751 VDD.n1438 VDD.n1383 51.0665
R6752 VDD.n1428 VDD.n1384 51.0665
R6753 VDD.n1416 VDD.n1385 51.0665
R6754 VDD.n1479 VDD.n1478 51.0665
R6755 VDD.n1725 VDD.n1038 51.0664
R6756 VDD.n1721 VDD.n1039 51.0664
R6757 VDD.n1717 VDD.n1040 51.0664
R6758 VDD.n1713 VDD.n1041 51.0664
R6759 VDD.n1709 VDD.n1042 51.0664
R6760 VDD.n1885 VDD.n1036 51.0664
R6761 VDD.n1886 VDD.n1885 51.0664
R6762 VDD.n1706 VDD.n1042 51.0664
R6763 VDD.n1710 VDD.n1041 51.0664
R6764 VDD.n1714 VDD.n1040 51.0664
R6765 VDD.n1718 VDD.n1039 51.0664
R6766 VDD.n1722 VDD.n1038 51.0664
R6767 VDD.n8366 VDD.n8365 50.7006
R6768 VDD.n8863 VDD.n8486 50.7006
R6769 VDD.n8764 VDD.n8477 50.7006
R6770 VDD.n7511 VDD.n7510 50.7006
R6771 VDD.n8008 VDD.n7631 50.7006
R6772 VDD.n7909 VDD.n7622 50.7006
R6773 VDD.n6657 VDD.n6656 50.7006
R6774 VDD.n7154 VDD.n6777 50.7006
R6775 VDD.n7055 VDD.n6768 50.7006
R6776 VDD.n5802 VDD.n5801 50.7006
R6777 VDD.n6299 VDD.n5922 50.7006
R6778 VDD.n6200 VDD.n5913 50.7006
R6779 VDD.n1856 VDD.n1061 50.7006
R6780 VDD.n925 VDD.n924 50.7006
R6781 VDD.n1095 VDD.n1094 50.7006
R6782 VDD.n8338 VDD.n8337 50.6999
R6783 VDD.n8999 VDD.n8273 50.6999
R6784 VDD.n8999 VDD.n8998 50.6999
R6785 VDD.n8641 VDD.n8637 50.6999
R6786 VDD.n8639 VDD.n8638 50.6999
R6787 VDD.n8865 VDD.n8467 50.6999
R6788 VDD.n8845 VDD.n8480 50.6999
R6789 VDD.n7483 VDD.n7482 50.6999
R6790 VDD.n8144 VDD.n7418 50.6999
R6791 VDD.n8144 VDD.n8143 50.6999
R6792 VDD.n7786 VDD.n7782 50.6999
R6793 VDD.n7784 VDD.n7783 50.6999
R6794 VDD.n8010 VDD.n7612 50.6999
R6795 VDD.n7990 VDD.n7625 50.6999
R6796 VDD.n6629 VDD.n6628 50.6999
R6797 VDD.n7290 VDD.n6564 50.6999
R6798 VDD.n7290 VDD.n7289 50.6999
R6799 VDD.n6932 VDD.n6928 50.6999
R6800 VDD.n6930 VDD.n6929 50.6999
R6801 VDD.n7156 VDD.n6758 50.6999
R6802 VDD.n7136 VDD.n6771 50.6999
R6803 VDD.n5774 VDD.n5773 50.6999
R6804 VDD.n6435 VDD.n5709 50.6999
R6805 VDD.n6435 VDD.n6434 50.6999
R6806 VDD.n6077 VDD.n6073 50.6999
R6807 VDD.n6075 VDD.n6074 50.6999
R6808 VDD.n6301 VDD.n5903 50.6999
R6809 VDD.n6281 VDD.n5916 50.6999
R6810 VDD.n1087 VDD.n1086 50.6999
R6811 VDD.n924 VDD.n920 50.6999
R6812 VDD.n1167 VDD.n1166 50.6999
R6813 VDD.n4018 VDD.n2464 50.6999
R6814 VDD.n4019 VDD.n4018 50.6999
R6815 VDD.n1861 VDD.n1059 50.6672
R6816 VDD.n8803 VDD.n8802 49.0945
R6817 VDD.n8806 VDD.n8797 49.0945
R6818 VDD.n8808 VDD.n8807 49.0945
R6819 VDD.n8378 VDD.n8295 49.0945
R6820 VDD.n8375 VDD.n8294 49.0945
R6821 VDD.n8378 VDD.n8294 49.0945
R6822 VDD.n8296 VDD.n8295 49.0945
R6823 VDD.n8354 VDD.n8353 49.0945
R6824 VDD.n8350 VDD.n8343 49.0945
R6825 VDD.n8349 VDD.n8348 49.0945
R6826 VDD.n8350 VDD.n8349 49.0945
R6827 VDD.n8353 VDD.n8343 49.0945
R6828 VDD.n8355 VDD.n8354 49.0945
R6829 VDD.n8807 VDD.n8806 49.0945
R6830 VDD.n8803 VDD.n8797 49.0945
R6831 VDD.n8802 VDD.n8801 49.0945
R6832 VDD.n7948 VDD.n7947 49.0945
R6833 VDD.n7951 VDD.n7942 49.0945
R6834 VDD.n7953 VDD.n7952 49.0945
R6835 VDD.n7523 VDD.n7440 49.0945
R6836 VDD.n7520 VDD.n7439 49.0945
R6837 VDD.n7523 VDD.n7439 49.0945
R6838 VDD.n7441 VDD.n7440 49.0945
R6839 VDD.n7499 VDD.n7498 49.0945
R6840 VDD.n7495 VDD.n7488 49.0945
R6841 VDD.n7494 VDD.n7493 49.0945
R6842 VDD.n7495 VDD.n7494 49.0945
R6843 VDD.n7498 VDD.n7488 49.0945
R6844 VDD.n7500 VDD.n7499 49.0945
R6845 VDD.n7952 VDD.n7951 49.0945
R6846 VDD.n7948 VDD.n7942 49.0945
R6847 VDD.n7947 VDD.n7946 49.0945
R6848 VDD.n7094 VDD.n7093 49.0945
R6849 VDD.n7097 VDD.n7088 49.0945
R6850 VDD.n7099 VDD.n7098 49.0945
R6851 VDD.n6669 VDD.n6586 49.0945
R6852 VDD.n6666 VDD.n6585 49.0945
R6853 VDD.n6669 VDD.n6585 49.0945
R6854 VDD.n6587 VDD.n6586 49.0945
R6855 VDD.n6645 VDD.n6644 49.0945
R6856 VDD.n6641 VDD.n6634 49.0945
R6857 VDD.n6640 VDD.n6639 49.0945
R6858 VDD.n6641 VDD.n6640 49.0945
R6859 VDD.n6644 VDD.n6634 49.0945
R6860 VDD.n6646 VDD.n6645 49.0945
R6861 VDD.n7098 VDD.n7097 49.0945
R6862 VDD.n7094 VDD.n7088 49.0945
R6863 VDD.n7093 VDD.n7092 49.0945
R6864 VDD.n6239 VDD.n6238 49.0945
R6865 VDD.n6242 VDD.n6233 49.0945
R6866 VDD.n6244 VDD.n6243 49.0945
R6867 VDD.n5814 VDD.n5731 49.0945
R6868 VDD.n5811 VDD.n5730 49.0945
R6869 VDD.n5814 VDD.n5730 49.0945
R6870 VDD.n5732 VDD.n5731 49.0945
R6871 VDD.n5790 VDD.n5789 49.0945
R6872 VDD.n5786 VDD.n5779 49.0945
R6873 VDD.n5785 VDD.n5784 49.0945
R6874 VDD.n5786 VDD.n5785 49.0945
R6875 VDD.n5789 VDD.n5779 49.0945
R6876 VDD.n5791 VDD.n5790 49.0945
R6877 VDD.n6243 VDD.n6242 49.0945
R6878 VDD.n6239 VDD.n6233 49.0945
R6879 VDD.n6238 VDD.n6237 49.0945
R6880 VDD.n1481 VDD.n1375 49.0838
R6881 VDD.n1486 VDD.n1484 49.0838
R6882 VDD.n1485 VDD.n1369 49.0838
R6883 VDD.n1497 VDD.n1496 49.0838
R6884 VDD.n1500 VDD.n1364 49.0838
R6885 VDD.n1502 VDD.n1501 49.0838
R6886 VDD.n1512 VDD.n1358 49.0838
R6887 VDD.n1513 VDD.n1353 49.0838
R6888 VDD.n1518 VDD.n1516 49.0838
R6889 VDD.n1517 VDD.n1347 49.0838
R6890 VDD.n1530 VDD.n1528 49.0838
R6891 VDD.n1529 VDD.n1341 49.0838
R6892 VDD.n1541 VDD.n1540 49.0838
R6893 VDD.n1544 VDD.n1336 49.0838
R6894 VDD.n1546 VDD.n1545 49.0838
R6895 VDD.n1556 VDD.n1330 49.0838
R6896 VDD.n1557 VDD.n1325 49.0838
R6897 VDD.n1562 VDD.n1560 49.0838
R6898 VDD.n1561 VDD.n1318 49.0838
R6899 VDD.n1572 VDD.n1571 49.0838
R6900 VDD.n1575 VDD.n1313 49.0838
R6901 VDD.n1577 VDD.n1576 49.0838
R6902 VDD.n1587 VDD.n1307 49.0838
R6903 VDD.n1588 VDD.n1302 49.0838
R6904 VDD.n1593 VDD.n1591 49.0838
R6905 VDD.n1592 VDD.n1296 49.0838
R6906 VDD.n1605 VDD.n1603 49.0838
R6907 VDD.n1604 VDD.n1290 49.0838
R6908 VDD.n1617 VDD.n1615 49.0838
R6909 VDD.n1616 VDD.n1276 49.0838
R6910 VDD.n1814 VDD.n1277 49.0838
R6911 VDD.n1805 VDD.n1622 49.0838
R6912 VDD.n1804 VDD.n1623 49.0838
R6913 VDD.n1801 VDD.n1800 49.0838
R6914 VDD.n1637 VDD.n1628 49.0838
R6915 VDD.n1790 VDD.n1638 49.0838
R6916 VDD.n1789 VDD.n1639 49.0838
R6917 VDD.n1786 VDD.n1785 49.0838
R6918 VDD.n1653 VDD.n1645 49.0838
R6919 VDD.n1776 VDD.n1654 49.0838
R6920 VDD.n1775 VDD.n1655 49.0838
R6921 VDD.n1772 VDD.n1771 49.0838
R6922 VDD.n1670 VDD.n1661 49.0838
R6923 VDD.n1761 VDD.n1671 49.0838
R6924 VDD.n1760 VDD.n1672 49.0838
R6925 VDD.n1757 VDD.n1756 49.0838
R6926 VDD.n1687 VDD.n1678 49.0838
R6927 VDD.n1746 VDD.n1688 49.0838
R6928 VDD.n1745 VDD.n1689 49.0838
R6929 VDD.n1742 VDD.n1741 49.0838
R6930 VDD.n1726 VDD.n1695 49.0838
R6931 VDD.n1731 VDD.n1727 49.0838
R6932 VDD.n2351 VDD.n2344 48.3613
R6933 VDD.n8390 VDD.n8389 48.0774
R6934 VDD.n7535 VDD.n7534 48.0774
R6935 VDD.n6681 VDD.n6680 48.0774
R6936 VDD.n5826 VDD.n5825 48.0774
R6937 VDD.n2289 VDD.n2213 46.4193
R6938 VDD.n3587 VDD.n3586 46.104
R6939 VDD.n3143 VDD.n3142 46.104
R6940 VDD.n3787 VDD.n3768 46.104
R6941 VDD.n2939 VDD.n2938 46.104
R6942 VDD.n63 VDD.n54 46.104
R6943 VDD.n5581 VDD.n5580 46.104
R6944 VDD.n209 VDD.n182 46.104
R6945 VDD.n3610 VDD.n2635 44.9671
R6946 VDD.n3169 VDD.n3093 44.9671
R6947 VDD.n8366 VDD.n8274 44.7682
R6948 VDD.n8864 VDD.n8477 44.7682
R6949 VDD.n8864 VDD.n8863 44.7682
R6950 VDD.n7511 VDD.n7419 44.7682
R6951 VDD.n8009 VDD.n7622 44.7682
R6952 VDD.n8009 VDD.n8008 44.7682
R6953 VDD.n6657 VDD.n6565 44.7682
R6954 VDD.n7155 VDD.n6768 44.7682
R6955 VDD.n7155 VDD.n7154 44.7682
R6956 VDD.n5802 VDD.n5710 44.7682
R6957 VDD.n6300 VDD.n5913 44.7682
R6958 VDD.n6300 VDD.n6299 44.7682
R6959 VDD.n1061 VDD.n1059 44.7682
R6960 VDD.n925 VDD.n921 44.7682
R6961 VDD.n1094 VDD.n1032 44.7682
R6962 VDD.n8337 VDD.n8274 44.768
R6963 VDD.n8274 VDD.n8273 44.768
R6964 VDD.n8998 VDD.n8274 44.768
R6965 VDD.n8637 VDD.n8502 44.768
R6966 VDD.n8638 VDD.n8502 44.768
R6967 VDD.n8865 VDD.n8864 44.768
R6968 VDD.n8864 VDD.n8480 44.768
R6969 VDD.n7482 VDD.n7419 44.768
R6970 VDD.n7419 VDD.n7418 44.768
R6971 VDD.n8143 VDD.n7419 44.768
R6972 VDD.n7782 VDD.n7647 44.768
R6973 VDD.n7783 VDD.n7647 44.768
R6974 VDD.n8010 VDD.n8009 44.768
R6975 VDD.n8009 VDD.n7625 44.768
R6976 VDD.n6628 VDD.n6565 44.768
R6977 VDD.n6565 VDD.n6564 44.768
R6978 VDD.n7289 VDD.n6565 44.768
R6979 VDD.n6928 VDD.n6793 44.768
R6980 VDD.n6929 VDD.n6793 44.768
R6981 VDD.n7156 VDD.n7155 44.768
R6982 VDD.n7155 VDD.n6771 44.768
R6983 VDD.n5773 VDD.n5710 44.768
R6984 VDD.n5710 VDD.n5709 44.768
R6985 VDD.n6434 VDD.n5710 44.768
R6986 VDD.n6073 VDD.n5938 44.768
R6987 VDD.n6074 VDD.n5938 44.768
R6988 VDD.n6301 VDD.n6300 44.768
R6989 VDD.n6300 VDD.n5916 44.768
R6990 VDD.n4020 VDD.n2464 44.768
R6991 VDD.n1087 VDD.n1059 44.768
R6992 VDD.n921 VDD.n920 44.768
R6993 VDD.n1166 VDD.n1032 44.768
R6994 VDD.n4020 VDD.n4019 44.768
R6995 VDD.n3950 VDD.n2473 44.4161
R6996 VDD.n2620 VDD.n2603 44.4161
R6997 VDD.n8400 VDD.n8286 43.5902
R6998 VDD.n7545 VDD.n7431 43.5902
R6999 VDD.n6691 VDD.n6577 43.5902
R7000 VDD.n5836 VDD.n5722 43.5902
R7001 VDD.n8960 VDD.n8959 41.7887
R7002 VDD.n8901 VDD.n8900 41.7887
R7003 VDD.n8105 VDD.n8104 41.7887
R7004 VDD.n8046 VDD.n8045 41.7887
R7005 VDD.n7251 VDD.n7250 41.7887
R7006 VDD.n7192 VDD.n7191 41.7887
R7007 VDD.n6396 VDD.n6395 41.7887
R7008 VDD.n6337 VDD.n6336 41.7887
R7009 VDD.n4355 VDD.n4354 41.7222
R7010 VDD.n2290 VDD.n2237 41.7221
R7011 VDD.n8388 VDD.n8387 41.6217
R7012 VDD.n8356 VDD.n8267 41.6217
R7013 VDD.n8800 VDD.n8709 41.6217
R7014 VDD.n7533 VDD.n7532 41.6217
R7015 VDD.n7501 VDD.n7412 41.6217
R7016 VDD.n7945 VDD.n7854 41.6217
R7017 VDD.n6679 VDD.n6678 41.6217
R7018 VDD.n6647 VDD.n6558 41.6217
R7019 VDD.n7091 VDD.n7000 41.6217
R7020 VDD.n5824 VDD.n5823 41.6217
R7021 VDD.n5792 VDD.n5703 41.6217
R7022 VDD.n6236 VDD.n6145 41.6217
R7023 VDD.n8388 VDD.n8293 41.6215
R7024 VDD.n8347 VDD.n8267 41.6215
R7025 VDD.n8809 VDD.n8709 41.6215
R7026 VDD.n7533 VDD.n7438 41.6215
R7027 VDD.n7492 VDD.n7412 41.6215
R7028 VDD.n7954 VDD.n7854 41.6215
R7029 VDD.n6679 VDD.n6584 41.6215
R7030 VDD.n6638 VDD.n6558 41.6215
R7031 VDD.n7100 VDD.n7000 41.6215
R7032 VDD.n5824 VDD.n5729 41.6215
R7033 VDD.n5783 VDD.n5703 41.6215
R7034 VDD.n6245 VDD.n6145 41.6215
R7035 VDD.n1884 VDD.n1037 41.1672
R7036 VDD.n3503 VDD.n3491 40.9783
R7037 VDD.n3514 VDD.n3505 40.9783
R7038 VDD.n3205 VDD.n3193 40.9783
R7039 VDD.n3216 VDD.n3207 40.9783
R7040 VDD.n3753 VDD.n3741 40.9783
R7041 VDD.n3831 VDD.n3738 40.9783
R7042 VDD.n3851 VDD.n3734 40.9783
R7043 VDD.n3884 VDD.n3875 40.9783
R7044 VDD.n3854 VDD.n3711 40.9783
R7045 VDD.n3873 VDD.n3706 40.9783
R7046 VDD.n2833 VDD.n2821 40.9783
R7047 VDD.n2975 VDD.n2963 40.9783
R7048 VDD.n8640 VDD.n8639 40.8219
R7049 VDD.n8857 VDD.n8485 40.8219
R7050 VDD.n8679 VDD.n8484 40.8219
R7051 VDD.n8690 VDD.n8483 40.8219
R7052 VDD.n8848 VDD.n8482 40.8219
R7053 VDD.n8845 VDD.n8481 40.8219
R7054 VDD.n8766 VDD.n8476 40.8219
R7055 VDD.n8770 VDD.n8475 40.8219
R7056 VDD.n8754 VDD.n8474 40.8219
R7057 VDD.n8776 VDD.n8473 40.8219
R7058 VDD.n8752 VDD.n8472 40.8219
R7059 VDD.n8782 VDD.n8471 40.8219
R7060 VDD.n8785 VDD.n8470 40.8219
R7061 VDD.n8469 VDD.n8467 40.8219
R7062 VDD.n8341 VDD.n8340 40.8219
R7063 VDD.n8339 VDD.n8338 40.8219
R7064 VDD.n8340 VDD.n8339 40.8219
R7065 VDD.n8365 VDD.n8341 40.8219
R7066 VDD.n8641 VDD.n8640 40.8219
R7067 VDD.n8764 VDD.n8476 40.8219
R7068 VDD.n8766 VDD.n8475 40.8219
R7069 VDD.n8770 VDD.n8474 40.8219
R7070 VDD.n8754 VDD.n8473 40.8219
R7071 VDD.n8776 VDD.n8472 40.8219
R7072 VDD.n8752 VDD.n8471 40.8219
R7073 VDD.n8782 VDD.n8470 40.8219
R7074 VDD.n8785 VDD.n8469 40.8219
R7075 VDD.n8486 VDD.n8485 40.8219
R7076 VDD.n8857 VDD.n8484 40.8219
R7077 VDD.n8679 VDD.n8483 40.8219
R7078 VDD.n8690 VDD.n8482 40.8219
R7079 VDD.n8848 VDD.n8481 40.8219
R7080 VDD.n7785 VDD.n7784 40.8219
R7081 VDD.n8002 VDD.n7630 40.8219
R7082 VDD.n7824 VDD.n7629 40.8219
R7083 VDD.n7835 VDD.n7628 40.8219
R7084 VDD.n7993 VDD.n7627 40.8219
R7085 VDD.n7990 VDD.n7626 40.8219
R7086 VDD.n7911 VDD.n7621 40.8219
R7087 VDD.n7915 VDD.n7620 40.8219
R7088 VDD.n7899 VDD.n7619 40.8219
R7089 VDD.n7921 VDD.n7618 40.8219
R7090 VDD.n7897 VDD.n7617 40.8219
R7091 VDD.n7927 VDD.n7616 40.8219
R7092 VDD.n7930 VDD.n7615 40.8219
R7093 VDD.n7614 VDD.n7612 40.8219
R7094 VDD.n7486 VDD.n7485 40.8219
R7095 VDD.n7484 VDD.n7483 40.8219
R7096 VDD.n7485 VDD.n7484 40.8219
R7097 VDD.n7510 VDD.n7486 40.8219
R7098 VDD.n7786 VDD.n7785 40.8219
R7099 VDD.n7909 VDD.n7621 40.8219
R7100 VDD.n7911 VDD.n7620 40.8219
R7101 VDD.n7915 VDD.n7619 40.8219
R7102 VDD.n7899 VDD.n7618 40.8219
R7103 VDD.n7921 VDD.n7617 40.8219
R7104 VDD.n7897 VDD.n7616 40.8219
R7105 VDD.n7927 VDD.n7615 40.8219
R7106 VDD.n7930 VDD.n7614 40.8219
R7107 VDD.n7631 VDD.n7630 40.8219
R7108 VDD.n8002 VDD.n7629 40.8219
R7109 VDD.n7824 VDD.n7628 40.8219
R7110 VDD.n7835 VDD.n7627 40.8219
R7111 VDD.n7993 VDD.n7626 40.8219
R7112 VDD.n6931 VDD.n6930 40.8219
R7113 VDD.n7148 VDD.n6776 40.8219
R7114 VDD.n6970 VDD.n6775 40.8219
R7115 VDD.n6981 VDD.n6774 40.8219
R7116 VDD.n7139 VDD.n6773 40.8219
R7117 VDD.n7136 VDD.n6772 40.8219
R7118 VDD.n7057 VDD.n6767 40.8219
R7119 VDD.n7061 VDD.n6766 40.8219
R7120 VDD.n7045 VDD.n6765 40.8219
R7121 VDD.n7067 VDD.n6764 40.8219
R7122 VDD.n7043 VDD.n6763 40.8219
R7123 VDD.n7073 VDD.n6762 40.8219
R7124 VDD.n7076 VDD.n6761 40.8219
R7125 VDD.n6760 VDD.n6758 40.8219
R7126 VDD.n6632 VDD.n6631 40.8219
R7127 VDD.n6630 VDD.n6629 40.8219
R7128 VDD.n6631 VDD.n6630 40.8219
R7129 VDD.n6656 VDD.n6632 40.8219
R7130 VDD.n6932 VDD.n6931 40.8219
R7131 VDD.n7055 VDD.n6767 40.8219
R7132 VDD.n7057 VDD.n6766 40.8219
R7133 VDD.n7061 VDD.n6765 40.8219
R7134 VDD.n7045 VDD.n6764 40.8219
R7135 VDD.n7067 VDD.n6763 40.8219
R7136 VDD.n7043 VDD.n6762 40.8219
R7137 VDD.n7073 VDD.n6761 40.8219
R7138 VDD.n7076 VDD.n6760 40.8219
R7139 VDD.n6777 VDD.n6776 40.8219
R7140 VDD.n7148 VDD.n6775 40.8219
R7141 VDD.n6970 VDD.n6774 40.8219
R7142 VDD.n6981 VDD.n6773 40.8219
R7143 VDD.n7139 VDD.n6772 40.8219
R7144 VDD.n6076 VDD.n6075 40.8219
R7145 VDD.n6293 VDD.n5921 40.8219
R7146 VDD.n6115 VDD.n5920 40.8219
R7147 VDD.n6126 VDD.n5919 40.8219
R7148 VDD.n6284 VDD.n5918 40.8219
R7149 VDD.n6281 VDD.n5917 40.8219
R7150 VDD.n6202 VDD.n5912 40.8219
R7151 VDD.n6206 VDD.n5911 40.8219
R7152 VDD.n6190 VDD.n5910 40.8219
R7153 VDD.n6212 VDD.n5909 40.8219
R7154 VDD.n6188 VDD.n5908 40.8219
R7155 VDD.n6218 VDD.n5907 40.8219
R7156 VDD.n6221 VDD.n5906 40.8219
R7157 VDD.n5905 VDD.n5903 40.8219
R7158 VDD.n5777 VDD.n5776 40.8219
R7159 VDD.n5775 VDD.n5774 40.8219
R7160 VDD.n5776 VDD.n5775 40.8219
R7161 VDD.n5801 VDD.n5777 40.8219
R7162 VDD.n6077 VDD.n6076 40.8219
R7163 VDD.n6200 VDD.n5912 40.8219
R7164 VDD.n6202 VDD.n5911 40.8219
R7165 VDD.n6206 VDD.n5910 40.8219
R7166 VDD.n6190 VDD.n5909 40.8219
R7167 VDD.n6212 VDD.n5908 40.8219
R7168 VDD.n6188 VDD.n5907 40.8219
R7169 VDD.n6218 VDD.n5906 40.8219
R7170 VDD.n6221 VDD.n5905 40.8219
R7171 VDD.n5922 VDD.n5921 40.8219
R7172 VDD.n6293 VDD.n5920 40.8219
R7173 VDD.n6115 VDD.n5919 40.8219
R7174 VDD.n6126 VDD.n5918 40.8219
R7175 VDD.n6284 VDD.n5917 40.8219
R7176 VDD.n1855 VDD.n1854 40.8219
R7177 VDD.n1067 VDD.n1063 40.8219
R7178 VDD.n1847 VDD.n1068 40.8219
R7179 VDD.n1846 VDD.n1845 40.8219
R7180 VDD.n1073 VDD.n1069 40.8219
R7181 VDD.n1838 VDD.n1074 40.8219
R7182 VDD.n1837 VDD.n1836 40.8219
R7183 VDD.n1835 VDD.n1834 40.8219
R7184 VDD.n1080 VDD.n1075 40.8219
R7185 VDD.n1827 VDD.n1081 40.8219
R7186 VDD.n1826 VDD.n1825 40.8219
R7187 VDD.n1086 VDD.n1082 40.8219
R7188 VDD.n1262 VDD.n1096 40.8219
R7189 VDD.n1261 VDD.n1260 40.8219
R7190 VDD.n1101 VDD.n1097 40.8219
R7191 VDD.n1253 VDD.n1102 40.8219
R7192 VDD.n1252 VDD.n1251 40.8219
R7193 VDD.n1107 VDD.n1103 40.8219
R7194 VDD.n1244 VDD.n1108 40.8219
R7195 VDD.n1243 VDD.n1242 40.8219
R7196 VDD.n1239 VDD.n1109 40.8219
R7197 VDD.n1238 VDD.n1237 40.8219
R7198 VDD.n1236 VDD.n1235 40.8219
R7199 VDD.n1118 VDD.n1112 40.8219
R7200 VDD.n1228 VDD.n1119 40.8219
R7201 VDD.n1227 VDD.n1226 40.8219
R7202 VDD.n1124 VDD.n1120 40.8219
R7203 VDD.n1219 VDD.n1125 40.8219
R7204 VDD.n1218 VDD.n1217 40.8219
R7205 VDD.n1130 VDD.n1126 40.8219
R7206 VDD.n1210 VDD.n1131 40.8219
R7207 VDD.n1209 VDD.n1208 40.8219
R7208 VDD.n1136 VDD.n1132 40.8219
R7209 VDD.n1201 VDD.n1137 40.8219
R7210 VDD.n1200 VDD.n1199 40.8219
R7211 VDD.n1142 VDD.n1138 40.8219
R7212 VDD.n1192 VDD.n1143 40.8219
R7213 VDD.n1191 VDD.n1190 40.8219
R7214 VDD.n1187 VDD.n1144 40.8219
R7215 VDD.n1186 VDD.n1185 40.8219
R7216 VDD.n1184 VDD.n1183 40.8219
R7217 VDD.n1153 VDD.n1147 40.8219
R7218 VDD.n1176 VDD.n1154 40.8219
R7219 VDD.n1175 VDD.n1174 40.8219
R7220 VDD.n1159 VDD.n1155 40.8219
R7221 VDD.n1167 VDD.n1160 40.8219
R7222 VDD.n1825 VDD.n1082 40.8219
R7223 VDD.n1827 VDD.n1826 40.8219
R7224 VDD.n1081 VDD.n1080 40.8219
R7225 VDD.n1834 VDD.n1075 40.8219
R7226 VDD.n1836 VDD.n1835 40.8219
R7227 VDD.n1838 VDD.n1837 40.8219
R7228 VDD.n1074 VDD.n1073 40.8219
R7229 VDD.n1845 VDD.n1069 40.8219
R7230 VDD.n1847 VDD.n1846 40.8219
R7231 VDD.n1068 VDD.n1067 40.8219
R7232 VDD.n1854 VDD.n1063 40.8219
R7233 VDD.n1856 VDD.n1855 40.8219
R7234 VDD.n1096 VDD.n1095 40.8219
R7235 VDD.n1262 VDD.n1261 40.8219
R7236 VDD.n1260 VDD.n1097 40.8219
R7237 VDD.n1102 VDD.n1101 40.8219
R7238 VDD.n1253 VDD.n1252 40.8219
R7239 VDD.n1251 VDD.n1103 40.8219
R7240 VDD.n1108 VDD.n1107 40.8219
R7241 VDD.n1244 VDD.n1243 40.8219
R7242 VDD.n1242 VDD.n1109 40.8219
R7243 VDD.n1239 VDD.n1238 40.8219
R7244 VDD.n1237 VDD.n1236 40.8219
R7245 VDD.n1235 VDD.n1112 40.8219
R7246 VDD.n1119 VDD.n1118 40.8219
R7247 VDD.n1228 VDD.n1227 40.8219
R7248 VDD.n1226 VDD.n1120 40.8219
R7249 VDD.n1125 VDD.n1124 40.8219
R7250 VDD.n1219 VDD.n1218 40.8219
R7251 VDD.n1217 VDD.n1126 40.8219
R7252 VDD.n1131 VDD.n1130 40.8219
R7253 VDD.n1210 VDD.n1209 40.8219
R7254 VDD.n1208 VDD.n1132 40.8219
R7255 VDD.n1137 VDD.n1136 40.8219
R7256 VDD.n1201 VDD.n1200 40.8219
R7257 VDD.n1199 VDD.n1138 40.8219
R7258 VDD.n1143 VDD.n1142 40.8219
R7259 VDD.n1192 VDD.n1191 40.8219
R7260 VDD.n1190 VDD.n1144 40.8219
R7261 VDD.n1187 VDD.n1186 40.8219
R7262 VDD.n1185 VDD.n1184 40.8219
R7263 VDD.n1183 VDD.n1147 40.8219
R7264 VDD.n1154 VDD.n1153 40.8219
R7265 VDD.n1176 VDD.n1175 40.8219
R7266 VDD.n1174 VDD.n1155 40.8219
R7267 VDD.n1160 VDD.n1159 40.8219
R7268 VDD.n1481 VDD.n1480 39.5838
R7269 VDD.n3596 VDD.n3595 39.5177
R7270 VDD.n3152 VDD.n3151 39.5177
R7271 VDD.n3781 VDD.n3642 39.5177
R7272 VDD.n2930 VDD.n2914 39.5177
R7273 VDD.n76 VDD.n50 39.5177
R7274 VDD.n5566 VDD.n5531 39.5177
R7275 VDD.n222 VDD.n179 39.5177
R7276 VDD.n4578 VDD.n4577 39.2068
R7277 VDD.n8746 VDD.n8723 38.7994
R7278 VDD.n8741 VDD.n8722 38.7994
R7279 VDD.n8738 VDD.n8721 38.7994
R7280 VDD.n8855 VDD.n8854 38.7994
R7281 VDD.n8397 VDD.n8396 38.7994
R7282 VDD.n8331 VDD.n8307 38.7994
R7283 VDD.n8330 VDD.n8308 38.7994
R7284 VDD.n8322 VDD.n8321 38.7994
R7285 VDD.n7891 VDD.n7868 38.7994
R7286 VDD.n7886 VDD.n7867 38.7994
R7287 VDD.n7883 VDD.n7866 38.7994
R7288 VDD.n8000 VDD.n7999 38.7994
R7289 VDD.n7542 VDD.n7541 38.7994
R7290 VDD.n7476 VDD.n7452 38.7994
R7291 VDD.n7475 VDD.n7453 38.7994
R7292 VDD.n7467 VDD.n7466 38.7994
R7293 VDD.n7037 VDD.n7014 38.7994
R7294 VDD.n7032 VDD.n7013 38.7994
R7295 VDD.n7029 VDD.n7012 38.7994
R7296 VDD.n7146 VDD.n7145 38.7994
R7297 VDD.n6688 VDD.n6687 38.7994
R7298 VDD.n6622 VDD.n6598 38.7994
R7299 VDD.n6621 VDD.n6599 38.7994
R7300 VDD.n6613 VDD.n6612 38.7994
R7301 VDD.n6182 VDD.n6159 38.7994
R7302 VDD.n6177 VDD.n6158 38.7994
R7303 VDD.n6174 VDD.n6157 38.7994
R7304 VDD.n6291 VDD.n6290 38.7994
R7305 VDD.n5833 VDD.n5832 38.7994
R7306 VDD.n5767 VDD.n5743 38.7994
R7307 VDD.n5766 VDD.n5744 38.7994
R7308 VDD.n5758 VDD.n5757 38.7994
R7309 VDD.n8739 VDD.n8722 38.7989
R7310 VDD.n8735 VDD.n8721 38.7989
R7311 VDD.n8746 VDD.n8745 38.7989
R7312 VDD.n8854 VDD.n8682 38.7989
R7313 VDD.n8397 VDD.n8287 38.7989
R7314 VDD.n8321 VDD.n8285 38.7989
R7315 VDD.n8320 VDD.n8308 38.7989
R7316 VDD.n8307 VDD.n8288 38.7989
R7317 VDD.n7884 VDD.n7867 38.7989
R7318 VDD.n7880 VDD.n7866 38.7989
R7319 VDD.n7891 VDD.n7890 38.7989
R7320 VDD.n7999 VDD.n7827 38.7989
R7321 VDD.n7542 VDD.n7432 38.7989
R7322 VDD.n7466 VDD.n7430 38.7989
R7323 VDD.n7465 VDD.n7453 38.7989
R7324 VDD.n7452 VDD.n7433 38.7989
R7325 VDD.n7030 VDD.n7013 38.7989
R7326 VDD.n7026 VDD.n7012 38.7989
R7327 VDD.n7037 VDD.n7036 38.7989
R7328 VDD.n7145 VDD.n6973 38.7989
R7329 VDD.n6688 VDD.n6578 38.7989
R7330 VDD.n6612 VDD.n6576 38.7989
R7331 VDD.n6611 VDD.n6599 38.7989
R7332 VDD.n6598 VDD.n6579 38.7989
R7333 VDD.n6175 VDD.n6158 38.7989
R7334 VDD.n6171 VDD.n6157 38.7989
R7335 VDD.n6182 VDD.n6181 38.7989
R7336 VDD.n6290 VDD.n6118 38.7989
R7337 VDD.n5833 VDD.n5723 38.7989
R7338 VDD.n5757 VDD.n5721 38.7989
R7339 VDD.n5756 VDD.n5744 38.7989
R7340 VDD.n5743 VDD.n5724 38.7989
R7341 VDD.n8852 VDD.n8688 38.7987
R7342 VDD.n8839 VDD.n8687 38.7987
R7343 VDD.n8852 VDD.n8851 38.7987
R7344 VDD.n8843 VDD.n8687 38.7987
R7345 VDD.n8773 VDD.n8686 38.7987
R7346 VDD.n8779 VDD.n8685 38.7987
R7347 VDD.n8788 VDD.n8684 38.7987
R7348 VDD.n8780 VDD.n8684 38.7987
R7349 VDD.n8774 VDD.n8685 38.7987
R7350 VDD.n8768 VDD.n8686 38.7987
R7351 VDD.n7997 VDD.n7833 38.7987
R7352 VDD.n7984 VDD.n7832 38.7987
R7353 VDD.n7997 VDD.n7996 38.7987
R7354 VDD.n7988 VDD.n7832 38.7987
R7355 VDD.n7918 VDD.n7831 38.7987
R7356 VDD.n7924 VDD.n7830 38.7987
R7357 VDD.n7933 VDD.n7829 38.7987
R7358 VDD.n7925 VDD.n7829 38.7987
R7359 VDD.n7919 VDD.n7830 38.7987
R7360 VDD.n7913 VDD.n7831 38.7987
R7361 VDD.n7143 VDD.n6979 38.7987
R7362 VDD.n7130 VDD.n6978 38.7987
R7363 VDD.n7143 VDD.n7142 38.7987
R7364 VDD.n7134 VDD.n6978 38.7987
R7365 VDD.n7064 VDD.n6977 38.7987
R7366 VDD.n7070 VDD.n6976 38.7987
R7367 VDD.n7079 VDD.n6975 38.7987
R7368 VDD.n7071 VDD.n6975 38.7987
R7369 VDD.n7065 VDD.n6976 38.7987
R7370 VDD.n7059 VDD.n6977 38.7987
R7371 VDD.n6288 VDD.n6124 38.7987
R7372 VDD.n6275 VDD.n6123 38.7987
R7373 VDD.n6288 VDD.n6287 38.7987
R7374 VDD.n6279 VDD.n6123 38.7987
R7375 VDD.n6209 VDD.n6122 38.7987
R7376 VDD.n6215 VDD.n6121 38.7987
R7377 VDD.n6224 VDD.n6120 38.7987
R7378 VDD.n6216 VDD.n6120 38.7987
R7379 VDD.n6210 VDD.n6121 38.7987
R7380 VDD.n6204 VDD.n6122 38.7987
R7381 VDD.n1724 VDD.n1705 38.777
R7382 VDD.n2459 VDD.n2458 38.4005
R7383 VDD.n8837 VDD.n8836 36.539
R7384 VDD.n8829 VDD.n8702 36.539
R7385 VDD.n7982 VDD.n7981 36.539
R7386 VDD.n7974 VDD.n7847 36.539
R7387 VDD.n7128 VDD.n7127 36.539
R7388 VDD.n7120 VDD.n6993 36.539
R7389 VDD.n6273 VDD.n6272 36.539
R7390 VDD.n6265 VDD.n6138 36.539
R7391 VDD.n2982 VDD.n2956 36.2246
R7392 VDD.n2458 VDD.n2442 36.2136
R7393 VDD.n5663 VDD.n5647 36.1417
R7394 VDD.n5663 VDD.n5662 36.1417
R7395 VDD.n5662 VDD.n5651 36.1417
R7396 VDD.n5658 VDD.n5651 36.1417
R7397 VDD.n5628 VDD.n5620 36.1417
R7398 VDD.n5639 VDD.n5620 36.1417
R7399 VDD.n5639 VDD.n5616 36.1417
R7400 VDD.n5670 VDD.n5616 36.1417
R7401 VDD.n6514 VDD.n6509 36.1417
R7402 VDD.n6514 VDD.n6513 36.1417
R7403 VDD.n6513 VDD.n6468 36.1417
R7404 VDD.n6519 VDD.n6468 36.1417
R7405 VDD.n6486 VDD.n6477 36.1417
R7406 VDD.n6491 VDD.n6477 36.1417
R7407 VDD.n6491 VDD.n6472 36.1417
R7408 VDD.n6502 VDD.n6472 36.1417
R7409 VDD.n7372 VDD.n7356 36.1417
R7410 VDD.n7372 VDD.n7371 36.1417
R7411 VDD.n7371 VDD.n7360 36.1417
R7412 VDD.n7367 VDD.n7360 36.1417
R7413 VDD.n7337 VDD.n7329 36.1417
R7414 VDD.n7348 VDD.n7329 36.1417
R7415 VDD.n7348 VDD.n7325 36.1417
R7416 VDD.n7379 VDD.n7325 36.1417
R7417 VDD.n8223 VDD.n8218 36.1417
R7418 VDD.n8223 VDD.n8222 36.1417
R7419 VDD.n8222 VDD.n8177 36.1417
R7420 VDD.n8228 VDD.n8177 36.1417
R7421 VDD.n8195 VDD.n8186 36.1417
R7422 VDD.n8200 VDD.n8186 36.1417
R7423 VDD.n8200 VDD.n8181 36.1417
R7424 VDD.n8211 VDD.n8181 36.1417
R7425 VDD.n8955 VDD.n8954 35.9626
R7426 VDD.n8100 VDD.n8099 35.9626
R7427 VDD.n7246 VDD.n7245 35.9626
R7428 VDD.n6391 VDD.n6390 35.9626
R7429 VDD.n8864 VDD.n8468 35.2569
R7430 VDD.n8009 VDD.n7613 35.2569
R7431 VDD.n7155 VDD.n6759 35.2569
R7432 VDD.n6300 VDD.n5904 35.2569
R7433 VDD.n5447 VDD.n5446 34.6359
R7434 VDD.n8994 VDD.n8274 34.6159
R7435 VDD.n8139 VDD.n7419 34.6159
R7436 VDD.n7285 VDD.n6565 34.6159
R7437 VDD.n6430 VDD.n5710 34.6159
R7438 VDD.n4721 VDD.n919 34.3808
R7439 VDD.n5160 VDD.n5159 34.3388
R7440 VDD.n1060 VDD.n1057 34.2989
R7441 VDD.n1472 VDD.n1471 33.9026
R7442 VDD.n4356 VDD.n4355 33.8538
R7443 VDD.n4356 VDD.n2237 33.8536
R7444 VDD.n8453 VDD.n8450 33.4435
R7445 VDD.n8964 VDD.n8963 33.4435
R7446 VDD.n8314 VDD.n8280 33.4435
R7447 VDD.n8310 VDD.n8305 33.4435
R7448 VDD.n8327 VDD.n8326 33.4435
R7449 VDD.n8313 VDD.n8312 33.4435
R7450 VDD.n8383 VDD.n8382 33.4435
R7451 VDD.n8302 VDD.n8299 33.4435
R7452 VDD.n8372 VDD.n8303 33.4435
R7453 VDD.n8535 VDD.n8533 33.4435
R7454 VDD.n8577 VDD.n8576 33.4435
R7455 VDD.n8646 VDD.n8645 33.4435
R7456 VDD.n7598 VDD.n7595 33.4435
R7457 VDD.n8109 VDD.n8108 33.4435
R7458 VDD.n7459 VDD.n7425 33.4435
R7459 VDD.n7455 VDD.n7450 33.4435
R7460 VDD.n7472 VDD.n7471 33.4435
R7461 VDD.n7458 VDD.n7457 33.4435
R7462 VDD.n7528 VDD.n7527 33.4435
R7463 VDD.n7447 VDD.n7444 33.4435
R7464 VDD.n7517 VDD.n7448 33.4435
R7465 VDD.n7680 VDD.n7678 33.4435
R7466 VDD.n7722 VDD.n7721 33.4435
R7467 VDD.n7791 VDD.n7790 33.4435
R7468 VDD.n6744 VDD.n6741 33.4435
R7469 VDD.n7255 VDD.n7254 33.4435
R7470 VDD.n6605 VDD.n6571 33.4435
R7471 VDD.n6601 VDD.n6596 33.4435
R7472 VDD.n6618 VDD.n6617 33.4435
R7473 VDD.n6604 VDD.n6603 33.4435
R7474 VDD.n6674 VDD.n6673 33.4435
R7475 VDD.n6593 VDD.n6590 33.4435
R7476 VDD.n6663 VDD.n6594 33.4435
R7477 VDD.n6826 VDD.n6824 33.4435
R7478 VDD.n6868 VDD.n6867 33.4435
R7479 VDD.n6937 VDD.n6936 33.4435
R7480 VDD.n5889 VDD.n5886 33.4435
R7481 VDD.n6400 VDD.n6399 33.4435
R7482 VDD.n5750 VDD.n5716 33.4435
R7483 VDD.n5746 VDD.n5741 33.4435
R7484 VDD.n5763 VDD.n5762 33.4435
R7485 VDD.n5749 VDD.n5748 33.4435
R7486 VDD.n5819 VDD.n5818 33.4435
R7487 VDD.n5738 VDD.n5735 33.4435
R7488 VDD.n5808 VDD.n5739 33.4435
R7489 VDD.n5971 VDD.n5969 33.4435
R7490 VDD.n6013 VDD.n6012 33.4435
R7491 VDD.n6082 VDD.n6081 33.4435
R7492 VDD.n2469 VDD.n2465 33.4435
R7493 VDD.n4021 VDD.n2463 33.4435
R7494 VDD.n1473 VDD.n1399 33.4435
R7495 VDD.n1400 VDD.n1392 33.4435
R7496 VDD.n1460 VDD.n1393 33.4435
R7497 VDD.n1450 VDD.n1394 33.4435
R7498 VDD.n1442 VDD.n1395 33.4435
R7499 VDD.n1432 VDD.n1396 33.4435
R7500 VDD.n1424 VDD.n1397 33.4435
R7501 VDD.n1472 VDD.n1398 33.4435
R7502 VDD.n1860 VDD.n1060 33.4435
R7503 VDD.n451 VDD.n393 33.4435
R7504 VDD.n5160 VDD.n677 33.4435
R7505 VDD.n4716 VDD.n919 33.4435
R7506 VDD.n8450 VDD.n8449 33.4431
R7507 VDD.n8963 VDD.n8962 33.4431
R7508 VDD.n8315 VDD.n8314 33.4431
R7509 VDD.n8316 VDD.n8313 33.4431
R7510 VDD.n8326 VDD.n8325 33.4431
R7511 VDD.n8311 VDD.n8310 33.4431
R7512 VDD.n8368 VDD.n8303 33.4431
R7513 VDD.n8373 VDD.n8302 33.4431
R7514 VDD.n8382 VDD.n8381 33.4431
R7515 VDD.n8576 VDD.n8575 33.4431
R7516 VDD.n8578 VDD.n8535 33.4431
R7517 VDD.n8645 VDD.n8505 33.4431
R7518 VDD.n7595 VDD.n7594 33.4431
R7519 VDD.n8108 VDD.n8107 33.4431
R7520 VDD.n7460 VDD.n7459 33.4431
R7521 VDD.n7461 VDD.n7458 33.4431
R7522 VDD.n7471 VDD.n7470 33.4431
R7523 VDD.n7456 VDD.n7455 33.4431
R7524 VDD.n7513 VDD.n7448 33.4431
R7525 VDD.n7518 VDD.n7447 33.4431
R7526 VDD.n7527 VDD.n7526 33.4431
R7527 VDD.n7721 VDD.n7720 33.4431
R7528 VDD.n7723 VDD.n7680 33.4431
R7529 VDD.n7790 VDD.n7650 33.4431
R7530 VDD.n6741 VDD.n6740 33.4431
R7531 VDD.n7254 VDD.n7253 33.4431
R7532 VDD.n6606 VDD.n6605 33.4431
R7533 VDD.n6607 VDD.n6604 33.4431
R7534 VDD.n6617 VDD.n6616 33.4431
R7535 VDD.n6602 VDD.n6601 33.4431
R7536 VDD.n6659 VDD.n6594 33.4431
R7537 VDD.n6664 VDD.n6593 33.4431
R7538 VDD.n6673 VDD.n6672 33.4431
R7539 VDD.n6867 VDD.n6866 33.4431
R7540 VDD.n6869 VDD.n6826 33.4431
R7541 VDD.n6936 VDD.n6796 33.4431
R7542 VDD.n5886 VDD.n5885 33.4431
R7543 VDD.n6399 VDD.n6398 33.4431
R7544 VDD.n5751 VDD.n5750 33.4431
R7545 VDD.n5752 VDD.n5749 33.4431
R7546 VDD.n5762 VDD.n5761 33.4431
R7547 VDD.n5747 VDD.n5746 33.4431
R7548 VDD.n5804 VDD.n5739 33.4431
R7549 VDD.n5809 VDD.n5738 33.4431
R7550 VDD.n5818 VDD.n5817 33.4431
R7551 VDD.n6012 VDD.n6011 33.4431
R7552 VDD.n6014 VDD.n5971 33.4431
R7553 VDD.n6081 VDD.n5941 33.4431
R7554 VDD.n5447 VDD.n282 33.4431
R7555 VDD.n2466 VDD.n2465 33.4431
R7556 VDD.n4022 VDD.n4021 33.4431
R7557 VDD.n1461 VDD.n1392 33.4431
R7558 VDD.n1449 VDD.n1393 33.4431
R7559 VDD.n1443 VDD.n1394 33.4431
R7560 VDD.n1431 VDD.n1395 33.4431
R7561 VDD.n1425 VDD.n1396 33.4431
R7562 VDD.n1397 VDD.n1389 33.4431
R7563 VDD.n1060 VDD.n1058 33.4431
R7564 VDD.n456 VDD.n451 33.4431
R7565 VDD.n5161 VDD.n5160 33.4431
R7566 VDD.n4719 VDD.n919 33.4431
R7567 VDD.n8761 VDD.n8478 33.4428
R7568 VDD.n8758 VDD.n8478 33.4428
R7569 VDD.n7906 VDD.n7623 33.4428
R7570 VDD.n7903 VDD.n7623 33.4428
R7571 VDD.n7052 VDD.n6769 33.4428
R7572 VDD.n7049 VDD.n6769 33.4428
R7573 VDD.n6197 VDD.n5914 33.4428
R7574 VDD.n6194 VDD.n5914 33.4428
R7575 VDD.n5448 VDD.n279 33.4428
R7576 VDD.n5450 VDD.n280 33.4428
R7577 VDD.n5439 VDD.n295 33.4428
R7578 VDD.n5428 VDD.n294 33.4428
R7579 VDD.n5419 VDD.n293 33.4428
R7580 VDD.n5416 VDD.n292 33.4428
R7581 VDD.n5407 VDD.n291 33.4428
R7582 VDD.n5404 VDD.n290 33.4428
R7583 VDD.n313 VDD.n289 33.4428
R7584 VDD.n5396 VDD.n288 33.4428
R7585 VDD.n5387 VDD.n287 33.4428
R7586 VDD.n5384 VDD.n286 33.4428
R7587 VDD.n5375 VDD.n285 33.4428
R7588 VDD.n5372 VDD.n284 33.4428
R7589 VDD.n328 VDD.n283 33.4428
R7590 VDD.n457 VDD.n447 33.4428
R7591 VDD.n468 VDD.n466 33.4428
R7592 VDD.n475 VDD.n443 33.4428
R7593 VDD.n476 VDD.n439 33.4428
R7594 VDD.n487 VDD.n486 33.4428
R7595 VDD.n488 VDD.n435 33.4428
R7596 VDD.n499 VDD.n497 33.4428
R7597 VDD.n506 VDD.n431 33.4428
R7598 VDD.n507 VDD.n427 33.4428
R7599 VDD.n518 VDD.n516 33.4428
R7600 VDD.n525 VDD.n423 33.4428
R7601 VDD.n526 VDD.n419 33.4428
R7602 VDD.n538 VDD.n535 33.4428
R7603 VDD.n536 VDD.n415 33.4428
R7604 VDD.n549 VDD.n547 33.4428
R7605 VDD.n556 VDD.n411 33.4428
R7606 VDD.n557 VDD.n407 33.4428
R7607 VDD.n568 VDD.n566 33.4428
R7608 VDD.n575 VDD.n403 33.4428
R7609 VDD.n576 VDD.n397 33.4428
R7610 VDD.n5371 VDD.n283 33.4428
R7611 VDD.n5376 VDD.n284 33.4428
R7612 VDD.n5383 VDD.n285 33.4428
R7613 VDD.n5388 VDD.n286 33.4428
R7614 VDD.n5395 VDD.n287 33.4428
R7615 VDD.n314 VDD.n288 33.4428
R7616 VDD.n5403 VDD.n289 33.4428
R7617 VDD.n5408 VDD.n290 33.4428
R7618 VDD.n5415 VDD.n291 33.4428
R7619 VDD.n5420 VDD.n292 33.4428
R7620 VDD.n5427 VDD.n293 33.4428
R7621 VDD.n5431 VDD.n294 33.4428
R7622 VDD.n5439 VDD.n5438 33.4428
R7623 VDD.n5451 VDD.n5450 33.4428
R7624 VDD.n458 VDD.n457 33.4428
R7625 VDD.n466 VDD.n465 33.4428
R7626 VDD.n467 VDD.n443 33.4428
R7627 VDD.n477 VDD.n476 33.4428
R7628 VDD.n486 VDD.n485 33.4428
R7629 VDD.n489 VDD.n488 33.4428
R7630 VDD.n497 VDD.n496 33.4428
R7631 VDD.n498 VDD.n431 33.4428
R7632 VDD.n508 VDD.n507 33.4428
R7633 VDD.n516 VDD.n515 33.4428
R7634 VDD.n517 VDD.n423 33.4428
R7635 VDD.n527 VDD.n526 33.4428
R7636 VDD.n535 VDD.n534 33.4428
R7637 VDD.n537 VDD.n536 33.4428
R7638 VDD.n547 VDD.n546 33.4428
R7639 VDD.n548 VDD.n411 33.4428
R7640 VDD.n558 VDD.n557 33.4428
R7641 VDD.n566 VDD.n565 33.4428
R7642 VDD.n567 VDD.n403 33.4428
R7643 VDD.n577 VDD.n576 33.4428
R7644 VDD.n8897 VDD.n8446 32.9658
R7645 VDD.n8042 VDD.n7591 32.9658
R7646 VDD.n7188 VDD.n6737 32.9658
R7647 VDD.n6333 VDD.n5882 32.9658
R7648 VDD.n2657 VDD.n2656 32.9315
R7649 VDD.n3126 VDD.n3125 32.9315
R7650 VDD.n2998 VDD.n2915 32.9315
R7651 VDD.n88 VDD.n85 32.9315
R7652 VDD.n5593 VDD.n5592 32.9315
R7653 VDD.n234 VDD.n233 32.9315
R7654 VDD.n8645 VDD.n8644 32.6607
R7655 VDD.n7790 VDD.n7789 32.6607
R7656 VDD.n6936 VDD.n6935 32.6607
R7657 VDD.n6081 VDD.n6080 32.6607
R7658 VDD.n8390 VDD.n8388 30.1287
R7659 VDD.n7535 VDD.n7533 30.1287
R7660 VDD.n6681 VDD.n6679 30.1287
R7661 VDD.n5826 VDD.n5824 30.1287
R7662 VDD.n8744 VDD.n8731 30.1181
R7663 VDD.n8359 VDD.n8358 30.1181
R7664 VDD.n8345 VDD.n8256 30.1181
R7665 VDD.n8820 VDD.n8712 30.1181
R7666 VDD.n8812 VDD.n8811 30.1181
R7667 VDD.n7889 VDD.n7876 30.1181
R7668 VDD.n7504 VDD.n7503 30.1181
R7669 VDD.n7490 VDD.n7401 30.1181
R7670 VDD.n7965 VDD.n7857 30.1181
R7671 VDD.n7957 VDD.n7956 30.1181
R7672 VDD.n7035 VDD.n7022 30.1181
R7673 VDD.n6650 VDD.n6649 30.1181
R7674 VDD.n6636 VDD.n6547 30.1181
R7675 VDD.n7111 VDD.n7003 30.1181
R7676 VDD.n7103 VDD.n7102 30.1181
R7677 VDD.n6180 VDD.n6167 30.1181
R7678 VDD.n5795 VDD.n5794 30.1181
R7679 VDD.n5781 VDD.n5692 30.1181
R7680 VDD.n6256 VDD.n6148 30.1181
R7681 VDD.n6248 VDD.n6247 30.1181
R7682 VDD.n8387 VDD.n8386 30.0704
R7683 VDD.n8357 VDD.n8356 30.0704
R7684 VDD.n8800 VDD.n8799 30.0704
R7685 VDD.n7532 VDD.n7531 30.0704
R7686 VDD.n7502 VDD.n7501 30.0704
R7687 VDD.n7945 VDD.n7944 30.0704
R7688 VDD.n6678 VDD.n6677 30.0704
R7689 VDD.n6648 VDD.n6647 30.0704
R7690 VDD.n7091 VDD.n7090 30.0704
R7691 VDD.n5823 VDD.n5822 30.0704
R7692 VDD.n5793 VDD.n5792 30.0704
R7693 VDD.n6236 VDD.n6235 30.0704
R7694 VDD.n8810 VDD.n8809 30.0702
R7695 VDD.n8300 VDD.n8293 30.0702
R7696 VDD.n8347 VDD.n8346 30.0702
R7697 VDD.n7955 VDD.n7954 30.0702
R7698 VDD.n7445 VDD.n7438 30.0702
R7699 VDD.n7492 VDD.n7491 30.0702
R7700 VDD.n7101 VDD.n7100 30.0702
R7701 VDD.n6591 VDD.n6584 30.0702
R7702 VDD.n6638 VDD.n6637 30.0702
R7703 VDD.n6246 VDD.n6245 30.0702
R7704 VDD.n5736 VDD.n5729 30.0702
R7705 VDD.n5783 VDD.n5782 30.0702
R7706 VDD.n3608 VDD.n2639 29.6384
R7707 VDD.n3167 VDD.n3096 29.6384
R7708 VDD.n2987 VDD.n2951 29.6384
R7709 VDD.n98 VDD.n97 29.6384
R7710 VDD.n5556 VDD.n5555 29.6384
R7711 VDD.n197 VDD.n196 29.6384
R7712 VDD.n8898 VDD.n8450 29.5303
R7713 VDD.n8963 VDD.n8418 29.5303
R7714 VDD.n8310 VDD.n8274 29.5303
R7715 VDD.n8326 VDD.n8274 29.5303
R7716 VDD.n8313 VDD.n8274 29.5303
R7717 VDD.n8314 VDD.n8274 29.5303
R7718 VDD.n8382 VDD.n8274 29.5303
R7719 VDD.n8302 VDD.n8274 29.5303
R7720 VDD.n8303 VDD.n8274 29.5303
R7721 VDD.n8536 VDD.n8535 29.5303
R7722 VDD.n8576 VDD.n8536 29.5303
R7723 VDD.n8043 VDD.n7595 29.5303
R7724 VDD.n8108 VDD.n7563 29.5303
R7725 VDD.n7455 VDD.n7419 29.5303
R7726 VDD.n7471 VDD.n7419 29.5303
R7727 VDD.n7458 VDD.n7419 29.5303
R7728 VDD.n7459 VDD.n7419 29.5303
R7729 VDD.n7527 VDD.n7419 29.5303
R7730 VDD.n7447 VDD.n7419 29.5303
R7731 VDD.n7448 VDD.n7419 29.5303
R7732 VDD.n7681 VDD.n7680 29.5303
R7733 VDD.n7721 VDD.n7681 29.5303
R7734 VDD.n7189 VDD.n6741 29.5303
R7735 VDD.n7254 VDD.n6709 29.5303
R7736 VDD.n6601 VDD.n6565 29.5303
R7737 VDD.n6617 VDD.n6565 29.5303
R7738 VDD.n6604 VDD.n6565 29.5303
R7739 VDD.n6605 VDD.n6565 29.5303
R7740 VDD.n6673 VDD.n6565 29.5303
R7741 VDD.n6593 VDD.n6565 29.5303
R7742 VDD.n6594 VDD.n6565 29.5303
R7743 VDD.n6827 VDD.n6826 29.5303
R7744 VDD.n6867 VDD.n6827 29.5303
R7745 VDD.n6334 VDD.n5886 29.5303
R7746 VDD.n6399 VDD.n5854 29.5303
R7747 VDD.n5746 VDD.n5710 29.5303
R7748 VDD.n5762 VDD.n5710 29.5303
R7749 VDD.n5749 VDD.n5710 29.5303
R7750 VDD.n5750 VDD.n5710 29.5303
R7751 VDD.n5818 VDD.n5710 29.5303
R7752 VDD.n5738 VDD.n5710 29.5303
R7753 VDD.n5739 VDD.n5710 29.5303
R7754 VDD.n5972 VDD.n5971 29.5303
R7755 VDD.n6012 VDD.n5972 29.5303
R7756 VDD.n4020 VDD.n2465 29.5303
R7757 VDD.n4021 VDD.n4020 29.5303
R7758 VDD.n1474 VDD.n1392 29.5303
R7759 VDD.n1474 VDD.n1393 29.5303
R7760 VDD.n1474 VDD.n1394 29.5303
R7761 VDD.n1474 VDD.n1395 29.5303
R7762 VDD.n1474 VDD.n1396 29.5303
R7763 VDD.n1474 VDD.n1397 29.5303
R7764 VDD.n1474 VDD.n1473 29.5303
R7765 VDD.n451 VDD.n395 29.5303
R7766 VDD.n8864 VDD.n8478 29.5301
R7767 VDD.n8009 VDD.n7623 29.5301
R7768 VDD.n7155 VDD.n6769 29.5301
R7769 VDD.n6300 VDD.n5914 29.5301
R7770 VDD.n5449 VDD.n283 29.5301
R7771 VDD.n5449 VDD.n284 29.5301
R7772 VDD.n5449 VDD.n285 29.5301
R7773 VDD.n5449 VDD.n286 29.5301
R7774 VDD.n5449 VDD.n287 29.5301
R7775 VDD.n5449 VDD.n288 29.5301
R7776 VDD.n5449 VDD.n289 29.5301
R7777 VDD.n5449 VDD.n290 29.5301
R7778 VDD.n5449 VDD.n291 29.5301
R7779 VDD.n5449 VDD.n292 29.5301
R7780 VDD.n5449 VDD.n293 29.5301
R7781 VDD.n5449 VDD.n294 29.5301
R7782 VDD.n5449 VDD.n5439 29.5301
R7783 VDD.n5450 VDD.n5449 29.5301
R7784 VDD.n5449 VDD.n5448 29.5301
R7785 VDD.n457 VDD.n395 29.5301
R7786 VDD.n466 VDD.n395 29.5301
R7787 VDD.n443 VDD.n395 29.5301
R7788 VDD.n476 VDD.n395 29.5301
R7789 VDD.n486 VDD.n395 29.5301
R7790 VDD.n488 VDD.n395 29.5301
R7791 VDD.n497 VDD.n395 29.5301
R7792 VDD.n431 VDD.n395 29.5301
R7793 VDD.n507 VDD.n395 29.5301
R7794 VDD.n516 VDD.n395 29.5301
R7795 VDD.n423 VDD.n395 29.5301
R7796 VDD.n526 VDD.n395 29.5301
R7797 VDD.n535 VDD.n395 29.5301
R7798 VDD.n536 VDD.n395 29.5301
R7799 VDD.n547 VDD.n395 29.5301
R7800 VDD.n411 VDD.n395 29.5301
R7801 VDD.n557 VDD.n395 29.5301
R7802 VDD.n566 VDD.n395 29.5301
R7803 VDD.n403 VDD.n395 29.5301
R7804 VDD.n576 VDD.n395 29.5301
R7805 VDD.n9017 VDD.n8251 29.4877
R7806 VDD.n9011 VDD.n8259 29.4877
R7807 VDD.n8162 VDD.n7396 29.4877
R7808 VDD.n8156 VDD.n7404 29.4877
R7809 VDD.n7308 VDD.n6542 29.4877
R7810 VDD.n7302 VDD.n6550 29.4877
R7811 VDD.n6453 VDD.n5687 29.4877
R7812 VDD.n6447 VDD.n5695 29.4877
R7813 VDD.n2618 VDD.n2617 29.4133
R7814 VDD.n2617 VDD.n2475 29.4133
R7815 VDD.t156 VDD.n8708 28.8467
R7816 VDD.t72 VDD.n8749 28.8467
R7817 VDD.t28 VDD.n8260 28.8467
R7818 VDD.t34 VDD.n7853 28.8467
R7819 VDD.t85 VDD.n7894 28.8467
R7820 VDD.t151 VDD.n7405 28.8467
R7821 VDD.t2 VDD.n6999 28.8467
R7822 VDD.t87 VDD.n7040 28.8467
R7823 VDD.t132 VDD.n6551 28.8467
R7824 VDD.t12 VDD.n6144 28.8467
R7825 VDD.t139 VDD.n6185 28.8467
R7826 VDD.t58 VDD.n5696 28.8467
R7827 VDD.n2471 VDD.n2468 28.5972
R7828 VDD.n2468 VDD.n2467 28.5972
R7829 VDD.n2467 VDD.n2462 28.5972
R7830 VDD.n4023 VDD.n2462 28.5972
R7831 VDD.n4287 VDD.n2367 28.5972
R7832 VDD.n4287 VDD.n4286 28.5972
R7833 VDD.n4286 VDD.n4285 28.5972
R7834 VDD.n4285 VDD.n2368 28.5972
R7835 VDD.n4276 VDD.n2368 28.5972
R7836 VDD.n4275 VDD.n4274 28.5972
R7837 VDD.n4274 VDD.n2375 28.5972
R7838 VDD.n4265 VDD.n2375 28.5972
R7839 VDD.n4265 VDD.n4264 28.5972
R7840 VDD.n4264 VDD.n4263 28.5972
R7841 VDD.n4263 VDD.n2384 28.5972
R7842 VDD.n4254 VDD.n4253 28.5972
R7843 VDD.n4253 VDD.n4252 28.5972
R7844 VDD.n4252 VDD.n2393 28.5972
R7845 VDD.n4243 VDD.n2393 28.5972
R7846 VDD.n4243 VDD.n4242 28.5972
R7847 VDD.n4242 VDD.n4241 28.5972
R7848 VDD.n2412 VDD.n2411 28.5972
R7849 VDD.n4231 VDD.n2412 28.5972
R7850 VDD.n4231 VDD.n4230 28.5972
R7851 VDD.n4230 VDD.n4229 28.5972
R7852 VDD.n4229 VDD.n2413 28.5972
R7853 VDD.n4220 VDD.n2413 28.5972
R7854 VDD.n4219 VDD.n4218 28.5972
R7855 VDD.n4218 VDD.n2422 28.5972
R7856 VDD.n4209 VDD.n2422 28.5972
R7857 VDD.n4209 VDD.n4208 28.5972
R7858 VDD.n4208 VDD.n4207 28.5972
R7859 VDD.n4207 VDD.n2431 28.5972
R7860 VDD.n4198 VDD.n2431 28.5972
R7861 VDD.n4082 VDD.n2440 28.5972
R7862 VDD.n4094 VDD.n4082 28.5972
R7863 VDD.n4095 VDD.n4094 28.5972
R7864 VDD.n4096 VDD.n4095 28.5972
R7865 VDD.n4096 VDD.n4075 28.5972
R7866 VDD.n4107 VDD.n4075 28.5972
R7867 VDD.n4109 VDD.n4108 28.5972
R7868 VDD.n4109 VDD.n4068 28.5972
R7869 VDD.n4120 VDD.n4068 28.5972
R7870 VDD.n4121 VDD.n4120 28.5972
R7871 VDD.n4123 VDD.n4121 28.5972
R7872 VDD.n4123 VDD.n4122 28.5972
R7873 VDD.n4135 VDD.n4134 28.5972
R7874 VDD.n4136 VDD.n4135 28.5972
R7875 VDD.n4136 VDD.n4056 28.5972
R7876 VDD.n4146 VDD.n4056 28.5972
R7877 VDD.n4147 VDD.n4146 28.5972
R7878 VDD.n4148 VDD.n4048 28.5972
R7879 VDD.n4158 VDD.n4048 28.5972
R7880 VDD.n4159 VDD.n4158 28.5972
R7881 VDD.n4160 VDD.n4159 28.5972
R7882 VDD.n4160 VDD.n4041 28.5972
R7883 VDD.n4171 VDD.n4041 28.5972
R7884 VDD.n4172 VDD.n4171 28.5972
R7885 VDD.n4173 VDD.n4172 28.5972
R7886 VDD.n4184 VDD.n4034 28.5972
R7887 VDD.n4185 VDD.n4184 28.5972
R7888 VDD.n4187 VDD.n4185 28.5972
R7889 VDD.n4187 VDD.n4186 28.5972
R7890 VDD.n5459 VDD.n270 28.5972
R7891 VDD.n5442 VDD.n270 28.5972
R7892 VDD.n5443 VDD.n5442 28.5972
R7893 VDD.n4134 VDD.t52 28.1767
R7894 VDD.n4186 VDD.n245 28.1767
R7895 VDD.n5667 VDD.t89 28.1564
R7896 VDD.t36 VDD.n6505 28.1564
R7897 VDD.n7376 VDD.t18 28.1564
R7898 VDD.t73 VDD.n8214 28.1564
R7899 VDD.n8583 VDD.n8532 28.0793
R7900 VDD.n7728 VDD.n7677 28.0793
R7901 VDD.n6874 VDD.n6823 28.0793
R7902 VDD.n6019 VDD.n5968 28.0793
R7903 VDD.n8244 VDD.t155 27.6955
R7904 VDD.n8244 VDD.t157 27.6955
R7905 VDD.n8243 VDD.t27 27.6955
R7906 VDD.n8243 VDD.t29 27.6955
R7907 VDD.n7389 VDD.t33 27.6955
R7908 VDD.n7389 VDD.t35 27.6955
R7909 VDD.n7388 VDD.t150 27.6955
R7910 VDD.n7388 VDD.t152 27.6955
R7911 VDD.n6535 VDD.t1 27.6955
R7912 VDD.n6535 VDD.t3 27.6955
R7913 VDD.n6534 VDD.t130 27.6955
R7914 VDD.n6534 VDD.t133 27.6955
R7915 VDD.n5680 VDD.t11 27.6955
R7916 VDD.n5680 VDD.t13 27.6955
R7917 VDD.n5679 VDD.t62 27.6955
R7918 VDD.n5679 VDD.t59 27.6955
R7919 VDD.n8747 VDD.n8722 26.8524
R7920 VDD.n8747 VDD.n8721 26.8524
R7921 VDD.n8747 VDD.n8746 26.8524
R7922 VDD.n8854 VDD.n8853 26.8524
R7923 VDD.n8398 VDD.n8397 26.8524
R7924 VDD.n8308 VDD.n8278 26.8524
R7925 VDD.n8321 VDD.n8278 26.8524
R7926 VDD.n8307 VDD.n8278 26.8524
R7927 VDD.n7892 VDD.n7867 26.8524
R7928 VDD.n7892 VDD.n7866 26.8524
R7929 VDD.n7892 VDD.n7891 26.8524
R7930 VDD.n7999 VDD.n7998 26.8524
R7931 VDD.n7543 VDD.n7542 26.8524
R7932 VDD.n7453 VDD.n7423 26.8524
R7933 VDD.n7466 VDD.n7423 26.8524
R7934 VDD.n7452 VDD.n7423 26.8524
R7935 VDD.n7038 VDD.n7013 26.8524
R7936 VDD.n7038 VDD.n7012 26.8524
R7937 VDD.n7038 VDD.n7037 26.8524
R7938 VDD.n7145 VDD.n7144 26.8524
R7939 VDD.n6689 VDD.n6688 26.8524
R7940 VDD.n6599 VDD.n6569 26.8524
R7941 VDD.n6612 VDD.n6569 26.8524
R7942 VDD.n6598 VDD.n6569 26.8524
R7943 VDD.n6183 VDD.n6158 26.8524
R7944 VDD.n6183 VDD.n6157 26.8524
R7945 VDD.n6183 VDD.n6182 26.8524
R7946 VDD.n6290 VDD.n6289 26.8524
R7947 VDD.n5834 VDD.n5833 26.8524
R7948 VDD.n5744 VDD.n5714 26.8524
R7949 VDD.n5757 VDD.n5714 26.8524
R7950 VDD.n5743 VDD.n5714 26.8524
R7951 VDD.n8853 VDD.n8852 26.8521
R7952 VDD.n8853 VDD.n8687 26.8521
R7953 VDD.n8853 VDD.n8684 26.8521
R7954 VDD.n8853 VDD.n8685 26.8521
R7955 VDD.n8853 VDD.n8686 26.8521
R7956 VDD.n7998 VDD.n7997 26.8521
R7957 VDD.n7998 VDD.n7832 26.8521
R7958 VDD.n7998 VDD.n7829 26.8521
R7959 VDD.n7998 VDD.n7830 26.8521
R7960 VDD.n7998 VDD.n7831 26.8521
R7961 VDD.n7144 VDD.n7143 26.8521
R7962 VDD.n7144 VDD.n6978 26.8521
R7963 VDD.n7144 VDD.n6975 26.8521
R7964 VDD.n7144 VDD.n6976 26.8521
R7965 VDD.n7144 VDD.n6977 26.8521
R7966 VDD.n6289 VDD.n6288 26.8521
R7967 VDD.n6289 VDD.n6123 26.8521
R7968 VDD.n6289 VDD.n6120 26.8521
R7969 VDD.n6289 VDD.n6121 26.8521
R7970 VDD.n6289 VDD.n6122 26.8521
R7971 VDD.n3950 VDD.n2497 26.6499
R7972 VDD.n2502 VDD.n2497 26.6499
R7973 VDD.n3982 VDD.n2502 26.6499
R7974 VDD.n3982 VDD.n2503 26.6499
R7975 VDD.n3947 VDD.n2501 26.6499
R7976 VDD.n3952 VDD.n2501 26.6499
R7977 VDD.n3953 VDD.n2496 26.6499
R7978 VDD.n2620 VDD.n2606 26.6499
R7979 VDD.n2624 VDD.n2597 26.6499
R7980 VDD.n5474 VDD.n269 26.6499
R7981 VDD.n5472 VDD.n269 26.6499
R7982 VDD.n5472 VDD.n5460 26.6499
R7983 VDD.n5460 VDD.n250 26.6499
R7984 VDD.n5501 VDD.n5500 26.6499
R7985 VDD.n5503 VDD.n246 26.6499
R7986 VDD.n2448 VDD.n2446 26.6499
R7987 VDD.n4009 VDD.n2478 26.6499
R7988 VDD.n2481 VDD.n2478 26.6499
R7989 VDD.n2483 VDD.n2481 26.6499
R7990 VDD.n4007 VDD.n2483 26.6499
R7991 VDD.n3999 VDD.n2489 26.6499
R7992 VDD.n3995 VDD.n3993 26.6499
R7993 VDD.t40 VDD.n4219 26.4945
R7994 VDD.n8736 VDD.n8713 26.3534
R7995 VDD.n7881 VDD.n7858 26.3534
R7996 VDD.n7027 VDD.n7004 26.3534
R7997 VDD.n6172 VDD.n6149 26.3534
R7998 VDD.n2349 VDD.n2344 26.3534
R7999 VDD.n2650 VDD.n2639 26.3453
R8000 VDD.n3122 VDD.n3096 26.3453
R8001 VDD.n2991 VDD.n2951 26.3453
R8002 VDD.n97 VDD.n47 26.3453
R8003 VDD.n5555 VDD.n5548 26.3453
R8004 VDD.n196 VDD.n192 26.3453
R8005 VDD.n3497 VDD.n3496 26.3366
R8006 VDD.n3512 VDD.n3509 26.3366
R8007 VDD.n3199 VDD.n3198 26.3366
R8008 VDD.n3214 VDD.n3211 26.3366
R8009 VDD.n3747 VDD.n3746 26.3366
R8010 VDD.n3840 VDD.n3839 26.3366
R8011 VDD.n3843 VDD.n3840 26.3366
R8012 VDD.n3882 VDD.n3879 26.3366
R8013 VDD.n3866 VDD.n3862 26.3366
R8014 VDD.n3866 VDD.n3865 26.3366
R8015 VDD.n2826 VDD.n2823 26.3366
R8016 VDD.n2968 VDD.n2965 26.3366
R8017 VDD.n2352 VDD.n2348 25.9875
R8018 VDD.n8648 VDD.n8647 25.7394
R8019 VDD.n7793 VDD.n7792 25.7394
R8020 VDD.n6939 VDD.n6938 25.7394
R8021 VDD.n6084 VDD.n6083 25.7394
R8022 VDD.n8744 VDD.n8743 25.6005
R8023 VDD.n8743 VDD.n8742 25.6005
R8024 VDD.n8742 VDD.n8740 25.6005
R8025 VDD.n8740 VDD.n8737 25.6005
R8026 VDD.n8737 VDD.n8736 25.6005
R8027 VDD.n8967 VDD.n8966 25.6005
R8028 VDD.n8966 VDD.n8965 25.6005
R8029 VDD.n8965 VDD.n8417 25.6005
R8030 VDD.n8960 VDD.n8417 25.6005
R8031 VDD.n8902 VDD.n8901 25.6005
R8032 VDD.n8902 VDD.n8444 25.6005
R8033 VDD.n8908 VDD.n8444 25.6005
R8034 VDD.n8909 VDD.n8908 25.6005
R8035 VDD.n8910 VDD.n8909 25.6005
R8036 VDD.n8910 VDD.n8440 25.6005
R8037 VDD.n8916 VDD.n8440 25.6005
R8038 VDD.n8917 VDD.n8916 25.6005
R8039 VDD.n8918 VDD.n8917 25.6005
R8040 VDD.n8918 VDD.n8436 25.6005
R8041 VDD.n8924 VDD.n8436 25.6005
R8042 VDD.n8925 VDD.n8924 25.6005
R8043 VDD.n8926 VDD.n8925 25.6005
R8044 VDD.n8926 VDD.n8432 25.6005
R8045 VDD.n8932 VDD.n8432 25.6005
R8046 VDD.n8933 VDD.n8932 25.6005
R8047 VDD.n8934 VDD.n8933 25.6005
R8048 VDD.n8934 VDD.n8428 25.6005
R8049 VDD.n8940 VDD.n8428 25.6005
R8050 VDD.n8941 VDD.n8940 25.6005
R8051 VDD.n8942 VDD.n8941 25.6005
R8052 VDD.n8942 VDD.n8424 25.6005
R8053 VDD.n8948 VDD.n8424 25.6005
R8054 VDD.n8949 VDD.n8948 25.6005
R8055 VDD.n8950 VDD.n8949 25.6005
R8056 VDD.n8950 VDD.n8420 25.6005
R8057 VDD.n8958 VDD.n8420 25.6005
R8058 VDD.n8959 VDD.n8958 25.6005
R8059 VDD.n8894 VDD.n8892 25.6005
R8060 VDD.n8894 VDD.n8893 25.6005
R8061 VDD.n8893 VDD.n8448 25.6005
R8062 VDD.n8900 VDD.n8448 25.6005
R8063 VDD.n8358 VDD.n8342 25.6005
R8064 VDD.n8352 VDD.n8342 25.6005
R8065 VDD.n8352 VDD.n8351 25.6005
R8066 VDD.n8351 VDD.n8344 25.6005
R8067 VDD.n8345 VDD.n8344 25.6005
R8068 VDD.n8798 VDD.n8712 25.6005
R8069 VDD.n8804 VDD.n8798 25.6005
R8070 VDD.n8805 VDD.n8804 25.6005
R8071 VDD.n8805 VDD.n8796 25.6005
R8072 VDD.n8811 VDD.n8796 25.6005
R8073 VDD.n7889 VDD.n7888 25.6005
R8074 VDD.n7888 VDD.n7887 25.6005
R8075 VDD.n7887 VDD.n7885 25.6005
R8076 VDD.n7885 VDD.n7882 25.6005
R8077 VDD.n7882 VDD.n7881 25.6005
R8078 VDD.n8112 VDD.n8111 25.6005
R8079 VDD.n8111 VDD.n8110 25.6005
R8080 VDD.n8110 VDD.n7562 25.6005
R8081 VDD.n8105 VDD.n7562 25.6005
R8082 VDD.n8047 VDD.n8046 25.6005
R8083 VDD.n8047 VDD.n7589 25.6005
R8084 VDD.n8053 VDD.n7589 25.6005
R8085 VDD.n8054 VDD.n8053 25.6005
R8086 VDD.n8055 VDD.n8054 25.6005
R8087 VDD.n8055 VDD.n7585 25.6005
R8088 VDD.n8061 VDD.n7585 25.6005
R8089 VDD.n8062 VDD.n8061 25.6005
R8090 VDD.n8063 VDD.n8062 25.6005
R8091 VDD.n8063 VDD.n7581 25.6005
R8092 VDD.n8069 VDD.n7581 25.6005
R8093 VDD.n8070 VDD.n8069 25.6005
R8094 VDD.n8071 VDD.n8070 25.6005
R8095 VDD.n8071 VDD.n7577 25.6005
R8096 VDD.n8077 VDD.n7577 25.6005
R8097 VDD.n8078 VDD.n8077 25.6005
R8098 VDD.n8079 VDD.n8078 25.6005
R8099 VDD.n8079 VDD.n7573 25.6005
R8100 VDD.n8085 VDD.n7573 25.6005
R8101 VDD.n8086 VDD.n8085 25.6005
R8102 VDD.n8087 VDD.n8086 25.6005
R8103 VDD.n8087 VDD.n7569 25.6005
R8104 VDD.n8093 VDD.n7569 25.6005
R8105 VDD.n8094 VDD.n8093 25.6005
R8106 VDD.n8095 VDD.n8094 25.6005
R8107 VDD.n8095 VDD.n7565 25.6005
R8108 VDD.n8103 VDD.n7565 25.6005
R8109 VDD.n8104 VDD.n8103 25.6005
R8110 VDD.n8039 VDD.n8037 25.6005
R8111 VDD.n8039 VDD.n8038 25.6005
R8112 VDD.n8038 VDD.n7593 25.6005
R8113 VDD.n8045 VDD.n7593 25.6005
R8114 VDD.n7503 VDD.n7487 25.6005
R8115 VDD.n7497 VDD.n7487 25.6005
R8116 VDD.n7497 VDD.n7496 25.6005
R8117 VDD.n7496 VDD.n7489 25.6005
R8118 VDD.n7490 VDD.n7489 25.6005
R8119 VDD.n7943 VDD.n7857 25.6005
R8120 VDD.n7949 VDD.n7943 25.6005
R8121 VDD.n7950 VDD.n7949 25.6005
R8122 VDD.n7950 VDD.n7941 25.6005
R8123 VDD.n7956 VDD.n7941 25.6005
R8124 VDD.n7035 VDD.n7034 25.6005
R8125 VDD.n7034 VDD.n7033 25.6005
R8126 VDD.n7033 VDD.n7031 25.6005
R8127 VDD.n7031 VDD.n7028 25.6005
R8128 VDD.n7028 VDD.n7027 25.6005
R8129 VDD.n7258 VDD.n7257 25.6005
R8130 VDD.n7257 VDD.n7256 25.6005
R8131 VDD.n7256 VDD.n6708 25.6005
R8132 VDD.n7251 VDD.n6708 25.6005
R8133 VDD.n7193 VDD.n7192 25.6005
R8134 VDD.n7193 VDD.n6735 25.6005
R8135 VDD.n7199 VDD.n6735 25.6005
R8136 VDD.n7200 VDD.n7199 25.6005
R8137 VDD.n7201 VDD.n7200 25.6005
R8138 VDD.n7201 VDD.n6731 25.6005
R8139 VDD.n7207 VDD.n6731 25.6005
R8140 VDD.n7208 VDD.n7207 25.6005
R8141 VDD.n7209 VDD.n7208 25.6005
R8142 VDD.n7209 VDD.n6727 25.6005
R8143 VDD.n7215 VDD.n6727 25.6005
R8144 VDD.n7216 VDD.n7215 25.6005
R8145 VDD.n7217 VDD.n7216 25.6005
R8146 VDD.n7217 VDD.n6723 25.6005
R8147 VDD.n7223 VDD.n6723 25.6005
R8148 VDD.n7224 VDD.n7223 25.6005
R8149 VDD.n7225 VDD.n7224 25.6005
R8150 VDD.n7225 VDD.n6719 25.6005
R8151 VDD.n7231 VDD.n6719 25.6005
R8152 VDD.n7232 VDD.n7231 25.6005
R8153 VDD.n7233 VDD.n7232 25.6005
R8154 VDD.n7233 VDD.n6715 25.6005
R8155 VDD.n7239 VDD.n6715 25.6005
R8156 VDD.n7240 VDD.n7239 25.6005
R8157 VDD.n7241 VDD.n7240 25.6005
R8158 VDD.n7241 VDD.n6711 25.6005
R8159 VDD.n7249 VDD.n6711 25.6005
R8160 VDD.n7250 VDD.n7249 25.6005
R8161 VDD.n7185 VDD.n7183 25.6005
R8162 VDD.n7185 VDD.n7184 25.6005
R8163 VDD.n7184 VDD.n6739 25.6005
R8164 VDD.n7191 VDD.n6739 25.6005
R8165 VDD.n6649 VDD.n6633 25.6005
R8166 VDD.n6643 VDD.n6633 25.6005
R8167 VDD.n6643 VDD.n6642 25.6005
R8168 VDD.n6642 VDD.n6635 25.6005
R8169 VDD.n6636 VDD.n6635 25.6005
R8170 VDD.n7089 VDD.n7003 25.6005
R8171 VDD.n7095 VDD.n7089 25.6005
R8172 VDD.n7096 VDD.n7095 25.6005
R8173 VDD.n7096 VDD.n7087 25.6005
R8174 VDD.n7102 VDD.n7087 25.6005
R8175 VDD.n6180 VDD.n6179 25.6005
R8176 VDD.n6179 VDD.n6178 25.6005
R8177 VDD.n6178 VDD.n6176 25.6005
R8178 VDD.n6176 VDD.n6173 25.6005
R8179 VDD.n6173 VDD.n6172 25.6005
R8180 VDD.n6403 VDD.n6402 25.6005
R8181 VDD.n6402 VDD.n6401 25.6005
R8182 VDD.n6401 VDD.n5853 25.6005
R8183 VDD.n6396 VDD.n5853 25.6005
R8184 VDD.n6338 VDD.n6337 25.6005
R8185 VDD.n6338 VDD.n5880 25.6005
R8186 VDD.n6344 VDD.n5880 25.6005
R8187 VDD.n6345 VDD.n6344 25.6005
R8188 VDD.n6346 VDD.n6345 25.6005
R8189 VDD.n6346 VDD.n5876 25.6005
R8190 VDD.n6352 VDD.n5876 25.6005
R8191 VDD.n6353 VDD.n6352 25.6005
R8192 VDD.n6354 VDD.n6353 25.6005
R8193 VDD.n6354 VDD.n5872 25.6005
R8194 VDD.n6360 VDD.n5872 25.6005
R8195 VDD.n6361 VDD.n6360 25.6005
R8196 VDD.n6362 VDD.n6361 25.6005
R8197 VDD.n6362 VDD.n5868 25.6005
R8198 VDD.n6368 VDD.n5868 25.6005
R8199 VDD.n6369 VDD.n6368 25.6005
R8200 VDD.n6370 VDD.n6369 25.6005
R8201 VDD.n6370 VDD.n5864 25.6005
R8202 VDD.n6376 VDD.n5864 25.6005
R8203 VDD.n6377 VDD.n6376 25.6005
R8204 VDD.n6378 VDD.n6377 25.6005
R8205 VDD.n6378 VDD.n5860 25.6005
R8206 VDD.n6384 VDD.n5860 25.6005
R8207 VDD.n6385 VDD.n6384 25.6005
R8208 VDD.n6386 VDD.n6385 25.6005
R8209 VDD.n6386 VDD.n5856 25.6005
R8210 VDD.n6394 VDD.n5856 25.6005
R8211 VDD.n6395 VDD.n6394 25.6005
R8212 VDD.n6330 VDD.n6328 25.6005
R8213 VDD.n6330 VDD.n6329 25.6005
R8214 VDD.n6329 VDD.n5884 25.6005
R8215 VDD.n6336 VDD.n5884 25.6005
R8216 VDD.n5794 VDD.n5778 25.6005
R8217 VDD.n5788 VDD.n5778 25.6005
R8218 VDD.n5788 VDD.n5787 25.6005
R8219 VDD.n5787 VDD.n5780 25.6005
R8220 VDD.n5781 VDD.n5780 25.6005
R8221 VDD.n6234 VDD.n6148 25.6005
R8222 VDD.n6240 VDD.n6234 25.6005
R8223 VDD.n6241 VDD.n6240 25.6005
R8224 VDD.n6241 VDD.n6232 25.6005
R8225 VDD.n6247 VDD.n6232 25.6005
R8226 VDD.n1724 VDD.n1723 25.6005
R8227 VDD.n1723 VDD.n1720 25.6005
R8228 VDD.n1720 VDD.n1719 25.6005
R8229 VDD.n1719 VDD.n1716 25.6005
R8230 VDD.n1716 VDD.n1715 25.6005
R8231 VDD.n1715 VDD.n1712 25.6005
R8232 VDD.n1712 VDD.n1711 25.6005
R8233 VDD.n1711 VDD.n1708 25.6005
R8234 VDD.n1708 VDD.n1707 25.6005
R8235 VDD.n1707 VDD.n1035 25.6005
R8236 VDD.n1887 VDD.n1035 25.6005
R8237 VDD.n1888 VDD.n1887 25.6005
R8238 VDD.n1890 VDD.n1888 25.6005
R8239 VDD.n1890 VDD.n1889 25.6005
R8240 VDD.n1889 VDD.n1015 25.6005
R8241 VDD.n4568 VDD.n1015 25.6005
R8242 VDD.n4568 VDD.n4567 25.6005
R8243 VDD.n4567 VDD.n4566 25.6005
R8244 VDD.n4566 VDD.n1016 25.6005
R8245 VDD.n1919 VDD.n1016 25.6005
R8246 VDD.n4549 VDD.n1919 25.6005
R8247 VDD.n4549 VDD.n4548 25.6005
R8248 VDD.n4548 VDD.n4547 25.6005
R8249 VDD.n4547 VDD.n1920 25.6005
R8250 VDD.n1950 VDD.n1920 25.6005
R8251 VDD.n4530 VDD.n1950 25.6005
R8252 VDD.n4530 VDD.n4529 25.6005
R8253 VDD.n4529 VDD.n4528 25.6005
R8254 VDD.n4528 VDD.n1951 25.6005
R8255 VDD.n1988 VDD.n1951 25.6005
R8256 VDD.n1990 VDD.n1988 25.6005
R8257 VDD.n1991 VDD.n1990 25.6005
R8258 VDD.n4505 VDD.n1991 25.6005
R8259 VDD.n4505 VDD.n4504 25.6005
R8260 VDD.n4504 VDD.n4503 25.6005
R8261 VDD.n4503 VDD.n1992 25.6005
R8262 VDD.n2024 VDD.n1992 25.6005
R8263 VDD.n4486 VDD.n2024 25.6005
R8264 VDD.n4486 VDD.n4485 25.6005
R8265 VDD.n4485 VDD.n4484 25.6005
R8266 VDD.n4484 VDD.n2025 25.6005
R8267 VDD.n2054 VDD.n2025 25.6005
R8268 VDD.n4467 VDD.n2054 25.6005
R8269 VDD.n4467 VDD.n4466 25.6005
R8270 VDD.n4466 VDD.n4465 25.6005
R8271 VDD.n4465 VDD.n2055 25.6005
R8272 VDD.n4452 VDD.n2055 25.6005
R8273 VDD.n4452 VDD.n4451 25.6005
R8274 VDD.n4451 VDD.n4450 25.6005
R8275 VDD.n4450 VDD.n2072 25.6005
R8276 VDD.n2108 VDD.n2072 25.6005
R8277 VDD.n4433 VDD.n2108 25.6005
R8278 VDD.n4433 VDD.n4432 25.6005
R8279 VDD.n4432 VDD.n4431 25.6005
R8280 VDD.n4431 VDD.n2109 25.6005
R8281 VDD.n2139 VDD.n2109 25.6005
R8282 VDD.n4414 VDD.n2139 25.6005
R8283 VDD.n4414 VDD.n4413 25.6005
R8284 VDD.n4413 VDD.n4412 25.6005
R8285 VDD.n4412 VDD.n2140 25.6005
R8286 VDD.n2170 VDD.n2140 25.6005
R8287 VDD.n4395 VDD.n2170 25.6005
R8288 VDD.n4395 VDD.n4394 25.6005
R8289 VDD.n4394 VDD.n4393 25.6005
R8290 VDD.n4393 VDD.n2171 25.6005
R8291 VDD.n2209 VDD.n2171 25.6005
R8292 VDD.n2211 VDD.n2209 25.6005
R8293 VDD.n2212 VDD.n2211 25.6005
R8294 VDD.n4370 VDD.n2212 25.6005
R8295 VDD.n4370 VDD.n4369 25.6005
R8296 VDD.n4369 VDD.n4368 25.6005
R8297 VDD.n4368 VDD.n2213 25.6005
R8298 VDD.n8367 VDD.n8366 25.3507
R8299 VDD.n8863 VDD.n8862 25.3507
R8300 VDD.n8762 VDD.n8477 25.3507
R8301 VDD.n7512 VDD.n7511 25.3507
R8302 VDD.n8008 VDD.n8007 25.3507
R8303 VDD.n7907 VDD.n7622 25.3507
R8304 VDD.n6658 VDD.n6657 25.3507
R8305 VDD.n7154 VDD.n7153 25.3507
R8306 VDD.n7053 VDD.n6768 25.3507
R8307 VDD.n5803 VDD.n5802 25.3507
R8308 VDD.n6299 VDD.n6298 25.3507
R8309 VDD.n6198 VDD.n5913 25.3507
R8310 VDD.n1859 VDD.n1061 25.3507
R8311 VDD.n926 VDD.n925 25.3507
R8312 VDD.n1094 VDD.n1088 25.3507
R8313 VDD.n8637 VDD.n8504 25.3505
R8314 VDD.n8638 VDD.n8501 25.3505
R8315 VDD.n8841 VDD.n8480 25.3505
R8316 VDD.n8866 VDD.n8865 25.3505
R8317 VDD.n8998 VDD.n8997 25.3505
R8318 VDD.n8298 VDD.n8273 25.3505
R8319 VDD.n8337 VDD.n8336 25.3505
R8320 VDD.n7782 VDD.n7649 25.3505
R8321 VDD.n7783 VDD.n7646 25.3505
R8322 VDD.n7986 VDD.n7625 25.3505
R8323 VDD.n8011 VDD.n8010 25.3505
R8324 VDD.n8143 VDD.n8142 25.3505
R8325 VDD.n7443 VDD.n7418 25.3505
R8326 VDD.n7482 VDD.n7481 25.3505
R8327 VDD.n6928 VDD.n6795 25.3505
R8328 VDD.n6929 VDD.n6792 25.3505
R8329 VDD.n7132 VDD.n6771 25.3505
R8330 VDD.n7157 VDD.n7156 25.3505
R8331 VDD.n7289 VDD.n7288 25.3505
R8332 VDD.n6589 VDD.n6564 25.3505
R8333 VDD.n6628 VDD.n6627 25.3505
R8334 VDD.n6073 VDD.n5940 25.3505
R8335 VDD.n6074 VDD.n5937 25.3505
R8336 VDD.n6277 VDD.n5916 25.3505
R8337 VDD.n6302 VDD.n6301 25.3505
R8338 VDD.n6434 VDD.n6433 25.3505
R8339 VDD.n5734 VDD.n5709 25.3505
R8340 VDD.n5773 VDD.n5772 25.3505
R8341 VDD.n4019 VDD.n2233 25.3505
R8342 VDD.n2470 VDD.n2464 25.3505
R8343 VDD.n1818 VDD.n1087 25.3505
R8344 VDD.n1166 VDD.n1165 25.3505
R8345 VDD.n4720 VDD.n920 25.3505
R8346 VDD.n4276 VDD.t41 24.8124
R8347 VDD.n4016 VDD.n2471 23.9713
R8348 VDD.n5652 VDD.t92 23.5572
R8349 VDD.n6521 VDD.t39 23.5572
R8350 VDD.n7361 VDD.t21 23.5572
R8351 VDD.n8230 VDD.t76 23.5572
R8352 VDD.n2350 VDD.n2348 23.4711
R8353 VDD.n4028 VDD.n267 23.2949
R8354 VDD.n3990 VDD.n3989 23.2817
R8355 VDD.n3987 VDD.n3986 23.2817
R8356 VDD.n8720 VDD.n8709 23.0774
R8357 VDD.n8816 VDD.n8747 23.0774
R8358 VDD.n8389 VDD.n8267 23.0774
R8359 VDD.n7865 VDD.n7854 23.0774
R8360 VDD.n7961 VDD.n7892 23.0774
R8361 VDD.n7534 VDD.n7412 23.0774
R8362 VDD.n7011 VDD.n7000 23.0774
R8363 VDD.n7107 VDD.n7038 23.0774
R8364 VDD.n6680 VDD.n6558 23.0774
R8365 VDD.n6156 VDD.n6145 23.0774
R8366 VDD.n6252 VDD.n6183 23.0774
R8367 VDD.n5825 VDD.n5703 23.0774
R8368 VDD.n2656 VDD.n2649 23.0522
R8369 VDD.n3125 VDD.n3123 23.0522
R8370 VDD.n2992 VDD.n2915 23.0522
R8371 VDD.n89 VDD.n88 23.0522
R8372 VDD.n5593 VDD.n5530 23.0522
R8373 VDD.n234 VDD.n178 23.0522
R8374 VDD.n5449 VDD.n281 22.7097
R8375 VDD.t6 VDD.n4034 22.2891
R8376 VDD.n3809 VDD.n3808 22.1478
R8377 VDD.n2809 VDD.n2807 22.1478
R8378 VDD.n3023 VDD.n2889 22.1478
R8379 VDD.n3665 VDD.n3664 22.1478
R8380 VDD.n3690 VDD.n3671 22.1478
R8381 VDD.n8701 VDD.t24 21.7954
R8382 VDD.n8395 VDD.t25 21.7954
R8383 VDD.t25 VDD.n8286 21.7954
R8384 VDD.n7846 VDD.t32 21.7954
R8385 VDD.n7540 VDD.t153 21.7954
R8386 VDD.t153 VDD.n7431 21.7954
R8387 VDD.n6992 VDD.t0 21.7954
R8388 VDD.n6686 VDD.t131 21.7954
R8389 VDD.t131 VDD.n6577 21.7954
R8390 VDD.n6137 VDD.t10 21.7954
R8391 VDD.n5831 VDD.t60 21.7954
R8392 VDD.t60 VDD.n5722 21.7954
R8393 VDD.n5474 VDD.n267 21.468
R8394 VDD.t50 VDD.n4147 21.448
R8395 VDD.n123 VDD.n122 21.2396
R8396 VDD.n119 VDD.n118 21.1681
R8397 VDD.n5648 VDD.n5643 21.1346
R8398 VDD.n6510 VDD.n6506 21.1346
R8399 VDD.n7357 VDD.n7352 21.1346
R8400 VDD.n8219 VDD.n8215 21.1346
R8401 VDD.n1480 VDD.n1381 20.7186
R8402 VDD.n1480 VDD.n1382 20.7186
R8403 VDD.n1480 VDD.n1383 20.7186
R8404 VDD.n1480 VDD.n1384 20.7186
R8405 VDD.n1480 VDD.n1385 20.7186
R8406 VDD.n1480 VDD.n1479 20.7186
R8407 VDD.n1885 VDD.n1884 20.7183
R8408 VDD.n1884 VDD.n1042 20.7183
R8409 VDD.n1884 VDD.n1041 20.7183
R8410 VDD.n1884 VDD.n1040 20.7183
R8411 VDD.n1884 VDD.n1039 20.7183
R8412 VDD.n1884 VDD.n1038 20.7183
R8413 VDD.n4108 VDD.t48 20.607
R8414 VDD.n8967 VDD.n8413 20.6044
R8415 VDD.n8112 VDD.n7558 20.6044
R8416 VDD.n7258 VDD.n6704 20.6044
R8417 VDD.n6403 VDD.n5849 20.6044
R8418 VDD.n3498 VDD.n3493 20.5156
R8419 VDD.n3200 VDD.n3195 20.5156
R8420 VDD.n3748 VDD.n3743 20.5156
R8421 VDD.n3511 VDD.n3510 20.5153
R8422 VDD.n3213 VDD.n3212 20.5153
R8423 VDD.n3881 VDD.n3880 20.5153
R8424 VDD.n2828 VDD.n2827 20.5152
R8425 VDD.n2970 VDD.n2969 20.5152
R8426 VDD.n8823 VDD.n8709 20.5133
R8427 VDD.n8750 VDD.n8747 20.5133
R8428 VDD.n9005 VDD.n8267 20.5133
R8429 VDD.n7968 VDD.n7854 20.5133
R8430 VDD.n7895 VDD.n7892 20.5133
R8431 VDD.n8150 VDD.n7412 20.5133
R8432 VDD.n7114 VDD.n7000 20.5133
R8433 VDD.n7041 VDD.n7038 20.5133
R8434 VDD.n7296 VDD.n6558 20.5133
R8435 VDD.n6259 VDD.n6145 20.5133
R8436 VDD.n6186 VDD.n6183 20.5133
R8437 VDD.n6441 VDD.n5703 20.5133
R8438 VDD.n3845 VDD.n3737 19.9534
R8439 VDD.n3845 VDD.n3844 19.9534
R8440 VDD.n3867 VDD.n3709 19.9534
R8441 VDD.n3867 VDD.n3710 19.9534
R8442 VDD.n3990 VDD.n2491 19.9425
R8443 VDD.n3986 VDD.n2495 19.9425
R8444 VDD.n3555 VDD.n2676 19.7698
R8445 VDD.n3548 VDD.n2674 19.7698
R8446 VDD.n3257 VDD.n3082 19.7698
R8447 VDD.n3250 VDD.n3080 19.7698
R8448 VDD.n3610 VDD.n3609 19.7591
R8449 VDD.n3169 VDD.n3168 19.7591
R8450 VDD.n2986 VDD.n2956 19.7591
R8451 VDD.n3560 VDD.n2677 19.7549
R8452 VDD.n3543 VDD.n2673 19.7549
R8453 VDD.n3262 VDD.n3083 19.7549
R8454 VDD.n3245 VDD.n3079 19.7549
R8455 VDD.n3565 VDD.n2669 19.7383
R8456 VDD.n3538 VDD.n2672 19.7383
R8457 VDD.n3267 VDD.n3075 19.7383
R8458 VDD.n3240 VDD.n3078 19.7383
R8459 VDD.n3571 VDD.n2679 19.7199
R8460 VDD.n3533 VDD.n2671 19.7199
R8461 VDD.n3460 VDD.n2695 19.7199
R8462 VDD.n3440 VDD.n3438 19.7199
R8463 VDD.n2725 VDD.n2720 19.7199
R8464 VDD.n3407 VDD.n3403 19.7199
R8465 VDD.n3386 VDD.n3384 19.7199
R8466 VDD.n3366 VDD.n3352 19.7199
R8467 VDD.n3295 VDD.n3294 19.7199
R8468 VDD.n3273 VDD.n3085 19.7199
R8469 VDD.n3235 VDD.n3077 19.7199
R8470 VDD.n3817 VDD.n3759 19.7199
R8471 VDD.n3720 VDD.n3661 19.7199
R8472 VDD.n3903 VDD.n3675 19.7199
R8473 VDD.n2848 VDD.n2847 19.7199
R8474 VDD.n3580 VDD.n3579 19.6997
R8475 VDD.n3528 VDD.n2670 19.6997
R8476 VDD.n3468 VDD.n3467 19.6997
R8477 VDD.n3446 VDD.n3436 19.6997
R8478 VDD.n3428 VDD.n3427 19.6997
R8479 VDD.n3415 VDD.n3414 19.6997
R8480 VDD.n3392 VDD.n3382 19.6997
R8481 VDD.n3359 VDD.n3351 19.6997
R8482 VDD.n3287 VDD.n3072 19.6997
R8483 VDD.n3282 VDD.n3281 19.6997
R8484 VDD.n3230 VDD.n3076 19.6997
R8485 VDD.n3822 VDD.n3757 19.6997
R8486 VDD.n3725 VDD.n3666 19.6997
R8487 VDD.n3898 VDD.n3673 19.6997
R8488 VDD.n2842 VDD.n2810 19.6997
R8489 VDD.n3523 VDD.n2678 19.6777
R8490 VDD.n3225 VDD.n3084 19.6777
R8491 VDD.n3827 VDD.n3755 19.6777
R8492 VDD.n3730 VDD.n3667 19.6777
R8493 VDD.n3893 VDD.n3674 19.6777
R8494 VDD.n2837 VDD.n2811 19.6777
R8495 VDD.n2925 VDD.n2923 19.3601
R8496 VDD.n65 VDD.n64 19.3601
R8497 VDD.n5570 VDD.n5569 19.3601
R8498 VDD.n3582 VDD.n2667 19.3599
R8499 VDD.n3138 VDD.n3136 19.3599
R8500 VDD.n3791 VDD.n3764 19.3599
R8501 VDD.n211 VDD.n210 19.3599
R8502 VDD.n5497 VDD.n251 19.2933
R8503 VDD.n46 VDD.n43 19.131
R8504 VDD.n5547 VDD.n5546 19.131
R8505 VDD.n191 VDD.n188 19.131
R8506 VDD.n3503 VDD.n3502 19.0069
R8507 VDD.n3517 VDD.n3505 19.0069
R8508 VDD.n3205 VDD.n3204 19.0069
R8509 VDD.n3219 VDD.n3207 19.0069
R8510 VDD.n3753 VDD.n3752 19.0069
R8511 VDD.n3831 VDD.n3739 19.0069
R8512 VDD.n3851 VDD.n3850 19.0069
R8513 VDD.n3887 VDD.n3875 19.0069
R8514 VDD.n3854 VDD.n3712 19.0069
R8515 VDD.n3873 VDD.n3872 19.0069
R8516 VDD.n2833 VDD.n2832 19.0069
R8517 VDD.n2975 VDD.n2974 19.0069
R8518 VDD.n2888 VDD.n2887 18.986
R8519 VDD.n2411 VDD.t80 18.9248
R8520 VDD.n2981 VDD.n2980 18.9099
R8521 VDD.n8892 VDD.n8891 18.7439
R8522 VDD.n8037 VDD.n8036 18.7439
R8523 VDD.n7183 VDD.n7182 18.7439
R8524 VDD.n6328 VDD.n6327 18.7439
R8525 VDD.n5497 VDD.n5496 17.9019
R8526 VDD.n5652 VDD.t154 17.8272
R8527 VDD.n6521 VDD.t129 17.8272
R8528 VDD.n7361 VDD.t93 17.8272
R8529 VDD.n8230 VDD.t97 17.8272
R8530 VDD.n5285 VDD.n395 17.8254
R8531 VDD.n3937 VDD.n3936 17.6125
R8532 VDD.n2565 VDD.n2517 17.3826
R8533 VDD.n5658 VDD.n5644 17.2489
R8534 VDD.n6519 VDD.n6518 17.2489
R8535 VDD.n7367 VDD.n7353 17.2489
R8536 VDD.n8228 VDD.n8227 17.2489
R8537 VDD.n4025 VDD.n4023 17.2426
R8538 VDD.t79 VDD.n2384 17.2426
R8539 VDD.n2576 VDD.n2575 16.6542
R8540 VDD.n3597 VDD.n3596 16.466
R8541 VDD.n3153 VDD.n3152 16.466
R8542 VDD.n3938 VDD.n3642 16.466
R8543 VDD.n2999 VDD.n2914 16.466
R8544 VDD.n84 VDD.n50 16.466
R8545 VDD.n5591 VDD.n5531 16.466
R8546 VDD.n232 VDD.n179 16.466
R8547 VDD.n2579 VDD.n2578 15.9242
R8548 VDD.n8814 VDD.n8812 15.6165
R8549 VDD.n9013 VDD.n8256 15.6165
R8550 VDD.n7959 VDD.n7957 15.6165
R8551 VDD.n8158 VDD.n7401 15.6165
R8552 VDD.n7105 VDD.n7103 15.6165
R8553 VDD.n7304 VDD.n6547 15.6165
R8554 VDD.n6250 VDD.n6248 15.6165
R8555 VDD.n6449 VDD.n5692 15.6165
R8556 VDD.n5285 VDD.n5284 15.0799
R8557 VDD.n121 VDD.n28 15.056
R8558 VDD.n2611 VDD.n2610 14.8411
R8559 VDD.t24 VDD.n8695 14.7441
R8560 VDD.n8823 VDD.t156 14.7441
R8561 VDD.n8750 VDD.t72 14.7441
R8562 VDD.t26 VDD.n8252 14.7441
R8563 VDD.n8258 VDD.t26 14.7441
R8564 VDD.n9005 VDD.t28 14.7441
R8565 VDD.t32 VDD.n7840 14.7441
R8566 VDD.n7968 VDD.t34 14.7441
R8567 VDD.n7895 VDD.t85 14.7441
R8568 VDD.t86 VDD.n7397 14.7441
R8569 VDD.n7403 VDD.t86 14.7441
R8570 VDD.n8150 VDD.t151 14.7441
R8571 VDD.t0 VDD.n6986 14.7441
R8572 VDD.n7114 VDD.t2 14.7441
R8573 VDD.n7041 VDD.t87 14.7441
R8574 VDD.t88 VDD.n6543 14.7441
R8575 VDD.n6549 VDD.t88 14.7441
R8576 VDD.n7296 VDD.t132 14.7441
R8577 VDD.t10 VDD.n6131 14.7441
R8578 VDD.n6259 VDD.t12 14.7441
R8579 VDD.n6186 VDD.t139 14.7441
R8580 VDD.t61 VDD.n5688 14.7441
R8581 VDD.n5694 VDD.t61 14.7441
R8582 VDD.n6441 VDD.t58 14.7441
R8583 VDD.n131 VDD.n130 14.6773
R8584 VDD.n1480 VDD.n1380 14.2505
R8585 VDD.n8812 VDD.n8795 14.2085
R8586 VDD.n8392 VDD.n8256 14.2085
R8587 VDD.n7957 VDD.n7940 14.2085
R8588 VDD.n7537 VDD.n7401 14.2085
R8589 VDD.n7103 VDD.n7086 14.2085
R8590 VDD.n6683 VDD.n6547 14.2085
R8591 VDD.n6248 VDD.n6231 14.2085
R8592 VDD.n5828 VDD.n5692 14.2085
R8593 VDD.n8749 VDD.n8251 14.1031
R8594 VDD.n9017 VDD.n8252 14.1031
R8595 VDD.n8259 VDD.n8258 14.1031
R8596 VDD.n9011 VDD.n8260 14.1031
R8597 VDD.n7894 VDD.n7396 14.1031
R8598 VDD.n8162 VDD.n7397 14.1031
R8599 VDD.n7404 VDD.n7403 14.1031
R8600 VDD.n8156 VDD.n7405 14.1031
R8601 VDD.n7040 VDD.n6542 14.1031
R8602 VDD.n7308 VDD.n6543 14.1031
R8603 VDD.n6550 VDD.n6549 14.1031
R8604 VDD.n7302 VDD.n6551 14.1031
R8605 VDD.n6185 VDD.n5687 14.1031
R8606 VDD.n6453 VDD.n5688 14.1031
R8607 VDD.n5695 VDD.n5694 14.1031
R8608 VDD.n6447 VDD.n5696 14.1031
R8609 VDD.n4198 VDD.t67 13.8783
R8610 VDD.n268 VDD.n248 13.8783
R8611 VDD.n5473 VDD.n247 13.8783
R8612 VDD.n2684 VDD.n2638 13.5534
R8613 VDD.n2652 VDD.n2651 13.5534
R8614 VDD.n3600 VDD.n2646 13.5534
R8615 VDD.n3594 VDD.n3593 13.5534
R8616 VDD.n2663 VDD.n2661 13.5534
R8617 VDD.n3098 VDD.n3095 13.5534
R8618 VDD.n3162 VDD.n3104 13.5534
R8619 VDD.n3156 VDD.n3119 13.5534
R8620 VDD.n3150 VDD.n3149 13.5534
R8621 VDD.n3132 VDD.n3130 13.5534
R8622 VDD.n3811 VDD.n3763 13.5534
R8623 VDD.n3928 VDD.n3927 13.5534
R8624 VDD.n3909 VDD.n3676 13.5534
R8625 VDD.n3786 VDD.n3773 13.5534
R8626 VDD.n2859 VDD.n2858 13.5534
R8627 VDD.n2941 VDD.n2940 13.5534
R8628 VDD.n2997 VDD.n2916 13.5534
R8629 VDD.n2990 VDD.n2952 13.5534
R8630 VDD.n2985 VDD.n2957 13.5534
R8631 VDD.n95 VDD.n94 13.5534
R8632 VDD.n77 VDD.n53 13.5534
R8633 VDD.n71 VDD.n60 13.5534
R8634 VDD.n5553 VDD.n5552 13.5534
R8635 VDD.n5585 VDD.n5563 13.5534
R8636 VDD.n5579 VDD.n5578 13.5534
R8637 VDD.n194 VDD.n170 13.5534
R8638 VDD.n223 VDD.n181 13.5534
R8639 VDD.n217 VDD.n206 13.5534
R8640 VDD.n8395 VDD.n8388 13.462
R8641 VDD.n7540 VDD.n7533 13.462
R8642 VDD.n6686 VDD.n6679 13.462
R8643 VDD.n5831 VDD.n5824 13.462
R8644 VDD.n2455 VDD.n2443 13.3252
R8645 VDD.t54 VDD.n2440 13.0372
R8646 VDD.n3805 VDD.n3648 12.8005
R8647 VDD.n3925 VDD.n3917 12.8005
R8648 VDD.n3688 VDD.n3672 12.8005
R8649 VDD.n3780 VDD.n3779 12.8005
R8650 VDD.n2856 VDD.n2855 12.8005
R8651 VDD.n2878 VDD.n2875 12.8005
R8652 VDD.n2929 VDD.n2896 12.8005
R8653 VDD.n86 VDD.n35 12.8005
R8654 VDD.n5534 VDD.n5529 12.8005
R8655 VDD.n226 VDD.n177 12.8005
R8656 VDD.t68 VDD.n5618 12.789
R8657 VDD.n6488 VDD.t144 12.789
R8658 VDD.t14 VDD.n7327 12.789
R8659 VDD.n8197 VDD.t65 12.789
R8660 VDD.n3581 VDD.n2680 12.6901
R8661 VDD.n2694 VDD.n2691 12.6901
R8662 VDD.n3445 VDD.n3435 12.6901
R8663 VDD.n2714 VDD.n2711 12.6901
R8664 VDD.n3416 VDD.n3404 12.6901
R8665 VDD.n3391 VDD.n3381 12.6901
R8666 VDD.n3283 VDD.n3086 12.6901
R8667 VDD.n1884 VDD.n1883 12.6672
R8668 VDD.n3360 VDD.n3354 12.2367
R8669 VDD.n3288 VDD.n3074 12.2367
R8670 VDD.n2353 VDD.n2352 12.1342
R8671 VDD.n5164 VDD.n5163 12.064
R8672 VDD.n8790 VDD.n8466 12.0325
R8673 VDD.n8403 VDD.n8402 12.0325
R8674 VDD.n7935 VDD.n7611 12.0325
R8675 VDD.n7548 VDD.n7547 12.0325
R8676 VDD.n7081 VDD.n6757 12.0325
R8677 VDD.n6694 VDD.n6693 12.0325
R8678 VDD.n6226 VDD.n5902 12.0325
R8679 VDD.n5839 VDD.n5838 12.0325
R8680 VDD.n4016 VDD.t142 11.8979
R8681 VDD.n4005 VDD.n4004 11.7802
R8682 VDD.n3945 VDD.n2506 11.7802
R8683 VDD.n2537 VDD.n2518 11.6711
R8684 VDD.n4012 VDD.n4011 11.5947
R8685 VDD.n4025 VDD.n2367 11.3551
R8686 VDD.n4254 VDD.t79 11.3551
R8687 VDD.n2346 VDD.n2345 11.1178
R8688 VDD.n2480 VDD.n2479 10.8935
R8689 VDD.n4008 VDD.n2482 10.8935
R8690 VDD.n8731 VDD.n8706 10.4112
R8691 VDD.n8731 VDD.n8730 10.4112
R8692 VDD.n7876 VDD.n7851 10.4112
R8693 VDD.n7876 VDD.n7875 10.4112
R8694 VDD.n7022 VDD.n6997 10.4112
R8695 VDD.n7022 VDD.n7021 10.4112
R8696 VDD.n6167 VDD.n6142 10.4112
R8697 VDD.n6167 VDD.n6166 10.4112
R8698 VDD.n3587 VDD.n2658 9.87981
R8699 VDD.n3143 VDD.n3127 9.87981
R8700 VDD.n3782 VDD.n3768 9.87981
R8701 VDD.n2938 VDD.n2931 9.87981
R8702 VDD.n75 VDD.n54 9.87981
R8703 VDD.n5582 VDD.n5581 9.87981
R8704 VDD.n221 VDD.n182 9.87981
R8705 VDD.n4241 VDD.t80 9.67292
R8706 VDD.n5443 VDD.n281 9.67292
R8707 VDD.n2666 VDD.n2664 9.3005
R8708 VDD.n3591 VDD.n2659 9.3005
R8709 VDD.n3601 VDD.n3600 9.3005
R8710 VDD.n3584 VDD.n3583 9.3005
R8711 VDD.n3585 VDD.n3584 9.3005
R8712 VDD.n2663 VDD.n2660 9.3005
R8713 VDD.n3590 VDD.n3589 9.3005
R8714 VDD.n3589 VDD.n2658 9.3005
R8715 VDD.n3593 VDD.n3592 9.3005
R8716 VDD.n3598 VDD.n2648 9.3005
R8717 VDD.n3598 VDD.n3597 9.3005
R8718 VDD.n3599 VDD.n2645 9.3005
R8719 VDD.n2685 VDD.n2684 9.3005
R8720 VDD.n3607 VDD.n3606 9.3005
R8721 VDD.n3608 VDD.n3607 9.3005
R8722 VDD.n2652 VDD.n2643 9.3005
R8723 VDD.n2654 VDD.n2644 9.3005
R8724 VDD.n2654 VDD.n2649 9.3005
R8725 VDD.n3613 VDD.n3612 9.3005
R8726 VDD.n3516 VDD.n3506 9.3005
R8727 VDD.n3518 VDD.n3517 9.3005
R8728 VDD.n3515 VDD.n3508 9.3005
R8729 VDD.n3515 VDD.n3514 9.3005
R8730 VDD.n3502 VDD.n3490 9.3005
R8731 VDD.n3501 VDD.n3500 9.3005
R8732 VDD.n3499 VDD.n3492 9.3005
R8733 VDD.n3492 VDD.n3491 9.3005
R8734 VDD.n3524 VDD.n3489 9.3005
R8735 VDD.n3529 VDD.n3488 9.3005
R8736 VDD.n3534 VDD.n3487 9.3005
R8737 VDD.n3539 VDD.n3486 9.3005
R8738 VDD.n3544 VDD.n3485 9.3005
R8739 VDD.n3549 VDD.n3484 9.3005
R8740 VDD.n3554 VDD.n3483 9.3005
R8741 VDD.n3559 VDD.n3482 9.3005
R8742 VDD.n3564 VDD.n3481 9.3005
R8743 VDD.n3566 VDD.n3565 9.3005
R8744 VDD.n3563 VDD.n3562 9.3005
R8745 VDD.n3561 VDD.n3560 9.3005
R8746 VDD.n3558 VDD.n3557 9.3005
R8747 VDD.n3556 VDD.n3555 9.3005
R8748 VDD.n3553 VDD.n3552 9.3005
R8749 VDD.n3551 VDD.n3550 9.3005
R8750 VDD.n3548 VDD.n3547 9.3005
R8751 VDD.n3546 VDD.n3545 9.3005
R8752 VDD.n3543 VDD.n3542 9.3005
R8753 VDD.n3541 VDD.n3540 9.3005
R8754 VDD.n3538 VDD.n3537 9.3005
R8755 VDD.n3536 VDD.n3535 9.3005
R8756 VDD.n3533 VDD.n3532 9.3005
R8757 VDD.n3531 VDD.n3530 9.3005
R8758 VDD.n3528 VDD.n3527 9.3005
R8759 VDD.n3526 VDD.n3525 9.3005
R8760 VDD.n3523 VDD.n3522 9.3005
R8761 VDD.n3579 VDD.n3578 9.3005
R8762 VDD.n3575 VDD.n3574 9.3005
R8763 VDD.n3572 VDD.n3571 9.3005
R8764 VDD.n3568 VDD.n3479 9.3005
R8765 VDD.n3474 VDD.n2681 9.3005
R8766 VDD.n3467 VDD.n3466 9.3005
R8767 VDD.n3464 VDD.n3463 9.3005
R8768 VDD.n3457 VDD.n2699 9.3005
R8769 VDD.n3461 VDD.n3460 9.3005
R8770 VDD.n3470 VDD.n3469 9.3005
R8771 VDD.n3443 VDD.n3442 9.3005
R8772 VDD.n3440 VDD.n3439 9.3005
R8773 VDD.n3437 VDD.n2705 9.3005
R8774 VDD.n3436 VDD.n2702 9.3005
R8775 VDD.n3448 VDD.n3447 9.3005
R8776 VDD.n3427 VDD.n3426 9.3005
R8777 VDD.n2719 VDD.n2716 9.3005
R8778 VDD.n2726 VDD.n2725 9.3005
R8779 VDD.n2723 VDD.n2722 9.3005
R8780 VDD.n3430 VDD.n3429 9.3005
R8781 VDD.n3414 VDD.n2732 9.3005
R8782 VDD.n3419 VDD.n3418 9.3005
R8783 VDD.n3408 VDD.n3407 9.3005
R8784 VDD.n3406 VDD.n3405 9.3005
R8785 VDD.n3413 VDD.n3412 9.3005
R8786 VDD.n3389 VDD.n3388 9.3005
R8787 VDD.n3386 VDD.n3385 9.3005
R8788 VDD.n3383 VDD.n2741 9.3005
R8789 VDD.n3382 VDD.n2738 9.3005
R8790 VDD.n3394 VDD.n3393 9.3005
R8791 VDD.n3351 VDD.n3328 9.3005
R8792 VDD.n3370 VDD.n3369 9.3005
R8793 VDD.n3367 VDD.n3366 9.3005
R8794 VDD.n3364 VDD.n3363 9.3005
R8795 VDD.n3358 VDD.n3357 9.3005
R8796 VDD.n3072 VDD.n3071 9.3005
R8797 VDD.n3297 VDD.n3296 9.3005
R8798 VDD.n3294 VDD.n3066 9.3005
R8799 VDD.n3292 VDD.n3291 9.3005
R8800 VDD.n3286 VDD.n3285 9.3005
R8801 VDD.n3218 VDD.n3208 9.3005
R8802 VDD.n3220 VDD.n3219 9.3005
R8803 VDD.n3217 VDD.n3210 9.3005
R8804 VDD.n3217 VDD.n3216 9.3005
R8805 VDD.n3204 VDD.n3192 9.3005
R8806 VDD.n3203 VDD.n3202 9.3005
R8807 VDD.n3201 VDD.n3194 9.3005
R8808 VDD.n3194 VDD.n3193 9.3005
R8809 VDD.n3226 VDD.n3191 9.3005
R8810 VDD.n3231 VDD.n3190 9.3005
R8811 VDD.n3236 VDD.n3189 9.3005
R8812 VDD.n3241 VDD.n3188 9.3005
R8813 VDD.n3246 VDD.n3187 9.3005
R8814 VDD.n3251 VDD.n3186 9.3005
R8815 VDD.n3256 VDD.n3185 9.3005
R8816 VDD.n3261 VDD.n3184 9.3005
R8817 VDD.n3266 VDD.n3183 9.3005
R8818 VDD.n3268 VDD.n3267 9.3005
R8819 VDD.n3265 VDD.n3264 9.3005
R8820 VDD.n3263 VDD.n3262 9.3005
R8821 VDD.n3260 VDD.n3259 9.3005
R8822 VDD.n3258 VDD.n3257 9.3005
R8823 VDD.n3255 VDD.n3254 9.3005
R8824 VDD.n3253 VDD.n3252 9.3005
R8825 VDD.n3250 VDD.n3249 9.3005
R8826 VDD.n3248 VDD.n3247 9.3005
R8827 VDD.n3245 VDD.n3244 9.3005
R8828 VDD.n3243 VDD.n3242 9.3005
R8829 VDD.n3240 VDD.n3239 9.3005
R8830 VDD.n3238 VDD.n3237 9.3005
R8831 VDD.n3235 VDD.n3234 9.3005
R8832 VDD.n3233 VDD.n3232 9.3005
R8833 VDD.n3230 VDD.n3229 9.3005
R8834 VDD.n3228 VDD.n3227 9.3005
R8835 VDD.n3225 VDD.n3224 9.3005
R8836 VDD.n3281 VDD.n3280 9.3005
R8837 VDD.n3277 VDD.n3276 9.3005
R8838 VDD.n3274 VDD.n3273 9.3005
R8839 VDD.n3270 VDD.n3181 9.3005
R8840 VDD.n3176 VDD.n3087 9.3005
R8841 VDD.n3155 VDD.n3118 9.3005
R8842 VDD.n3147 VDD.n3128 9.3005
R8843 VDD.n3135 VDD.n3133 9.3005
R8844 VDD.n3140 VDD.n3139 9.3005
R8845 VDD.n3141 VDD.n3140 9.3005
R8846 VDD.n3132 VDD.n3129 9.3005
R8847 VDD.n3146 VDD.n3145 9.3005
R8848 VDD.n3145 VDD.n3127 9.3005
R8849 VDD.n3149 VDD.n3148 9.3005
R8850 VDD.n3154 VDD.n3121 9.3005
R8851 VDD.n3154 VDD.n3153 9.3005
R8852 VDD.n3157 VDD.n3156 9.3005
R8853 VDD.n3098 VDD.n3097 9.3005
R8854 VDD.n3166 VDD.n3165 9.3005
R8855 VDD.n3167 VDD.n3166 9.3005
R8856 VDD.n3159 VDD.n3105 9.3005
R8857 VDD.n3123 VDD.n3105 9.3005
R8858 VDD.n3163 VDD.n3162 9.3005
R8859 VDD.n3172 VDD.n3171 9.3005
R8860 VDD.n3658 VDD.n3655 9.3005
R8861 VDD.n3914 VDD.n3911 9.3005
R8862 VDD.n3913 VDD.n3912 9.3005
R8863 VDD.n3916 VDD.n3915 9.3005
R8864 VDD.n3922 VDD.n3921 9.3005
R8865 VDD.n3719 VDD.n3715 9.3005
R8866 VDD.n3724 VDD.n3714 9.3005
R8867 VDD.n3729 VDD.n3713 9.3005
R8868 VDD.n3731 VDD.n3730 9.3005
R8869 VDD.n3728 VDD.n3727 9.3005
R8870 VDD.n3726 VDD.n3725 9.3005
R8871 VDD.n3723 VDD.n3722 9.3005
R8872 VDD.n3721 VDD.n3720 9.3005
R8873 VDD.n3718 VDD.n3717 9.3005
R8874 VDD.n3682 VDD.n3681 9.3005
R8875 VDD.n3693 VDD.n3691 9.3005
R8876 VDD.n3692 VDD.n3687 9.3005
R8877 VDD.n3695 VDD.n3694 9.3005
R8878 VDD.n3684 VDD.n3683 9.3005
R8879 VDD.n3904 VDD.n3702 9.3005
R8880 VDD.n3903 VDD.n3902 9.3005
R8881 VDD.n3894 VDD.n3704 9.3005
R8882 VDD.n3901 VDD.n3900 9.3005
R8883 VDD.n3896 VDD.n3895 9.3005
R8884 VDD.n3893 VDD.n3892 9.3005
R8885 VDD.n3898 VDD.n3897 9.3005
R8886 VDD.n3899 VDD.n3703 9.3005
R8887 VDD.n3906 VDD.n3905 9.3005
R8888 VDD.n3858 VDD.n3857 9.3005
R8889 VDD.n3871 VDD.n3870 9.3005
R8890 VDD.n3856 VDD.n3712 9.3005
R8891 VDD.n3859 VDD.n3708 9.3005
R8892 VDD.n3859 VDD.n3711 9.3005
R8893 VDD.n3869 VDD.n3707 9.3005
R8894 VDD.n3707 VDD.n3706 9.3005
R8895 VDD.n3872 VDD.n3705 9.3005
R8896 VDD.n3886 VDD.n3876 9.3005
R8897 VDD.n3888 VDD.n3887 9.3005
R8898 VDD.n3885 VDD.n3878 9.3005
R8899 VDD.n3885 VDD.n3884 9.3005
R8900 VDD.n3850 VDD.n3733 9.3005
R8901 VDD.n3833 VDD.n3739 9.3005
R8902 VDD.n3752 VDD.n3740 9.3005
R8903 VDD.n3751 VDD.n3750 9.3005
R8904 VDD.n3749 VDD.n3742 9.3005
R8905 VDD.n3742 VDD.n3741 9.3005
R8906 VDD.n3835 VDD.n3834 9.3005
R8907 VDD.n3836 VDD.n3736 9.3005
R8908 VDD.n3836 VDD.n3738 9.3005
R8909 VDD.n3849 VDD.n3848 9.3005
R8910 VDD.n3847 VDD.n3735 9.3005
R8911 VDD.n3735 VDD.n3734 9.3005
R8912 VDD.n3826 VDD.n3756 9.3005
R8913 VDD.n3821 VDD.n3758 9.3005
R8914 VDD.n3816 VDD.n3760 9.3005
R8915 VDD.n3828 VDD.n3827 9.3005
R8916 VDD.n3825 VDD.n3824 9.3005
R8917 VDD.n3823 VDD.n3822 9.3005
R8918 VDD.n3820 VDD.n3819 9.3005
R8919 VDD.n3818 VDD.n3817 9.3005
R8920 VDD.n3815 VDD.n3814 9.3005
R8921 VDD.n3795 VDD.n3794 9.3005
R8922 VDD.n3793 VDD.n3647 9.3005
R8923 VDD.n3802 VDD.n3801 9.3005
R8924 VDD.n3800 VDD.n3799 9.3005
R8925 VDD.n3797 VDD.n3796 9.3005
R8926 VDD.n3769 VDD.n3766 9.3005
R8927 VDD.n3773 VDD.n3772 9.3005
R8928 VDD.n3789 VDD.n3767 9.3005
R8929 VDD.n3789 VDD.n3788 9.3005
R8930 VDD.n3776 VDD.n3774 9.3005
R8931 VDD.n3778 VDD.n3777 9.3005
R8932 VDD.n3641 VDD.n3639 9.3005
R8933 VDD.n3940 VDD.n3939 9.3005
R8934 VDD.n3939 VDD.n3938 9.3005
R8935 VDD.n3783 VDD.n3775 9.3005
R8936 VDD.n3783 VDD.n3782 9.3005
R8937 VDD.n2831 VDD.n2830 9.3005
R8938 VDD.n2829 VDD.n2822 9.3005
R8939 VDD.n2822 VDD.n2821 9.3005
R8940 VDD.n2832 VDD.n2820 9.3005
R8941 VDD.n2818 VDD.n2813 9.3005
R8942 VDD.n2847 VDD.n2846 9.3005
R8943 VDD.n2838 VDD.n2819 9.3005
R8944 VDD.n2845 VDD.n2812 9.3005
R8945 VDD.n2840 VDD.n2839 9.3005
R8946 VDD.n2837 VDD.n2836 9.3005
R8947 VDD.n2842 VDD.n2841 9.3005
R8948 VDD.n2844 VDD.n2843 9.3005
R8949 VDD.n2817 VDD.n2816 9.3005
R8950 VDD.n2860 VDD.n2802 9.3005
R8951 VDD.n2852 VDD.n2849 9.3005
R8952 VDD.n2851 VDD.n2850 9.3005
R8953 VDD.n2854 VDD.n2853 9.3005
R8954 VDD.n2862 VDD.n2861 9.3005
R8955 VDD.n2881 VDD.n2877 9.3005
R8956 VDD.n2880 VDD.n2879 9.3005
R8957 VDD.n2886 VDD.n2885 9.3005
R8958 VDD.n2876 VDD.n2874 9.3005
R8959 VDD.n2883 VDD.n2882 9.3005
R8960 VDD.n2919 VDD.n2918 9.3005
R8961 VDD.n2927 VDD.n2926 9.3005
R8962 VDD.n2928 VDD.n2927 9.3005
R8963 VDD.n2942 VDD.n2941 9.3005
R8964 VDD.n2973 VDD.n2972 9.3005
R8965 VDD.n2971 VDD.n2964 9.3005
R8966 VDD.n2964 VDD.n2963 9.3005
R8967 VDD.n2974 VDD.n2962 9.3005
R8968 VDD.n2978 VDD.n2958 9.3005
R8969 VDD.n2959 VDD.n2953 9.3005
R8970 VDD.n2950 VDD.n2949 9.3005
R8971 VDD.n2954 VDD.n2952 9.3005
R8972 VDD.n2988 VDD.n2955 9.3005
R8973 VDD.n2988 VDD.n2987 9.3005
R8974 VDD.n2960 VDD.n2957 9.3005
R8975 VDD.n2983 VDD.n2961 9.3005
R8976 VDD.n2983 VDD.n2982 9.3005
R8977 VDD.n2980 VDD.n2979 9.3005
R8978 VDD.n2994 VDD.n2993 9.3005
R8979 VDD.n2993 VDD.n2992 9.3005
R8980 VDD.n2913 VDD.n2911 9.3005
R8981 VDD.n2934 VDD.n2933 9.3005
R8982 VDD.n2936 VDD.n2935 9.3005
R8983 VDD.n2936 VDD.n2931 9.3005
R8984 VDD.n2932 VDD.n2895 9.3005
R8985 VDD.n3001 VDD.n3000 9.3005
R8986 VDD.n3000 VDD.n2999 9.3005
R8987 VDD.n70 VDD.n59 9.3005
R8988 VDD.n69 VDD.n62 9.3005
R8989 VDD.n69 VDD.n68 9.3005
R8990 VDD.n72 VDD.n71 9.3005
R8991 VDD.n74 VDD.n73 9.3005
R8992 VDD.n75 VDD.n74 9.3005
R8993 VDD.n58 VDD.n55 9.3005
R8994 VDD.n51 VDD.n36 9.3005
R8995 VDD.n45 VDD.n44 9.3005
R8996 VDD.n93 VDD.n92 9.3005
R8997 VDD.n43 VDD.n41 9.3005
R8998 VDD.n91 VDD.n90 9.3005
R8999 VDD.n90 VDD.n89 9.3005
R9000 VDD.n99 VDD.n42 9.3005
R9001 VDD.n99 VDD.n98 9.3005
R9002 VDD.n57 VDD.n53 9.3005
R9003 VDD.n83 VDD.n82 9.3005
R9004 VDD.n84 VDD.n83 9.3005
R9005 VDD.n80 VDD.n52 9.3005
R9006 VDD.n114 VDD.n29 9.3005
R9007 VDD.n127 VDD.n125 9.3005
R9008 VDD.n113 VDD.n112 9.3005
R9009 VDD.n118 VDD.n110 9.3005
R9010 VDD.n134 VDD.n133 9.3005
R9011 VDD.n133 VDD.n132 9.3005
R9012 VDD.n126 VDD.n117 9.3005
R9013 VDD.n132 VDD.n117 9.3005
R9014 VDD.n129 VDD.n128 9.3005
R9015 VDD.n116 VDD.n115 9.3005
R9016 VDD.n132 VDD.n116 9.3005
R9017 VDD.n5576 VDD.n5568 9.3005
R9018 VDD.n5575 VDD.n5574 9.3005
R9019 VDD.n5574 VDD.n5567 9.3005
R9020 VDD.n5578 VDD.n5577 9.3005
R9021 VDD.n5583 VDD.n5565 9.3005
R9022 VDD.n5583 VDD.n5582 9.3005
R9023 VDD.n5584 VDD.n5561 9.3005
R9024 VDD.n5536 VDD.n5535 9.3005
R9025 VDD.n5545 VDD.n5544 9.3005
R9026 VDD.n5551 VDD.n5550 9.3005
R9027 VDD.n5546 VDD.n5542 9.3005
R9028 VDD.n5528 VDD.n164 9.3005
R9029 VDD.n5530 VDD.n5528 9.3005
R9030 VDD.n5558 VDD.n5557 9.3005
R9031 VDD.n5557 VDD.n5556 9.3005
R9032 VDD.n5586 VDD.n5585 9.3005
R9033 VDD.n5590 VDD.n5589 9.3005
R9034 VDD.n5591 VDD.n5590 9.3005
R9035 VDD.n5537 VDD.n5532 9.3005
R9036 VDD.n204 VDD.n183 9.3005
R9037 VDD.n216 VDD.n205 9.3005
R9038 VDD.n220 VDD.n219 9.3005
R9039 VDD.n221 VDD.n220 9.3005
R9040 VDD.n215 VDD.n208 9.3005
R9041 VDD.n215 VDD.n214 9.3005
R9042 VDD.n218 VDD.n217 9.3005
R9043 VDD.n229 VDD.n180 9.3005
R9044 VDD.n175 VDD.n171 9.3005
R9045 VDD.n203 VDD.n181 9.3005
R9046 VDD.n190 VDD.n189 9.3005
R9047 VDD.n188 VDD.n186 9.3005
R9048 VDD.n198 VDD.n187 9.3005
R9049 VDD.n198 VDD.n197 9.3005
R9050 VDD.n176 VDD.n173 9.3005
R9051 VDD.n178 VDD.n176 9.3005
R9052 VDD.n231 VDD.n230 9.3005
R9053 VDD.n232 VDD.n231 9.3005
R9054 VDD.n228 VDD.n227 9.3005
R9055 VDD.n5496 VDD.n5495 9.3005
R9056 VDD.n5473 VDD.n250 9.3005
R9057 VDD.n5474 VDD.n5473 9.3005
R9058 VDD.n5473 VDD.n5472 9.3005
R9059 VDD.n5494 VDD.n249 9.3005
R9060 VDD.n4008 VDD.n4007 9.3005
R9061 VDD.n4008 VDD.n2481 9.3005
R9062 VDD.n4009 VDD.n4008 9.3005
R9063 VDD.n3983 VDD.n2496 9.3005
R9064 VDD.n3950 VDD.n2015 9.3005
R9065 VDD.n2503 VDD.n2015 9.3005
R9066 VDD.n2502 VDD.n2015 9.3005
R9067 VDD.n2581 VDD.n2511 9.3005
R9068 VDD.n2586 VDD.n2585 9.3005
R9069 VDD.n2529 VDD.n2528 9.3005
R9070 VDD.n2526 VDD.n2515 9.3005
R9071 VDD.n2568 VDD.n2567 9.3005
R9072 VDD.n2566 VDD.n2533 9.3005
R9073 VDD.n2557 VDD.n2536 9.3005
R9074 VDD.n2559 VDD.n2558 9.3005
R9075 VDD.n2556 VDD.n2555 9.3005
R9076 VDD.n2547 VDD.n2546 9.3005
R9077 VDD.n2544 VDD.n2540 9.3005
R9078 VDD.n2543 VDD.n2542 9.3005
R9079 VDD.n2521 VDD.n2520 9.3005
R9080 VDD.n2583 VDD.n2582 9.3005
R9081 VDD.n3926 VDD.n3663 9.1381
R9082 VDD.n3910 VDD.n3670 9.1381
R9083 VDD.n3810 VDD.n3798 9.1381
R9084 VDD.n2857 VDD.n2805 9.1381
R9085 VDD.n3024 VDD.n2884 9.1381
R9086 VDD.n3926 VDD.n3662 9.12656
R9087 VDD.n3910 VDD.n3669 9.12656
R9088 VDD.n3810 VDD.n3803 9.12656
R9089 VDD.n2857 VDD.n2803 9.12656
R9090 VDD.n3025 VDD.n3024 9.12656
R9091 VDD.n3926 VDD.n3660 9.11505
R9092 VDD.n3910 VDD.n3668 9.11505
R9093 VDD.n3810 VDD.n3761 9.11505
R9094 VDD.n2857 VDD.n2806 9.11505
R9095 VDD.n2456 VDD.n2455 9.01711
R9096 VDD.n4017 VDD.n2235 8.99396
R9097 VDD.n8860 VDD.n8678 8.9605
R9098 VDD.n9002 VDD.n9001 8.9605
R9099 VDD.n8005 VDD.n7823 8.9605
R9100 VDD.n8147 VDD.n8146 8.9605
R9101 VDD.n7151 VDD.n6969 8.9605
R9102 VDD.n7293 VDD.n7292 8.9605
R9103 VDD.n6296 VDD.n6114 8.9605
R9104 VDD.n6438 VDD.n6437 8.9605
R9105 VDD.n3581 VDD.n2676 8.90247
R9106 VDD.n3581 VDD.n2674 8.90247
R9107 VDD.n3283 VDD.n3082 8.90247
R9108 VDD.n3283 VDD.n3080 8.90247
R9109 VDD.n3581 VDD.n2677 8.89163
R9110 VDD.n3581 VDD.n2673 8.89163
R9111 VDD.n3283 VDD.n3083 8.89163
R9112 VDD.n3283 VDD.n3079 8.89163
R9113 VDD.n3581 VDD.n2672 8.88085
R9114 VDD.n3581 VDD.n2669 8.88085
R9115 VDD.n3283 VDD.n3078 8.88085
R9116 VDD.n3283 VDD.n3075 8.88085
R9117 VDD.n3581 VDD.n2679 8.87012
R9118 VDD.n3581 VDD.n2671 8.87012
R9119 VDD.n2695 VDD.n2694 8.87012
R9120 VDD.n3445 VDD.n3438 8.87012
R9121 VDD.n2720 VDD.n2714 8.87012
R9122 VDD.n3416 VDD.n3403 8.87012
R9123 VDD.n3391 VDD.n3384 8.87012
R9124 VDD.n3360 VDD.n3352 8.87012
R9125 VDD.n3295 VDD.n3288 8.87012
R9126 VDD.n3283 VDD.n3085 8.87012
R9127 VDD.n3283 VDD.n3077 8.87012
R9128 VDD.n3926 VDD.n3661 8.87012
R9129 VDD.n3910 VDD.n3675 8.87012
R9130 VDD.n3810 VDD.n3759 8.87012
R9131 VDD.n2857 VDD.n2848 8.87012
R9132 VDD.n3581 VDD.n3580 8.85944
R9133 VDD.n3581 VDD.n2670 8.85944
R9134 VDD.n3468 VDD.n2694 8.85944
R9135 VDD.n3446 VDD.n3445 8.85944
R9136 VDD.n3428 VDD.n2714 8.85944
R9137 VDD.n3416 VDD.n3415 8.85944
R9138 VDD.n3392 VDD.n3391 8.85944
R9139 VDD.n3360 VDD.n3359 8.85944
R9140 VDD.n3288 VDD.n3287 8.85944
R9141 VDD.n3283 VDD.n3282 8.85944
R9142 VDD.n3283 VDD.n3076 8.85944
R9143 VDD.n3926 VDD.n3666 8.85944
R9144 VDD.n3910 VDD.n3673 8.85944
R9145 VDD.n3810 VDD.n3757 8.85944
R9146 VDD.n2857 VDD.n2810 8.85944
R9147 VDD.n5647 VDD.n5646 8.85536
R9148 VDD.n5664 VDD.n5663 8.85536
R9149 VDD.n5662 VDD.n5645 8.85536
R9150 VDD.n5651 VDD.n5650 8.85536
R9151 VDD.n5628 VDD.n5627 8.85536
R9152 VDD.n5620 VDD.n5619 8.85536
R9153 VDD.n5619 VDD.n5618 8.85536
R9154 VDD.n5640 VDD.n5639 8.85536
R9155 VDD.n5641 VDD.n5640 8.85536
R9156 VDD.n5617 VDD.n5616 8.85536
R9157 VDD.n5642 VDD.n5617 8.85536
R9158 VDD.n5670 VDD.n5669 8.85536
R9159 VDD.n5669 VDD.n5668 8.85536
R9160 VDD.n6509 VDD.n6508 8.85536
R9161 VDD.n6515 VDD.n6514 8.85536
R9162 VDD.n6513 VDD.n6507 8.85536
R9163 VDD.n6469 VDD.n6468 8.85536
R9164 VDD.n6487 VDD.n6486 8.85536
R9165 VDD.n6478 VDD.n6477 8.85536
R9166 VDD.n6488 VDD.n6478 8.85536
R9167 VDD.n6491 VDD.n6490 8.85536
R9168 VDD.n6490 VDD.n6489 8.85536
R9169 VDD.n6472 VDD.n6471 8.85536
R9170 VDD.n6471 VDD.n6470 8.85536
R9171 VDD.n6503 VDD.n6502 8.85536
R9172 VDD.n6504 VDD.n6503 8.85536
R9173 VDD.n7356 VDD.n7355 8.85536
R9174 VDD.n7373 VDD.n7372 8.85536
R9175 VDD.n7371 VDD.n7354 8.85536
R9176 VDD.n7360 VDD.n7359 8.85536
R9177 VDD.n7337 VDD.n7336 8.85536
R9178 VDD.n7329 VDD.n7328 8.85536
R9179 VDD.n7328 VDD.n7327 8.85536
R9180 VDD.n7349 VDD.n7348 8.85536
R9181 VDD.n7350 VDD.n7349 8.85536
R9182 VDD.n7326 VDD.n7325 8.85536
R9183 VDD.n7351 VDD.n7326 8.85536
R9184 VDD.n7379 VDD.n7378 8.85536
R9185 VDD.n7378 VDD.n7377 8.85536
R9186 VDD.n8218 VDD.n8217 8.85536
R9187 VDD.n8224 VDD.n8223 8.85536
R9188 VDD.n8222 VDD.n8216 8.85536
R9189 VDD.n8178 VDD.n8177 8.85536
R9190 VDD.n8196 VDD.n8195 8.85536
R9191 VDD.n8187 VDD.n8186 8.85536
R9192 VDD.n8197 VDD.n8187 8.85536
R9193 VDD.n8200 VDD.n8199 8.85536
R9194 VDD.n8199 VDD.n8198 8.85536
R9195 VDD.n8181 VDD.n8180 8.85536
R9196 VDD.n8180 VDD.n8179 8.85536
R9197 VDD.n8212 VDD.n8211 8.85536
R9198 VDD.n8213 VDD.n8212 8.85536
R9199 VDD.n2578 VDD.n2577 8.85412
R9200 VDD.n3581 VDD.n2678 8.84881
R9201 VDD.n3283 VDD.n3084 8.84881
R9202 VDD.n3810 VDD.n3755 8.84881
R9203 VDD.n3926 VDD.n3667 8.84881
R9204 VDD.n3910 VDD.n3674 8.84881
R9205 VDD.n2857 VDD.n2811 8.84881
R9206 VDD.n2577 VDD.n2576 8.84352
R9207 VDD.n2577 VDD.n2517 8.83298
R9208 VDD.n3993 VDD.n3992 8.78757
R9209 VDD.n5500 VDD.n5499 8.77128
R9210 VDD.n3867 VDD.n3866 8.76429
R9211 VDD.n3845 VDD.n3840 8.76429
R9212 VDD.n8791 VDD.n8790 8.7045
R9213 VDD.n8792 VDD.n8791 8.7045
R9214 VDD.n8795 VDD.n8792 8.7045
R9215 VDD.n8814 VDD.n8813 8.7045
R9216 VDD.n8813 VDD.n8255 8.7045
R9217 VDD.n9015 VDD.n8255 8.7045
R9218 VDD.n9015 VDD.n9014 8.7045
R9219 VDD.n9014 VDD.n9013 8.7045
R9220 VDD.n8393 VDD.n8392 8.7045
R9221 VDD.n8393 VDD.n8283 8.7045
R9222 VDD.n8402 VDD.n8283 8.7045
R9223 VDD.n7936 VDD.n7935 8.7045
R9224 VDD.n7937 VDD.n7936 8.7045
R9225 VDD.n7940 VDD.n7937 8.7045
R9226 VDD.n7959 VDD.n7958 8.7045
R9227 VDD.n7958 VDD.n7400 8.7045
R9228 VDD.n8160 VDD.n7400 8.7045
R9229 VDD.n8160 VDD.n8159 8.7045
R9230 VDD.n8159 VDD.n8158 8.7045
R9231 VDD.n7538 VDD.n7537 8.7045
R9232 VDD.n7538 VDD.n7428 8.7045
R9233 VDD.n7547 VDD.n7428 8.7045
R9234 VDD.n7082 VDD.n7081 8.7045
R9235 VDD.n7083 VDD.n7082 8.7045
R9236 VDD.n7086 VDD.n7083 8.7045
R9237 VDD.n7105 VDD.n7104 8.7045
R9238 VDD.n7104 VDD.n6546 8.7045
R9239 VDD.n7306 VDD.n6546 8.7045
R9240 VDD.n7306 VDD.n7305 8.7045
R9241 VDD.n7305 VDD.n7304 8.7045
R9242 VDD.n6684 VDD.n6683 8.7045
R9243 VDD.n6684 VDD.n6574 8.7045
R9244 VDD.n6693 VDD.n6574 8.7045
R9245 VDD.n6227 VDD.n6226 8.7045
R9246 VDD.n6228 VDD.n6227 8.7045
R9247 VDD.n6231 VDD.n6228 8.7045
R9248 VDD.n6250 VDD.n6249 8.7045
R9249 VDD.n6249 VDD.n5691 8.7045
R9250 VDD.n6451 VDD.n5691 8.7045
R9251 VDD.n6451 VDD.n6450 8.7045
R9252 VDD.n6450 VDD.n6449 8.7045
R9253 VDD.n5829 VDD.n5828 8.7045
R9254 VDD.n5829 VDD.n5719 8.7045
R9255 VDD.n5838 VDD.n5719 8.7045
R9256 VDD.n2620 VDD.n2604 8.65557
R9257 VDD.n3947 VDD.n2499 8.65557
R9258 VDD.n4357 VDD.n4356 8.46493
R9259 VDD.n2455 VDD.n2454 8.45089
R9260 VDD.n2622 VDD.n2598 8.45089
R9261 VDD.n3993 VDD.n2491 8.45089
R9262 VDD.n3997 VDD.n2489 8.45089
R9263 VDD.n2446 VDD.n2444 8.45089
R9264 VDD.n5504 VDD.n5503 8.45089
R9265 VDD.n5500 VDD.n249 8.45089
R9266 VDD.n2626 VDD.n2597 8.45089
R9267 VDD.n2620 VDD.n2619 8.45089
R9268 VDD.n4001 VDD.n2487 8.45089
R9269 VDD.n3955 VDD.n3952 8.45089
R9270 VDD.n3948 VDD.n3947 8.45089
R9271 VDD.n2496 VDD.n2495 8.45089
R9272 VDD.n268 VDD.n250 8.40959
R9273 VDD.n5474 VDD.n268 8.40959
R9274 VDD.n5472 VDD.n268 8.40959
R9275 VDD.n4007 VDD.n2479 8.40959
R9276 VDD.n2481 VDD.n2479 8.40959
R9277 VDD.n4009 VDD.n2479 8.40959
R9278 VDD.n3951 VDD.n3950 8.40959
R9279 VDD.n3951 VDD.n2503 8.40959
R9280 VDD.n3951 VDD.n2502 8.40959
R9281 VDD.n5665 VDD.n5645 8.39408
R9282 VDD.n5665 VDD.n5664 8.39408
R9283 VDD.n5650 VDD.n5644 8.39408
R9284 VDD.n6516 VDD.n6507 8.39408
R9285 VDD.n6516 VDD.n6515 8.39408
R9286 VDD.n6518 VDD.n6469 8.39408
R9287 VDD.n7374 VDD.n7354 8.39408
R9288 VDD.n7374 VDD.n7373 8.39408
R9289 VDD.n7359 VDD.n7353 8.39408
R9290 VDD.n8225 VDD.n8216 8.39408
R9291 VDD.n8225 VDD.n8224 8.39408
R9292 VDD.n8227 VDD.n8178 8.39408
R9293 VDD.n5646 VDD.n5643 8.39405
R9294 VDD.n6508 VDD.n6506 8.39405
R9295 VDD.n7355 VDD.n7352 8.39405
R9296 VDD.n8217 VDD.n8215 8.39405
R9297 VDD.n2588 VDD.n2509 8.08763
R9298 VDD.n4011 VDD.n2476 8.07007
R9299 VDD.n1816 VDD.n1030 8.06816
R9300 VDD.n1011 VDD.n1002 8.06816
R9301 VDD.n4570 VDD.n1012 8.06816
R9302 VDD.n4555 VDD.n1910 8.06816
R9303 VDD.n4554 VDD.n1911 8.06816
R9304 VDD.n4551 VDD.n1917 8.06816
R9305 VDD.n1923 VDD.n1922 8.06816
R9306 VDD.n4545 VDD.n1924 8.06816
R9307 VDD.n4535 VDD.n1942 8.06816
R9308 VDD.n4532 VDD.n1948 8.06816
R9309 VDD.n4526 VDD.n1954 8.06816
R9310 VDD.n4520 VDD.n1962 8.06816
R9311 VDD.n4519 VDD.n1963 8.06816
R9312 VDD.n4511 VDD.n1979 8.06816
R9313 VDD.n4510 VDD.n1980 8.06816
R9314 VDD.n4507 VDD.n1986 8.06816
R9315 VDD.n1995 VDD.n1994 8.06816
R9316 VDD.n4501 VDD.n1996 8.06816
R9317 VDD.n4488 VDD.n2022 8.06816
R9318 VDD.n2028 VDD.n2027 8.06816
R9319 VDD.n4482 VDD.n2029 8.06816
R9320 VDD.n4473 VDD.n2046 8.06816
R9321 VDD.n4472 VDD.n2047 8.06816
R9322 VDD.n2089 VDD.n2057 8.06816
R9323 VDD.n4463 VDD.n2058 8.06816
R9324 VDD.n2069 VDD.n2068 8.06816
R9325 VDD.n4454 VDD.n2070 8.06816
R9326 VDD.n2075 VDD.n2074 8.06816
R9327 VDD.n4448 VDD.n2076 8.06816
R9328 VDD.n4439 VDD.n2099 8.06816
R9329 VDD.n4438 VDD.n2100 8.06816
R9330 VDD.n4435 VDD.n2106 8.06816
R9331 VDD.n2112 VDD.n2111 8.06816
R9332 VDD.n4429 VDD.n2113 8.06816
R9333 VDD.n4420 VDD.n2130 8.06816
R9334 VDD.n4416 VDD.n2137 8.06816
R9335 VDD.n2143 VDD.n2142 8.06816
R9336 VDD.n4410 VDD.n2144 8.06816
R9337 VDD.n4401 VDD.n2161 8.06816
R9338 VDD.n4400 VDD.n2162 8.06816
R9339 VDD.n4397 VDD.n2168 8.06816
R9340 VDD.n4391 VDD.n2175 8.06816
R9341 VDD.n4385 VDD.n2183 8.06816
R9342 VDD.n4384 VDD.n2184 8.06816
R9343 VDD.n4376 VDD.n2200 8.06816
R9344 VDD.n4375 VDD.n2201 8.06816
R9345 VDD.n4372 VDD.n2207 8.06816
R9346 VDD.n4366 VDD.n2217 8.06816
R9347 VDD.n4357 VDD.n2234 8.06816
R9348 VDD.t48 VDD.n4107 7.99076
R9349 VDD.n2543 VDD.n2518 7.52991
R9350 VDD.n3496 VDD.n3495 7.45411
R9351 VDD.n3513 VDD.n3512 7.45411
R9352 VDD.n3198 VDD.n3197 7.45411
R9353 VDD.n3215 VDD.n3214 7.45411
R9354 VDD.n3746 VDD.n3745 7.45411
R9355 VDD.n3839 VDD.n3838 7.45411
R9356 VDD.n3843 VDD.n3842 7.45411
R9357 VDD.n3883 VDD.n3882 7.45411
R9358 VDD.n3862 VDD.n3861 7.45411
R9359 VDD.n3865 VDD.n3864 7.45411
R9360 VDD.n2826 VDD.n2825 7.45411
R9361 VDD.n2968 VDD.n2967 7.45411
R9362 VDD.n3355 VDD.n3354 7.33876
R9363 VDD.n3284 VDD.n3074 7.33876
R9364 VDD.n4148 VDD.t50 7.14968
R9365 VDD.n8245 VDD.n8244 7.09014
R9366 VDD.n9022 VDD.n8243 7.09014
R9367 VDD.n7390 VDD.n7389 7.09014
R9368 VDD.n8167 VDD.n7388 7.09014
R9369 VDD.n6536 VDD.n6535 7.09014
R9370 VDD.n7313 VDD.n6534 7.09014
R9371 VDD.n5681 VDD.n5680 7.09014
R9372 VDD.n6458 VDD.n5679 7.09014
R9373 VDD.n8635 VDD.n8506 7.07692
R9374 VDD.n8629 VDD.n8506 7.07692
R9375 VDD.n8629 VDD.n8628 7.07692
R9376 VDD.n8628 VDD.n8627 7.07692
R9377 VDD.n8627 VDD.n8510 7.07692
R9378 VDD.n8621 VDD.n8510 7.07692
R9379 VDD.n8621 VDD.n8620 7.07692
R9380 VDD.n8620 VDD.n8619 7.07692
R9381 VDD.n8619 VDD.n8514 7.07692
R9382 VDD.n8613 VDD.n8514 7.07692
R9383 VDD.n8613 VDD.n8612 7.07692
R9384 VDD.n8612 VDD.n8611 7.07692
R9385 VDD.n8611 VDD.n8518 7.07692
R9386 VDD.n8605 VDD.n8518 7.07692
R9387 VDD.n8605 VDD.n8604 7.07692
R9388 VDD.n8604 VDD.n8603 7.07692
R9389 VDD.n8603 VDD.n8522 7.07692
R9390 VDD.n8597 VDD.n8522 7.07692
R9391 VDD.n8597 VDD.n8596 7.07692
R9392 VDD.n8596 VDD.n8595 7.07692
R9393 VDD.n8595 VDD.n8526 7.07692
R9394 VDD.n8589 VDD.n8526 7.07692
R9395 VDD.n8589 VDD.n8588 7.07692
R9396 VDD.n8588 VDD.n8587 7.07692
R9397 VDD.n8587 VDD.n8530 7.07692
R9398 VDD.n7780 VDD.n7651 7.07692
R9399 VDD.n7774 VDD.n7651 7.07692
R9400 VDD.n7774 VDD.n7773 7.07692
R9401 VDD.n7773 VDD.n7772 7.07692
R9402 VDD.n7772 VDD.n7655 7.07692
R9403 VDD.n7766 VDD.n7655 7.07692
R9404 VDD.n7766 VDD.n7765 7.07692
R9405 VDD.n7765 VDD.n7764 7.07692
R9406 VDD.n7764 VDD.n7659 7.07692
R9407 VDD.n7758 VDD.n7659 7.07692
R9408 VDD.n7758 VDD.n7757 7.07692
R9409 VDD.n7757 VDD.n7756 7.07692
R9410 VDD.n7756 VDD.n7663 7.07692
R9411 VDD.n7750 VDD.n7663 7.07692
R9412 VDD.n7750 VDD.n7749 7.07692
R9413 VDD.n7749 VDD.n7748 7.07692
R9414 VDD.n7748 VDD.n7667 7.07692
R9415 VDD.n7742 VDD.n7667 7.07692
R9416 VDD.n7742 VDD.n7741 7.07692
R9417 VDD.n7741 VDD.n7740 7.07692
R9418 VDD.n7740 VDD.n7671 7.07692
R9419 VDD.n7734 VDD.n7671 7.07692
R9420 VDD.n7734 VDD.n7733 7.07692
R9421 VDD.n7733 VDD.n7732 7.07692
R9422 VDD.n7732 VDD.n7675 7.07692
R9423 VDD.n6926 VDD.n6797 7.07692
R9424 VDD.n6920 VDD.n6797 7.07692
R9425 VDD.n6920 VDD.n6919 7.07692
R9426 VDD.n6919 VDD.n6918 7.07692
R9427 VDD.n6918 VDD.n6801 7.07692
R9428 VDD.n6912 VDD.n6801 7.07692
R9429 VDD.n6912 VDD.n6911 7.07692
R9430 VDD.n6911 VDD.n6910 7.07692
R9431 VDD.n6910 VDD.n6805 7.07692
R9432 VDD.n6904 VDD.n6805 7.07692
R9433 VDD.n6904 VDD.n6903 7.07692
R9434 VDD.n6903 VDD.n6902 7.07692
R9435 VDD.n6902 VDD.n6809 7.07692
R9436 VDD.n6896 VDD.n6809 7.07692
R9437 VDD.n6896 VDD.n6895 7.07692
R9438 VDD.n6895 VDD.n6894 7.07692
R9439 VDD.n6894 VDD.n6813 7.07692
R9440 VDD.n6888 VDD.n6813 7.07692
R9441 VDD.n6888 VDD.n6887 7.07692
R9442 VDD.n6887 VDD.n6886 7.07692
R9443 VDD.n6886 VDD.n6817 7.07692
R9444 VDD.n6880 VDD.n6817 7.07692
R9445 VDD.n6880 VDD.n6879 7.07692
R9446 VDD.n6879 VDD.n6878 7.07692
R9447 VDD.n6878 VDD.n6821 7.07692
R9448 VDD.n6071 VDD.n5942 7.07692
R9449 VDD.n6065 VDD.n5942 7.07692
R9450 VDD.n6065 VDD.n6064 7.07692
R9451 VDD.n6064 VDD.n6063 7.07692
R9452 VDD.n6063 VDD.n5946 7.07692
R9453 VDD.n6057 VDD.n5946 7.07692
R9454 VDD.n6057 VDD.n6056 7.07692
R9455 VDD.n6056 VDD.n6055 7.07692
R9456 VDD.n6055 VDD.n5950 7.07692
R9457 VDD.n6049 VDD.n5950 7.07692
R9458 VDD.n6049 VDD.n6048 7.07692
R9459 VDD.n6048 VDD.n6047 7.07692
R9460 VDD.n6047 VDD.n5954 7.07692
R9461 VDD.n6041 VDD.n5954 7.07692
R9462 VDD.n6041 VDD.n6040 7.07692
R9463 VDD.n6040 VDD.n6039 7.07692
R9464 VDD.n6039 VDD.n5958 7.07692
R9465 VDD.n6033 VDD.n5958 7.07692
R9466 VDD.n6033 VDD.n6032 7.07692
R9467 VDD.n6032 VDD.n6031 7.07692
R9468 VDD.n6031 VDD.n5962 7.07692
R9469 VDD.n6025 VDD.n5962 7.07692
R9470 VDD.n6025 VDD.n6024 7.07692
R9471 VDD.n6024 VDD.n6023 7.07692
R9472 VDD.n6023 VDD.n5966 7.07692
R9473 VDD.n8837 VDD.n8683 7.05178
R9474 VDD.n8836 VDD.n8695 7.05178
R9475 VDD.n8829 VDD.n8701 7.05178
R9476 VDD.n8708 VDD.n8702 7.05178
R9477 VDD.n7982 VDD.n7828 7.05178
R9478 VDD.n7981 VDD.n7840 7.05178
R9479 VDD.n7974 VDD.n7846 7.05178
R9480 VDD.n7853 VDD.n7847 7.05178
R9481 VDD.n7128 VDD.n6974 7.05178
R9482 VDD.n7127 VDD.n6986 7.05178
R9483 VDD.n7120 VDD.n6992 7.05178
R9484 VDD.n6999 VDD.n6993 7.05178
R9485 VDD.n6273 VDD.n6119 7.05178
R9486 VDD.n6272 VDD.n6131 7.05178
R9487 VDD.n6265 VDD.n6137 7.05178
R9488 VDD.n6144 VDD.n6138 7.05178
R9489 VDD.n3952 VDD.n2500 6.89484
R9490 VDD.n2605 VDD.n2597 6.89484
R9491 VDD.n2623 VDD.n2622 6.89484
R9492 VDD.n2446 VDD.n2445 6.89484
R9493 VDD.n5503 VDD.n5502 6.89484
R9494 VDD.n4001 VDD.n4000 6.89484
R9495 VDD.n3994 VDD.n2489 6.89484
R9496 VDD.n3498 VDD.n3497 6.80334
R9497 VDD.n3200 VDD.n3199 6.80334
R9498 VDD.n3748 VDD.n3747 6.80334
R9499 VDD.n2828 VDD.n2823 6.80105
R9500 VDD.n2970 VDD.n2965 6.80105
R9501 VDD.n3510 VDD.n3509 6.80104
R9502 VDD.n3212 VDD.n3211 6.80104
R9503 VDD.n3880 VDD.n3879 6.80104
R9504 VDD.n8580 VDD.n8579 6.59444
R9505 VDD.n8579 VDD.n8534 6.59444
R9506 VDD.n8574 VDD.n8534 6.59444
R9507 VDD.n8574 VDD.n8573 6.59444
R9508 VDD.n8573 VDD.n8572 6.59444
R9509 VDD.n8572 VDD.n8538 6.59444
R9510 VDD.n8566 VDD.n8538 6.59444
R9511 VDD.n8566 VDD.n8565 6.59444
R9512 VDD.n8565 VDD.n8564 6.59444
R9513 VDD.n8564 VDD.n8543 6.59444
R9514 VDD.n8558 VDD.n8543 6.59444
R9515 VDD.n8558 VDD.n8557 6.59444
R9516 VDD.n8557 VDD.n8556 6.59444
R9517 VDD.n8556 VDD.n8547 6.59444
R9518 VDD.n8550 VDD.n8547 6.59444
R9519 VDD.n8550 VDD.n8549 6.59444
R9520 VDD.n8549 VDD.n8276 6.59444
R9521 VDD.n7725 VDD.n7724 6.59444
R9522 VDD.n7724 VDD.n7679 6.59444
R9523 VDD.n7719 VDD.n7679 6.59444
R9524 VDD.n7719 VDD.n7718 6.59444
R9525 VDD.n7718 VDD.n7717 6.59444
R9526 VDD.n7717 VDD.n7683 6.59444
R9527 VDD.n7711 VDD.n7683 6.59444
R9528 VDD.n7711 VDD.n7710 6.59444
R9529 VDD.n7710 VDD.n7709 6.59444
R9530 VDD.n7709 VDD.n7688 6.59444
R9531 VDD.n7703 VDD.n7688 6.59444
R9532 VDD.n7703 VDD.n7702 6.59444
R9533 VDD.n7702 VDD.n7701 6.59444
R9534 VDD.n7701 VDD.n7692 6.59444
R9535 VDD.n7695 VDD.n7692 6.59444
R9536 VDD.n7695 VDD.n7694 6.59444
R9537 VDD.n7694 VDD.n7421 6.59444
R9538 VDD.n6871 VDD.n6870 6.59444
R9539 VDD.n6870 VDD.n6825 6.59444
R9540 VDD.n6865 VDD.n6825 6.59444
R9541 VDD.n6865 VDD.n6864 6.59444
R9542 VDD.n6864 VDD.n6863 6.59444
R9543 VDD.n6863 VDD.n6829 6.59444
R9544 VDD.n6857 VDD.n6829 6.59444
R9545 VDD.n6857 VDD.n6856 6.59444
R9546 VDD.n6856 VDD.n6855 6.59444
R9547 VDD.n6855 VDD.n6834 6.59444
R9548 VDD.n6849 VDD.n6834 6.59444
R9549 VDD.n6849 VDD.n6848 6.59444
R9550 VDD.n6848 VDD.n6847 6.59444
R9551 VDD.n6847 VDD.n6838 6.59444
R9552 VDD.n6841 VDD.n6838 6.59444
R9553 VDD.n6841 VDD.n6840 6.59444
R9554 VDD.n6840 VDD.n6567 6.59444
R9555 VDD.n6016 VDD.n6015 6.59444
R9556 VDD.n6015 VDD.n5970 6.59444
R9557 VDD.n6010 VDD.n5970 6.59444
R9558 VDD.n6010 VDD.n6009 6.59444
R9559 VDD.n6009 VDD.n6008 6.59444
R9560 VDD.n6008 VDD.n5974 6.59444
R9561 VDD.n6002 VDD.n5974 6.59444
R9562 VDD.n6002 VDD.n6001 6.59444
R9563 VDD.n6001 VDD.n6000 6.59444
R9564 VDD.n6000 VDD.n5979 6.59444
R9565 VDD.n5994 VDD.n5979 6.59444
R9566 VDD.n5994 VDD.n5993 6.59444
R9567 VDD.n5993 VDD.n5992 6.59444
R9568 VDD.n5992 VDD.n5983 6.59444
R9569 VDD.n5986 VDD.n5983 6.59444
R9570 VDD.n5986 VDD.n5985 6.59444
R9571 VDD.n5985 VDD.n5712 6.59444
R9572 VDD.n2216 VDD.t77 6.48108
R9573 VDD.n4419 VDD.t81 6.34882
R9574 VDD.n2723 VDD.n2721 6.31678
R9575 VDD.n3418 VDD.n3417 6.31678
R9576 VDD.n3364 VDD.n3361 6.31678
R9577 VDD.n3292 VDD.n3289 6.31678
R9578 VDD.n3455 VDD.n2699 6.31678
R9579 VDD.n3444 VDD.n3443 6.31678
R9580 VDD.n3390 VDD.n3389 6.31678
R9581 VDD.n2547 VDD.n2516 6.31321
R9582 VDD.n4173 VDD.t6 6.3086
R9583 VDD.n2619 VDD.n2618 6.30775
R9584 VDD.n3620 VDD.n2475 6.30775
R9585 VDD.n8868 VDD.n8867 6.17355
R9586 VDD.n8869 VDD.n8868 6.17355
R9587 VDD.n8869 VDD.n8462 6.17355
R9588 VDD.n8875 VDD.n8462 6.17355
R9589 VDD.n8876 VDD.n8875 6.17355
R9590 VDD.n8877 VDD.n8876 6.17355
R9591 VDD.n8877 VDD.n8458 6.17355
R9592 VDD.n8883 VDD.n8458 6.17355
R9593 VDD.n8884 VDD.n8883 6.17355
R9594 VDD.n8885 VDD.n8884 6.17355
R9595 VDD.n8885 VDD.n8454 6.17355
R9596 VDD.n8891 VDD.n8454 6.17355
R9597 VDD.n8013 VDD.n8012 6.17355
R9598 VDD.n8014 VDD.n8013 6.17355
R9599 VDD.n8014 VDD.n7607 6.17355
R9600 VDD.n8020 VDD.n7607 6.17355
R9601 VDD.n8021 VDD.n8020 6.17355
R9602 VDD.n8022 VDD.n8021 6.17355
R9603 VDD.n8022 VDD.n7603 6.17355
R9604 VDD.n8028 VDD.n7603 6.17355
R9605 VDD.n8029 VDD.n8028 6.17355
R9606 VDD.n8030 VDD.n8029 6.17355
R9607 VDD.n8030 VDD.n7599 6.17355
R9608 VDD.n8036 VDD.n7599 6.17355
R9609 VDD.n7159 VDD.n7158 6.17355
R9610 VDD.n7160 VDD.n7159 6.17355
R9611 VDD.n7160 VDD.n6753 6.17355
R9612 VDD.n7166 VDD.n6753 6.17355
R9613 VDD.n7167 VDD.n7166 6.17355
R9614 VDD.n7168 VDD.n7167 6.17355
R9615 VDD.n7168 VDD.n6749 6.17355
R9616 VDD.n7174 VDD.n6749 6.17355
R9617 VDD.n7175 VDD.n7174 6.17355
R9618 VDD.n7176 VDD.n7175 6.17355
R9619 VDD.n7176 VDD.n6745 6.17355
R9620 VDD.n7182 VDD.n6745 6.17355
R9621 VDD.n6304 VDD.n6303 6.17355
R9622 VDD.n6305 VDD.n6304 6.17355
R9623 VDD.n6305 VDD.n5898 6.17355
R9624 VDD.n6311 VDD.n5898 6.17355
R9625 VDD.n6312 VDD.n6311 6.17355
R9626 VDD.n6313 VDD.n6312 6.17355
R9627 VDD.n6313 VDD.n5894 6.17355
R9628 VDD.n6319 VDD.n5894 6.17355
R9629 VDD.n6320 VDD.n6319 6.17355
R9630 VDD.n6321 VDD.n6320 6.17355
R9631 VDD.n6321 VDD.n5890 6.17355
R9632 VDD.n6327 VDD.n5890 6.17355
R9633 VDD.n4577 VDD.n4576 6.08431
R9634 VDD.n2664 VDD.n2663 6.02403
R9635 VDD.n2667 VDD.n2665 6.02403
R9636 VDD.n3555 VDD.n3554 6.02403
R9637 VDD.n3549 VDD.n3548 6.02403
R9638 VDD.n3257 VDD.n3256 6.02403
R9639 VDD.n3251 VDD.n3250 6.02403
R9640 VDD.n3133 VDD.n3132 6.02403
R9641 VDD.n3136 VDD.n3134 6.02403
R9642 VDD.n3791 VDD.n3790 6.02403
R9643 VDD.n3773 VDD.n3766 6.02403
R9644 VDD.n2923 VDD.n2922 6.02403
R9645 VDD.n2941 VDD.n2919 6.02403
R9646 VDD.n71 VDD.n70 6.02403
R9647 VDD.n65 VDD.n61 6.02403
R9648 VDD.n5578 VDD.n5568 6.02403
R9649 VDD.n5573 VDD.n5570 6.02403
R9650 VDD.n217 VDD.n216 6.02403
R9651 VDD.n211 VDD.n207 6.02403
R9652 VDD.n1271 VDD.n1270 5.96815
R9653 VDD.n4536 VDD.t46 5.95205
R9654 VDD.n2090 VDD.t106 5.95205
R9655 VDD.n8705 VDD.n8678 5.80317
R9656 VDD.n8827 VDD.n8705 5.80317
R9657 VDD.n8827 VDD.n8826 5.80317
R9658 VDD.n8826 VDD.n8825 5.80317
R9659 VDD.n8825 VDD.n8706 5.80317
R9660 VDD.n8730 VDD.n8725 5.80317
R9661 VDD.n8726 VDD.n8725 5.80317
R9662 VDD.n8726 VDD.n8270 5.80317
R9663 VDD.n9003 VDD.n8270 5.80317
R9664 VDD.n9003 VDD.n9002 5.80317
R9665 VDD.n7850 VDD.n7823 5.80317
R9666 VDD.n7972 VDD.n7850 5.80317
R9667 VDD.n7972 VDD.n7971 5.80317
R9668 VDD.n7971 VDD.n7970 5.80317
R9669 VDD.n7970 VDD.n7851 5.80317
R9670 VDD.n7875 VDD.n7870 5.80317
R9671 VDD.n7871 VDD.n7870 5.80317
R9672 VDD.n7871 VDD.n7415 5.80317
R9673 VDD.n8148 VDD.n7415 5.80317
R9674 VDD.n8148 VDD.n8147 5.80317
R9675 VDD.n6996 VDD.n6969 5.80317
R9676 VDD.n7118 VDD.n6996 5.80317
R9677 VDD.n7118 VDD.n7117 5.80317
R9678 VDD.n7117 VDD.n7116 5.80317
R9679 VDD.n7116 VDD.n6997 5.80317
R9680 VDD.n7021 VDD.n7016 5.80317
R9681 VDD.n7017 VDD.n7016 5.80317
R9682 VDD.n7017 VDD.n6561 5.80317
R9683 VDD.n7294 VDD.n6561 5.80317
R9684 VDD.n7294 VDD.n7293 5.80317
R9685 VDD.n6141 VDD.n6114 5.80317
R9686 VDD.n6263 VDD.n6141 5.80317
R9687 VDD.n6263 VDD.n6262 5.80317
R9688 VDD.n6262 VDD.n6261 5.80317
R9689 VDD.n6261 VDD.n6142 5.80317
R9690 VDD.n6166 VDD.n6161 5.80317
R9691 VDD.n6162 VDD.n6161 5.80317
R9692 VDD.n6162 VDD.n5706 5.80317
R9693 VDD.n6439 VDD.n5706 5.80317
R9694 VDD.n6439 VDD.n6438 5.80317
R9695 VDD.n2981 VDD.n2977 5.73742
R9696 VDD.n3494 VDD.n3493 5.64756
R9697 VDD.n3502 VDD.n3501 5.64756
R9698 VDD.n3517 VDD.n3516 5.64756
R9699 VDD.n3511 VDD.n3507 5.64756
R9700 VDD.n3196 VDD.n3195 5.64756
R9701 VDD.n3204 VDD.n3203 5.64756
R9702 VDD.n3219 VDD.n3218 5.64756
R9703 VDD.n3213 VDD.n3209 5.64756
R9704 VDD.n3744 VDD.n3743 5.64756
R9705 VDD.n3752 VDD.n3751 5.64756
R9706 VDD.n3835 VDD.n3739 5.64756
R9707 VDD.n3837 VDD.n3737 5.64756
R9708 VDD.n3844 VDD.n3841 5.64756
R9709 VDD.n3850 VDD.n3849 5.64756
R9710 VDD.n3887 VDD.n3886 5.64756
R9711 VDD.n3881 VDD.n3877 5.64756
R9712 VDD.n3858 VDD.n3712 5.64756
R9713 VDD.n3860 VDD.n3709 5.64756
R9714 VDD.n3863 VDD.n3710 5.64756
R9715 VDD.n3872 VDD.n3871 5.64756
R9716 VDD.n2827 VDD.n2824 5.64756
R9717 VDD.n2832 VDD.n2831 5.64756
R9718 VDD.n2969 VDD.n2966 5.64756
R9719 VDD.n2974 VDD.n2973 5.64756
R9720 VDD.n100 VDD.n99 5.64756
R9721 VDD.n133 VDD.n111 5.64756
R9722 VDD.n5557 VDD.n5543 5.64756
R9723 VDD.n199 VDD.n198 5.64756
R9724 VDD.n2544 VDD.n2543 5.64756
R9725 VDD.n2548 VDD.n2547 5.64756
R9726 VDD.n2681 VDD.n2680 5.63005
R9727 VDD.n3469 VDD.n2691 5.63005
R9728 VDD.n3447 VDD.n3435 5.63005
R9729 VDD.n3429 VDD.n2711 5.63005
R9730 VDD.n3413 VDD.n3404 5.63005
R9731 VDD.n3393 VDD.n3381 5.63005
R9732 VDD.n3087 VDD.n3086 5.63005
R9733 VDD.n8991 VDD.n8404 5.61598
R9734 VDD.n8991 VDD.n8990 5.61598
R9735 VDD.n8990 VDD.n8989 5.61598
R9736 VDD.n8989 VDD.n8405 5.61598
R9737 VDD.n8983 VDD.n8405 5.61598
R9738 VDD.n8983 VDD.n8982 5.61598
R9739 VDD.n8982 VDD.n8981 5.61598
R9740 VDD.n8981 VDD.n8409 5.61598
R9741 VDD.n8975 VDD.n8409 5.61598
R9742 VDD.n8975 VDD.n8974 5.61598
R9743 VDD.n8974 VDD.n8973 5.61598
R9744 VDD.n8973 VDD.n8413 5.61598
R9745 VDD.n8136 VDD.n7549 5.61598
R9746 VDD.n8136 VDD.n8135 5.61598
R9747 VDD.n8135 VDD.n8134 5.61598
R9748 VDD.n8134 VDD.n7550 5.61598
R9749 VDD.n8128 VDD.n7550 5.61598
R9750 VDD.n8128 VDD.n8127 5.61598
R9751 VDD.n8127 VDD.n8126 5.61598
R9752 VDD.n8126 VDD.n7554 5.61598
R9753 VDD.n8120 VDD.n7554 5.61598
R9754 VDD.n8120 VDD.n8119 5.61598
R9755 VDD.n8119 VDD.n8118 5.61598
R9756 VDD.n8118 VDD.n7558 5.61598
R9757 VDD.n7282 VDD.n6695 5.61598
R9758 VDD.n7282 VDD.n7281 5.61598
R9759 VDD.n7281 VDD.n7280 5.61598
R9760 VDD.n7280 VDD.n6696 5.61598
R9761 VDD.n7274 VDD.n6696 5.61598
R9762 VDD.n7274 VDD.n7273 5.61598
R9763 VDD.n7273 VDD.n7272 5.61598
R9764 VDD.n7272 VDD.n6700 5.61598
R9765 VDD.n7266 VDD.n6700 5.61598
R9766 VDD.n7266 VDD.n7265 5.61598
R9767 VDD.n7265 VDD.n7264 5.61598
R9768 VDD.n7264 VDD.n6704 5.61598
R9769 VDD.n6427 VDD.n5840 5.61598
R9770 VDD.n6427 VDD.n6426 5.61598
R9771 VDD.n6426 VDD.n6425 5.61598
R9772 VDD.n6425 VDD.n5841 5.61598
R9773 VDD.n6419 VDD.n5841 5.61598
R9774 VDD.n6419 VDD.n6418 5.61598
R9775 VDD.n6418 VDD.n6417 5.61598
R9776 VDD.n6417 VDD.n5845 5.61598
R9777 VDD.n6411 VDD.n5845 5.61598
R9778 VDD.n6411 VDD.n6410 5.61598
R9779 VDD.n6410 VDD.n6409 5.61598
R9780 VDD.n6409 VDD.n5849 5.61598
R9781 VDD.n3173 VDD.n3093 5.57349
R9782 VDD.n3614 VDD.n2635 5.57349
R9783 VDD.t107 VDD.n3581 5.5395
R9784 VDD.n3581 VDD.t124 5.5395
R9785 VDD.n2694 VDD.t124 5.5395
R9786 VDD.n2694 VDD.t82 5.5395
R9787 VDD.n3445 VDD.t95 5.5395
R9788 VDD.n3445 VDD.t78 5.5395
R9789 VDD.n2714 VDD.t143 5.5395
R9790 VDD.n2714 VDD.t158 5.5395
R9791 VDD.n3416 VDD.t159 5.5395
R9792 VDD.n3416 VDD.t84 5.5395
R9793 VDD.n3391 VDD.t128 5.5395
R9794 VDD.n3391 VDD.t45 5.5395
R9795 VDD.n3360 VDD.t136 5.5395
R9796 VDD.n3360 VDD.t138 5.5395
R9797 VDD.n3288 VDD.t137 5.5395
R9798 VDD.n3288 VDD.t122 5.5395
R9799 VDD.t122 VDD.n3283 5.5395
R9800 VDD.n3283 VDD.t116 5.5395
R9801 VDD.n3810 VDD.t109 5.5395
R9802 VDD.n3810 VDD.t104 5.5395
R9803 VDD.n3926 VDD.t104 5.5395
R9804 VDD.n3926 VDD.t113 5.5395
R9805 VDD.t113 VDD.n3910 5.5395
R9806 VDD.n3910 VDD.t111 5.5395
R9807 VDD.n2857 VDD.t127 5.5395
R9808 VDD.n2857 VDD.t5 5.5395
R9809 VDD.n3024 VDD.t9 5.5395
R9810 VDD.n3024 VDD.t119 5.5395
R9811 VDD.n132 VDD.t49 5.5395
R9812 VDD.n132 VDD.t53 5.5395
R9813 VDD.n2014 VDD.n2013 5.42303
R9814 VDD.n3553 VDD.n2675 5.39401
R9815 VDD.n3255 VDD.n3081 5.39401
R9816 VDD.n3550 VDD.n2675 5.39321
R9817 VDD.n3252 VDD.n3081 5.39321
R9818 VDD.n6524 VDD 5.2805
R9819 VDD.n8233 VDD 5.2805
R9820 VDD.n4298 VDD.t96 5.27719
R9821 VDD.n3593 VDD.n2659 5.27109
R9822 VDD.n3588 VDD.n2661 5.27109
R9823 VDD.n3560 VDD.n3559 5.27109
R9824 VDD.n3544 VDD.n3543 5.27109
R9825 VDD.n3262 VDD.n3261 5.27109
R9826 VDD.n3246 VDD.n3245 5.27109
R9827 VDD.n3149 VDD.n3128 5.27109
R9828 VDD.n3144 VDD.n3130 5.27109
R9829 VDD.n55 VDD.n53 5.27109
R9830 VDD.n60 VDD.n56 5.27109
R9831 VDD.n5585 VDD.n5584 5.27109
R9832 VDD.n5579 VDD.n5564 5.27109
R9833 VDD.n183 VDD.n181 5.27109
R9834 VDD.n206 VDD.n184 5.27109
R9835 VDD.n46 VDD.n40 5.25364
R9836 VDD.n5547 VDD.n5541 5.25364
R9837 VDD.n191 VDD.n185 5.25364
R9838 VDD.n8757 VDD.n8756 5.2318
R9839 VDD.n7902 VDD.n7901 5.2318
R9840 VDD.n7048 VDD.n7047 5.2318
R9841 VDD.n6193 VDD.n6192 5.2318
R9842 VDD.n2615 VDD.n2607 5.15851
R9843 VDD.n2835 VDD.n2811 4.96787
R9844 VDD.n3521 VDD.n2678 4.95584
R9845 VDD.n3223 VDD.n3084 4.95584
R9846 VDD.n3829 VDD.n3755 4.95584
R9847 VDD.n3732 VDD.n3667 4.95584
R9848 VDD.n3891 VDD.n3674 4.95584
R9849 VDD.n315 VDD.n310 4.91801
R9850 VDD.n5348 VDD.n341 4.91801
R9851 VDD.n380 VDD.n377 4.91801
R9852 VDD.n490 VDD.n438 4.91801
R9853 VDD.n545 VDD.n544 4.91801
R9854 VDD.n593 VDD.n590 4.91801
R9855 VDD.n5222 VDD.n632 4.91801
R9856 VDD.n5172 VDD.n5171 4.91801
R9857 VDD.n3786 VDD.n3785 4.89462
R9858 VDD.n2940 VDD.n2920 4.89462
R9859 VDD.n2584 VDD.n2583 4.89462
R9860 VDD.n2557 VDD.n2556 4.89462
R9861 VDD.n2621 VDD.n2602 4.894
R9862 VDD.n5440 VDD.n274 4.89039
R9863 VDD.n5445 VDD.n5440 4.89039
R9864 VDD.n5402 VDD.n5401 4.8457
R9865 VDD.n5354 VDD.n337 4.8457
R9866 VDD.n5304 VDD.n5303 4.8457
R9867 VDD.n484 VDD.n483 4.8457
R9868 VDD.n543 VDD.n416 4.8457
R9869 VDD.n5271 VDD.n5270 4.8457
R9870 VDD.n5223 VDD.n629 4.8457
R9871 VDD.n671 VDD.n670 4.8457
R9872 VDD.n2585 VDD.n2509 4.78705
R9873 VDD.n8819 VDD.n8818 4.78659
R9874 VDD.n7964 VDD.n7963 4.78659
R9875 VDD.n7110 VDD.n7109 4.78659
R9876 VDD.n6255 VDD.n6254 4.78659
R9877 VDD.n1484 VDD.n1375 4.7505
R9878 VDD.n1486 VDD.n1485 4.7505
R9879 VDD.n1496 VDD.n1369 4.7505
R9880 VDD.n1497 VDD.n1364 4.7505
R9881 VDD.n1502 VDD.n1500 4.7505
R9882 VDD.n1501 VDD.n1358 4.7505
R9883 VDD.n1513 VDD.n1512 4.7505
R9884 VDD.n1516 VDD.n1353 4.7505
R9885 VDD.n1518 VDD.n1517 4.7505
R9886 VDD.n1528 VDD.n1347 4.7505
R9887 VDD.n1530 VDD.n1529 4.7505
R9888 VDD.n1540 VDD.n1341 4.7505
R9889 VDD.n1541 VDD.n1336 4.7505
R9890 VDD.n1546 VDD.n1544 4.7505
R9891 VDD.n1545 VDD.n1330 4.7505
R9892 VDD.n1557 VDD.n1556 4.7505
R9893 VDD.n1560 VDD.n1325 4.7505
R9894 VDD.n1562 VDD.n1561 4.7505
R9895 VDD.n1571 VDD.n1318 4.7505
R9896 VDD.n1572 VDD.n1313 4.7505
R9897 VDD.n1577 VDD.n1575 4.7505
R9898 VDD.n1576 VDD.n1307 4.7505
R9899 VDD.n1588 VDD.n1587 4.7505
R9900 VDD.n1591 VDD.n1302 4.7505
R9901 VDD.n1593 VDD.n1592 4.7505
R9902 VDD.n1603 VDD.n1296 4.7505
R9903 VDD.n1605 VDD.n1604 4.7505
R9904 VDD.n1615 VDD.n1290 4.7505
R9905 VDD.n1617 VDD.n1616 4.7505
R9906 VDD.n1622 VDD.n1277 4.7505
R9907 VDD.n1805 VDD.n1804 4.7505
R9908 VDD.n1801 VDD.n1623 4.7505
R9909 VDD.n1800 VDD.n1628 4.7505
R9910 VDD.n1638 VDD.n1637 4.7505
R9911 VDD.n1790 VDD.n1789 4.7505
R9912 VDD.n1786 VDD.n1639 4.7505
R9913 VDD.n1785 VDD.n1645 4.7505
R9914 VDD.n1654 VDD.n1653 4.7505
R9915 VDD.n1776 VDD.n1775 4.7505
R9916 VDD.n1772 VDD.n1655 4.7505
R9917 VDD.n1771 VDD.n1661 4.7505
R9918 VDD.n1671 VDD.n1670 4.7505
R9919 VDD.n1761 VDD.n1760 4.7505
R9920 VDD.n1757 VDD.n1672 4.7505
R9921 VDD.n1756 VDD.n1678 4.7505
R9922 VDD.n1688 VDD.n1687 4.7505
R9923 VDD.n1746 VDD.n1745 4.7505
R9924 VDD.n1742 VDD.n1689 4.7505
R9925 VDD.n1741 VDD.n1695 4.7505
R9926 VDD.n1727 VDD.n1726 4.7505
R9927 VDD.n1731 VDD.n1730 4.7505
R9928 VDD.n3504 VDD.n3503 4.73575
R9929 VDD.n3519 VDD.n3505 4.73575
R9930 VDD.n3206 VDD.n3205 4.73575
R9931 VDD.n3221 VDD.n3207 4.73575
R9932 VDD.n3754 VDD.n3753 4.73575
R9933 VDD.n3832 VDD.n3831 4.73575
R9934 VDD.n3852 VDD.n3851 4.73575
R9935 VDD.n3889 VDD.n3875 4.73575
R9936 VDD.n3855 VDD.n3854 4.73575
R9937 VDD.n3874 VDD.n3873 4.73575
R9938 VDD.n2834 VDD.n2833 4.73575
R9939 VDD.n2976 VDD.n2975 4.73575
R9940 VDD.n8643 VDD.n8642 4.73093
R9941 VDD.n8642 VDD.n8636 4.73093
R9942 VDD.n8636 VDD.n8500 4.73093
R9943 VDD.n8651 VDD.n8500 4.73093
R9944 VDD.n8652 VDD.n8651 4.73093
R9945 VDD.n8653 VDD.n8652 4.73093
R9946 VDD.n8653 VDD.n8496 4.73093
R9947 VDD.n8659 VDD.n8496 4.73093
R9948 VDD.n8660 VDD.n8659 4.73093
R9949 VDD.n8661 VDD.n8660 4.73093
R9950 VDD.n8661 VDD.n8492 4.73093
R9951 VDD.n8667 VDD.n8492 4.73093
R9952 VDD.n8668 VDD.n8667 4.73093
R9953 VDD.n8669 VDD.n8668 4.73093
R9954 VDD.n8669 VDD.n8488 4.73093
R9955 VDD.n8676 VDD.n8488 4.73093
R9956 VDD.n8677 VDD.n8676 4.73093
R9957 VDD.n7788 VDD.n7787 4.73093
R9958 VDD.n7787 VDD.n7781 4.73093
R9959 VDD.n7781 VDD.n7645 4.73093
R9960 VDD.n7796 VDD.n7645 4.73093
R9961 VDD.n7797 VDD.n7796 4.73093
R9962 VDD.n7798 VDD.n7797 4.73093
R9963 VDD.n7798 VDD.n7641 4.73093
R9964 VDD.n7804 VDD.n7641 4.73093
R9965 VDD.n7805 VDD.n7804 4.73093
R9966 VDD.n7806 VDD.n7805 4.73093
R9967 VDD.n7806 VDD.n7637 4.73093
R9968 VDD.n7812 VDD.n7637 4.73093
R9969 VDD.n7813 VDD.n7812 4.73093
R9970 VDD.n7814 VDD.n7813 4.73093
R9971 VDD.n7814 VDD.n7633 4.73093
R9972 VDD.n7821 VDD.n7633 4.73093
R9973 VDD.n7822 VDD.n7821 4.73093
R9974 VDD.n6934 VDD.n6933 4.73093
R9975 VDD.n6933 VDD.n6927 4.73093
R9976 VDD.n6927 VDD.n6791 4.73093
R9977 VDD.n6942 VDD.n6791 4.73093
R9978 VDD.n6943 VDD.n6942 4.73093
R9979 VDD.n6944 VDD.n6943 4.73093
R9980 VDD.n6944 VDD.n6787 4.73093
R9981 VDD.n6950 VDD.n6787 4.73093
R9982 VDD.n6951 VDD.n6950 4.73093
R9983 VDD.n6952 VDD.n6951 4.73093
R9984 VDD.n6952 VDD.n6783 4.73093
R9985 VDD.n6958 VDD.n6783 4.73093
R9986 VDD.n6959 VDD.n6958 4.73093
R9987 VDD.n6960 VDD.n6959 4.73093
R9988 VDD.n6960 VDD.n6779 4.73093
R9989 VDD.n6967 VDD.n6779 4.73093
R9990 VDD.n6968 VDD.n6967 4.73093
R9991 VDD.n6079 VDD.n6078 4.73093
R9992 VDD.n6078 VDD.n6072 4.73093
R9993 VDD.n6072 VDD.n5936 4.73093
R9994 VDD.n6087 VDD.n5936 4.73093
R9995 VDD.n6088 VDD.n6087 4.73093
R9996 VDD.n6089 VDD.n6088 4.73093
R9997 VDD.n6089 VDD.n5932 4.73093
R9998 VDD.n6095 VDD.n5932 4.73093
R9999 VDD.n6096 VDD.n6095 4.73093
R10000 VDD.n6097 VDD.n6096 4.73093
R10001 VDD.n6097 VDD.n5928 4.73093
R10002 VDD.n6103 VDD.n5928 4.73093
R10003 VDD.n6104 VDD.n6103 4.73093
R10004 VDD.n6105 VDD.n6104 4.73093
R10005 VDD.n6105 VDD.n5924 4.73093
R10006 VDD.n6112 VDD.n5924 4.73093
R10007 VDD.n6113 VDD.n6112 4.73093
R10008 VDD.n1876 VDD.n1050 4.70536
R10009 VDD.n5398 VDD.n5397 4.70106
R10010 VDD.n5347 VDD.n342 4.70106
R10011 VDD.n5300 VDD.n5299 4.70106
R10012 VDD.n491 VDD.n436 4.70106
R10013 VDD.n550 VDD.n414 4.70106
R10014 VDD.n5267 VDD.n5266 4.70106
R10015 VDD.n5216 VDD.n636 4.70106
R10016 VDD.n5170 VDD.n672 4.70106
R10017 VDD.n5629 VDD.n5628 4.6533
R10018 VDD.n6486 VDD.n6485 4.6533
R10019 VDD.n7338 VDD.n7337 4.6533
R10020 VDD.n8195 VDD.n8194 4.6533
R10021 VDD.n5663 VDD.n5649 4.6505
R10022 VDD.n5662 VDD.n5661 4.6505
R10023 VDD.n5660 VDD.n5651 4.6505
R10024 VDD.n5659 VDD.n5658 4.6505
R10025 VDD.n5632 VDD.n5620 4.6505
R10026 VDD.n5639 VDD.n5638 4.6505
R10027 VDD.n5623 VDD.n5616 4.6505
R10028 VDD VDD.n5670 4.6505
R10029 VDD.n5622 VDD.n5615 4.6505
R10030 VDD.n5625 VDD.n5622 4.6505
R10031 VDD.n5631 VDD.n5630 4.6505
R10032 VDD.n6514 VDD.n6511 4.6505
R10033 VDD.n6513 VDD.n6512 4.6505
R10034 VDD.n6468 VDD.n6467 4.6505
R10035 VDD.n6520 VDD.n6519 4.6505
R10036 VDD.n6481 VDD.n6477 4.6505
R10037 VDD.n6492 VDD.n6491 4.6505
R10038 VDD.n6498 VDD.n6472 4.6505
R10039 VDD.n6502 VDD 4.6505
R10040 VDD.n6501 VDD.n6500 4.6505
R10041 VDD.n6500 VDD.n6474 4.6505
R10042 VDD.n6480 VDD.n6479 4.6505
R10043 VDD.n7372 VDD.n7358 4.6505
R10044 VDD.n7371 VDD.n7370 4.6505
R10045 VDD.n7369 VDD.n7360 4.6505
R10046 VDD.n7368 VDD.n7367 4.6505
R10047 VDD.n7341 VDD.n7329 4.6505
R10048 VDD.n7348 VDD.n7347 4.6505
R10049 VDD.n7332 VDD.n7325 4.6505
R10050 VDD VDD.n7379 4.6505
R10051 VDD.n7331 VDD.n7324 4.6505
R10052 VDD.n7334 VDD.n7331 4.6505
R10053 VDD.n7340 VDD.n7339 4.6505
R10054 VDD.n8223 VDD.n8220 4.6505
R10055 VDD.n8222 VDD.n8221 4.6505
R10056 VDD.n8177 VDD.n8176 4.6505
R10057 VDD.n8229 VDD.n8228 4.6505
R10058 VDD.n8190 VDD.n8186 4.6505
R10059 VDD.n8201 VDD.n8200 4.6505
R10060 VDD.n8207 VDD.n8181 4.6505
R10061 VDD.n8211 VDD 4.6505
R10062 VDD.n8210 VDD.n8209 4.6505
R10063 VDD.n8209 VDD.n8183 4.6505
R10064 VDD.n8189 VDD.n8188 4.6505
R10065 VDD.n3868 VDD.n3867 4.6505
R10066 VDD.n3846 VDD.n3845 4.6505
R10067 VDD.n2355 VDD.n2344 4.6505
R10068 VDD.n5456 VDD.n5455 4.6505
R10069 VDD.n4291 VDD.n4290 4.6505
R10070 VDD.n2370 VDD.n2363 4.6505
R10071 VDD.n4282 VDD.n4281 4.6505
R10072 VDD.n4280 VDD.n4279 4.6505
R10073 VDD.n2373 VDD.n2372 4.6505
R10074 VDD.n2380 VDD.n2378 4.6505
R10075 VDD.n4271 VDD.n4270 4.6505
R10076 VDD.n4269 VDD.n4268 4.6505
R10077 VDD.n2382 VDD.n2381 4.6505
R10078 VDD.n2389 VDD.n2387 4.6505
R10079 VDD.n4260 VDD.n4259 4.6505
R10080 VDD.n4258 VDD.n4257 4.6505
R10081 VDD.n2391 VDD.n2390 4.6505
R10082 VDD.n2398 VDD.n2396 4.6505
R10083 VDD.n4249 VDD.n4248 4.6505
R10084 VDD.n4247 VDD.n4246 4.6505
R10085 VDD.n2400 VDD.n2399 4.6505
R10086 VDD.n2406 VDD.n2404 4.6505
R10087 VDD.n4237 VDD.n4236 4.6505
R10088 VDD.n4235 VDD.n4234 4.6505
R10089 VDD.n2408 VDD.n2407 4.6505
R10090 VDD.n2418 VDD.n2416 4.6505
R10091 VDD.n4226 VDD.n4225 4.6505
R10092 VDD.n4224 VDD.n4223 4.6505
R10093 VDD.n2420 VDD.n2419 4.6505
R10094 VDD.n2427 VDD.n2425 4.6505
R10095 VDD.n4215 VDD.n4214 4.6505
R10096 VDD.n4213 VDD.n4212 4.6505
R10097 VDD.n2429 VDD.n2428 4.6505
R10098 VDD.n2436 VDD.n2434 4.6505
R10099 VDD.n4204 VDD.n4203 4.6505
R10100 VDD.n4202 VDD.n4201 4.6505
R10101 VDD.n4085 VDD.n2437 4.6505
R10102 VDD.n4088 VDD.n4087 4.6505
R10103 VDD.n4090 VDD.n4089 4.6505
R10104 VDD.n4080 VDD.n4079 4.6505
R10105 VDD.n4101 VDD.n4100 4.6505
R10106 VDD.n4102 VDD.n4077 4.6505
R10107 VDD.n4104 VDD.n4103 4.6505
R10108 VDD.n4073 VDD.n4072 4.6505
R10109 VDD.n4114 VDD.n4113 4.6505
R10110 VDD.n4115 VDD.n4070 4.6505
R10111 VDD.n4117 VDD.n4116 4.6505
R10112 VDD.n4066 VDD.n4065 4.6505
R10113 VDD.n4128 VDD.n4127 4.6505
R10114 VDD.n4129 VDD.n4063 4.6505
R10115 VDD.n4131 VDD.n4130 4.6505
R10116 VDD.n4060 VDD.n4059 4.6505
R10117 VDD.n4140 VDD.n4139 4.6505
R10118 VDD.n4142 VDD.n4141 4.6505
R10119 VDD.n4143 VDD.n4052 4.6505
R10120 VDD.n4152 VDD.n4151 4.6505
R10121 VDD.n4153 VDD.n4050 4.6505
R10122 VDD.n4155 VDD.n4154 4.6505
R10123 VDD.n4046 VDD.n4045 4.6505
R10124 VDD.n4165 VDD.n4164 4.6505
R10125 VDD.n4166 VDD.n4043 4.6505
R10126 VDD.n4168 VDD.n4167 4.6505
R10127 VDD.n4039 VDD.n4038 4.6505
R10128 VDD.n4178 VDD.n4177 4.6505
R10129 VDD.n4179 VDD.n4036 4.6505
R10130 VDD.n4181 VDD.n4180 4.6505
R10131 VDD.n4031 VDD.n4030 4.6505
R10132 VDD.n4191 VDD.n4190 4.6505
R10133 VDD.n4193 VDD.n4192 4.6505
R10134 VDD.n275 VDD.n273 4.6505
R10135 VDD.n4293 VDD.n2362 4.6505
R10136 VDD.n1466 VDD.n1465 4.6505
R10137 VDD.n1464 VDD.n1463 4.6505
R10138 VDD.n1406 VDD.n1402 4.6505
R10139 VDD.n1455 VDD.n1454 4.6505
R10140 VDD.n1453 VDD.n1452 4.6505
R10141 VDD.n1445 VDD.n1408 4.6505
R10142 VDD.n1413 VDD.n1411 4.6505
R10143 VDD.n1437 VDD.n1436 4.6505
R10144 VDD.n1435 VDD.n1434 4.6505
R10145 VDD.n1427 VDD.n1414 4.6505
R10146 VDD.n1420 VDD.n1419 4.6505
R10147 VDD.n1418 VDD.n1387 4.6505
R10148 VDD.n1388 VDD.n1027 4.6505
R10149 VDD.n1898 VDD.n1897 4.6505
R10150 VDD.n1899 VDD.n1005 4.6505
R10151 VDD.n1900 VDD.n1006 4.6505
R10152 VDD.n1902 VDD.n1901 4.6505
R10153 VDD.n1903 VDD.n1023 4.6505
R10154 VDD.n4561 VDD.n4560 4.6505
R10155 VDD.n4559 VDD.n4558 4.6505
R10156 VDD.n1914 VDD.n1024 4.6505
R10157 VDD.n1933 VDD.n1932 4.6505
R10158 VDD.n1934 VDD.n1928 4.6505
R10159 VDD.n4542 VDD.n4541 4.6505
R10160 VDD.n4540 VDD.n4539 4.6505
R10161 VDD.n1945 VDD.n1929 4.6505
R10162 VDD.n1968 VDD.n1967 4.6505
R10163 VDD.n1973 VDD.n1972 4.6505
R10164 VDD.n1974 VDD.n1957 4.6505
R10165 VDD.n4517 VDD.n4516 4.6505
R10166 VDD.n4515 VDD.n4514 4.6505
R10167 VDD.n1983 VDD.n1975 4.6505
R10168 VDD.n2005 VDD.n2004 4.6505
R10169 VDD.n2006 VDD.n2000 4.6505
R10170 VDD.n4498 VDD.n4497 4.6505
R10171 VDD.n4496 VDD.n4495 4.6505
R10172 VDD.n2018 VDD.n2001 4.6505
R10173 VDD.n2038 VDD.n2037 4.6505
R10174 VDD.n2039 VDD.n2033 4.6505
R10175 VDD.n4479 VDD.n4478 4.6505
R10176 VDD.n4477 VDD.n4476 4.6505
R10177 VDD.n2050 VDD.n2034 4.6505
R10178 VDD.n2085 VDD.n2084 4.6505
R10179 VDD.n2086 VDD.n2062 4.6505
R10180 VDD.n4460 VDD.n4459 4.6505
R10181 VDD.n4458 VDD.n4457 4.6505
R10182 VDD.n2078 VDD.n2063 4.6505
R10183 VDD.n4445 VDD.n4444 4.6505
R10184 VDD.n4443 VDD.n4442 4.6505
R10185 VDD.n2103 VDD.n2081 4.6505
R10186 VDD.n2122 VDD.n2121 4.6505
R10187 VDD.n2123 VDD.n2117 4.6505
R10188 VDD.n4426 VDD.n4425 4.6505
R10189 VDD.n4424 VDD.n4423 4.6505
R10190 VDD.n2133 VDD.n2118 4.6505
R10191 VDD.n2153 VDD.n2152 4.6505
R10192 VDD.n2154 VDD.n2148 4.6505
R10193 VDD.n4407 VDD.n4406 4.6505
R10194 VDD.n4405 VDD.n4404 4.6505
R10195 VDD.n2165 VDD.n2149 4.6505
R10196 VDD.n2189 VDD.n2188 4.6505
R10197 VDD.n2194 VDD.n2193 4.6505
R10198 VDD.n2195 VDD.n2178 4.6505
R10199 VDD.n4382 VDD.n4381 4.6505
R10200 VDD.n4380 VDD.n4379 4.6505
R10201 VDD.n2204 VDD.n2196 4.6505
R10202 VDD.n2226 VDD.n2225 4.6505
R10203 VDD.n2227 VDD.n2221 4.6505
R10204 VDD.n4363 VDD.n4362 4.6505
R10205 VDD.n4361 VDD.n4360 4.6505
R10206 VDD.n2224 VDD.n2222 4.6505
R10207 VDD.n1491 VDD.n1490 4.6505
R10208 VDD.n1493 VDD.n1492 4.6505
R10209 VDD.n1366 VDD.n1361 4.6505
R10210 VDD.n1507 VDD.n1506 4.6505
R10211 VDD.n1509 VDD.n1508 4.6505
R10212 VDD.n1356 VDD.n1350 4.6505
R10213 VDD.n1522 VDD.n1521 4.6505
R10214 VDD.n1524 VDD.n1523 4.6505
R10215 VDD.n1345 VDD.n1344 4.6505
R10216 VDD.n1535 VDD.n1534 4.6505
R10217 VDD.n1537 VDD.n1536 4.6505
R10218 VDD.n1338 VDD.n1333 4.6505
R10219 VDD.n1551 VDD.n1550 4.6505
R10220 VDD.n1553 VDD.n1552 4.6505
R10221 VDD.n1328 VDD.n1321 4.6505
R10222 VDD.n1566 VDD.n1565 4.6505
R10223 VDD.n1568 VDD.n1567 4.6505
R10224 VDD.n1316 VDD.n1310 4.6505
R10225 VDD.n1582 VDD.n1581 4.6505
R10226 VDD.n1584 VDD.n1583 4.6505
R10227 VDD.n1305 VDD.n1299 4.6505
R10228 VDD.n1597 VDD.n1596 4.6505
R10229 VDD.n1599 VDD.n1598 4.6505
R10230 VDD.n1294 VDD.n1293 4.6505
R10231 VDD.n1610 VDD.n1609 4.6505
R10232 VDD.n1612 VDD.n1611 4.6505
R10233 VDD.n1287 VDD.n1282 4.6505
R10234 VDD.n1811 VDD.n1810 4.6505
R10235 VDD.n1809 VDD.n1808 4.6505
R10236 VDD.n1625 VDD.n1283 4.6505
R10237 VDD.n1632 VDD.n1630 4.6505
R10238 VDD.n1796 VDD.n1795 4.6505
R10239 VDD.n1794 VDD.n1793 4.6505
R10240 VDD.n1643 VDD.n1633 4.6505
R10241 VDD.n1782 VDD.n1781 4.6505
R10242 VDD.n1780 VDD.n1779 4.6505
R10243 VDD.n1658 VDD.n1648 4.6505
R10244 VDD.n1665 VDD.n1663 4.6505
R10245 VDD.n1767 VDD.n1766 4.6505
R10246 VDD.n1765 VDD.n1764 4.6505
R10247 VDD.n1675 VDD.n1666 4.6505
R10248 VDD.n1682 VDD.n1680 4.6505
R10249 VDD.n1752 VDD.n1751 4.6505
R10250 VDD.n1750 VDD.n1749 4.6505
R10251 VDD.n1692 VDD.n1683 4.6505
R10252 VDD.n1699 VDD.n1697 4.6505
R10253 VDD.n1737 VDD.n1736 4.6505
R10254 VDD.n1735 VDD.n1734 4.6505
R10255 VDD.n1703 VDD.n1700 4.6505
R10256 VDD.n1048 VDD.n1046 4.6505
R10257 VDD.n1377 VDD.n1372 4.6505
R10258 VDD.n1880 VDD.n1879 4.6505
R10259 VDD.n1878 VDD.n1877 4.6505
R10260 VDD.n1054 VDD.n1049 4.6505
R10261 VDD.n1869 VDD.n1868 4.6505
R10262 VDD.n1867 VDD.n1866 4.6505
R10263 VDD.n1062 VDD.n1056 4.6505
R10264 VDD.n1852 VDD.n1851 4.6505
R10265 VDD.n1850 VDD.n1849 4.6505
R10266 VDD.n1066 VDD.n1065 4.6505
R10267 VDD.n1843 VDD.n1842 4.6505
R10268 VDD.n1841 VDD.n1840 4.6505
R10269 VDD.n1076 VDD.n1071 4.6505
R10270 VDD.n1832 VDD.n1831 4.6505
R10271 VDD.n1830 VDD.n1829 4.6505
R10272 VDD.n1079 VDD.n1078 4.6505
R10273 VDD.n1823 VDD.n1822 4.6505
R10274 VDD.n1821 VDD.n1820 4.6505
R10275 VDD.n1085 VDD.n1084 4.6505
R10276 VDD.n1274 VDD.n1273 4.6505
R10277 VDD.n1272 VDD.n1089 4.6505
R10278 VDD.n1269 VDD.n1090 4.6505
R10279 VDD.n1267 VDD.n1266 4.6505
R10280 VDD.n1265 VDD.n1264 4.6505
R10281 VDD.n1093 VDD.n1092 4.6505
R10282 VDD.n1258 VDD.n1257 4.6505
R10283 VDD.n1256 VDD.n1255 4.6505
R10284 VDD.n1100 VDD.n1099 4.6505
R10285 VDD.n1249 VDD.n1248 4.6505
R10286 VDD.n1247 VDD.n1246 4.6505
R10287 VDD.n1106 VDD.n1105 4.6505
R10288 VDD.n1240 VDD.n1111 4.6505
R10289 VDD.n1115 VDD.n1113 4.6505
R10290 VDD.n1233 VDD.n1232 4.6505
R10291 VDD.n1231 VDD.n1230 4.6505
R10292 VDD.n1117 VDD.n1116 4.6505
R10293 VDD.n1224 VDD.n1223 4.6505
R10294 VDD.n1222 VDD.n1221 4.6505
R10295 VDD.n1123 VDD.n1122 4.6505
R10296 VDD.n1215 VDD.n1214 4.6505
R10297 VDD.n1213 VDD.n1212 4.6505
R10298 VDD.n1129 VDD.n1128 4.6505
R10299 VDD.n1206 VDD.n1205 4.6505
R10300 VDD.n1204 VDD.n1203 4.6505
R10301 VDD.n1135 VDD.n1134 4.6505
R10302 VDD.n1197 VDD.n1196 4.6505
R10303 VDD.n1195 VDD.n1194 4.6505
R10304 VDD.n1141 VDD.n1140 4.6505
R10305 VDD.n1188 VDD.n1146 4.6505
R10306 VDD.n1150 VDD.n1148 4.6505
R10307 VDD.n1181 VDD.n1180 4.6505
R10308 VDD.n1179 VDD.n1178 4.6505
R10309 VDD.n1152 VDD.n1151 4.6505
R10310 VDD.n1172 VDD.n1171 4.6505
R10311 VDD.n1170 VDD.n1169 4.6505
R10312 VDD.n1158 VDD.n1157 4.6505
R10313 VDD.n1163 VDD.n1162 4.6505
R10314 VDD.n999 VDD.n998 4.6505
R10315 VDD.n4584 VDD.n4583 4.6505
R10316 VDD.n4585 VDD.n996 4.6505
R10317 VDD.n4587 VDD.n4586 4.6505
R10318 VDD.n992 VDD.n991 4.6505
R10319 VDD.n4596 VDD.n4595 4.6505
R10320 VDD.n4598 VDD.n4597 4.6505
R10321 VDD.n4599 VDD.n984 4.6505
R10322 VDD.n4607 VDD.n4606 4.6505
R10323 VDD.n4608 VDD.n982 4.6505
R10324 VDD.n4610 VDD.n4609 4.6505
R10325 VDD.n978 VDD.n977 4.6505
R10326 VDD.n4620 VDD.n4619 4.6505
R10327 VDD.n4621 VDD.n975 4.6505
R10328 VDD.n4623 VDD.n4622 4.6505
R10329 VDD.n971 VDD.n970 4.6505
R10330 VDD.n4633 VDD.n4632 4.6505
R10331 VDD.n4634 VDD.n968 4.6505
R10332 VDD.n4636 VDD.n4635 4.6505
R10333 VDD.n964 VDD.n963 4.6505
R10334 VDD.n4646 VDD.n4645 4.6505
R10335 VDD.n4647 VDD.n961 4.6505
R10336 VDD.n4649 VDD.n4648 4.6505
R10337 VDD.n957 VDD.n956 4.6505
R10338 VDD.n4658 VDD.n4657 4.6505
R10339 VDD.n4660 VDD.n4659 4.6505
R10340 VDD.n950 VDD.n949 4.6505
R10341 VDD.n4669 VDD.n4668 4.6505
R10342 VDD.n4670 VDD.n947 4.6505
R10343 VDD.n4672 VDD.n4671 4.6505
R10344 VDD.n943 VDD.n942 4.6505
R10345 VDD.n4682 VDD.n4681 4.6505
R10346 VDD.n4683 VDD.n940 4.6505
R10347 VDD.n4685 VDD.n4684 4.6505
R10348 VDD.n936 VDD.n935 4.6505
R10349 VDD.n4695 VDD.n4694 4.6505
R10350 VDD.n4696 VDD.n933 4.6505
R10351 VDD.n4698 VDD.n4697 4.6505
R10352 VDD.n929 VDD.n928 4.6505
R10353 VDD.n4707 VDD.n4706 4.6505
R10354 VDD.n4709 VDD.n4708 4.6505
R10355 VDD.n4711 VDD.n917 4.6505
R10356 VDD.n5157 VDD.n5156 4.6505
R10357 VDD.n5155 VDD.n5154 4.6505
R10358 VDD.n5145 VDD.n682 4.6505
R10359 VDD.n5144 VDD.n5143 4.6505
R10360 VDD.n5142 VDD.n5141 4.6505
R10361 VDD.n690 VDD.n689 4.6505
R10362 VDD.n5133 VDD.n5132 4.6505
R10363 VDD.n5131 VDD.n694 4.6505
R10364 VDD.n5130 VDD.n5129 4.6505
R10365 VDD.n697 VDD.n696 4.6505
R10366 VDD.n5120 VDD.n5119 4.6505
R10367 VDD.n5118 VDD.n701 4.6505
R10368 VDD.n5117 VDD.n5116 4.6505
R10369 VDD.n704 VDD.n703 4.6505
R10370 VDD.n5107 VDD.n5106 4.6505
R10371 VDD.n5105 VDD.n708 4.6505
R10372 VDD.n5104 VDD.n5103 4.6505
R10373 VDD.n711 VDD.n710 4.6505
R10374 VDD.n5094 VDD.n5093 4.6505
R10375 VDD.n5092 VDD.n5091 4.6505
R10376 VDD.n718 VDD.n717 4.6505
R10377 VDD.n5083 VDD.n5082 4.6505
R10378 VDD.n5081 VDD.n722 4.6505
R10379 VDD.n5080 VDD.n5079 4.6505
R10380 VDD.n725 VDD.n724 4.6505
R10381 VDD.n5070 VDD.n5069 4.6505
R10382 VDD.n5068 VDD.n729 4.6505
R10383 VDD.n5067 VDD.n5066 4.6505
R10384 VDD.n732 VDD.n731 4.6505
R10385 VDD.n5057 VDD.n5056 4.6505
R10386 VDD.n5055 VDD.n736 4.6505
R10387 VDD.n5054 VDD.n5053 4.6505
R10388 VDD.n739 VDD.n738 4.6505
R10389 VDD.n5044 VDD.n5043 4.6505
R10390 VDD.n5042 VDD.n743 4.6505
R10391 VDD.n5041 VDD.n5040 4.6505
R10392 VDD.n5031 VDD.n745 4.6505
R10393 VDD.n5030 VDD.n5029 4.6505
R10394 VDD.n5028 VDD.n5027 4.6505
R10395 VDD.n752 VDD.n751 4.6505
R10396 VDD.n5019 VDD.n5018 4.6505
R10397 VDD.n5017 VDD.n756 4.6505
R10398 VDD.n5016 VDD.n5015 4.6505
R10399 VDD.n759 VDD.n758 4.6505
R10400 VDD.n5006 VDD.n5005 4.6505
R10401 VDD.n5004 VDD.n763 4.6505
R10402 VDD.n5003 VDD.n5002 4.6505
R10403 VDD.n766 VDD.n765 4.6505
R10404 VDD.n4993 VDD.n4992 4.6505
R10405 VDD.n4991 VDD.n770 4.6505
R10406 VDD.n4990 VDD.n4989 4.6505
R10407 VDD.n773 VDD.n772 4.6505
R10408 VDD.n4980 VDD.n4979 4.6505
R10409 VDD.n4978 VDD.n4977 4.6505
R10410 VDD.n780 VDD.n779 4.6505
R10411 VDD.n4969 VDD.n4968 4.6505
R10412 VDD.n4967 VDD.n784 4.6505
R10413 VDD.n4966 VDD.n4965 4.6505
R10414 VDD.n787 VDD.n786 4.6505
R10415 VDD.n4956 VDD.n4955 4.6505
R10416 VDD.n4954 VDD.n791 4.6505
R10417 VDD.n4953 VDD.n4952 4.6505
R10418 VDD.n794 VDD.n793 4.6505
R10419 VDD.n4943 VDD.n4942 4.6505
R10420 VDD.n4941 VDD.n798 4.6505
R10421 VDD.n4940 VDD.n4939 4.6505
R10422 VDD.n801 VDD.n800 4.6505
R10423 VDD.n4930 VDD.n4929 4.6505
R10424 VDD.n4928 VDD.n805 4.6505
R10425 VDD.n4927 VDD.n4926 4.6505
R10426 VDD.n4917 VDD.n807 4.6505
R10427 VDD.n4916 VDD.n4915 4.6505
R10428 VDD.n4914 VDD.n4913 4.6505
R10429 VDD.n814 VDD.n813 4.6505
R10430 VDD.n4905 VDD.n4904 4.6505
R10431 VDD.n4903 VDD.n818 4.6505
R10432 VDD.n4902 VDD.n4901 4.6505
R10433 VDD.n821 VDD.n820 4.6505
R10434 VDD.n4892 VDD.n4891 4.6505
R10435 VDD.n4890 VDD.n825 4.6505
R10436 VDD.n4889 VDD.n4888 4.6505
R10437 VDD.n828 VDD.n827 4.6505
R10438 VDD.n4879 VDD.n4878 4.6505
R10439 VDD.n4877 VDD.n832 4.6505
R10440 VDD.n4876 VDD.n4875 4.6505
R10441 VDD.n835 VDD.n834 4.6505
R10442 VDD.n4866 VDD.n4865 4.6505
R10443 VDD.n4864 VDD.n4863 4.6505
R10444 VDD.n842 VDD.n841 4.6505
R10445 VDD.n4855 VDD.n4854 4.6505
R10446 VDD.n4853 VDD.n846 4.6505
R10447 VDD.n4852 VDD.n4851 4.6505
R10448 VDD.n849 VDD.n848 4.6505
R10449 VDD.n4842 VDD.n4841 4.6505
R10450 VDD.n4840 VDD.n853 4.6505
R10451 VDD.n4839 VDD.n4838 4.6505
R10452 VDD.n856 VDD.n855 4.6505
R10453 VDD.n4829 VDD.n4828 4.6505
R10454 VDD.n4827 VDD.n860 4.6505
R10455 VDD.n4826 VDD.n4825 4.6505
R10456 VDD.n863 VDD.n862 4.6505
R10457 VDD.n4816 VDD.n4815 4.6505
R10458 VDD.n4814 VDD.n867 4.6505
R10459 VDD.n4813 VDD.n4812 4.6505
R10460 VDD.n4803 VDD.n869 4.6505
R10461 VDD.n4802 VDD.n4801 4.6505
R10462 VDD.n4800 VDD.n4799 4.6505
R10463 VDD.n876 VDD.n875 4.6505
R10464 VDD.n4791 VDD.n4790 4.6505
R10465 VDD.n4789 VDD.n880 4.6505
R10466 VDD.n4788 VDD.n4787 4.6505
R10467 VDD.n883 VDD.n882 4.6505
R10468 VDD.n4778 VDD.n4777 4.6505
R10469 VDD.n4776 VDD.n887 4.6505
R10470 VDD.n4775 VDD.n4774 4.6505
R10471 VDD.n890 VDD.n889 4.6505
R10472 VDD.n4765 VDD.n4764 4.6505
R10473 VDD.n4763 VDD.n894 4.6505
R10474 VDD.n4762 VDD.n4761 4.6505
R10475 VDD.n897 VDD.n896 4.6505
R10476 VDD.n4752 VDD.n4751 4.6505
R10477 VDD.n4750 VDD.n4749 4.6505
R10478 VDD.n904 VDD.n903 4.6505
R10479 VDD.n4741 VDD.n4740 4.6505
R10480 VDD.n4739 VDD.n908 4.6505
R10481 VDD.n4738 VDD.n4737 4.6505
R10482 VDD.n911 VDD.n910 4.6505
R10483 VDD.n4728 VDD.n4727 4.6505
R10484 VDD.n4726 VDD.n915 4.6505
R10485 VDD.n4725 VDD.n4724 4.6505
R10486 VDD.n278 VDD.n276 4.6505
R10487 VDD.n299 VDD.n297 4.6505
R10488 VDD.n5436 VDD.n5435 4.6505
R10489 VDD.n5434 VDD.n5433 4.6505
R10490 VDD.n5430 VDD.n300 4.6505
R10491 VDD.n303 VDD.n301 4.6505
R10492 VDD.n5425 VDD.n5424 4.6505
R10493 VDD.n5423 VDD.n5422 4.6505
R10494 VDD.n5418 VDD.n304 4.6505
R10495 VDD.n307 VDD.n305 4.6505
R10496 VDD.n5413 VDD.n5412 4.6505
R10497 VDD.n5411 VDD.n5410 4.6505
R10498 VDD.n5406 VDD.n308 4.6505
R10499 VDD.n311 VDD.n309 4.6505
R10500 VDD.n5401 VDD.n5400 4.6505
R10501 VDD.n5399 VDD.n5398 4.6505
R10502 VDD.n316 VDD.n312 4.6505
R10503 VDD.n5393 VDD.n5392 4.6505
R10504 VDD.n5391 VDD.n5390 4.6505
R10505 VDD.n5386 VDD.n318 4.6505
R10506 VDD.n321 VDD.n319 4.6505
R10507 VDD.n5381 VDD.n5380 4.6505
R10508 VDD.n5379 VDD.n5378 4.6505
R10509 VDD.n5374 VDD.n322 4.6505
R10510 VDD.n325 VDD.n323 4.6505
R10511 VDD.n5369 VDD.n5368 4.6505
R10512 VDD.n5367 VDD.n5366 4.6505
R10513 VDD.n327 VDD.n326 4.6505
R10514 VDD.n335 VDD.n333 4.6505
R10515 VDD.n5358 VDD.n5357 4.6505
R10516 VDD.n5356 VDD.n5355 4.6505
R10517 VDD.n337 VDD.n336 4.6505
R10518 VDD.n5347 VDD.n5346 4.6505
R10519 VDD.n5345 VDD.n5344 4.6505
R10520 VDD.n344 VDD.n343 4.6505
R10521 VDD.n351 VDD.n349 4.6505
R10522 VDD.n5336 VDD.n5335 4.6505
R10523 VDD.n5334 VDD.n5333 4.6505
R10524 VDD.n353 VDD.n352 4.6505
R10525 VDD.n360 VDD.n358 4.6505
R10526 VDD.n5325 VDD.n5324 4.6505
R10527 VDD.n5323 VDD.n5322 4.6505
R10528 VDD.n362 VDD.n361 4.6505
R10529 VDD.n369 VDD.n367 4.6505
R10530 VDD.n5314 VDD.n5313 4.6505
R10531 VDD.n5312 VDD.n5311 4.6505
R10532 VDD.n371 VDD.n370 4.6505
R10533 VDD.n378 VDD.n376 4.6505
R10534 VDD.n5303 VDD.n5302 4.6505
R10535 VDD.n5301 VDD.n5300 4.6505
R10536 VDD.n381 VDD.n379 4.6505
R10537 VDD.n390 VDD.n388 4.6505
R10538 VDD.n5292 VDD.n5291 4.6505
R10539 VDD.n5290 VDD.n5289 4.6505
R10540 VDD.n392 VDD.n391 4.6505
R10541 VDD.n454 VDD.n453 4.6505
R10542 VDD.n450 VDD.n449 4.6505
R10543 VDD.n461 VDD.n460 4.6505
R10544 VDD.n463 VDD.n462 4.6505
R10545 VDD.n446 VDD.n445 4.6505
R10546 VDD.n471 VDD.n470 4.6505
R10547 VDD.n473 VDD.n472 4.6505
R10548 VDD.n442 VDD.n441 4.6505
R10549 VDD.n480 VDD.n479 4.6505
R10550 VDD.n482 VDD.n481 4.6505
R10551 VDD.n483 VDD.n437 4.6505
R10552 VDD.n492 VDD.n491 4.6505
R10553 VDD.n494 VDD.n493 4.6505
R10554 VDD.n434 VDD.n433 4.6505
R10555 VDD.n502 VDD.n501 4.6505
R10556 VDD.n504 VDD.n503 4.6505
R10557 VDD.n430 VDD.n429 4.6505
R10558 VDD.n511 VDD.n510 4.6505
R10559 VDD.n513 VDD.n512 4.6505
R10560 VDD.n426 VDD.n425 4.6505
R10561 VDD.n521 VDD.n520 4.6505
R10562 VDD.n523 VDD.n522 4.6505
R10563 VDD.n422 VDD.n421 4.6505
R10564 VDD.n530 VDD.n529 4.6505
R10565 VDD.n532 VDD.n531 4.6505
R10566 VDD.n418 VDD.n417 4.6505
R10567 VDD.n541 VDD.n540 4.6505
R10568 VDD.n543 VDD.n542 4.6505
R10569 VDD.n414 VDD.n413 4.6505
R10570 VDD.n552 VDD.n551 4.6505
R10571 VDD.n554 VDD.n553 4.6505
R10572 VDD.n410 VDD.n409 4.6505
R10573 VDD.n561 VDD.n560 4.6505
R10574 VDD.n563 VDD.n562 4.6505
R10575 VDD.n406 VDD.n405 4.6505
R10576 VDD.n571 VDD.n570 4.6505
R10577 VDD.n573 VDD.n572 4.6505
R10578 VDD.n402 VDD.n401 4.6505
R10579 VDD.n581 VDD.n580 4.6505
R10580 VDD.n582 VDD.n399 4.6505
R10581 VDD.n5281 VDD.n5280 4.6505
R10582 VDD.n5279 VDD.n5278 4.6505
R10583 VDD.n584 VDD.n583 4.6505
R10584 VDD.n591 VDD.n589 4.6505
R10585 VDD.n5270 VDD.n5269 4.6505
R10586 VDD.n5268 VDD.n5267 4.6505
R10587 VDD.n594 VDD.n592 4.6505
R10588 VDD.n603 VDD.n601 4.6505
R10589 VDD.n5259 VDD.n5258 4.6505
R10590 VDD.n5257 VDD.n5256 4.6505
R10591 VDD.n605 VDD.n604 4.6505
R10592 VDD.n612 VDD.n610 4.6505
R10593 VDD.n5248 VDD.n5247 4.6505
R10594 VDD.n5246 VDD.n5245 4.6505
R10595 VDD.n614 VDD.n613 4.6505
R10596 VDD.n621 VDD.n619 4.6505
R10597 VDD.n5237 VDD.n5236 4.6505
R10598 VDD.n5235 VDD.n5234 4.6505
R10599 VDD.n623 VDD.n622 4.6505
R10600 VDD.n630 VDD.n628 4.6505
R10601 VDD.n5226 VDD.n5225 4.6505
R10602 VDD.n5224 VDD.n5223 4.6505
R10603 VDD.n636 VDD.n631 4.6505
R10604 VDD.n5215 VDD.n5214 4.6505
R10605 VDD.n5213 VDD.n5212 4.6505
R10606 VDD.n639 VDD.n638 4.6505
R10607 VDD.n646 VDD.n644 4.6505
R10608 VDD.n5204 VDD.n5203 4.6505
R10609 VDD.n5202 VDD.n5201 4.6505
R10610 VDD.n648 VDD.n647 4.6505
R10611 VDD.n655 VDD.n653 4.6505
R10612 VDD.n5193 VDD.n5192 4.6505
R10613 VDD.n5191 VDD.n5190 4.6505
R10614 VDD.n657 VDD.n656 4.6505
R10615 VDD.n664 VDD.n662 4.6505
R10616 VDD.n5182 VDD.n5181 4.6505
R10617 VDD.n5180 VDD.n5179 4.6505
R10618 VDD.n666 VDD.n665 4.6505
R10619 VDD.n5454 VDD.n5453 4.6505
R10620 VDD.n5170 VDD.n5169 4.6505
R10621 VDD.n5168 VDD.n5167 4.6505
R10622 VDD.n675 VDD.n674 4.6505
R10623 VDD.n673 VDD.n671 4.6505
R10624 VDD.n1877 VDD.n1047 4.63618
R10625 VDD.n4753 VDD.n901 4.60579
R10626 VDD.n4810 VDD.n870 4.60579
R10627 VDD.n4867 VDD.n839 4.60579
R10628 VDD.n4924 VDD.n808 4.60579
R10629 VDD.n4981 VDD.n777 4.60579
R10630 VDD.n5038 VDD.n746 4.60579
R10631 VDD.n5095 VDD.n715 4.60579
R10632 VDD.n5153 VDD.n683 4.60579
R10633 VDD.n1241 VDD.n1240 4.58155
R10634 VDD.n1240 VDD.n1110 4.58155
R10635 VDD.n1189 VDD.n1188 4.58155
R10636 VDD.n1188 VDD.n1145 4.58155
R10637 VDD.n4606 VDD.n985 4.58155
R10638 VDD.n4606 VDD.n986 4.58155
R10639 VDD.n4660 VDD.n954 4.58155
R10640 VDD.n4660 VDD.n955 4.58155
R10641 VDD.n4710 VDD.n918 4.58155
R10642 VDD.n5405 VDD.n309 4.55643
R10643 VDD.n5355 VDD.n334 4.55643
R10644 VDD.n376 VDD.n375 4.55643
R10645 VDD.n482 VDD.n440 4.55643
R10646 VDD.n540 VDD.n539 4.55643
R10647 VDD.n589 VDD.n588 4.55643
R10648 VDD.n5227 VDD.n5226 4.55643
R10649 VDD.n5178 VDD.n666 4.55643
R10650 VDD.n3630 VDD.n3624 4.53566
R10651 VDD.n3979 VDD.n2631 4.53566
R10652 VDD.n2545 VDD.n2539 4.5337
R10653 VDD.n3972 VDD.n3618 4.53087
R10654 VDD.n3964 VDD.n3963 4.52784
R10655 VDD.n5476 VDD.n263 4.52055
R10656 VDD.n3600 VDD.n3599 4.51815
R10657 VDD.n3594 VDD.n2647 4.51815
R10658 VDD.n3565 VDD.n3564 4.51815
R10659 VDD.n3539 VDD.n3538 4.51815
R10660 VDD.n3267 VDD.n3266 4.51815
R10661 VDD.n3241 VDD.n3240 4.51815
R10662 VDD.n3156 VDD.n3155 4.51815
R10663 VDD.n3150 VDD.n3120 4.51815
R10664 VDD.n3799 VDD.n3763 4.51815
R10665 VDD.n3928 VDD.n3658 4.51815
R10666 VDD.n3682 VDD.n3676 4.51815
R10667 VDD.n3936 VDD.n3641 4.51815
R10668 VDD.n2860 VDD.n2859 4.51815
R10669 VDD.n2887 VDD.n2886 4.51815
R10670 VDD.n2916 VDD.n2913 4.51815
R10671 VDD.n94 VDD.n93 4.51815
R10672 VDD.n78 VDD.n77 4.51815
R10673 VDD.n114 VDD.n28 4.51815
R10674 VDD.n5552 VDD.n5551 4.51815
R10675 VDD.n5563 VDD.n5562 4.51815
R10676 VDD.n175 VDD.n170 4.51815
R10677 VDD.n224 VDD.n223 4.51815
R10678 VDD.n1274 VDD.n1089 4.51815
R10679 VDD.n1270 VDD.n1089 4.51815
R10680 VDD.n2528 VDD.n2527 4.51815
R10681 VDD.n3604 VDD.n3602 4.51417
R10682 VDD.n3567 VDD.n3477 4.51417
R10683 VDD.n3456 VDD.n2697 4.51417
R10684 VDD.n3450 VDD.n2706 4.51417
R10685 VDD.n2728 VDD.n2717 4.51417
R10686 VDD.n3410 VDD.n3402 4.51417
R10687 VDD.n3396 VDD.n2742 4.51417
R10688 VDD.n3269 VDD.n3179 4.51417
R10689 VDD.n3158 VDD.n3102 4.51417
R10690 VDD.n3716 VDD.n3659 4.5005
R10691 VDD.n3908 VDD.n3907 4.5005
R10692 VDD.n3813 VDD.n3812 4.5005
R10693 VDD.n3942 VDD.n3634 4.5005
R10694 VDD.n3935 VDD.n3934 4.5005
R10695 VDD.n3698 VDD.n3689 4.5005
R10696 VDD.n3689 VDD.n3686 4.5005
R10697 VDD.n3698 VDD.n3688 4.5005
R10698 VDD.n3698 VDD.n3697 4.5005
R10699 VDD.n3697 VDD.n3686 4.5005
R10700 VDD.n3686 VDD.n3685 4.5005
R10701 VDD.n3929 VDD.n3656 4.5005
R10702 VDD.n3930 VDD.n3654 4.5005
R10703 VDD.n3664 VDD.n3654 4.5005
R10704 VDD.n3696 VDD.n3690 4.5005
R10705 VDD.n3697 VDD.n3696 4.5005
R10706 VDD.n3933 VDD.n3645 4.5005
R10707 VDD.n3931 VDD.n3646 4.5005
R10708 VDD.n3933 VDD.n3646 4.5005
R10709 VDD.n3933 VDD.n3932 4.5005
R10710 VDD.n3932 VDD.n3648 4.5005
R10711 VDD.n3932 VDD.n3931 4.5005
R10712 VDD.n3931 VDD.n3651 4.5005
R10713 VDD.n3934 VDD.n3633 4.5005
R10714 VDD.n3779 VDD.n3633 4.5005
R10715 VDD.n3942 VDD.n3633 4.5005
R10716 VDD.n3942 VDD.n3941 4.5005
R10717 VDD.n3941 VDD.n3637 4.5005
R10718 VDD.n3804 VDD.n3651 4.5005
R10719 VDD.n3808 VDD.n3645 4.5005
R10720 VDD.n3656 VDD.n3654 4.5005
R10721 VDD.n3656 VDD.n3652 4.5005
R10722 VDD.n3917 VDD.n3652 4.5005
R10723 VDD.n3930 VDD.n3652 4.5005
R10724 VDD.n3930 VDD.n3929 4.5005
R10725 VDD.n3924 VDD.n3923 4.5005
R10726 VDD.n3923 VDD.n3656 4.5005
R10727 VDD.n3689 VDD.n3677 4.5005
R10728 VDD.n3785 VDD.n3634 4.5005
R10729 VDD.n3934 VDD.n3634 4.5005
R10730 VDD.n3631 VDD.n3630 4.5005
R10731 VDD.n3631 VDD.n3623 4.5005
R10732 VDD.n3957 VDD.n3623 4.5005
R10733 VDD.n3957 VDD.n3956 4.5005
R10734 VDD.n3956 VDD.n3631 4.5005
R10735 VDD.n2815 VDD.n2804 4.5005
R10736 VDD.n2996 VDD.n2995 4.5005
R10737 VDD.n3003 VDD.n2894 4.5005
R10738 VDD.n3005 VDD.n2894 4.5005
R10739 VDD.n3028 VDD.n2869 4.5005
R10740 VDD.n2873 VDD.n2869 4.5005
R10741 VDD.n3005 VDD.n2892 4.5005
R10742 VDD.n2920 VDD.n2892 4.5005
R10743 VDD.n2907 VDD.n2899 4.5005
R10744 VDD.n2906 VDD.n2905 4.5005
R10745 VDD.n2907 VDD.n2906 4.5005
R10746 VDD.n2905 VDD.n2899 4.5005
R10747 VDD.n3028 VDD.n2871 4.5005
R10748 VDD.n3028 VDD.n2868 4.5005
R10749 VDD.n3028 VDD.n3027 4.5005
R10750 VDD.n2878 VDD.n2868 4.5005
R10751 VDD.n2873 VDD.n2868 4.5005
R10752 VDD.n3027 VDD.n2873 4.5005
R10753 VDD.n3027 VDD.n3026 4.5005
R10754 VDD.n2864 VDD.n2796 4.5005
R10755 VDD.n2800 VDD.n2796 4.5005
R10756 VDD.n2864 VDD.n2797 4.5005
R10757 VDD.n2807 VDD.n2795 4.5005
R10758 VDD.n2864 VDD.n2795 4.5005
R10759 VDD.n2800 VDD.n2795 4.5005
R10760 VDD.n2855 VDD.n2797 4.5005
R10761 VDD.n2800 VDD.n2797 4.5005
R10762 VDD.n2863 VDD.n2799 4.5005
R10763 VDD.n2864 VDD.n2863 4.5005
R10764 VDD.n2889 VDD.n2871 4.5005
R10765 VDD.n3003 VDD.n2892 4.5005
R10766 VDD.n3004 VDD.n3003 4.5005
R10767 VDD.n3004 VDD.n2896 4.5005
R10768 VDD.n3005 VDD.n3004 4.5005
R10769 VDD.n3002 VDD.n2910 4.5005
R10770 VDD.n3003 VDD.n3002 4.5005
R10771 VDD.n101 VDD.n100 4.5005
R10772 VDD.n135 VDD.n111 4.5005
R10773 VDD.n4295 VDD.n2358 4.5005
R10774 VDD.n5559 VDD.n5543 4.5005
R10775 VDD.n200 VDD.n199 4.5005
R10776 VDD.n5510 VDD.n168 4.5005
R10777 VDD.n5510 VDD.n166 4.5005
R10778 VDD.n5588 VDD.n5533 4.5005
R10779 VDD.n5588 VDD.n5526 4.5005
R10780 VDD.n5597 VDD.n161 4.5005
R10781 VDD.n5534 VDD.n161 4.5005
R10782 VDD.n5597 VDD.n163 4.5005
R10783 VDD.n5597 VDD.n160 4.5005
R10784 VDD.n5596 VDD.n5595 4.5005
R10785 VDD.n5526 VDD.n161 4.5005
R10786 VDD.n139 VDD.n138 4.5005
R10787 VDD.n138 VDD.n106 4.5005
R10788 VDD.n138 VDD.n24 4.5005
R10789 VDD.n140 VDD.n25 4.5005
R10790 VDD.n81 VDD.n37 4.5005
R10791 VDD.n81 VDD.n79 4.5005
R10792 VDD.n104 VDD.n35 4.5005
R10793 VDD.n37 VDD.n33 4.5005
R10794 VDD.n37 VDD.n32 4.5005
R10795 VDD.n49 VDD.n31 4.5005
R10796 VDD.n105 VDD.n32 4.5005
R10797 VDD.n140 VDD.n26 4.5005
R10798 VDD.n138 VDD.n26 4.5005
R10799 VDD.n120 VDD.n26 4.5005
R10800 VDD.n5596 VDD.n5526 4.5005
R10801 VDD.n5526 VDD.n160 4.5005
R10802 VDD.n5526 VDD.n163 4.5005
R10803 VDD.n5549 VDD.n163 4.5005
R10804 VDD.n5510 VDD.n5509 4.5005
R10805 VDD.n5508 VDD.n237 4.5005
R10806 VDD.n5508 VDD.n165 4.5005
R10807 VDD.n193 VDD.n165 4.5005
R10808 VDD.n5510 VDD.n165 4.5005
R10809 VDD.n237 VDD.n236 4.5005
R10810 VDD.n5509 VDD.n5508 4.5005
R10811 VDD.n48 VDD.n33 4.5005
R10812 VDD.n105 VDD.n33 4.5005
R10813 VDD.n105 VDD.n31 4.5005
R10814 VDD.n105 VDD.n104 4.5005
R10815 VDD.n37 VDD.n31 4.5005
R10816 VDD.n122 VDD.n25 4.5005
R10817 VDD.n130 VDD.n24 4.5005
R10818 VDD.n140 VDD.n24 4.5005
R10819 VDD.n124 VDD.n106 4.5005
R10820 VDD.n140 VDD.n139 4.5005
R10821 VDD.n5597 VDD.n5596 4.5005
R10822 VDD.n225 VDD.n166 4.5005
R10823 VDD.n226 VDD.n168 4.5005
R10824 VDD.n5508 VDD.n168 4.5005
R10825 VDD.n5507 VDD.n238 4.5005
R10826 VDD.n5490 VDD.n253 4.5005
R10827 VDD.n5505 VDD.n242 4.5005
R10828 VDD.n254 VDD.n252 4.5005
R10829 VDD.n5483 VDD.n5482 4.5005
R10830 VDD.n5481 VDD.n257 4.5005
R10831 VDD.n5465 VDD.n5464 4.5005
R10832 VDD.n5467 VDD.n5466 4.5005
R10833 VDD.n5469 VDD.n258 4.5005
R10834 VDD.n5463 VDD.n5462 4.5005
R10835 VDD.n242 VDD.n238 4.5005
R10836 VDD.n2453 VDD.n2452 4.5005
R10837 VDD.n5493 VDD.n5492 4.5005
R10838 VDD.n2589 VDD.n2588 4.5005
R10839 VDD.n2523 VDD.n2512 4.5005
R10840 VDD.n2571 VDD.n2570 4.5005
R10841 VDD.n2549 VDD.n2548 4.5005
R10842 VDD.n2553 VDD.n2552 4.5005
R10843 VDD.n2565 VDD.n2564 4.5005
R10844 VDD.n2551 VDD.n2538 4.5005
R10845 VDD.n2554 VDD.n2537 4.5005
R10846 VDD.n2561 VDD.n2560 4.5005
R10847 VDD.n2562 VDD.n2534 4.5005
R10848 VDD.n2541 VDD.n2539 4.5005
R10849 VDD.n2572 VDD.n2522 4.5005
R10850 VDD.n2575 VDD.n2574 4.5005
R10851 VDD.n2530 VDD.n2527 4.5005
R10852 VDD.n2525 VDD.n2524 4.5005
R10853 VDD.n2580 VDD.n2579 4.5005
R10854 VDD.n2584 VDD.n2510 4.5005
R10855 VDD.n2587 VDD.n2508 4.5005
R10856 VDD.n3174 VDD.n3173 4.5005
R10857 VDD.n3271 VDD.n3068 4.5005
R10858 VDD.n3272 VDD.n3271 4.5005
R10859 VDD.n3302 VDD.n3301 4.5005
R10860 VDD.n3069 VDD.n3061 4.5005
R10861 VDD.n3069 VDD.n3064 4.5005
R10862 VDD.n3293 VDD.n3069 4.5005
R10863 VDD.n3300 VDD.n3069 4.5005
R10864 VDD.n3299 VDD.n3061 4.5005
R10865 VDD.n3299 VDD.n3064 4.5005
R10866 VDD.n3299 VDD.n3298 4.5005
R10867 VDD.n3373 VDD.n3327 4.5005
R10868 VDD.n3399 VDD.n3398 4.5005
R10869 VDD.n3398 VDD.n2740 4.5005
R10870 VDD.n3177 VDD.n3175 4.5005
R10871 VDD.n3279 VDD.n3175 4.5005
R10872 VDD.n3279 VDD.n3068 4.5005
R10873 VDD.n3174 VDD.n3090 4.5005
R10874 VDD.n3099 VDD.n3090 4.5005
R10875 VDD.n3117 VDD.n3090 4.5005
R10876 VDD.n3160 VDD.n3117 4.5005
R10877 VDD.n3116 VDD.n2486 4.5005
R10878 VDD.n3114 VDD.n2486 4.5005
R10879 VDD.n3116 VDD.n3115 4.5005
R10880 VDD.n3115 VDD.n3114 4.5005
R10881 VDD.n3103 VDD.n3102 4.5005
R10882 VDD.n3161 VDD.n3160 4.5005
R10883 VDD.n3279 VDD.n3088 4.5005
R10884 VDD.n3301 VDD.n3063 4.5005
R10885 VDD.n3067 VDD.n3061 4.5005
R10886 VDD.n3284 VDD.n3067 4.5005
R10887 VDD.n3300 VDD.n3067 4.5005
R10888 VDD.n3348 VDD.n2766 4.5005
R10889 VDD.n3355 VDD.n2766 4.5005
R10890 VDD.n3373 VDD.n2766 4.5005
R10891 VDD.n3373 VDD.n3372 4.5005
R10892 VDD.n3372 VDD.n3371 4.5005
R10893 VDD.n3327 VDD.n2765 4.5005
R10894 VDD.n3365 VDD.n3327 4.5005
R10895 VDD.n3348 VDD.n3327 4.5005
R10896 VDD.n3423 VDD.n2731 4.5005
R10897 VDD.n3420 VDD.n3401 4.5005
R10898 VDD.n3399 VDD.n2736 4.5005
R10899 VDD.n3387 VDD.n2736 4.5005
R10900 VDD.n3379 VDD.n2736 4.5005
R10901 VDD.n3432 VDD.n2710 4.5005
R10902 VDD.n2724 VDD.n2710 4.5005
R10903 VDD.n3424 VDD.n2710 4.5005
R10904 VDD.n3425 VDD.n2715 4.5005
R10905 VDD.n3423 VDD.n3422 4.5005
R10906 VDD.n3422 VDD.n2733 4.5005
R10907 VDD.n3422 VDD.n3421 4.5005
R10908 VDD.n3453 VDD.n3452 4.5005
R10909 VDD.n3452 VDD.n2704 4.5005
R10910 VDD.n3432 VDD.n3431 4.5005
R10911 VDD.n3472 VDD.n3471 4.5005
R10912 VDD.n3569 VDD.n2688 4.5005
R10913 VDD.n3570 VDD.n3569 4.5005
R10914 VDD.n3615 VDD.n2634 4.5005
R10915 VDD.n2653 VDD.n2634 4.5005
R10916 VDD.n2687 VDD.n2634 4.5005
R10917 VDD.n2686 VDD.n2640 4.5005
R10918 VDD.n3617 VDD.n2630 4.5005
R10919 VDD.n3978 VDD.n3617 4.5005
R10920 VDD.n3977 VDD.n2630 4.5005
R10921 VDD.n2595 VDD.n2592 4.5005
R10922 VDD.n2628 VDD.n2592 4.5005
R10923 VDD.n2627 VDD.n2595 4.5005
R10924 VDD.n2628 VDD.n2591 4.5005
R10925 VDD.n2628 VDD.n2627 4.5005
R10926 VDD.n3475 VDD.n3473 4.5005
R10927 VDD.n3577 VDD.n3473 4.5005
R10928 VDD.n3577 VDD.n2688 4.5005
R10929 VDD.n3472 VDD.n2689 4.5005
R10930 VDD.n3465 VDD.n2689 4.5005
R10931 VDD.n3454 VDD.n2689 4.5005
R10932 VDD.n3458 VDD.n3454 4.5005
R10933 VDD.n3453 VDD.n2700 4.5005
R10934 VDD.n3441 VDD.n2700 4.5005
R10935 VDD.n3433 VDD.n2700 4.5005
R10936 VDD.n2698 VDD.n2697 4.5005
R10937 VDD.n3459 VDD.n3458 4.5005
R10938 VDD.n3577 VDD.n2682 4.5005
R10939 VDD.n3615 VDD.n3614 4.5005
R10940 VDD.n3979 VDD.n3978 4.5005
R10941 VDD.n3979 VDD.n2630 4.5005
R10942 VDD.n2595 VDD.n2591 4.5005
R10943 VDD.n3978 VDD.n3977 4.5005
R10944 VDD.n3604 VDD.n2642 4.5005
R10945 VDD.n2687 VDD.n2686 4.5005
R10946 VDD.n3478 VDD.n3477 4.5005
R10947 VDD.n3434 VDD.n3433 4.5005
R10948 VDD.n3451 VDD.n3450 4.5005
R10949 VDD.n2729 VDD.n2728 4.5005
R10950 VDD.n3425 VDD.n3424 4.5005
R10951 VDD.n3410 VDD.n3400 4.5005
R10952 VDD.n3421 VDD.n3420 4.5005
R10953 VDD.n3380 VDD.n3379 4.5005
R10954 VDD.n3397 VDD.n3396 4.5005
R10955 VDD.n3301 VDD.n3062 4.5005
R10956 VDD.n3300 VDD.n3299 4.5005
R10957 VDD.n3180 VDD.n3179 4.5005
R10958 VDD.n1870 VDD.n1054 4.4978
R10959 VDD.n2354 VDD.n2353 4.48249
R10960 VDD.n4749 VDD.n4748 4.47034
R10961 VDD.n4752 VDD.n902 4.47034
R10962 VDD.n4804 VDD.n4803 4.47034
R10963 VDD.n4812 VDD.n4811 4.47034
R10964 VDD.n4863 VDD.n4862 4.47034
R10965 VDD.n4866 VDD.n840 4.47034
R10966 VDD.n4918 VDD.n4917 4.47034
R10967 VDD.n4926 VDD.n4925 4.47034
R10968 VDD.n4977 VDD.n4976 4.47034
R10969 VDD.n4980 VDD.n778 4.47034
R10970 VDD.n5032 VDD.n5031 4.47034
R10971 VDD.n5040 VDD.n5039 4.47034
R10972 VDD.n5091 VDD.n5090 4.47034
R10973 VDD.n5094 VDD.n716 4.47034
R10974 VDD.n5146 VDD.n5145 4.47034
R10975 VDD.n5154 VDD.n681 4.47034
R10976 VDD.n5453 VDD.n5452 4.4118
R10977 VDD.n5394 VDD.n316 4.4118
R10978 VDD.n5344 VDD.n5343 4.4118
R10979 VDD.n387 VDD.n381 4.4118
R10980 VDD.n495 VDD.n494 4.4118
R10981 VDD.n551 VDD.n412 4.4118
R10982 VDD.n600 VDD.n594 4.4118
R10983 VDD.n5215 VDD.n637 4.4118
R10984 VDD.n5167 VDD.n5166 4.4118
R10985 VDD.n1032 VDD.n1031 4.36497
R10986 VDD.n132 VDD.n119 4.35817
R10987 VDD.n1881 VDD.n1880 4.3536
R10988 VDD.n251 VDD.n250 4.31361
R10989 VDD.n5475 VDD.n5474 4.31361
R10990 VDD.n5472 VDD.n5471 4.31361
R10991 VDD.n4007 VDD.n4006 4.31361
R10992 VDD.n3110 VDD.n2481 4.31361
R10993 VDD.n4009 VDD.n2476 4.31361
R10994 VDD.n3950 VDD.n3620 4.31361
R10995 VDD.n3980 VDD.n2503 4.31361
R10996 VDD.n2504 VDD.n2502 4.31361
R10997 VDD.n2452 VDD.n2442 4.31327
R10998 VDD.n1245 VDD.n1106 4.31208
R10999 VDD.n1234 VDD.n1113 4.31208
R11000 VDD.n1193 VDD.n1141 4.31208
R11001 VDD.n1182 VDD.n1148 4.31208
R11002 VDD.n4600 VDD.n4599 4.31208
R11003 VDD.n4611 VDD.n982 4.31208
R11004 VDD.n4657 VDD.n4656 4.31208
R11005 VDD.n4666 VDD.n950 4.31208
R11006 VDD.n4712 VDD.n4711 4.31208
R11007 VDD.n1468 VDD.n1379 4.30941
R11008 VDD.n1858 VDD.n1857 4.26717
R11009 VDD.n1839 VDD.n1072 4.26717
R11010 VDD.n5409 VDD.n5406 4.26717
R11011 VDD.n5359 VDD.n5358 4.26717
R11012 VDD.n5310 VDD.n371 4.26717
R11013 VDD.n479 VDD.n478 4.26717
R11014 VDD.n533 VDD.n418 4.26717
R11015 VDD.n5277 VDD.n584 4.26717
R11016 VDD.n628 VDD.n627 4.26717
R11017 VDD.n5179 VDD.n663 4.26717
R11018 VDD.n4722 VDD.n918 4.24471
R11019 VDD.n3583 VDD.n3582 4.23768
R11020 VDD.n3139 VDD.n3138 4.23768
R11021 VDD.n3767 VDD.n3764 4.23768
R11022 VDD.n210 VDD.n208 4.23768
R11023 VDD.n2926 VDD.n2925 4.23684
R11024 VDD.n64 VDD.n62 4.23684
R11025 VDD.n5575 VDD.n5569 4.23684
R11026 VDD.n1869 VDD.n1055 4.22104
R11027 VDD.n909 VDD.n904 4.19944
R11028 VDD.n4759 VDD.n897 4.19944
R11029 VDD.n4802 VDD.n874 4.19944
R11030 VDD.n4817 VDD.n867 4.19944
R11031 VDD.n847 VDD.n842 4.19944
R11032 VDD.n4873 VDD.n835 4.19944
R11033 VDD.n4916 VDD.n812 4.19944
R11034 VDD.n4931 VDD.n805 4.19944
R11035 VDD.n785 VDD.n780 4.19944
R11036 VDD.n4987 VDD.n773 4.19944
R11037 VDD.n5030 VDD.n750 4.19944
R11038 VDD.n5045 VDD.n743 4.19944
R11039 VDD.n723 VDD.n718 4.19944
R11040 VDD.n5101 VDD.n711 4.19944
R11041 VDD.n5144 VDD.n688 4.19944
R11042 VDD.n5158 VDD.n5157 4.19944
R11043 VDD.n2604 VDD.n2600 4.18565
R11044 VDD.n3951 VDD.n2499 4.18565
R11045 VDD.n8361 VDD.n8360 4.17441
R11046 VDD.n7506 VDD.n7505 4.17441
R11047 VDD.n6652 VDD.n6651 4.17441
R11048 VDD.n5797 VDD.n5796 4.17441
R11049 VDD.n3612 VDD.n3611 4.14168
R11050 VDD.n3525 VDD.n3524 4.14168
R11051 VDD.n3227 VDD.n3226 4.14168
R11052 VDD.n3171 VDD.n3170 4.14168
R11053 VDD.n3797 VDD.n3794 4.14168
R11054 VDD.n3805 VDD.n3804 4.14168
R11055 VDD.n3826 VDD.n3825 4.14168
R11056 VDD.n3912 VDD.n3911 4.14168
R11057 VDD.n3925 VDD.n3924 4.14168
R11058 VDD.n3729 VDD.n3728 4.14168
R11059 VDD.n3694 VDD.n3693 4.14168
R11060 VDD.n3685 VDD.n3672 4.14168
R11061 VDD.n3895 VDD.n3894 4.14168
R11062 VDD.n3783 VDD.n3774 4.14168
R11063 VDD.n3780 VDD.n3637 4.14168
R11064 VDD.n2850 VDD.n2849 4.14168
R11065 VDD.n2856 VDD.n2799 4.14168
R11066 VDD.n2839 VDD.n2838 4.14168
R11067 VDD.n2883 VDD.n2877 4.14168
R11068 VDD.n3026 VDD.n2875 4.14168
R11069 VDD.n2936 VDD.n2933 4.14168
R11070 VDD.n2929 VDD.n2910 4.14168
R11071 VDD.n2984 VDD.n2983 4.14168
R11072 VDD.n2983 VDD.n2958 4.14168
R11073 VDD.n83 VDD.n52 4.14168
R11074 VDD.n125 VDD.n117 4.14168
R11075 VDD.n5590 VDD.n5532 4.14168
R11076 VDD.n231 VDD.n180 4.14168
R11077 VDD.n1840 VDD.n1070 4.14168
R11078 VDD.n1833 VDD.n1076 4.14168
R11079 VDD.n1422 VDD.n1421 4.13172
R11080 VDD.n1477 VDD.n1476 4.13172
R11081 VDD.n1388 VDD.n1028 4.13172
R11082 VDD.n4524 VDD.n4523 4.13172
R11083 VDD.n1961 VDD.n1960 4.13172
R11084 VDD.n4517 VDD.n1966 4.13172
R11085 VDD.n2065 VDD.n2064 4.13172
R11086 VDD.n4456 VDD.n2066 4.13172
R11087 VDD.n2079 VDD.n2078 4.13172
R11088 VDD.n4389 VDD.n4388 4.13172
R11089 VDD.n2182 VDD.n2181 4.13172
R11090 VDD.n4382 VDD.n2187 4.13172
R11091 VDD.n296 VDD.n278 4.12253
R11092 VDD.n5393 VDD.n317 4.12253
R11093 VDD.n348 VDD.n344 4.12253
R11094 VDD.n5293 VDD.n388 4.12253
R11095 VDD.n500 VDD.n434 4.12253
R11096 VDD.n555 VDD.n554 4.12253
R11097 VDD.n5260 VDD.n601 4.12253
R11098 VDD.n5212 VDD.n5211 4.12253
R11099 VDD.n2174 VDD.t94 4.10046
R11100 VDD.n4195 VDD.n265 4.08166
R11101 VDD.n1420 VDD.n1417 4.06399
R11102 VDD.n1972 VDD.n1971 4.06399
R11103 VDD.n4461 VDD.n4460 4.06399
R11104 VDD.n2193 VDD.n2192 4.06399
R11105 VDD.n5446 VDD.n277 4.05022
R11106 VDD.n1246 VDD.n1104 4.04261
R11107 VDD.n1233 VDD.n1114 4.04261
R11108 VDD.n1194 VDD.n1139 4.04261
R11109 VDD.n1181 VDD.n1149 4.04261
R11110 VDD.n4598 VDD.n990 4.04261
R11111 VDD.n4610 VDD.n983 4.04261
R11112 VDD.n962 VDD.n957 4.04261
R11113 VDD.n4668 VDD.n4667 4.04261
R11114 VDD.n4709 VDD.n927 4.04261
R11115 VDD.n2356 VDD.n2342 4.03708
R11116 VDD.n2356 VDD.n2343 4.03708
R11117 VDD.n5410 VDD.n306 3.9779
R11118 VDD.n333 VDD.n332 3.9779
R11119 VDD.n5311 VDD.n368 3.9779
R11120 VDD.n474 VDD.n442 3.9779
R11121 VDD.n532 VDD.n420 3.9779
R11122 VDD.n5278 VDD.n400 3.9779
R11123 VDD.n5233 VDD.n623 3.9779
R11124 VDD.n5183 VDD.n5182 3.9779
R11125 VDD.t94 VDD.n2173 3.9682
R11126 VDD.n1866 VDD.n1865 3.94428
R11127 VDD.n1379 VDD.n1378 3.92921
R11128 VDD.n1488 VDD.n1373 3.92921
R11129 VDD.n1489 VDD.n1371 3.92921
R11130 VDD.n1323 VDD.n1320 3.92921
R11131 VDD.n1569 VDD.n1317 3.92921
R11132 VDD.n1315 VDD.n1311 3.92921
R11133 VDD.n1642 VDD.n1635 3.92921
R11134 VDD.n1783 VDD.n1644 3.92921
R11135 VDD.n1649 VDD.n1647 3.92921
R11136 VDD.n4742 VDD.n4741 3.92854
R11137 VDD.n4761 VDD.n4760 3.92854
R11138 VDD.n4799 VDD.n4798 3.92854
R11139 VDD.n4816 VDD.n868 3.92854
R11140 VDD.n4856 VDD.n4855 3.92854
R11141 VDD.n4875 VDD.n4874 3.92854
R11142 VDD.n4913 VDD.n4912 3.92854
R11143 VDD.n4930 VDD.n806 3.92854
R11144 VDD.n4970 VDD.n4969 3.92854
R11145 VDD.n4989 VDD.n4988 3.92854
R11146 VDD.n5027 VDD.n5026 3.92854
R11147 VDD.n5044 VDD.n744 3.92854
R11148 VDD.n5084 VDD.n5083 3.92854
R11149 VDD.n5103 VDD.n5102 3.92854
R11150 VDD.n5141 VDD.n5140 3.92854
R11151 VDD.n1844 VDD.n1843 3.8907
R11152 VDD.n1832 VDD.n1077 3.8907
R11153 VDD.n1897 VDD.n1896 3.86082
R11154 VDD.n4514 VDD.n4513 3.86082
R11155 VDD.n4445 VDD.n2080 3.86082
R11156 VDD.n4379 VDD.n4378 3.86082
R11157 VDD.n5437 VDD.n297 3.83327
R11158 VDD.n5390 VDD.n5389 3.83327
R11159 VDD.n5337 VDD.n349 3.83327
R11160 VDD.n5292 VDD.n389 3.83327
R11161 VDD.n501 VDD.n432 3.83327
R11162 VDD.n559 VDD.n410 3.83327
R11163 VDD.n5259 VDD.n602 3.83327
R11164 VDD.n643 VDD.n639 3.83327
R11165 VDD.n1430 VDD.n1427 3.79309
R11166 VDD.n1968 VDD.n1947 3.79309
R11167 VDD.n2087 VDD.n2086 3.79309
R11168 VDD.n2189 VDD.n2167 3.79309
R11169 VDD.n2354 VDD.n2346 3.79052
R11170 VDD.t41 VDD.n4275 3.78536
R11171 VDD.n8821 VDD.n8711 3.78485
R11172 VDD.n8718 VDD.n8717 3.78485
R11173 VDD.n9008 VDD.n8264 3.78485
R11174 VDD.n7966 VDD.n7856 3.78485
R11175 VDD.n7863 VDD.n7862 3.78485
R11176 VDD.n8153 VDD.n7409 3.78485
R11177 VDD.n7112 VDD.n7002 3.78485
R11178 VDD.n7009 VDD.n7008 3.78485
R11179 VDD.n7299 VDD.n6555 3.78485
R11180 VDD.n6257 VDD.n6147 3.78485
R11181 VDD.n6154 VDD.n6153 3.78485
R11182 VDD.n6444 VDD.n5700 3.78485
R11183 VDD.n1250 VDD.n1249 3.77313
R11184 VDD.n1230 VDD.n1229 3.77313
R11185 VDD.n1198 VDD.n1197 3.77313
R11186 VDD.n1178 VDD.n1177 3.77313
R11187 VDD.n4595 VDD.n4594 3.77313
R11188 VDD.n4617 VDD.n978 3.77313
R11189 VDD.n4650 VDD.n4649 3.77313
R11190 VDD.n4673 VDD.n947 3.77313
R11191 VDD.n4706 VDD.n4705 3.77313
R11192 VDD.n2653 VDD.n2652 3.76521
R11193 VDD.n2655 VDD.n2646 3.76521
R11194 VDD.n3571 VDD.n3570 3.76521
R11195 VDD.n3534 VDD.n3533 3.76521
R11196 VDD.n3460 VDD.n3459 3.76521
R11197 VDD.n3441 VDD.n3440 3.76521
R11198 VDD.n2725 VDD.n2724 3.76521
R11199 VDD.n3407 VDD.n3401 3.76521
R11200 VDD.n3387 VDD.n3386 3.76521
R11201 VDD.n3366 VDD.n3365 3.76521
R11202 VDD.n3294 VDD.n3293 3.76521
R11203 VDD.n3273 VDD.n3272 3.76521
R11204 VDD.n3236 VDD.n3235 3.76521
R11205 VDD.n3162 VDD.n3161 3.76521
R11206 VDD.n3124 VDD.n3119 3.76521
R11207 VDD.n87 VDD.n86 3.76521
R11208 VDD.n2353 VDD.n2347 3.76521
R11209 VDD.n5594 VDD.n5529 3.76521
R11210 VDD.n235 VDD.n177 3.76521
R11211 VDD.n1469 VDD.n1468 3.73911
R11212 VDD.n1493 VDD.n1368 3.73911
R11213 VDD.n1565 VDD.n1322 3.73911
R11214 VDD.n1581 VDD.n1580 3.73911
R11215 VDD.n1793 VDD.n1634 3.73911
R11216 VDD.n1779 VDD.n1778 3.73911
R11217 VDD.n1892 VDD.n1032 3.70369
R11218 VDD.n5414 VDD.n5413 3.68864
R11219 VDD.n5365 VDD.n327 3.68864
R11220 VDD.n5315 VDD.n5314 3.68864
R11221 VDD.n473 VDD.n444 3.68864
R11222 VDD.n529 VDD.n528 3.68864
R11223 VDD.n5282 VDD.n5281 3.68864
R11224 VDD.n5234 VDD.n620 3.68864
R11225 VDD.n662 VDD.n661 3.68864
R11226 VDD.n5648 VDD.n5647 3.67828
R11227 VDD.n6510 VDD.n6509 3.67828
R11228 VDD.n7357 VDD.n7356 3.67828
R11229 VDD.n8219 VDD.n8218 3.67828
R11230 VDD.n4736 VDD.n908 3.65764
R11231 VDD.n4766 VDD.n894 3.65764
R11232 VDD.n881 VDD.n876 3.65764
R11233 VDD.n4823 VDD.n863 3.65764
R11234 VDD.n4850 VDD.n846 3.65764
R11235 VDD.n4880 VDD.n832 3.65764
R11236 VDD.n819 VDD.n814 3.65764
R11237 VDD.n4937 VDD.n801 3.65764
R11238 VDD.n4964 VDD.n784 3.65764
R11239 VDD.n4994 VDD.n770 3.65764
R11240 VDD.n757 VDD.n752 3.65764
R11241 VDD.n5051 VDD.n739 3.65764
R11242 VDD.n5078 VDD.n722 3.65764
R11243 VDD.n5108 VDD.n708 3.65764
R11244 VDD.n695 VDD.n690 3.65764
R11245 VDD.n8644 VDD.n8635 3.64278
R11246 VDD.n7789 VDD.n7780 3.64278
R11247 VDD.n6935 VDD.n6926 3.64278
R11248 VDD.n6080 VDD.n6071 3.64278
R11249 VDD.n1848 VDD.n1066 3.63972
R11250 VDD.n1829 VDD.n1828 3.63972
R11251 VDD.n4574 VDD.n1005 3.58992
R11252 VDD.n1984 VDD.n1983 3.58992
R11253 VDD.n4442 VDD.n4441 3.58992
R11254 VDD.n2205 VDD.n2204 3.58992
R11255 VDD.n5436 VDD.n298 3.544
R11256 VDD.n5386 VDD.n5385 3.544
R11257 VDD.n5336 VDD.n350 3.544
R11258 VDD.n5289 VDD.n5288 3.544
R11259 VDD.n505 VDD.n504 3.544
R11260 VDD.n560 VDD.n408 3.544
R11261 VDD.n5256 VDD.n5255 3.544
R11262 VDD.n5205 VDD.n644 3.544
R11263 VDD.n1434 VDD.n1415 3.52219
R11264 VDD.n1945 VDD.n1931 3.52219
R11265 VDD.n2085 VDD.n2052 3.52219
R11266 VDD.n2165 VDD.n2151 3.52219
R11267 VDD.n1254 VDD.n1100 3.50366
R11268 VDD.n1225 VDD.n1117 3.50366
R11269 VDD.n1202 VDD.n1135 3.50366
R11270 VDD.n1173 VDD.n1152 3.50366
R11271 VDD.n997 VDD.n992 3.50366
R11272 VDD.n4619 VDD.n4618 3.50366
R11273 VDD.n4644 VDD.n961 3.50366
R11274 VDD.n4672 VDD.n948 3.50366
R11275 VDD.n934 VDD.n929 3.50366
R11276 VDD.n1366 VDD.n1362 3.48565
R11277 VDD.n1329 VDD.n1328 3.48565
R11278 VDD.n1585 VDD.n1584 3.48565
R11279 VDD.n1797 VDD.n1796 3.48565
R11280 VDD.n1659 VDD.n1658 3.48565
R11281 VDD.n1703 VDD.n1702 3.48565
R11282 VDD.n6527 VDD.n6520 3.43528
R11283 VDD.n8236 VDD.n8229 3.43528
R11284 VDD.n2829 VDD.n2828 3.42768
R11285 VDD.n2971 VDD.n2970 3.42768
R11286 VDD.n3510 VDD.n3508 3.42765
R11287 VDD.n3212 VDD.n3210 3.42765
R11288 VDD.n3880 VDD.n3878 3.42765
R11289 VDD.n3499 VDD.n3498 3.42683
R11290 VDD.n3201 VDD.n3200 3.42683
R11291 VDD.n3749 VDD.n3748 3.42683
R11292 VDD.n263 VDD.n255 3.42673
R11293 VDD.n3965 VDD.n3964 3.42318
R11294 VDD.n3960 VDD.n3624 3.42286
R11295 VDD.n8276 VDD.n8271 3.42221
R11296 VDD.n7421 VDD.n7416 3.42221
R11297 VDD.n6567 VDD.n6562 3.42221
R11298 VDD.n5712 VDD.n5707 3.42221
R11299 VDD.n5489 VDD.n5488 3.41892
R11300 VDD.n3966 VDD.n2631 3.41503
R11301 VDD.n3622 VDD.n3621 3.4105
R11302 VDD.n3959 VDD.n3958 3.4105
R11303 VDD.n3959 VDD.n3943 3.4105
R11304 VDD.n3944 VDD.n3943 3.4105
R11305 VDD.n3958 VDD.n3944 3.4105
R11306 VDD.n3943 VDD.n3628 3.4105
R11307 VDD.n3958 VDD.n3628 3.4105
R11308 VDD.n3961 VDD.n3960 3.4105
R11309 VDD.n3962 VDD.n3628 3.4105
R11310 VDD.n3963 VDD.n3962 3.4105
R11311 VDD.n5488 VDD.n5487 3.4105
R11312 VDD.n260 VDD.n256 3.4105
R11313 VDD.n256 VDD.n2 3.4105
R11314 VDD.n5479 VDD.n5478 3.4105
R11315 VDD.n5468 VDD.n2 3.4105
R11316 VDD.n260 VDD.n259 3.4105
R11317 VDD.n259 VDD.n2 3.4105
R11318 VDD.n5479 VDD.n262 3.4105
R11319 VDD.n5480 VDD.n5479 3.4105
R11320 VDD.n5479 VDD.n259 3.4105
R11321 VDD.n264 VDD.n259 3.4105
R11322 VDD.n5479 VDD.n256 3.4105
R11323 VDD.n5484 VDD.n256 3.4105
R11324 VDD.n3975 VDD.n3971 3.4105
R11325 VDD.n3975 VDD.n3974 3.4105
R11326 VDD.n3975 VDD.n3968 3.4105
R11327 VDD.n3974 VDD.n3616 3.4105
R11328 VDD.n3967 VDD.n2632 3.4105
R11329 VDD.n3303 VDD.n3302 3.4105
R11330 VDD.n3350 VDD.n2765 3.4105
R11331 VDD.n3303 VDD.n3063 3.4105
R11332 VDD.n3303 VDD.n3062 3.4105
R11333 VDD.n2762 VDD.n2753 3.4105
R11334 VDD.n2762 VDD.n2755 3.4105
R11335 VDD.n2762 VDD.n2754 3.4105
R11336 VDD.n3375 VDD.n2762 3.4105
R11337 VDD.n2762 VDD.n2749 3.4105
R11338 VDD.n2762 VDD.n2758 3.4105
R11339 VDD.n2762 VDD.n2750 3.4105
R11340 VDD.n2762 VDD.n2757 3.4105
R11341 VDD.n2762 VDD.n2746 3.4105
R11342 VDD.n2764 VDD.n2753 3.4105
R11343 VDD.n2764 VDD.n2755 3.4105
R11344 VDD.n2764 VDD.n2754 3.4105
R11345 VDD.n3375 VDD.n2764 3.4105
R11346 VDD.n2764 VDD.n2749 3.4105
R11347 VDD.n2764 VDD.n2758 3.4105
R11348 VDD.n2764 VDD.n2750 3.4105
R11349 VDD.n2764 VDD.n2757 3.4105
R11350 VDD.n2764 VDD.n2746 3.4105
R11351 VDD.n3375 VDD.n2761 3.4105
R11352 VDD.n2761 VDD.n2749 3.4105
R11353 VDD.n2761 VDD.n2758 3.4105
R11354 VDD.n2761 VDD.n2750 3.4105
R11355 VDD.n2761 VDD.n2757 3.4105
R11356 VDD.n3331 VDD.n2761 3.4105
R11357 VDD.n2761 VDD.n2746 3.4105
R11358 VDD.n2761 VDD.n2754 3.4105
R11359 VDD.n2761 VDD.n2755 3.4105
R11360 VDD.n2761 VDD.n2753 3.4105
R11361 VDD.n3376 VDD.n2754 3.4105
R11362 VDD.n3376 VDD.n2755 3.4105
R11363 VDD.n3376 VDD.n2753 3.4105
R11364 VDD.n2753 VDD.n2747 3.4105
R11365 VDD.n2755 VDD.n2747 3.4105
R11366 VDD.n2754 VDD.n2747 3.4105
R11367 VDD.n3375 VDD.n2747 3.4105
R11368 VDD.n2749 VDD.n2747 3.4105
R11369 VDD.n2758 VDD.n2747 3.4105
R11370 VDD.n2750 VDD.n2747 3.4105
R11371 VDD.n2757 VDD.n2747 3.4105
R11372 VDD.n3377 VDD.n2747 3.4105
R11373 VDD.n2752 VDD.n2747 3.4105
R11374 VDD.n2760 VDD.n2746 3.4105
R11375 VDD.n3331 VDD.n2760 3.4105
R11376 VDD.n2760 VDD.n2757 3.4105
R11377 VDD.n2760 VDD.n2750 3.4105
R11378 VDD.n2760 VDD.n2758 3.4105
R11379 VDD.n2760 VDD.n2749 3.4105
R11380 VDD.n3375 VDD.n2760 3.4105
R11381 VDD.n2760 VDD.n2754 3.4105
R11382 VDD.n2760 VDD.n2755 3.4105
R11383 VDD.n2760 VDD.n2753 3.4105
R11384 VDD.n3376 VDD.n2752 3.4105
R11385 VDD.n3377 VDD.n3376 3.4105
R11386 VDD.n3376 VDD.n2757 3.4105
R11387 VDD.n3376 VDD.n2750 3.4105
R11388 VDD.n3376 VDD.n2758 3.4105
R11389 VDD.n3376 VDD.n2749 3.4105
R11390 VDD.n3376 VDD.n3375 3.4105
R11391 VDD.n3305 VDD.n3057 3.4105
R11392 VDD.n3057 VDD.n2770 3.4105
R11393 VDD.n3308 VDD.n3307 3.4105
R11394 VDD.n3308 VDD.n2770 3.4105
R11395 VDD.n3045 VDD.n2784 3.4105
R11396 VDD.n2784 VDD.n2773 3.4105
R11397 VDD.n2784 VDD.n2782 3.4105
R11398 VDD.n2784 VDD.n2774 3.4105
R11399 VDD.n2784 VDD.n2781 3.4105
R11400 VDD.n2784 VDD.n2775 3.4105
R11401 VDD.n2784 VDD.n2780 3.4105
R11402 VDD.n2784 VDD.n2779 3.4105
R11403 VDD.n2784 VDD.n2778 3.4105
R11404 VDD.n2786 VDD.n2782 3.4105
R11405 VDD.n2786 VDD.n2774 3.4105
R11406 VDD.n2786 VDD.n2781 3.4105
R11407 VDD.n2786 VDD.n2775 3.4105
R11408 VDD.n2786 VDD.n2780 3.4105
R11409 VDD.n2786 VDD.n2776 3.4105
R11410 VDD.n2786 VDD.n2779 3.4105
R11411 VDD.n3042 VDD.n2786 3.4105
R11412 VDD.n2865 VDD.n2793 3.4105
R11413 VDD.n2865 VDD.n2789 3.4105
R11414 VDD.n3042 VDD.n2789 3.4105
R11415 VDD.n2789 VDD.n2779 3.4105
R11416 VDD.n2789 VDD.n2780 3.4105
R11417 VDD.n2789 VDD.n2775 3.4105
R11418 VDD.n2789 VDD.n2781 3.4105
R11419 VDD.n2789 VDD.n2774 3.4105
R11420 VDD.n2789 VDD.n2782 3.4105
R11421 VDD.n2789 VDD.n2773 3.4105
R11422 VDD.n2789 VDD.n2783 3.4105
R11423 VDD.n2789 VDD.n2785 3.4105
R11424 VDD.n3046 VDD.n2778 3.4105
R11425 VDD.n3046 VDD.n2779 3.4105
R11426 VDD.n3046 VDD.n2776 3.4105
R11427 VDD.n3046 VDD.n2780 3.4105
R11428 VDD.n3046 VDD.n2775 3.4105
R11429 VDD.n3046 VDD.n2781 3.4105
R11430 VDD.n3046 VDD.n2774 3.4105
R11431 VDD.n3046 VDD.n2782 3.4105
R11432 VDD.n3046 VDD.n2773 3.4105
R11433 VDD.n3046 VDD.n3045 3.4105
R11434 VDD.n2793 VDD.n2783 3.4105
R11435 VDD.n2793 VDD.n2782 3.4105
R11436 VDD.n2793 VDD.n2774 3.4105
R11437 VDD.n2793 VDD.n2781 3.4105
R11438 VDD.n2793 VDD.n2775 3.4105
R11439 VDD.n2793 VDD.n2780 3.4105
R11440 VDD.n2793 VDD.n2776 3.4105
R11441 VDD.n2793 VDD.n2779 3.4105
R11442 VDD.n2793 VDD.n2785 3.4105
R11443 VDD.n3043 VDD.n2773 3.4105
R11444 VDD.n3043 VDD.n2782 3.4105
R11445 VDD.n3043 VDD.n2774 3.4105
R11446 VDD.n3043 VDD.n2781 3.4105
R11447 VDD.n3043 VDD.n2775 3.4105
R11448 VDD.n3043 VDD.n2780 3.4105
R11449 VDD.n3043 VDD.n2776 3.4105
R11450 VDD.n3043 VDD.n2779 3.4105
R11451 VDD.n3043 VDD.n3042 3.4105
R11452 VDD.n3042 VDD.n2793 3.4105
R11453 VDD.n3307 VDD.n3050 3.4105
R11454 VDD.n3047 VDD.n2770 3.4105
R11455 VDD.n3310 VDD.n3047 3.4105
R11456 VDD.n3050 VDD.n2770 3.4105
R11457 VDD.n3307 VDD.n3047 3.4105
R11458 VDD.n3056 VDD.n2772 3.4105
R11459 VDD.n3310 VDD.n2772 3.4105
R11460 VDD.n2772 VDD.n2770 3.4105
R11461 VDD.n3306 VDD.n2770 3.4105
R11462 VDD.n3307 VDD.n3306 3.4105
R11463 VDD.n3306 VDD.n3305 3.4105
R11464 VDD.n3056 VDD.n3050 3.4105
R11465 VDD.n3043 VDD.n2778 3.4105
R11466 VDD.n2786 VDD.n2778 3.4105
R11467 VDD.n5602 VDD.n18 3.4105
R11468 VDD.n5600 VDD.n6 3.4105
R11469 VDD.n10 VDD.n6 3.4105
R11470 VDD.n148 VDD.n6 3.4105
R11471 VDD.n5603 VDD.n6 3.4105
R11472 VDD.n147 VDD.n6 3.4105
R11473 VDD.n11 VDD.n6 3.4105
R11474 VDD.n12 VDD.n1 3.4105
R11475 VDD.n147 VDD.n1 3.4105
R11476 VDD.n21 VDD.n1 3.4105
R11477 VDD.n13 VDD.n1 3.4105
R11478 VDD.n19 VDD.n1 3.4105
R11479 VDD.n18 VDD.n1 3.4105
R11480 VDD.n5600 VDD.n1 3.4105
R11481 VDD.n10 VDD.n1 3.4105
R11482 VDD.n148 VDD.n1 3.4105
R11483 VDD.n5603 VDD.n8 3.4105
R11484 VDD.n5602 VDD.n16 3.4105
R11485 VDD.n5512 VDD.n6 3.4105
R11486 VDD.n13 VDD.n6 3.4105
R11487 VDD.n19 VDD.n6 3.4105
R11488 VDD.n5602 VDD.n19 3.4105
R11489 VDD.n19 VDD.n4 3.4105
R11490 VDD.n13 VDD.n4 3.4105
R11491 VDD.n5602 VDD.n13 3.4105
R11492 VDD.n5602 VDD.n21 3.4105
R11493 VDD.n16 VDD.n4 3.4105
R11494 VDD.n15 VDD.n6 3.4105
R11495 VDD.n15 VDD.n8 3.4105
R11496 VDD.n5512 VDD.n8 3.4105
R11497 VDD.n21 VDD.n8 3.4105
R11498 VDD.n21 VDD.n5 3.4105
R11499 VDD.n13 VDD.n5 3.4105
R11500 VDD.n13 VDD.n8 3.4105
R11501 VDD.n19 VDD.n8 3.4105
R11502 VDD.n19 VDD.n5 3.4105
R11503 VDD.n18 VDD.n5 3.4105
R11504 VDD.n18 VDD.n8 3.4105
R11505 VDD.n10 VDD.n5 3.4105
R11506 VDD.n10 VDD.n8 3.4105
R11507 VDD.n148 VDD.n8 3.4105
R11508 VDD.n148 VDD.n5 3.4105
R11509 VDD.n5603 VDD.n5 3.4105
R11510 VDD.n5603 VDD.n1 3.4105
R11511 VDD.n147 VDD.n8 3.4105
R11512 VDD.n147 VDD.n5 3.4105
R11513 VDD.n12 VDD.n5 3.4105
R11514 VDD.n11 VDD.n8 3.4105
R11515 VDD.n12 VDD.n4 3.4105
R11516 VDD.n5602 VDD.n12 3.4105
R11517 VDD.n5602 VDD.n147 3.4105
R11518 VDD.n147 VDD.n4 3.4105
R11519 VDD.n5603 VDD.n4 3.4105
R11520 VDD.n5603 VDD.n5602 3.4105
R11521 VDD.n5602 VDD.n148 3.4105
R11522 VDD.n148 VDD.n4 3.4105
R11523 VDD.n10 VDD.n4 3.4105
R11524 VDD.n5602 VDD.n10 3.4105
R11525 VDD.n18 VDD.n4 3.4105
R11526 VDD.n18 VDD.n6 3.4105
R11527 VDD.n5417 VDD.n305 3.39937
R11528 VDD.n5366 VDD.n324 3.39937
R11529 VDD.n367 VDD.n366 3.39937
R11530 VDD.n470 VDD.n469 3.39937
R11531 VDD.n524 VDD.n422 3.39937
R11532 VDD.n579 VDD.n399 3.39937
R11533 VDD.n5238 VDD.n5237 3.39937
R11534 VDD.n5189 VDD.n657 3.39937
R11535 VDD.n8861 VDD.n8677 3.39504
R11536 VDD.n8006 VDD.n7822 3.39504
R11537 VDD.n7152 VDD.n6968 3.39504
R11538 VDD.n6297 VDD.n6113 3.39504
R11539 VDD.n3607 VDD.n2640 3.38874
R11540 VDD.n3607 VDD.n2641 3.38874
R11541 VDD.n3574 VDD.n2682 3.38874
R11542 VDD.n3530 VDD.n3529 3.38874
R11543 VDD.n3465 VDD.n3464 3.38874
R11544 VDD.n3437 VDD.n2704 3.38874
R11545 VDD.n2719 VDD.n2715 3.38874
R11546 VDD.n3405 VDD.n2733 3.38874
R11547 VDD.n3383 VDD.n2740 3.38874
R11548 VDD.n3371 VDD.n3370 3.38874
R11549 VDD.n3298 VDD.n3297 3.38874
R11550 VDD.n3276 VDD.n3088 3.38874
R11551 VDD.n3232 VDD.n3231 3.38874
R11552 VDD.n3166 VDD.n3099 3.38874
R11553 VDD.n3166 VDD.n3100 3.38874
R11554 VDD.n3812 VDD.n3811 3.38874
R11555 VDD.n3816 VDD.n3815 3.38874
R11556 VDD.n3821 VDD.n3820 3.38874
R11557 VDD.n3927 VDD.n3659 3.38874
R11558 VDD.n3719 VDD.n3718 3.38874
R11559 VDD.n3724 VDD.n3723 3.38874
R11560 VDD.n3909 VDD.n3908 3.38874
R11561 VDD.n3905 VDD.n3904 3.38874
R11562 VDD.n3900 VDD.n3899 3.38874
R11563 VDD.n2858 VDD.n2804 3.38874
R11564 VDD.n2816 VDD.n2813 3.38874
R11565 VDD.n2843 VDD.n2812 3.38874
R11566 VDD.n2997 VDD.n2996 3.38874
R11567 VDD.n2993 VDD.n2950 3.38874
R11568 VDD.n2989 VDD.n2988 3.38874
R11569 VDD.n2988 VDD.n2953 3.38874
R11570 VDD.n1849 VDD.n1064 3.38874
R11571 VDD.n1824 VDD.n1079 3.38874
R11572 VDD.n2567 VDD.n2566 3.38874
R11573 VDD.n4737 VDD.n4735 3.38674
R11574 VDD.n4765 VDD.n895 3.38674
R11575 VDD.n4792 VDD.n4791 3.38674
R11576 VDD.n4825 VDD.n4824 3.38674
R11577 VDD.n4851 VDD.n4849 3.38674
R11578 VDD.n4879 VDD.n833 3.38674
R11579 VDD.n4906 VDD.n4905 3.38674
R11580 VDD.n4939 VDD.n4938 3.38674
R11581 VDD.n4965 VDD.n4963 3.38674
R11582 VDD.n4993 VDD.n771 3.38674
R11583 VDD.n5020 VDD.n5019 3.38674
R11584 VDD.n5053 VDD.n5052 3.38674
R11585 VDD.n5079 VDD.n5077 3.38674
R11586 VDD.n5107 VDD.n709 3.38674
R11587 VDD.n5134 VDD.n5133 3.38674
R11588 VDD.n3109 VDD.n2476 3.33963
R11589 VDD.n3110 VDD.n3109 3.33963
R11590 VDD.n3110 VDD.n2485 3.33963
R11591 VDD.n4006 VDD.n2485 3.33963
R11592 VDD.n3998 VDD.n2487 3.33963
R11593 VDD.n3998 VDD.n3997 3.33963
R11594 VDD.n3997 VDD.n3996 3.33963
R11595 VDD.n3996 VDD.n2491 3.33963
R11596 VDD.n2619 VDD.n2596 3.33963
R11597 VDD.n2626 VDD.n2596 3.33963
R11598 VDD.n2626 VDD.n2625 3.33963
R11599 VDD.n2625 VDD.n2598 3.33963
R11600 VDD.n5475 VDD.n266 3.33963
R11601 VDD.n5471 VDD.n266 3.33963
R11602 VDD.n5471 VDD.n5461 3.33963
R11603 VDD.n5461 VDD.n251 3.33963
R11604 VDD.n5504 VDD.n243 3.33963
R11605 VDD.n5504 VDD.n244 3.33963
R11606 VDD.n2444 VDD.n244 3.33963
R11607 VDD.n2449 VDD.n2444 3.33963
R11608 VDD.n3620 VDD.n3619 3.33963
R11609 VDD.n3619 VDD.n2504 3.33963
R11610 VDD.n3981 VDD.n2504 3.33963
R11611 VDD.n3981 VDD.n3980 3.33963
R11612 VDD.n3949 VDD.n3948 3.33963
R11613 VDD.n3955 VDD.n3949 3.33963
R11614 VDD.n3955 VDD.n3954 3.33963
R11615 VDD.n3954 VDD.n2495 3.33963
R11616 VDD.n1009 VDD.n1006 3.31902
R11617 VDD.n2008 VDD.n2005 3.31902
R11618 VDD.n2104 VDD.n2103 3.31902
R11619 VDD.n2229 VDD.n2226 3.31902
R11620 VDD.n1705 VDD.n1704 3.29555
R11621 VDD.n3585 VDD.n2662 3.2936
R11622 VDD.n3141 VDD.n3131 3.2936
R11623 VDD.n3788 VDD.n3765 3.2936
R11624 VDD.n2928 VDD.n2921 3.2936
R11625 VDD.n68 VDD.n67 3.2936
R11626 VDD.n5572 VDD.n5567 3.2936
R11627 VDD.n214 VDD.n213 3.2936
R11628 VDD.n5433 VDD.n5432 3.25474
R11629 VDD.n5382 VDD.n319 3.25474
R11630 VDD.n5333 VDD.n5332 3.25474
R11631 VDD.n452 VDD.n392 3.25474
R11632 VDD.n509 VDD.n430 3.25474
R11633 VDD.n564 VDD.n563 3.25474
R11634 VDD.n609 VDD.n605 3.25474
R11635 VDD.n5204 VDD.n645 3.25474
R11636 VDD.n5457 VDD.n5456 3.25377
R11637 VDD.n1440 VDD.n1437 3.25129
R11638 VDD.n4539 VDD.n1930 3.25129
R11639 VDD.n2050 VDD.n2036 3.25129
R11640 VDD.n4404 VDD.n2150 3.25129
R11641 VDD.n1255 VDD.n1098 3.23418
R11642 VDD.n1224 VDD.n1121 3.23418
R11643 VDD.n1203 VDD.n1133 3.23418
R11644 VDD.n1172 VDD.n1156 3.23418
R11645 VDD.n4588 VDD.n4587 3.23418
R11646 VDD.n4624 VDD.n975 3.23418
R11647 VDD.n4645 VDD.n4643 3.23418
R11648 VDD.n4679 VDD.n943 3.23418
R11649 VDD.n4699 VDD.n4698 3.23418
R11650 VDD.n1506 VDD.n1505 3.23218
R11651 VDD.n1553 VDD.n1332 3.23218
R11652 VDD.n1305 VDD.n1304 3.23218
R11653 VDD.n1630 VDD.n1627 3.23218
R11654 VDD.n1769 VDD.n1663 3.23218
R11655 VDD.n1734 VDD.n1701 3.23218
R11656 VDD.n5659 VDD.n5657 3.20702
R11657 VDD.n7368 VDD.n7366 3.20702
R11658 VDD.n2621 VDD.n1018 3.17466
R11659 VDD.n2600 VDD.n2599 3.17466
R11660 VDD.n8834 VDD.n8694 3.17267
R11661 VDD.n8833 VDD.n8832 3.17267
R11662 VDD.n8831 VDD.n8699 3.17267
R11663 VDD.n7979 VDD.n7839 3.17267
R11664 VDD.n7978 VDD.n7977 3.17267
R11665 VDD.n7976 VDD.n7844 3.17267
R11666 VDD.n7125 VDD.n6985 3.17267
R11667 VDD.n7124 VDD.n7123 3.17267
R11668 VDD.n7122 VDD.n6990 3.17267
R11669 VDD.n6270 VDD.n6130 3.17267
R11670 VDD.n6269 VDD.n6268 3.17267
R11671 VDD.n6267 VDD.n6135 3.17267
R11672 VDD.n1815 VDD.n1276 3.16717
R11673 VDD.n5492 VDD.n243 3.15412
R11674 VDD.n1853 VDD.n1852 3.13775
R11675 VDD.n1823 VDD.n1083 3.13775
R11676 VDD.n916 VDD.n911 3.11584
R11677 VDD.n4772 VDD.n890 3.11584
R11678 VDD.n4786 VDD.n880 3.11584
R11679 VDD.n4830 VDD.n860 3.11584
R11680 VDD.n854 VDD.n849 3.11584
R11681 VDD.n4886 VDD.n828 3.11584
R11682 VDD.n4900 VDD.n818 3.11584
R11683 VDD.n4944 VDD.n798 3.11584
R11684 VDD.n792 VDD.n787 3.11584
R11685 VDD.n5000 VDD.n766 3.11584
R11686 VDD.n5014 VDD.n756 3.11584
R11687 VDD.n5058 VDD.n736 3.11584
R11688 VDD.n730 VDD.n725 3.11584
R11689 VDD.n5114 VDD.n704 3.11584
R11690 VDD.n5128 VDD.n694 3.11584
R11691 VDD.n5421 VDD.n5418 3.1101
R11692 VDD.n5370 VDD.n5369 3.1101
R11693 VDD.n5321 VDD.n362 3.1101
R11694 VDD.n464 VDD.n446 3.1101
R11695 VDD.n523 VDD.n424 3.1101
R11696 VDD.n580 VDD.n578 3.1101
R11697 VDD.n619 VDD.n618 3.1101
R11698 VDD.n5190 VDD.n654 3.1101
R11699 VDD.n2337 VDD.n2335 3.10907
R11700 VDD.n2335 VDD.n2333 3.10907
R11701 VDD.n2333 VDD.n2331 3.10907
R11702 VDD.n2331 VDD.n2329 3.10907
R11703 VDD.n2329 VDD.n2327 3.10907
R11704 VDD.n2327 VDD.n2325 3.10907
R11705 VDD.n2325 VDD.n2323 3.10907
R11706 VDD.n2323 VDD.n2321 3.10907
R11707 VDD.n2321 VDD.n2319 3.10907
R11708 VDD.n2319 VDD.n2317 3.10907
R11709 VDD.n2317 VDD.n2315 3.10907
R11710 VDD.n2315 VDD.n2313 3.10907
R11711 VDD.n2313 VDD.n2311 3.10907
R11712 VDD.n2311 VDD.n2309 3.10907
R11713 VDD.n2309 VDD.n2307 3.10907
R11714 VDD.n2307 VDD.n2305 3.10907
R11715 VDD.n2305 VDD.n2303 3.10907
R11716 VDD.n2303 VDD.n2301 3.10907
R11717 VDD.n2301 VDD.n2299 3.10907
R11718 VDD.n2299 VDD.n2297 3.10907
R11719 VDD.n2297 VDD.n2295 3.10907
R11720 VDD.n2295 VDD.n2293 3.10907
R11721 VDD.n2293 VDD.n2291 3.10907
R11722 VDD.n2291 VDD.n2289 3.10907
R11723 VDD.n5630 VDD.n5629 3.10102
R11724 VDD.n6485 VDD.n6479 3.10102
R11725 VDD.n7339 VDD.n7338 3.10102
R11726 VDD.n8194 VDD.n8188 3.10102
R11727 VDD.n5622 VDD.n5614 3.09792
R11728 VDD.n6500 VDD.n6499 3.09792
R11729 VDD.n7331 VDD.n7323 3.09792
R11730 VDD.n8209 VDD.n8208 3.09792
R11731 VDD.n1905 VDD.n1902 3.04812
R11732 VDD.n2006 VDD.n1998 3.04812
R11733 VDD.n2125 VDD.n2122 3.04812
R11734 VDD.n2227 VDD.n2219 3.04812
R11735 VDD.n3936 VDD.n3935 3.03311
R11736 VDD.n3763 VDD.n3646 3.03311
R11737 VDD.n3929 VDD.n3928 3.03311
R11738 VDD.n3677 VDD.n3676 3.03311
R11739 VDD.n2887 VDD.n2869 3.03311
R11740 VDD.n2859 VDD.n2796 3.03311
R11741 VDD.n2916 VDD.n2894 3.03311
R11742 VDD.n94 VDD.n32 3.03311
R11743 VDD.n5552 VDD.n160 3.03311
R11744 VDD.n5509 VDD.n170 3.03311
R11745 VDD.n139 VDD.n28 3.03311
R11746 VDD.n2444 VDD.n238 3.03311
R11747 VDD.n5505 VDD.n5504 3.03311
R11748 VDD.n5485 VDD.n251 3.03311
R11749 VDD.n5476 VDD.n5475 3.03311
R11750 VDD.n5471 VDD.n5470 3.03311
R11751 VDD.n2598 VDD.n2591 3.03311
R11752 VDD.n2906 VDD.n2491 3.03311
R11753 VDD.n3997 VDD.n2490 3.03311
R11754 VDD.n4006 VDD.n2486 3.03311
R11755 VDD.n2899 VDD.n2487 3.03311
R11756 VDD.n3956 VDD.n3955 3.03311
R11757 VDD.n3948 VDD.n3623 3.03311
R11758 VDD.n3630 VDD.n2495 3.03311
R11759 VDD.n3977 VDD.n3620 3.03311
R11760 VDD.n2569 VDD.n2519 3.03311
R11761 VDD.n3115 VDD.n3110 3.03311
R11762 VDD.n3617 VDD.n2504 3.03311
R11763 VDD.n2619 VDD.n2592 3.03311
R11764 VDD.n2627 VDD.n2626 3.03311
R11765 VDD.n3980 VDD.n3979 3.03311
R11766 VDD.n3112 VDD.n2476 3.03311
R11767 VDD.n2684 VDD.n2640 3.01226
R11768 VDD.n2651 VDD.n2641 3.01226
R11769 VDD.n3579 VDD.n2682 3.01226
R11770 VDD.n3529 VDD.n3528 3.01226
R11771 VDD.n3467 VDD.n3465 3.01226
R11772 VDD.n3436 VDD.n2704 3.01226
R11773 VDD.n3427 VDD.n2715 3.01226
R11774 VDD.n3414 VDD.n2733 3.01226
R11775 VDD.n3382 VDD.n2740 3.01226
R11776 VDD.n3358 VDD.n3355 3.01226
R11777 VDD.n3371 VDD.n3351 3.01226
R11778 VDD.n3286 VDD.n3284 3.01226
R11779 VDD.n3298 VDD.n3072 3.01226
R11780 VDD.n3281 VDD.n3088 3.01226
R11781 VDD.n3231 VDD.n3230 3.01226
R11782 VDD.n3099 VDD.n3098 3.01226
R11783 VDD.n3104 VDD.n3100 3.01226
R11784 VDD.n3817 VDD.n3816 3.01226
R11785 VDD.n3822 VDD.n3821 3.01226
R11786 VDD.n3720 VDD.n3719 3.01226
R11787 VDD.n3725 VDD.n3724 3.01226
R11788 VDD.n3904 VDD.n3903 3.01226
R11789 VDD.n3899 VDD.n3898 3.01226
R11790 VDD.n2847 VDD.n2813 3.01226
R11791 VDD.n2843 VDD.n2842 3.01226
R11792 VDD.n2952 VDD.n2950 3.01226
R11793 VDD.n2990 VDD.n2989 3.01226
R11794 VDD.n2957 VDD.n2953 3.01226
R11795 VDD.n96 VDD.n95 3.01226
R11796 VDD.n5554 VDD.n5553 3.01226
R11797 VDD.n195 VDD.n194 3.01226
R11798 VDD.n2575 VDD.n2520 3.01226
R11799 VDD.n2567 VDD.n2519 3.01226
R11800 VDD.n1411 VDD.n1410 2.98039
R11801 VDD.n4543 VDD.n4542 2.98039
R11802 VDD.n4476 VDD.n2035 2.98039
R11803 VDD.n4408 VDD.n4407 2.98039
R11804 VDD.n1510 VDD.n1509 2.97872
R11805 VDD.n1550 VDD.n1548 2.97872
R11806 VDD.n1596 VDD.n1595 2.97872
R11807 VDD.n1625 VDD.n1285 2.97872
R11808 VDD.n1767 VDD.n1664 2.97872
R11809 VDD.n1738 VDD.n1737 2.97872
R11810 VDD.n5430 VDD.n5429 2.96547
R11811 VDD.n5381 VDD.n320 2.96547
R11812 VDD.n357 VDD.n353 2.96547
R11813 VDD.n455 VDD.n454 2.96547
R11814 VDD.n510 VDD.n428 2.96547
R11815 VDD.n569 VDD.n406 2.96547
R11816 VDD.n5249 VDD.n610 2.96547
R11817 VDD.n5201 VDD.n5200 2.96547
R11818 VDD.n1259 VDD.n1258 2.96471
R11819 VDD.n1221 VDD.n1220 2.96471
R11820 VDD.n1207 VDD.n1206 2.96471
R11821 VDD.n1169 VDD.n1168 2.96471
R11822 VDD.n4582 VDD.n996 2.96471
R11823 VDD.n4623 VDD.n976 2.96471
R11824 VDD.n969 VDD.n964 2.96471
R11825 VDD.n4681 VDD.n4680 2.96471
R11826 VDD.n4693 VDD.n933 2.96471
R11827 VDD.n3812 VDD.n3761 2.96007
R11828 VDD.n3660 VDD.n3659 2.96007
R11829 VDD.n3908 VDD.n3668 2.96007
R11830 VDD.n2806 VDD.n2804 2.96007
R11831 VDD.n4289 VDD.n2364 2.91154
R11832 VDD.n4239 VDD.n4238 2.91154
R11833 VDD.n4092 VDD.n4091 2.91154
R11834 VDD.n4150 VDD.n4054 2.91154
R11835 VDD.n2615 VDD.n1953 2.91015
R11836 VDD.n1857 VDD.n1062 2.88677
R11837 VDD.n1820 VDD.n1819 2.88677
R11838 VDD.n2404 VDD.n2403 2.86873
R11839 VDD.n4090 VDD.n4084 2.86873
R11840 VDD.n4151 VDD.n4053 2.86873
R11841 VDD.n3024 VDD.n2888 2.85341
R11842 VDD.n4729 VDD.n4728 2.84494
R11843 VDD.n4774 VDD.n4773 2.84494
R11844 VDD.n4787 VDD.n4785 2.84494
R11845 VDD.n4829 VDD.n861 2.84494
R11846 VDD.n4843 VDD.n4842 2.84494
R11847 VDD.n4888 VDD.n4887 2.84494
R11848 VDD.n4901 VDD.n4899 2.84494
R11849 VDD.n4943 VDD.n799 2.84494
R11850 VDD.n4957 VDD.n4956 2.84494
R11851 VDD.n5002 VDD.n5001 2.84494
R11852 VDD.n5015 VDD.n5013 2.84494
R11853 VDD.n5057 VDD.n737 2.84494
R11854 VDD.n5071 VDD.n5070 2.84494
R11855 VDD.n5116 VDD.n5115 2.84494
R11856 VDD.n5129 VDD.n5127 2.84494
R11857 VDD.n5422 VDD.n302 2.82084
R11858 VDD.n5373 VDD.n323 2.82084
R11859 VDD.n5322 VDD.n359 2.82084
R11860 VDD.n463 VDD.n448 2.82084
R11861 VDD.n520 VDD.n519 2.82084
R11862 VDD.n574 VDD.n402 2.82084
R11863 VDD.n5244 VDD.n614 2.82084
R11864 VDD.n5194 VDD.n5193 2.82084
R11865 VDD.n4283 VDD.n2370 2.78311
R11866 VDD.n4237 VDD.n2405 2.78311
R11867 VDD.n4098 VDD.n4080 2.78311
R11868 VDD.n4156 VDD.n4050 2.78311
R11869 VDD.n1466 VDD.n1401 2.77722
R11870 VDD.n1903 VDD.n1021 2.77722
R11871 VDD.n4498 VDD.n1999 2.77722
R11872 VDD.n2123 VDD.n2115 2.77722
R11873 VDD.n4363 VDD.n2220 2.77722
R11874 VDD.n2577 VDD.t47 2.77
R11875 VDD.n2577 VDD.t101 2.77
R11876 VDD.n1356 VDD.n1355 2.72525
R11877 VDD.n1339 VDD.n1338 2.72525
R11878 VDD.n1600 VDD.n1599 2.72525
R11879 VDD.n1808 VDD.n1284 2.72525
R11880 VDD.n1764 VDD.n1763 2.72525
R11881 VDD.n1697 VDD.n1694 2.72525
R11882 VDD.n1448 VDD.n1445 2.70949
R11883 VDD.n1935 VDD.n1934 2.70949
R11884 VDD.n4480 VDD.n4479 2.70949
R11885 VDD.n2155 VDD.n2154 2.70949
R11886 VDD.n4245 VDD.n2400 2.69749
R11887 VDD.n4087 VDD.n4086 2.69749
R11888 VDD.n4144 VDD.n4143 2.69749
R11889 VDD.n1269 VDD.n1268 2.69524
R11890 VDD.n1263 VDD.n1093 2.69524
R11891 VDD.n1216 VDD.n1123 2.69524
R11892 VDD.n1211 VDD.n1129 2.69524
R11893 VDD.n1164 VDD.n1158 2.69524
R11894 VDD.n4583 VDD.n4581 2.69524
R11895 VDD.n4630 VDD.n971 2.69524
R11896 VDD.n4637 VDD.n4636 2.69524
R11897 VDD.n4686 VDD.n940 2.69524
R11898 VDD.n4694 VDD.n4692 2.69524
R11899 VDD.n5475 VDD.n265 2.69036
R11900 VDD.n5426 VDD.n301 2.67621
R11901 VDD.n5378 VDD.n5377 2.67621
R11902 VDD.n5326 VDD.n358 2.67621
R11903 VDD.n459 VDD.n450 2.67621
R11904 VDD.n514 VDD.n513 2.67621
R11905 VDD.n570 VDD.n404 2.67621
R11906 VDD.n5248 VDD.n611 2.67621
R11907 VDD.n652 VDD.n648 2.67621
R11908 VDD.n8317 VDD.n8282 2.64609
R11909 VDD.n7462 VDD.n7427 2.64609
R11910 VDD.n6608 VDD.n6573 2.64609
R11911 VDD.n5753 VDD.n5718 2.64609
R11912 VDD.n4492 VDD.n2014 2.64563
R11913 VDD.n3951 VDD.n2021 2.64563
R11914 VDD.n2654 VDD.n2653 2.63579
R11915 VDD.n2655 VDD.n2654 2.63579
R11916 VDD.n3570 VDD.n3479 2.63579
R11917 VDD.n3535 VDD.n3534 2.63579
R11918 VDD.n3459 VDD.n2699 2.63579
R11919 VDD.n3443 VDD.n3441 2.63579
R11920 VDD.n2724 VDD.n2723 2.63579
R11921 VDD.n3418 VDD.n3401 2.63579
R11922 VDD.n3389 VDD.n3387 2.63579
R11923 VDD.n3365 VDD.n3364 2.63579
R11924 VDD.n3293 VDD.n3292 2.63579
R11925 VDD.n3272 VDD.n3181 2.63579
R11926 VDD.n3237 VDD.n3236 2.63579
R11927 VDD.n3161 VDD.n3105 2.63579
R11928 VDD.n3124 VDD.n3105 2.63579
R11929 VDD.n2993 VDD.n2917 2.63579
R11930 VDD.n48 VDD.n45 2.63579
R11931 VDD.n120 VDD.n113 2.63579
R11932 VDD.n2349 VDD.n2347 2.63579
R11933 VDD.n5549 VDD.n5545 2.63579
R11934 VDD.n193 VDD.n190 2.63579
R11935 VDD.n1275 VDD.n1085 2.63579
R11936 VDD.n2579 VDD.n2511 2.63579
R11937 VDD.n4282 VDD.n2371 2.61187
R11938 VDD.n4234 VDD.n4233 2.61187
R11939 VDD.n4100 VDD.n4099 2.61187
R11940 VDD.n4155 VDD.n4051 2.61187
R11941 VDD.n4723 VDD.n915 2.57404
R11942 VDD.n4779 VDD.n887 2.57404
R11943 VDD.n888 VDD.n883 2.57404
R11944 VDD.n4836 VDD.n856 2.57404
R11945 VDD.n4837 VDD.n853 2.57404
R11946 VDD.n4893 VDD.n825 2.57404
R11947 VDD.n826 VDD.n821 2.57404
R11948 VDD.n4950 VDD.n794 2.57404
R11949 VDD.n4951 VDD.n791 2.57404
R11950 VDD.n5007 VDD.n763 2.57404
R11951 VDD.n764 VDD.n759 2.57404
R11952 VDD.n5064 VDD.n732 2.57404
R11953 VDD.n5065 VDD.n729 2.57404
R11954 VDD.n5121 VDD.n701 2.57404
R11955 VDD.n702 VDD.n697 2.57404
R11956 VDD.n8859 VDD.n8858 2.56805
R11957 VDD.n8759 VDD.n8692 2.56805
R11958 VDD.n8760 VDD.n8759 2.56805
R11959 VDD.n8765 VDD.n8763 2.56805
R11960 VDD.n8767 VDD.n8765 2.56805
R11961 VDD.n8786 VDD.n8784 2.56805
R11962 VDD.n8004 VDD.n8003 2.56805
R11963 VDD.n7904 VDD.n7837 2.56805
R11964 VDD.n7905 VDD.n7904 2.56805
R11965 VDD.n7910 VDD.n7908 2.56805
R11966 VDD.n7912 VDD.n7910 2.56805
R11967 VDD.n7931 VDD.n7929 2.56805
R11968 VDD.n7150 VDD.n7149 2.56805
R11969 VDD.n7050 VDD.n6983 2.56805
R11970 VDD.n7051 VDD.n7050 2.56805
R11971 VDD.n7056 VDD.n7054 2.56805
R11972 VDD.n7058 VDD.n7056 2.56805
R11973 VDD.n7077 VDD.n7075 2.56805
R11974 VDD.n6295 VDD.n6294 2.56805
R11975 VDD.n6195 VDD.n6128 2.56805
R11976 VDD.n6196 VDD.n6195 2.56805
R11977 VDD.n6201 VDD.n6199 2.56805
R11978 VDD.n6203 VDD.n6201 2.56805
R11979 VDD.n6222 VDD.n6220 2.56805
R11980 VDD.n119 VDD.n109 2.56676
R11981 VDD.n8262 VDD.n8248 2.5605
R11982 VDD.n9009 VDD.n8263 2.5605
R11983 VDD.n7407 VDD.n7393 2.5605
R11984 VDD.n8154 VDD.n7408 2.5605
R11985 VDD.n6553 VDD.n6539 2.5605
R11986 VDD.n7300 VDD.n6554 2.5605
R11987 VDD.n5698 VDD.n5684 2.5605
R11988 VDD.n6445 VDD.n5699 2.5605
R11989 VDD.n5426 VDD.n5425 2.53157
R11990 VDD.n5377 VDD.n5374 2.53157
R11991 VDD.n5326 VDD.n5325 2.53157
R11992 VDD.n460 VDD.n459 2.53157
R11993 VDD.n514 VDD.n426 2.53157
R11994 VDD.n573 VDD.n404 2.53157
R11995 VDD.n5245 VDD.n611 2.53157
R11996 VDD.n653 VDD.n652 2.53157
R11997 VDD.n4246 VDD.n2397 2.52625
R11998 VDD.n4142 VDD.n4058 2.52625
R11999 VDD.n9030 VDD 2.50745
R12000 VDD.n1463 VDD.n1462 2.50632
R12001 VDD.n4561 VDD.n1022 2.50632
R12002 VDD.n4495 VDD.n4494 2.50632
R12003 VDD.n4426 VDD.n2116 2.50632
R12004 VDD.n4360 VDD.n4359 2.50632
R12005 VDD.n1521 VDD.n1520 2.47179
R12006 VDD.n1538 VDD.n1537 2.47179
R12007 VDD.n1607 VDD.n1294 2.47179
R12008 VDD.n1812 VDD.n1811 2.47179
R12009 VDD.n1676 VDD.n1675 2.47179
R12010 VDD.n1692 VDD.n1685 2.47179
R12011 VDD.n4279 VDD.n4278 2.44063
R12012 VDD.n2415 VDD.n2408 2.44063
R12013 VDD.n4105 VDD.n4077 2.44063
R12014 VDD.n4162 VDD.n4046 2.44063
R12015 VDD.n1452 VDD.n1409 2.4386
R12016 VDD.n1933 VDD.n1916 2.4386
R12017 VDD.n2040 VDD.n2039 2.4386
R12018 VDD.n2153 VDD.n2135 2.4386
R12019 VDD.n8335 VDD.n8290 2.43651
R12020 VDD.n7480 VDD.n7435 2.43651
R12021 VDD.n6626 VDD.n6581 2.43651
R12022 VDD.n5771 VDD.n5726 2.43651
R12023 VDD.n1267 VDD.n1091 2.42576
R12024 VDD.n1264 VDD.n1091 2.42576
R12025 VDD.n1215 VDD.n1127 2.42576
R12026 VDD.n1212 VDD.n1127 2.42576
R12027 VDD.n1163 VDD.n1161 2.42576
R12028 VDD.n1161 VDD.n999 2.42576
R12029 VDD.n4632 VDD.n4631 2.42576
R12030 VDD.n4631 VDD.n968 2.42576
R12031 VDD.n4685 VDD.n941 2.42576
R12032 VDD.n941 VDD.n936 2.42576
R12033 VDD.n6523 VDD.n6522 2.42534
R12034 VDD.n8232 VDD.n8231 2.42534
R12035 VDD.n5425 VDD.n302 2.38694
R12036 VDD.n5374 VDD.n5373 2.38694
R12037 VDD.n5325 VDD.n359 2.38694
R12038 VDD.n460 VDD.n448 2.38694
R12039 VDD.n519 VDD.n426 2.38694
R12040 VDD.n574 VDD.n573 2.38694
R12041 VDD.n5245 VDD.n5244 2.38694
R12042 VDD.n5194 VDD.n653 2.38694
R12043 VDD.n5159 VDD.n675 2.38694
R12044 VDD.n2577 VDD.n2509 2.37942
R12045 VDD.n2356 VDD.n2355 2.3755
R12046 VDD.n4359 VDD.n2224 2.37087
R12047 VDD.n1270 VDD.n1269 2.35839
R12048 VDD.n4250 VDD.n4249 2.35502
R12049 VDD.n4201 VDD.n2435 2.35502
R12050 VDD.n4139 VDD.n4138 2.35502
R12051 VDD.n5634 VDD.n5626 2.30684
R12052 VDD.n6484 VDD.n6483 2.30684
R12053 VDD.n7343 VDD.n7335 2.30684
R12054 VDD.n8193 VDD.n8192 2.30684
R12055 VDD.n4724 VDD.n4723 2.30315
R12056 VDD.n4779 VDD.n4778 2.30315
R12057 VDD.n4778 VDD.n888 2.30315
R12058 VDD.n4838 VDD.n4836 2.30315
R12059 VDD.n4838 VDD.n4837 2.30315
R12060 VDD.n4893 VDD.n4892 2.30315
R12061 VDD.n4892 VDD.n826 2.30315
R12062 VDD.n4952 VDD.n4950 2.30315
R12063 VDD.n4952 VDD.n4951 2.30315
R12064 VDD.n5007 VDD.n5006 2.30315
R12065 VDD.n5006 VDD.n764 2.30315
R12066 VDD.n5066 VDD.n5064 2.30315
R12067 VDD.n5066 VDD.n5065 2.30315
R12068 VDD.n5121 VDD.n5120 2.30315
R12069 VDD.n5120 VDD.n702 2.30315
R12070 VDD.n102 VDD.n38 2.28225
R12071 VDD.n136 VDD.n108 2.28225
R12072 VDD.n5587 VDD.n5560 2.28225
R12073 VDD.n202 VDD.n201 2.28225
R12074 VDD.n2377 VDD.n2373 2.2694
R12075 VDD.n4227 VDD.n2416 2.2694
R12076 VDD.n4104 VDD.n4078 2.2694
R12077 VDD.n4164 VDD.n4163 2.2694
R12078 VDD.n3112 VDD.n3106 2.25953
R12079 VDD.n3611 VDD.n2638 2.25932
R12080 VDD.n3524 VDD.n3523 2.25932
R12081 VDD.n3226 VDD.n3225 2.25932
R12082 VDD.n3170 VDD.n3095 2.25932
R12083 VDD.n3794 VDD.n3793 2.25932
R12084 VDD.n3827 VDD.n3826 2.25932
R12085 VDD.n3916 VDD.n3911 2.25932
R12086 VDD.n3730 VDD.n3729 2.25932
R12087 VDD.n3693 VDD.n3692 2.25932
R12088 VDD.n3894 VDD.n3893 2.25932
R12089 VDD.n3778 VDD.n3774 2.25932
R12090 VDD.n2854 VDD.n2849 2.25932
R12091 VDD.n2838 VDD.n2837 2.25932
R12092 VDD.n2879 VDD.n2877 2.25932
R12093 VDD.n2933 VDD.n2932 2.25932
R12094 VDD.n2985 VDD.n2984 2.25932
R12095 VDD.n2980 VDD.n2958 2.25932
R12096 VDD.n90 VDD.n49 2.25932
R12097 VDD.n52 VDD.n51 2.25932
R12098 VDD.n124 VDD.n116 2.25932
R12099 VDD.n129 VDD.n125 2.25932
R12100 VDD.n5595 VDD.n5528 2.25932
R12101 VDD.n5535 VDD.n5532 2.25932
R12102 VDD.n236 VDD.n176 2.25932
R12103 VDD.n227 VDD.n180 2.25932
R12104 VDD.n2566 VDD.n2565 2.25932
R12105 VDD.n131 VDD.n124 2.25379
R12106 VDD.n3362 VDD.n2765 2.25051
R12107 VDD.n3290 VDD.n3064 2.25051
R12108 VDD.n5634 VDD.n5633 2.2505
R12109 VDD.n5635 VDD.n5621 2.2505
R12110 VDD.n5637 VDD.n5636 2.2505
R12111 VDD.n5624 VDD.n5613 2.2505
R12112 VDD.n5672 VDD.n5671 2.2505
R12113 VDD.n6483 VDD.n6482 2.2505
R12114 VDD.n6476 VDD.n6475 2.2505
R12115 VDD.n6494 VDD.n6493 2.2505
R12116 VDD.n6497 VDD.n6496 2.2505
R12117 VDD.n6495 VDD.n6473 2.2505
R12118 VDD.n7343 VDD.n7342 2.2505
R12119 VDD.n7344 VDD.n7330 2.2505
R12120 VDD.n7346 VDD.n7345 2.2505
R12121 VDD.n7333 VDD.n7322 2.2505
R12122 VDD.n7381 VDD.n7380 2.2505
R12123 VDD.n8192 VDD.n8191 2.2505
R12124 VDD.n8185 VDD.n8184 2.2505
R12125 VDD.n8203 VDD.n8202 2.2505
R12126 VDD.n8206 VDD.n8205 2.2505
R12127 VDD.n8204 VDD.n8182 2.2505
R12128 VDD.n3396 VDD.n2744 2.25002
R12129 VDD.n2728 VDD.n2718 2.25002
R12130 VDD.n3604 VDD.n3603 2.25002
R12131 VDD.n3450 VDD.n2708 2.25002
R12132 VDD.n3353 VDD.n2765 2.24905
R12133 VDD.n3073 VDD.n3064 2.24905
R12134 VDD.n3102 VDD.n3101 2.24807
R12135 VDD.n3278 VDD.n3179 2.24807
R12136 VDD.n3410 VDD.n2734 2.24807
R12137 VDD.n2697 VDD.n2696 2.24807
R12138 VDD.n3576 VDD.n3477 2.24807
R12139 VDD.n3935 VDD.n3635 2.24691
R12140 VDD.n3696 VDD.n3678 2.24691
R12141 VDD.n3651 VDD.n3644 2.24691
R12142 VDD.n3923 VDD.n3653 2.24691
R12143 VDD.n2900 VDD.n2490 2.24691
R12144 VDD.n2863 VDD.n2801 2.24691
R12145 VDD.n3002 VDD.n2893 2.24691
R12146 VDD.n5588 VDD.n162 2.24691
R12147 VDD.n137 VDD.n25 2.24691
R12148 VDD.n104 VDD.n103 2.24691
R12149 VDD.n237 VDD.n167 2.24691
R12150 VDD.n5506 VDD.n5505 2.24691
R12151 VDD.n3630 VDD.n3625 2.24691
R12152 VDD.n3178 VDD.n3177 2.24691
R12153 VDD.n3160 VDD.n3091 2.24691
R12154 VDD.n3372 VDD.n3349 2.24691
R12155 VDD.n3420 VDD.n2730 2.24691
R12156 VDD.n3380 VDD.n2737 2.24691
R12157 VDD.n3425 VDD.n2709 2.24691
R12158 VDD.n2686 VDD.n2633 2.24691
R12159 VDD.n3476 VDD.n3475 2.24691
R12160 VDD.n3458 VDD.n2690 2.24691
R12161 VDD.n3434 VDD.n2701 2.24691
R12162 VDD.n3679 VDD.n3677 2.24671
R12163 VDD.n3941 VDD.n3638 2.24671
R12164 VDD.n3650 VDD.n3645 2.24671
R12165 VDD.n2904 VDD.n2490 2.24671
R12166 VDD.n2891 VDD.n2871 2.24671
R12167 VDD.n172 VDD.n166 2.24671
R12168 VDD.n106 VDD.n23 2.24671
R12169 VDD.n81 VDD.n30 2.24671
R12170 VDD.n3113 VDD.n3112 2.24671
R12171 VDD.n3173 VDD.n3092 2.24671
R12172 VDD.n3271 VDD.n3182 2.24671
R12173 VDD.n3398 VDD.n2739 2.24671
R12174 VDD.n2735 VDD.n2731 2.24671
R12175 VDD.n3452 VDD.n2703 2.24671
R12176 VDD.n3431 VDD.n2712 2.24671
R12177 VDD.n3471 VDD.n2692 2.24671
R12178 VDD.n3569 VDD.n3480 2.24671
R12179 VDD.n3614 VDD.n2636 2.24671
R12180 VDD.n3700 VDD.n3680 2.24661
R12181 VDD.n3807 VDD.n3806 2.24661
R12182 VDD.n102 VDD.n40 2.24613
R12183 VDD.n136 VDD.n109 2.24613
R12184 VDD.n5560 VDD.n5541 2.24613
R12185 VDD.n201 VDD.n185 2.24613
R12186 VDD.n240 VDD.n239 2.24365
R12187 VDD.n5429 VDD.n301 2.24231
R12188 VDD.n5378 VDD.n320 2.24231
R12189 VDD.n358 VDD.n357 2.24231
R12190 VDD.n455 VDD.n450 2.24231
R12191 VDD.n513 VDD.n428 2.24231
R12192 VDD.n570 VDD.n569 2.24231
R12193 VDD.n5249 VDD.n5248 2.24231
R12194 VDD.n5200 VDD.n648 2.24231
R12195 VDD.n3275 VDD.n3179 2.23886
R12196 VDD.n3065 VDD.n3064 2.23886
R12197 VDD.n3070 VDD.n3064 2.23886
R12198 VDD.n3164 VDD.n3102 2.23886
R12199 VDD.n3410 VDD.n3409 2.23886
R12200 VDD.n3396 VDD.n2743 2.23886
R12201 VDD.n2728 VDD.n2727 2.23886
R12202 VDD.n3573 VDD.n3477 2.23886
R12203 VDD.n3605 VDD.n3604 2.23886
R12204 VDD.n3462 VDD.n2697 2.23886
R12205 VDD.n3450 VDD.n2707 2.23886
R12206 VDD.n1459 VDD.n1406 2.23542
R12207 VDD.n4558 VDD.n4557 2.23542
R12208 VDD.n2019 VDD.n2018 2.23542
R12209 VDD.n4423 VDD.n4422 2.23542
R12210 VDD.n3804 VDD.n3803 2.22452
R12211 VDD.n3924 VDD.n3662 2.22452
R12212 VDD.n3685 VDD.n3669 2.22452
R12213 VDD.n2803 VDD.n2799 2.22452
R12214 VDD.n3026 VDD.n3025 2.22452
R12215 VDD.n1525 VDD.n1524 2.21832
R12216 VDD.n1534 VDD.n1533 2.21832
R12217 VDD.n1609 VDD.n1292 2.21832
R12218 VDD.n1288 VDD.n1287 2.21832
R12219 VDD.n1754 VDD.n1680 2.21832
R12220 VDD.n1749 VDD.n1684 2.21832
R12221 VDD.n6525 VDD.n6524 2.19693
R12222 VDD.n8234 VDD.n8233 2.19693
R12223 VDD.n2396 VDD.n2395 2.18378
R12224 VDD.n4205 VDD.n4204 2.18378
R12225 VDD.n4064 VDD.n4060 2.18378
R12226 VDD.n4193 VDD.n4029 2.18378
R12227 VDD.n1458 VDD.n1455 2.1677
R12228 VDD.n1914 VDD.n1026 2.1677
R12229 VDD.n2038 VDD.n2020 2.1677
R12230 VDD.n2133 VDD.n2120 2.1677
R12231 VDD.n1268 VDD.n1267 2.15629
R12232 VDD.n1264 VDD.n1263 2.15629
R12233 VDD.n1216 VDD.n1215 2.15629
R12234 VDD.n1212 VDD.n1211 2.15629
R12235 VDD.n1164 VDD.n1163 2.15629
R12236 VDD.n4581 VDD.n999 2.15629
R12237 VDD.n4632 VDD.n4630 2.15629
R12238 VDD.n4637 VDD.n968 2.15629
R12239 VDD.n4686 VDD.n4685 2.15629
R12240 VDD.n4692 VDD.n936 2.15629
R12241 VDD.t46 VDD.n1941 2.11661
R12242 VDD.n4469 VDD.t106 2.11661
R12243 VDD.n3937 VDD.n3643 2.10401
R12244 VDD.n4220 VDD.t40 2.1032
R12245 VDD.n4272 VDD.n2378 2.09816
R12246 VDD.n4226 VDD.n2417 2.09816
R12247 VDD.n4111 VDD.n4073 2.09816
R12248 VDD.n4169 VDD.n4043 2.09816
R12249 VDD.n5422 VDD.n5421 2.09768
R12250 VDD.n5370 VDD.n323 2.09768
R12251 VDD.n5322 VDD.n5321 2.09768
R12252 VDD.n464 VDD.n463 2.09768
R12253 VDD.n520 VDD.n424 2.09768
R12254 VDD.n578 VDD.n402 2.09768
R12255 VDD.n618 VDD.n614 2.09768
R12256 VDD.n5193 VDD.n654 2.09768
R12257 VDD.n2339 VDD.n2337 2.07664
R12258 VDD.n5657 VDD.n5653 2.0723
R12259 VDD.n7366 VDD.n7362 2.0723
R12260 VDD.n4729 VDD.n915 2.03225
R12261 VDD.n4773 VDD.n887 2.03225
R12262 VDD.n4785 VDD.n883 2.03225
R12263 VDD.n861 VDD.n856 2.03225
R12264 VDD.n4843 VDD.n853 2.03225
R12265 VDD.n4887 VDD.n825 2.03225
R12266 VDD.n4899 VDD.n821 2.03225
R12267 VDD.n799 VDD.n794 2.03225
R12268 VDD.n4957 VDD.n791 2.03225
R12269 VDD.n5001 VDD.n763 2.03225
R12270 VDD.n5013 VDD.n759 2.03225
R12271 VDD.n737 VDD.n732 2.03225
R12272 VDD.n5071 VDD.n729 2.03225
R12273 VDD.n5115 VDD.n701 2.03225
R12274 VDD.n5127 VDD.n697 2.03225
R12275 VDD.n4256 VDD.n2391 2.01254
R12276 VDD.n2434 VDD.n2433 2.01254
R12277 VDD.n4132 VDD.n4131 2.01254
R12278 VDD.n4190 VDD.n4189 2.01254
R12279 VDD.n8820 VDD.n8819 2.00398
R12280 VDD.n8818 VDD.n8713 2.00398
R12281 VDD.n8360 VDD.n8359 2.00398
R12282 VDD.n7965 VDD.n7964 2.00398
R12283 VDD.n7963 VDD.n7858 2.00398
R12284 VDD.n7505 VDD.n7504 2.00398
R12285 VDD.n7111 VDD.n7110 2.00398
R12286 VDD.n7109 VDD.n7004 2.00398
R12287 VDD.n6651 VDD.n6650 2.00398
R12288 VDD.n6256 VDD.n6255 2.00398
R12289 VDD.n6254 VDD.n6149 2.00398
R12290 VDD.n5796 VDD.n5795 2.00398
R12291 VDD.n4577 VDD.n1001 1.98435
R12292 VDD.n8581 VDD.n8530 1.97774
R12293 VDD.n7726 VDD.n7675 1.97774
R12294 VDD.n6872 VDD.n6821 1.97774
R12295 VDD.n6017 VDD.n5966 1.97774
R12296 VDD.n1526 VDD.n1345 1.96486
R12297 VDD.n1532 VDD.n1345 1.96486
R12298 VDD.n1613 VDD.n1612 1.96486
R12299 VDD.n1612 VDD.n1289 1.96486
R12300 VDD.n1753 VDD.n1752 1.96486
R12301 VDD.n1752 VDD.n1681 1.96486
R12302 VDD.n1455 VDD.n1407 1.96452
R12303 VDD.n1915 VDD.n1914 1.96452
R12304 VDD.n2041 VDD.n2038 1.96452
R12305 VDD.n2134 VDD.n2133 1.96452
R12306 VDD.n8858 VDD.n8856 1.96392
R12307 VDD.n8689 VDD.n8680 1.96392
R12308 VDD.n8850 VDD.n8691 1.96392
R12309 VDD.n8849 VDD.n8847 1.96392
R12310 VDD.n8846 VDD.n8844 1.96392
R12311 VDD.n8842 VDD.n8840 1.96392
R12312 VDD.n8003 VDD.n8001 1.96392
R12313 VDD.n7834 VDD.n7825 1.96392
R12314 VDD.n7995 VDD.n7836 1.96392
R12315 VDD.n7994 VDD.n7992 1.96392
R12316 VDD.n7991 VDD.n7989 1.96392
R12317 VDD.n7987 VDD.n7985 1.96392
R12318 VDD.n7149 VDD.n7147 1.96392
R12319 VDD.n6980 VDD.n6971 1.96392
R12320 VDD.n7141 VDD.n6982 1.96392
R12321 VDD.n7140 VDD.n7138 1.96392
R12322 VDD.n7137 VDD.n7135 1.96392
R12323 VDD.n7133 VDD.n7131 1.96392
R12324 VDD.n6294 VDD.n6292 1.96392
R12325 VDD.n6125 VDD.n6116 1.96392
R12326 VDD.n6286 VDD.n6127 1.96392
R12327 VDD.n6285 VDD.n6283 1.96392
R12328 VDD.n6282 VDD.n6280 1.96392
R12329 VDD.n6278 VDD.n6276 1.96392
R12330 VDD.n5432 VDD.n5430 1.95304
R12331 VDD.n5382 VDD.n5381 1.95304
R12332 VDD.n5332 VDD.n353 1.95304
R12333 VDD.n454 VDD.n452 1.95304
R12334 VDD.n510 VDD.n509 1.95304
R12335 VDD.n564 VDD.n406 1.95304
R12336 VDD.n610 VDD.n609 1.95304
R12337 VDD.n5201 VDD.n645 1.95304
R12338 VDD.n8404 VDD.n8403 1.94579
R12339 VDD.n7549 VDD.n7548 1.94579
R12340 VDD.n6695 VDD.n6694 1.94579
R12341 VDD.n5840 VDD.n5839 1.94579
R12342 VDD.n3975 VDD.n3618 1.93951
R12343 VDD.n4271 VDD.n2379 1.92692
R12344 VDD.n4223 VDD.n4222 1.92692
R12345 VDD.n4113 VDD.n4112 1.92692
R12346 VDD.n4168 VDD.n4044 1.92692
R12347 VDD.n2361 VDD.n2287 1.90031
R12348 VDD.n1469 VDD.n1467 1.8968
R12349 VDD.n1406 VDD.n1405 1.8968
R12350 VDD.n4558 VDD.n1025 1.8968
R12351 VDD.n2018 VDD.n2003 1.8968
R12352 VDD.n4423 VDD.n2119 1.8968
R12353 VDD.n8867 VDD.n8466 1.88841
R12354 VDD.n8012 VDD.n7611 1.88841
R12355 VDD.n7158 VDD.n6757 1.88841
R12356 VDD.n6303 VDD.n5902 1.88841
R12357 VDD.n1259 VDD.n1093 1.88682
R12358 VDD.n1220 VDD.n1123 1.88682
R12359 VDD.n1207 VDD.n1129 1.88682
R12360 VDD.n1168 VDD.n1158 1.88682
R12361 VDD.n4583 VDD.n4582 1.88682
R12362 VDD.n976 VDD.n971 1.88682
R12363 VDD.n4636 VDD.n969 1.88682
R12364 VDD.n4680 VDD.n940 1.88682
R12365 VDD.n4694 VDD.n4693 1.88682
R12366 VDD.n3599 VDD.n3598 1.88285
R12367 VDD.n3598 VDD.n2647 1.88285
R12368 VDD.n3564 VDD.n3563 1.88285
R12369 VDD.n3540 VDD.n3539 1.88285
R12370 VDD.n3266 VDD.n3265 1.88285
R12371 VDD.n3242 VDD.n3241 1.88285
R12372 VDD.n3155 VDD.n3154 1.88285
R12373 VDD.n3154 VDD.n3120 1.88285
R12374 VDD.n3802 VDD.n3799 1.88285
R12375 VDD.n3921 VDD.n3658 1.88285
R12376 VDD.n3683 VDD.n3682 1.88285
R12377 VDD.n3939 VDD.n3640 1.88285
R12378 VDD.n3939 VDD.n3641 1.88285
R12379 VDD.n2861 VDD.n2860 1.88285
R12380 VDD.n2886 VDD.n2876 1.88285
R12381 VDD.n3000 VDD.n2912 1.88285
R12382 VDD.n3000 VDD.n2913 1.88285
R12383 VDD.n93 VDD.n90 1.88285
R12384 VDD.n116 VDD.n114 1.88285
R12385 VDD.n5551 VDD.n5528 1.88285
R12386 VDD.n176 VDD.n175 1.88285
R12387 VDD.n1275 VDD.n1274 1.88285
R12388 VDD.n121 VDD.n120 1.87949
R12389 VDD.n4020 VDD.n2360 1.85282
R12390 VDD.n4257 VDD.n2388 1.8413
R12391 VDD.n4211 VDD.n2429 1.8413
R12392 VDD.n4126 VDD.n4063 1.8413
R12393 VDD.n4037 VDD.n4031 1.8413
R12394 VDD.n1467 VDD.n1466 1.82907
R12395 VDD.n3581 VDD.n2675 1.81303
R12396 VDD.n3283 VDD.n3081 1.81303
R12397 VDD.n5418 VDD.n5417 1.80841
R12398 VDD.n5369 VDD.n324 1.80841
R12399 VDD.n366 VDD.n362 1.80841
R12400 VDD.n469 VDD.n446 1.80841
R12401 VDD.n524 VDD.n523 1.80841
R12402 VDD.n580 VDD.n579 1.80841
R12403 VDD.n5238 VDD.n619 1.80841
R12404 VDD.n5190 VDD.n5189 1.80841
R12405 VDD.n8821 VDD.n8820 1.78137
R12406 VDD.n8359 VDD.n8264 1.78137
R12407 VDD.n7966 VDD.n7965 1.78137
R12408 VDD.n7504 VDD.n7409 1.78137
R12409 VDD.n7112 VDD.n7111 1.78137
R12410 VDD.n6650 VDD.n6555 1.78137
R12411 VDD.n6257 VDD.n6256 1.78137
R12412 VDD.n5795 VDD.n5700 1.78137
R12413 VDD.n4728 VDD.n916 1.76135
R12414 VDD.n4774 VDD.n4772 1.76135
R12415 VDD.n4787 VDD.n4786 1.76135
R12416 VDD.n4830 VDD.n4829 1.76135
R12417 VDD.n4842 VDD.n854 1.76135
R12418 VDD.n4888 VDD.n4886 1.76135
R12419 VDD.n4901 VDD.n4900 1.76135
R12420 VDD.n4944 VDD.n4943 1.76135
R12421 VDD.n4956 VDD.n792 1.76135
R12422 VDD.n5002 VDD.n5000 1.76135
R12423 VDD.n5015 VDD.n5014 1.76135
R12424 VDD.n5058 VDD.n5057 1.76135
R12425 VDD.n5070 VDD.n730 1.76135
R12426 VDD.n5116 VDD.n5114 1.76135
R12427 VDD.n5129 VDD.n5128 1.76135
R12428 VDD.n4268 VDD.n4267 1.75568
R12429 VDD.n2424 VDD.n2420 1.75568
R12430 VDD.n4118 VDD.n4070 1.75568
R12431 VDD.n4175 VDD.n4039 1.75568
R12432 VDD.n8581 VDD.n8580 1.74595
R12433 VDD.n7726 VDD.n7725 1.74595
R12434 VDD.n6872 VDD.n6871 1.74595
R12435 VDD.n6017 VDD.n6016 1.74595
R12436 VDD.n2136 VDD.t81 1.71984
R12437 VDD.n3974 VDD.n3972 1.71462
R12438 VDD.n8334 VDD.n8333 1.71235
R12439 VDD.n8332 VDD.n8306 1.71235
R12440 VDD.n8329 VDD.n8328 1.71235
R12441 VDD.n8324 VDD.n8309 1.71235
R12442 VDD.n8323 VDD.n8319 1.71235
R12443 VDD.n8318 VDD.n8317 1.71235
R12444 VDD.n7479 VDD.n7478 1.71235
R12445 VDD.n7477 VDD.n7451 1.71235
R12446 VDD.n7474 VDD.n7473 1.71235
R12447 VDD.n7469 VDD.n7454 1.71235
R12448 VDD.n7468 VDD.n7464 1.71235
R12449 VDD.n7463 VDD.n7462 1.71235
R12450 VDD.n6625 VDD.n6624 1.71235
R12451 VDD.n6623 VDD.n6597 1.71235
R12452 VDD.n6620 VDD.n6619 1.71235
R12453 VDD.n6615 VDD.n6600 1.71235
R12454 VDD.n6614 VDD.n6610 1.71235
R12455 VDD.n6609 VDD.n6608 1.71235
R12456 VDD.n5770 VDD.n5769 1.71235
R12457 VDD.n5768 VDD.n5742 1.71235
R12458 VDD.n5765 VDD.n5764 1.71235
R12459 VDD.n5760 VDD.n5745 1.71235
R12460 VDD.n5759 VDD.n5755 1.71235
R12461 VDD.n5754 VDD.n5753 1.71235
R12462 VDD.n1524 VDD.n1349 1.71139
R12463 VDD.n1534 VDD.n1343 1.71139
R12464 VDD.n1609 VDD.n1608 1.71139
R12465 VDD.n1287 VDD.n1280 1.71139
R12466 VDD.n1680 VDD.n1677 1.71139
R12467 VDD.n1749 VDD.n1748 1.71139
R12468 VDD.n3304 VDD.n3058 1.71033
R12469 VDD.n2791 VDD.n2778 1.70907
R12470 VDD.n2792 VDD.n2773 1.70593
R12471 VDD.n3310 VDD.n3309 1.70593
R12472 VDD.n3307 VDD.n3054 1.70592
R12473 VDD.n2788 VDD.n2776 1.70592
R12474 VDD.n3331 VDD.n2751 1.70592
R12475 VDD.n21 VDD.n20 1.70591
R12476 VDD.n3331 VDD.n3330 1.70591
R12477 VDD.n5600 VDD.n150 1.7059
R12478 VDD.n3310 VDD.n3048 1.70583
R12479 VDD.n3042 VDD.n2777 1.70583
R12480 VDD.n3045 VDD.n3044 1.70582
R12481 VDD.n3305 VDD.n3051 1.70582
R12482 VDD.n3316 VDD.n2768 1.7058
R12483 VDD.n3316 VDD.n2769 1.70579
R12484 VDD.n16 VDD.n14 1.70578
R12485 VDD.n5601 VDD.n5600 1.70577
R12486 VDD.n5674 VDD.n5612 1.7055
R12487 VDD.n6529 VDD.n6528 1.7055
R12488 VDD.n7383 VDD.n7321 1.7055
R12489 VDD.n8238 VDD.n8237 1.7055
R12490 VDD.n2867 VDD.n2787 1.7055
R12491 VDD.n2945 VDD.n2898 1.7055
R12492 VDD.n3008 VDD.n3007 1.7055
R12493 VDD.n3011 VDD.n3010 1.7055
R12494 VDD.n3016 VDD.n3015 1.7055
R12495 VDD.n3019 VDD.n3018 1.7055
R12496 VDD.n3030 VDD.n3029 1.7055
R12497 VDD.n3033 VDD.n3032 1.7055
R12498 VDD.n3036 VDD.n3035 1.7055
R12499 VDD.n3040 VDD.n2790 1.7055
R12500 VDD.n145 VDD.n3 1.7055
R12501 VDD.n144 VDD.n22 1.7055
R12502 VDD.n5560 VDD.n5540 1.7055
R12503 VDD.n159 VDD.n149 1.7055
R12504 VDD.n5525 VDD.n5524 1.7055
R12505 VDD.n5517 VDD.n5516 1.7055
R12506 VDD.n5514 VDD.n5513 1.7055
R12507 VDD.n5522 VDD.n5521 1.7055
R12508 VDD.n5598 VDD.n151 1.7055
R12509 VDD.n157 VDD.n156 1.7055
R12510 VDD.n152 VDD.n7 1.7055
R12511 VDD.n5519 VDD.n5518 1.7055
R12512 VDD.n154 VDD.n153 1.7055
R12513 VDD.n3052 VDD.n3049 1.7055
R12514 VDD.n3312 VDD.n3311 1.7055
R12515 VDD.n3315 VDD.n3314 1.7055
R12516 VDD.n3318 VDD.n3317 1.7055
R12517 VDD.n3321 VDD.n3320 1.7055
R12518 VDD.n3324 VDD.n3323 1.7055
R12519 VDD.n3326 VDD.n2763 1.7055
R12520 VDD.n2748 VDD.n2745 1.7055
R12521 VDD.n3333 VDD.n3332 1.7055
R12522 VDD.n3336 VDD.n3335 1.7055
R12523 VDD.n3341 VDD.n3340 1.7055
R12524 VDD.n3344 VDD.n3343 1.7055
R12525 VDD.n3347 VDD.n3346 1.7055
R12526 VDD.n3059 VDD.n3055 1.7055
R12527 VDD.n3319 VDD.n2753 1.7055
R12528 VDD.n3322 VDD.n2755 1.7055
R12529 VDD.n3378 VDD.n3377 1.7055
R12530 VDD.n3331 VDD.n3329 1.7055
R12531 VDD.n3334 VDD.n2757 1.7055
R12532 VDD.n3339 VDD.n2750 1.7055
R12533 VDD.n3342 VDD.n2758 1.7055
R12534 VDD.n3345 VDD.n2749 1.7055
R12535 VDD.n3375 VDD.n3374 1.7055
R12536 VDD.n2866 VDD.n2865 1.7055
R12537 VDD.n2908 VDD.n2783 1.7055
R12538 VDD.n3006 VDD.n2773 1.7055
R12539 VDD.n3009 VDD.n2782 1.7055
R12540 VDD.n3014 VDD.n2774 1.7055
R12541 VDD.n3017 VDD.n2781 1.7055
R12542 VDD.n3031 VDD.n2780 1.7055
R12543 VDD.n3034 VDD.n2776 1.7055
R12544 VDD.n3039 VDD.n2779 1.7055
R12545 VDD.n3042 VDD.n3041 1.7055
R12546 VDD.n3307 VDD.n3053 1.7055
R12547 VDD.n3310 VDD.n2771 1.7055
R12548 VDD.n3313 VDD.n2770 1.7055
R12549 VDD.n3060 VDD.n3056 1.7055
R12550 VDD.n143 VDD.n142 1.7055
R12551 VDD.n5603 VDD.n9 1.7055
R12552 VDD.n5512 VDD.n5511 1.7055
R12553 VDD.n5515 VDD.n21 1.7055
R12554 VDD.n5520 VDD.n13 1.7055
R12555 VDD.n5523 VDD.n19 1.7055
R12556 VDD.n158 VDD.n10 1.7055
R12557 VDD.n155 VDD.n148 1.7055
R12558 VDD.n147 VDD.n146 1.7055
R12559 VDD.n5539 VDD.n18 1.7055
R12560 VDD.n3316 VDD.n2756 1.70519
R12561 VDD.n142 VDD.n141 1.70511
R12562 VDD.n3973 VDD.n2632 1.70413
R12563 VDD.n3961 VDD.n3632 1.70404
R12564 VDD.n3962 VDD.n3627 1.70006
R12565 VDD.n3970 VDD.n3616 1.70006
R12566 VDD.n1452 VDD.n1451 1.69362
R12567 VDD.n1936 VDD.n1933 1.69362
R12568 VDD.n2039 VDD.n2031 1.69362
R12569 VDD.n2156 VDD.n2153 1.69362
R12570 VDD.t67 VDD.t54 1.68266
R12571 VDD.n8362 VDD.n8361 1.67007
R12572 VDD.n7507 VDD.n7506 1.67007
R12573 VDD.n6653 VDD.n6652 1.67007
R12574 VDD.n5798 VDD.n5797 1.67007
R12575 VDD.n2450 VDD.n2449 1.67007
R12576 VDD.n4261 VDD.n4260 1.67007
R12577 VDD.n4212 VDD.n2426 1.67007
R12578 VDD.n4127 VDD.n4125 1.67007
R12579 VDD.n4182 VDD.n4181 1.67007
R12580 VDD.n5433 VDD.n298 1.66378
R12581 VDD.n5385 VDD.n319 1.66378
R12582 VDD.n5333 VDD.n350 1.66378
R12583 VDD.n5288 VDD.n392 1.66378
R12584 VDD.n505 VDD.n430 1.66378
R12585 VDD.n563 VDD.n408 1.66378
R12586 VDD.n5255 VDD.n605 1.66378
R12587 VDD.n5205 VDD.n5204 1.66378
R12588 VDD.n8771 VDD.n8769 1.66186
R12589 VDD.n8772 VDD.n8755 1.66186
R12590 VDD.n8777 VDD.n8775 1.66186
R12591 VDD.n8778 VDD.n8753 1.66186
R12592 VDD.n8783 VDD.n8781 1.66186
R12593 VDD.n8787 VDD.n8786 1.66186
R12594 VDD.n7916 VDD.n7914 1.66186
R12595 VDD.n7917 VDD.n7900 1.66186
R12596 VDD.n7922 VDD.n7920 1.66186
R12597 VDD.n7923 VDD.n7898 1.66186
R12598 VDD.n7928 VDD.n7926 1.66186
R12599 VDD.n7932 VDD.n7931 1.66186
R12600 VDD.n7062 VDD.n7060 1.66186
R12601 VDD.n7063 VDD.n7046 1.66186
R12602 VDD.n7068 VDD.n7066 1.66186
R12603 VDD.n7069 VDD.n7044 1.66186
R12604 VDD.n7074 VDD.n7072 1.66186
R12605 VDD.n7078 VDD.n7077 1.66186
R12606 VDD.n6207 VDD.n6205 1.66186
R12607 VDD.n6208 VDD.n6191 1.66186
R12608 VDD.n6213 VDD.n6211 1.66186
R12609 VDD.n6214 VDD.n6189 1.66186
R12610 VDD.n6219 VDD.n6217 1.66186
R12611 VDD.n6223 VDD.n6222 1.66186
R12612 VDD.n3926 VDD.n3665 1.64452
R12613 VDD.n3910 VDD.n3671 1.64452
R12614 VDD.n3810 VDD.n3809 1.64447
R12615 VDD.n2857 VDD.n2809 1.64446
R12616 VDD.n3024 VDD.n3023 1.64446
R12617 VDD.n1819 VDD.n1085 1.63187
R12618 VDD.n1463 VDD.n1404 1.6259
R12619 VDD.n4562 VDD.n4561 1.6259
R12620 VDD.n4495 VDD.n2002 1.6259
R12621 VDD.n4427 VDD.n4426 1.6259
R12622 VDD.n4360 VDD.n2223 1.6259
R12623 VDD.n2357 VDD.n2356 1.62066
R12624 VDD.n1258 VDD.n1098 1.61734
R12625 VDD.n1221 VDD.n1121 1.61734
R12626 VDD.n1206 VDD.n1133 1.61734
R12627 VDD.n1169 VDD.n1156 1.61734
R12628 VDD.n4588 VDD.n996 1.61734
R12629 VDD.n4624 VDD.n4623 1.61734
R12630 VDD.n4643 VDD.n964 1.61734
R12631 VDD.n4681 VDD.n4679 1.61734
R12632 VDD.n4699 VDD.n933 1.61734
R12633 VDD.n4353 VDD.n4352 1.61534
R12634 VDD.n4352 VDD.n4351 1.61534
R12635 VDD.n4351 VDD.n4349 1.61534
R12636 VDD.n4349 VDD.n4347 1.61534
R12637 VDD.n4347 VDD.n4345 1.61534
R12638 VDD.n4345 VDD.n4343 1.61534
R12639 VDD.n4343 VDD.n4341 1.61534
R12640 VDD.n4341 VDD.n4339 1.61534
R12641 VDD.n4339 VDD.n4337 1.61534
R12642 VDD.n4337 VDD.n4335 1.61534
R12643 VDD.n4335 VDD.n4333 1.61534
R12644 VDD.n4333 VDD.n4331 1.61534
R12645 VDD.n4328 VDD.n4326 1.61534
R12646 VDD.n4326 VDD.n4324 1.61534
R12647 VDD.n4324 VDD.n4322 1.61534
R12648 VDD.n4322 VDD.n4320 1.61534
R12649 VDD.n4320 VDD.n4318 1.61534
R12650 VDD.n4318 VDD.n4316 1.61534
R12651 VDD.n4316 VDD.n4314 1.61534
R12652 VDD.n4314 VDD.n4312 1.61534
R12653 VDD.n4312 VDD.n4310 1.61534
R12654 VDD.n4310 VDD.n4308 1.61534
R12655 VDD.n4308 VDD.n4306 1.61534
R12656 VDD.n4306 VDD.n4304 1.61534
R12657 VDD.n8718 VDD.n8716 1.61441
R12658 VDD.n7863 VDD.n7861 1.61441
R12659 VDD.n7009 VDD.n7007 1.61441
R12660 VDD.n6154 VDD.n6152 1.61441
R12661 VDD.t77 VDD.n2215 1.58758
R12662 VDD.n2386 VDD.n2382 1.58445
R12663 VDD.n4216 VDD.n2425 1.58445
R12664 VDD.n4200 VDD.n2438 1.58445
R12665 VDD.n4117 VDD.n4071 1.58445
R12666 VDD.n4177 VDD.n4176 1.58445
R12667 VDD.n1815 VDD.n1814 1.58383
R12668 VDD.n2453 VDD.n2450 1.57731
R12669 VDD.n4724 VDD.n4722 1.55817
R12670 VDD.n4294 VDD.n4293 1.5505
R12671 VDD.n5414 VDD.n305 1.51914
R12672 VDD.n5366 VDD.n5365 1.51914
R12673 VDD.n5315 VDD.n367 1.51914
R12674 VDD.n470 VDD.n444 1.51914
R12675 VDD.n528 VDD.n422 1.51914
R12676 VDD.n5282 VDD.n399 1.51914
R12677 VDD.n5237 VDD.n620 1.51914
R12678 VDD.n661 VDD.n657 1.51914
R12679 VDD.n102 VDD.n101 1.51334
R12680 VDD.n136 VDD.n135 1.51334
R12681 VDD.n5560 VDD.n5559 1.51334
R12682 VDD.n201 VDD.n200 1.51334
R12683 VDD.n83 VDD.n79 1.50638
R12684 VDD.n122 VDD.n117 1.50638
R12685 VDD.n5590 VDD.n5533 1.50638
R12686 VDD.n231 VDD.n225 1.50638
R12687 VDD.n2585 VDD.n2584 1.50638
R12688 VDD.n2558 VDD.n2557 1.50638
R12689 VDD.n2556 VDD.n2537 1.50638
R12690 VDD.n4293 VDD.n4292 1.5044
R12691 VDD.n132 VDD.n123 1.50148
R12692 VDD.n5486 VDD.n5485 1.5005
R12693 VDD.n5477 VDD.n5476 1.5005
R12694 VDD.n5493 VDD.n5491 1.5005
R12695 VDD.n2564 VDD.n2563 1.5005
R12696 VDD.n2554 VDD.n2535 1.5005
R12697 VDD.n2550 VDD.n2549 1.5005
R12698 VDD.n2569 VDD.n2532 1.5005
R12699 VDD.n2574 VDD.n2573 1.5005
R12700 VDD.n2531 VDD.n2530 1.5005
R12701 VDD.n2580 VDD.n2514 1.5005
R12702 VDD.n2513 VDD.n2510 1.5005
R12703 VDD.n2387 VDD.n2386 1.49883
R12704 VDD.n4216 VDD.n4215 1.49883
R12705 VDD.n4071 VDD.n4066 1.49883
R12706 VDD.n4176 VDD.n4036 1.49883
R12707 VDD.n102 VDD.n34 1.49119
R12708 VDD.n136 VDD.n107 1.49076
R12709 VDD.n201 VDD.n174 1.49076
R12710 VDD.n3770 VDD.n3636 1.49076
R12711 VDD.n3806 VDD.n3649 1.49076
R12712 VDD.n3920 VDD.n3919 1.49076
R12713 VDD.n2798 VDD.n2794 1.49076
R12714 VDD.n4735 VDD.n911 1.49045
R12715 VDD.n895 VDD.n890 1.49045
R12716 VDD.n4792 VDD.n880 1.49045
R12717 VDD.n4824 VDD.n860 1.49045
R12718 VDD.n4849 VDD.n849 1.49045
R12719 VDD.n833 VDD.n828 1.49045
R12720 VDD.n4906 VDD.n818 1.49045
R12721 VDD.n4938 VDD.n798 1.49045
R12722 VDD.n4963 VDD.n787 1.49045
R12723 VDD.n771 VDD.n766 1.49045
R12724 VDD.n5020 VDD.n756 1.49045
R12725 VDD.n5052 VDD.n736 1.49045
R12726 VDD.n5077 VDD.n725 1.49045
R12727 VDD.n709 VDD.n704 1.49045
R12728 VDD.n5134 VDD.n694 1.49045
R12729 VDD.n3919 VDD.n3918 1.4899
R12730 VDD.n3771 VDD.n3770 1.4899
R12731 VDD.n2808 VDD.n2794 1.4899
R12732 VDD.n3808 VDD.n3798 1.4871
R12733 VDD.n3664 VDD.n3663 1.4871
R12734 VDD.n3690 VDD.n3670 1.4871
R12735 VDD.n2807 VDD.n2805 1.4871
R12736 VDD.n2889 VDD.n2884 1.4871
R12737 VDD.n3102 VDD.n3094 1.48392
R12738 VDD.n3179 VDD.n3089 1.48392
R12739 VDD.n3411 VDD.n3410 1.48392
R12740 VDD.n2728 VDD.n2713 1.48392
R12741 VDD.n2697 VDD.n2693 1.48392
R12742 VDD.n3477 VDD.n2683 1.48392
R12743 VDD.n3604 VDD.n2637 1.48392
R12744 VDD.n3450 VDD.n3449 1.48392
R12745 VDD.n3396 VDD.n3395 1.48392
R12746 VDD.n3111 VDD.n3107 1.48264
R12747 VDD.n3362 VDD.n3361 1.47597
R12748 VDD.n3290 VDD.n3289 1.47597
R12749 VDD.n3456 VDD.n3455 1.46766
R12750 VDD.n3444 VDD.n2706 1.46766
R12751 VDD.n3390 VDD.n2742 1.46766
R12752 VDD.n2721 VDD.n2717 1.46766
R12753 VDD.n3417 VDD.n3402 1.46766
R12754 VDD.n9000 VDD.n8272 1.45846
R12755 VDD.n8369 VDD.n8304 1.45846
R12756 VDD.n8364 VDD.n8304 1.45846
R12757 VDD.n8145 VDD.n7417 1.45846
R12758 VDD.n7514 VDD.n7449 1.45846
R12759 VDD.n7509 VDD.n7449 1.45846
R12760 VDD.n7291 VDD.n6563 1.45846
R12761 VDD.n6660 VDD.n6595 1.45846
R12762 VDD.n6655 VDD.n6595 1.45846
R12763 VDD.n6436 VDD.n5708 1.45846
R12764 VDD.n5805 VDD.n5740 1.45846
R12765 VDD.n5800 VDD.n5740 1.45846
R12766 VDD.n1521 VDD.n1351 1.45793
R12767 VDD.n1537 VDD.n1340 1.45793
R12768 VDD.n1601 VDD.n1294 1.45793
R12769 VDD.n1811 VDD.n1281 1.45793
R12770 VDD.n1675 VDD.n1668 1.45793
R12771 VDD.n1693 VDD.n1692 1.45793
R12772 VDD.n4017 VDD.n4016 1.45532
R12773 VDD.n1445 VDD.n1444 1.42272
R12774 VDD.n1934 VDD.n1926 1.42272
R12775 VDD.n4479 VDD.n2032 1.42272
R12776 VDD.n2154 VDD.n2146 1.42272
R12777 VDD.n4261 VDD.n2387 1.41321
R12778 VDD.n4215 VDD.n2426 1.41321
R12779 VDD.n4125 VDD.n4066 1.41321
R12780 VDD.n4182 VDD.n4036 1.41321
R12781 VDD.n4195 VDD.n4194 1.41321
R12782 VDD.n5496 VDD.n249 1.3918
R12783 VDD.n1853 VDD.n1062 1.38089
R12784 VDD.n1820 VDD.n1083 1.38089
R12785 VDD.n5437 VDD.n5436 1.37451
R12786 VDD.n5389 VDD.n5386 1.37451
R12787 VDD.n5337 VDD.n5336 1.37451
R12788 VDD.n5289 VDD.n389 1.37451
R12789 VDD.n504 VDD.n432 1.37451
R12790 VDD.n560 VDD.n559 1.37451
R12791 VDD.n5256 VDD.n602 1.37451
R12792 VDD.n644 VDD.n643 1.37451
R12793 VDD.n1904 VDD.n1903 1.355
R12794 VDD.n4499 VDD.n4498 1.355
R12795 VDD.n2124 VDD.n2123 1.355
R12796 VDD.n4364 VDD.n4363 1.355
R12797 VDD.n8398 VDD.n8289 1.35125
R12798 VDD.n7543 VDD.n7434 1.35125
R12799 VDD.n6689 VDD.n6580 1.35125
R12800 VDD.n5834 VDD.n5725 1.35125
R12801 VDD.n1255 VDD.n1254 1.34787
R12802 VDD.n1225 VDD.n1224 1.34787
R12803 VDD.n1203 VDD.n1202 1.34787
R12804 VDD.n1173 VDD.n1172 1.34787
R12805 VDD.n4587 VDD.n997 1.34787
R12806 VDD.n4618 VDD.n975 1.34787
R12807 VDD.n4645 VDD.n4644 1.34787
R12808 VDD.n948 VDD.n943 1.34787
R12809 VDD.n4698 VDD.n934 1.34787
R12810 VDD.n2947 VDD.n2897 1.3466
R12811 VDD.n3022 VDD.n3021 1.3449
R12812 VDD.n3356 VDD.n2765 1.34458
R12813 VDD.n3368 VDD.n2765 1.34227
R12814 VDD.n9020 VDD.n9019 1.33615
R12815 VDD.n8165 VDD.n8164 1.33615
R12816 VDD.n7311 VDD.n7310 1.33615
R12817 VDD.n6456 VDD.n6455 1.33615
R12818 VDD.n4267 VDD.n2382 1.32759
R12819 VDD.n2425 VDD.n2424 1.32759
R12820 VDD.n4118 VDD.n4117 1.32759
R12821 VDD.n4177 VDD.n4175 1.32759
R12822 VDD.n8860 VDD.n8859 1.32203
R12823 VDD.n8763 VDD.n8757 1.32203
R12824 VDD.n8005 VDD.n8004 1.32203
R12825 VDD.n7908 VDD.n7902 1.32203
R12826 VDD.n7151 VDD.n7150 1.32203
R12827 VDD.n7054 VDD.n7048 1.32203
R12828 VDD.n6296 VDD.n6295 1.32203
R12829 VDD.n6199 VDD.n6193 1.32203
R12830 VDD.n4353 VDD.n2287 1.28287
R12831 VDD.n2545 VDD.n2516 1.26837
R12832 VDD.n8644 VDD.n8643 1.25267
R12833 VDD.n7789 VDD.n7788 1.25267
R12834 VDD.n6935 VDD.n6934 1.25267
R12835 VDD.n6080 VDD.n6079 1.25267
R12836 VDD.n8861 VDD.n8860 1.24652
R12837 VDD.n8760 VDD.n8757 1.24652
R12838 VDD.n8006 VDD.n8005 1.24652
R12839 VDD.n7905 VDD.n7902 1.24652
R12840 VDD.n7152 VDD.n7151 1.24652
R12841 VDD.n7051 VDD.n7048 1.24652
R12842 VDD.n6297 VDD.n6296 1.24652
R12843 VDD.n6196 VDD.n6193 1.24652
R12844 VDD.n4260 VDD.n2388 1.24197
R12845 VDD.n4212 VDD.n4211 1.24197
R12846 VDD.n4127 VDD.n4126 1.24197
R12847 VDD.n4181 VDD.n4037 1.24197
R12848 VDD.n5413 VDD.n306 1.22988
R12849 VDD.n332 VDD.n327 1.22988
R12850 VDD.n5314 VDD.n368 1.22988
R12851 VDD.n474 VDD.n473 1.22988
R12852 VDD.n529 VDD.n420 1.22988
R12853 VDD.n5281 VDD.n400 1.22988
R12854 VDD.n5234 VDD.n5233 1.22988
R12855 VDD.n5183 VDD.n662 1.22988
R12856 VDD.n8717 VDD.n8247 1.22485
R12857 VDD.n9020 VDD.n8247 1.22485
R12858 VDD.n9019 VDD.n8248 1.22485
R12859 VDD.n8263 VDD.n8262 1.22485
R12860 VDD.n9009 VDD.n9008 1.22485
R12861 VDD.n7862 VDD.n7392 1.22485
R12862 VDD.n8165 VDD.n7392 1.22485
R12863 VDD.n8164 VDD.n7393 1.22485
R12864 VDD.n7408 VDD.n7407 1.22485
R12865 VDD.n8154 VDD.n8153 1.22485
R12866 VDD.n7008 VDD.n6538 1.22485
R12867 VDD.n7311 VDD.n6538 1.22485
R12868 VDD.n7310 VDD.n6539 1.22485
R12869 VDD.n6554 VDD.n6553 1.22485
R12870 VDD.n7300 VDD.n7299 1.22485
R12871 VDD.n6153 VDD.n5683 1.22485
R12872 VDD.n6456 VDD.n5683 1.22485
R12873 VDD.n6455 VDD.n5684 1.22485
R12874 VDD.n5699 VDD.n5698 1.22485
R12875 VDD.n6445 VDD.n6444 1.22485
R12876 VDD.n4737 VDD.n4736 1.21955
R12877 VDD.n4766 VDD.n4765 1.21955
R12878 VDD.n4791 VDD.n881 1.21955
R12879 VDD.n4825 VDD.n4823 1.21955
R12880 VDD.n4851 VDD.n4850 1.21955
R12881 VDD.n4880 VDD.n4879 1.21955
R12882 VDD.n4905 VDD.n819 1.21955
R12883 VDD.n4939 VDD.n4937 1.21955
R12884 VDD.n4965 VDD.n4964 1.21955
R12885 VDD.n4994 VDD.n4993 1.21955
R12886 VDD.n5019 VDD.n757 1.21955
R12887 VDD.n5053 VDD.n5051 1.21955
R12888 VDD.n5079 VDD.n5078 1.21955
R12889 VDD.n5108 VDD.n5107 1.21955
R12890 VDD.n5133 VDD.n695 1.21955
R12891 VDD.n1357 VDD.n1356 1.20446
R12892 VDD.n1338 VDD.n1334 1.20446
R12893 VDD.n1599 VDD.n1298 1.20446
R12894 VDD.n1808 VDD.n1807 1.20446
R12895 VDD.n1764 VDD.n1667 1.20446
R12896 VDD.n1739 VDD.n1697 1.20446
R12897 VDD.n6495 VDD.n6466 1.20001
R12898 VDD.n8204 VDD.n8175 1.20001
R12899 VDD.n5673 VDD.n5672 1.1947
R12900 VDD.n7382 VDD.n7381 1.1947
R12901 VDD.n4268 VDD.n2379 1.15635
R12902 VDD.n4222 VDD.n2420 1.15635
R12903 VDD.n4112 VDD.n4070 1.15635
R12904 VDD.n4044 VDD.n4039 1.15635
R12905 VDD.n4300 VDD.n2357 1.15386
R12906 VDD.n1441 VDD.n1411 1.15182
R12907 VDD.n4542 VDD.n1927 1.15182
R12908 VDD.n4476 VDD.n4475 1.15182
R12909 VDD.n4407 VDD.n2147 1.15182
R12910 VDD.n3038 VDD.n3037 1.13717
R12911 VDD.n3021 VDD.n3020 1.13717
R12912 VDD.n3013 VDD.n3012 1.13717
R12913 VDD.n2947 VDD.n2946 1.13717
R12914 VDD.n2944 VDD.n2909 1.13717
R12915 VDD.n3304 VDD.n3303 1.13717
R12916 VDD.n3338 VDD.n3337 1.13717
R12917 VDD.n2765 VDD.n2759 1.13717
R12918 VDD.n5468 VDD.n261 1.13602
R12919 VDD.n3589 VDD.n2659 1.12991
R12920 VDD.n3589 VDD.n3588 1.12991
R12921 VDD.n3559 VDD.n3558 1.12991
R12922 VDD.n3545 VDD.n3544 1.12991
R12923 VDD.n3261 VDD.n3260 1.12991
R12924 VDD.n3247 VDD.n3246 1.12991
R12925 VDD.n3145 VDD.n3128 1.12991
R12926 VDD.n3145 VDD.n3144 1.12991
R12927 VDD.n3784 VDD.n3783 1.12991
R12928 VDD.n2937 VDD.n2936 1.12991
R12929 VDD.n74 VDD.n55 1.12991
R12930 VDD.n74 VDD.n56 1.12991
R12931 VDD.n5584 VDD.n5583 1.12991
R12932 VDD.n5583 VDD.n5564 1.12991
R12933 VDD.n220 VDD.n183 1.12991
R12934 VDD.n220 VDD.n184 1.12991
R12935 VDD.n1852 VDD.n1064 1.12991
R12936 VDD.n1824 VDD.n1823 1.12991
R12937 VDD.n2583 VDD.n2511 1.12991
R12938 VDD.n2528 VDD.n2520 1.12991
R12939 VDD.n8385 VDD.n8272 1.11541
R12940 VDD.n8384 VDD.n8297 1.11541
R12941 VDD.n8380 VDD.n8379 1.11541
R12942 VDD.n8377 VDD.n8376 1.11541
R12943 VDD.n8374 VDD.n8301 1.11541
R12944 VDD.n8371 VDD.n8370 1.11541
R12945 VDD.n7530 VDD.n7417 1.11541
R12946 VDD.n7529 VDD.n7442 1.11541
R12947 VDD.n7525 VDD.n7524 1.11541
R12948 VDD.n7522 VDD.n7521 1.11541
R12949 VDD.n7519 VDD.n7446 1.11541
R12950 VDD.n7516 VDD.n7515 1.11541
R12951 VDD.n6676 VDD.n6563 1.11541
R12952 VDD.n6675 VDD.n6588 1.11541
R12953 VDD.n6671 VDD.n6670 1.11541
R12954 VDD.n6668 VDD.n6667 1.11541
R12955 VDD.n6665 VDD.n6592 1.11541
R12956 VDD.n6662 VDD.n6661 1.11541
R12957 VDD.n5821 VDD.n5708 1.11541
R12958 VDD.n5820 VDD.n5733 1.11541
R12959 VDD.n5816 VDD.n5815 1.11541
R12960 VDD.n5813 VDD.n5812 1.11541
R12961 VDD.n5810 VDD.n5737 1.11541
R12962 VDD.n5807 VDD.n5806 1.11541
R12963 VDD.n241 VDD.n239 1.11031
R12964 VDD.n3700 VDD.n3699 1.10923
R12965 VDD.n136 VDD.n27 1.10918
R12966 VDD.n201 VDD.n169 1.10899
R12967 VDD.n102 VDD.n39 1.10899
R12968 VDD.n5657 VDD 1.09833
R12969 VDD.n7366 VDD 1.09833
R12970 VDD.n4298 VDD.n0 1.09663
R12971 VDD.n297 VDD.n296 1.08525
R12972 VDD.n5390 VDD.n317 1.08525
R12973 VDD.n349 VDD.n348 1.08525
R12974 VDD.n5293 VDD.n5292 1.08525
R12975 VDD.n501 VDD.n500 1.08525
R12976 VDD.n555 VDD.n410 1.08525
R12977 VDD.n5260 VDD.n5259 1.08525
R12978 VDD.n5211 VDD.n639 1.08525
R12979 VDD.n1902 VDD.n1010 1.0841
R12980 VDD.n2007 VDD.n2006 1.0841
R12981 VDD.n2122 VDD.n2105 1.0841
R12982 VDD.n2228 VDD.n2227 1.0841
R12983 VDD.n1250 VDD.n1100 1.07839
R12984 VDD.n1229 VDD.n1117 1.07839
R12985 VDD.n1198 VDD.n1135 1.07839
R12986 VDD.n1177 VDD.n1152 1.07839
R12987 VDD.n4594 VDD.n992 1.07839
R12988 VDD.n4619 VDD.n4617 1.07839
R12989 VDD.n4650 VDD.n961 1.07839
R12990 VDD.n4673 VDD.n4672 1.07839
R12991 VDD.n4705 VDD.n929 1.07839
R12992 VDD.n4290 VDD.n2361 1.07073
R12993 VDD.n4257 VDD.n4256 1.07073
R12994 VDD.n2433 VDD.n2429 1.07073
R12995 VDD.n4132 VDD.n4063 1.07073
R12996 VDD.n4189 VDD.n4031 1.07073
R12997 VDD.n4300 VDD.n4299 1.04401
R12998 VDD.n4301 VDD.n2341 1.04351
R12999 VDD.n5470 VDD.n5468 1.04225
R13000 VDD.n2947 VDD.n2943 1.02922
R13001 VDD.n5560 VDD.n5527 1.0272
R13002 VDD.n3021 VDD.n2872 1.02676
R13003 VDD.n5560 VDD.n5538 1.02649
R13004 VDD.n4304 VDD.n4302 1.02165
R13005 VDD.n4293 VDD.n2361 0.997903
R13006 VDD.n3495 VDD.n3491 0.994314
R13007 VDD.n3514 VDD.n3513 0.994314
R13008 VDD.n3197 VDD.n3193 0.994314
R13009 VDD.n3216 VDD.n3215 0.994314
R13010 VDD.n3745 VDD.n3741 0.994314
R13011 VDD.n3838 VDD.n3738 0.994314
R13012 VDD.n3842 VDD.n3734 0.994314
R13013 VDD.n3884 VDD.n3883 0.994314
R13014 VDD.n3861 VDD.n3711 0.994314
R13015 VDD.n3864 VDD.n3706 0.994314
R13016 VDD.n2825 VDD.n2821 0.994314
R13017 VDD.n2967 VDD.n2963 0.994314
R13018 VDD.n4272 VDD.n4271 0.985115
R13019 VDD.n4223 VDD.n2417 0.985115
R13020 VDD.n4113 VDD.n4111 0.985115
R13021 VDD.n4169 VDD.n4168 0.985115
R13022 VDD.n1509 VDD.n1360 0.950995
R13023 VDD.n1550 VDD.n1549 0.950995
R13024 VDD.n1596 VDD.n1300 0.950995
R13025 VDD.n1626 VDD.n1625 0.950995
R13026 VDD.n1768 VDD.n1767 0.950995
R13027 VDD.n1737 VDD.n1698 0.950995
R13028 VDD.n4742 VDD.n908 0.948648
R13029 VDD.n4760 VDD.n894 0.948648
R13030 VDD.n4798 VDD.n876 0.948648
R13031 VDD.n868 VDD.n863 0.948648
R13032 VDD.n4856 VDD.n846 0.948648
R13033 VDD.n4874 VDD.n832 0.948648
R13034 VDD.n4912 VDD.n814 0.948648
R13035 VDD.n806 VDD.n801 0.948648
R13036 VDD.n4970 VDD.n784 0.948648
R13037 VDD.n4988 VDD.n770 0.948648
R13038 VDD.n5026 VDD.n752 0.948648
R13039 VDD.n744 VDD.n739 0.948648
R13040 VDD.n5084 VDD.n722 0.948648
R13041 VDD.n5102 VDD.n708 0.948648
R13042 VDD.n5140 VDD.n690 0.948648
R13043 VDD.n4085 VDD.n2438 0.942306
R13044 VDD.n4195 VDD.n273 0.942306
R13045 VDD.n5410 VDD.n5409 0.940613
R13046 VDD.n5359 VDD.n333 0.940613
R13047 VDD.n5311 VDD.n5310 0.940613
R13048 VDD.n478 VDD.n442 0.940613
R13049 VDD.n533 VDD.n532 0.940613
R13050 VDD.n5278 VDD.n5277 0.940613
R13051 VDD.n627 VDD.n623 0.940613
R13052 VDD.n5182 VDD.n663 0.940613
R13053 VDD.n8335 VDD.n8334 0.934239
R13054 VDD.n8333 VDD.n8332 0.934239
R13055 VDD.n8329 VDD.n8306 0.934239
R13056 VDD.n8328 VDD.n8309 0.934239
R13057 VDD.n8324 VDD.n8323 0.934239
R13058 VDD.n8319 VDD.n8318 0.934239
R13059 VDD.n7480 VDD.n7479 0.934239
R13060 VDD.n7478 VDD.n7477 0.934239
R13061 VDD.n7474 VDD.n7451 0.934239
R13062 VDD.n7473 VDD.n7454 0.934239
R13063 VDD.n7469 VDD.n7468 0.934239
R13064 VDD.n7464 VDD.n7463 0.934239
R13065 VDD.n6626 VDD.n6625 0.934239
R13066 VDD.n6624 VDD.n6623 0.934239
R13067 VDD.n6620 VDD.n6597 0.934239
R13068 VDD.n6619 VDD.n6600 0.934239
R13069 VDD.n6615 VDD.n6614 0.934239
R13070 VDD.n6610 VDD.n6609 0.934239
R13071 VDD.n5771 VDD.n5770 0.934239
R13072 VDD.n5769 VDD.n5768 0.934239
R13073 VDD.n5765 VDD.n5742 0.934239
R13074 VDD.n5764 VDD.n5745 0.934239
R13075 VDD.n5760 VDD.n5759 0.934239
R13076 VDD.n5755 VDD.n5754 0.934239
R13077 VDD.n1816 VDD.n1815 0.926297
R13078 VDD.n1892 VDD.n1030 0.926297
R13079 VDD.n1031 VDD.n1001 0.926297
R13080 VDD.n4576 VDD.n1002 0.926297
R13081 VDD.n4570 VDD.n1011 0.926297
R13082 VDD.n2602 VDD.n1012 0.926297
R13083 VDD.n4564 VDD.n1018 0.926297
R13084 VDD.n2599 VDD.n1910 0.926297
R13085 VDD.n4555 VDD.n4554 0.926297
R13086 VDD.n4551 VDD.n1911 0.926297
R13087 VDD.n1922 VDD.n1917 0.926297
R13088 VDD.n4545 VDD.n1923 0.926297
R13089 VDD.n1941 VDD.n1924 0.926297
R13090 VDD.n4536 VDD.n4535 0.926297
R13091 VDD.n4532 VDD.n1942 0.926297
R13092 VDD.n2607 VDD.n1948 0.926297
R13093 VDD.n4526 VDD.n1953 0.926297
R13094 VDD.n1962 VDD.n1954 0.926297
R13095 VDD.n4520 VDD.n4519 0.926297
R13096 VDD.n4511 VDD.n4510 0.926297
R13097 VDD.n4507 VDD.n1980 0.926297
R13098 VDD.n1994 VDD.n1986 0.926297
R13099 VDD.n4501 VDD.n1995 0.926297
R13100 VDD.n2013 VDD.n1996 0.926297
R13101 VDD.n4492 VDD.n4491 0.926297
R13102 VDD.n4488 VDD.n2021 0.926297
R13103 VDD.n2027 VDD.n2022 0.926297
R13104 VDD.n4482 VDD.n2028 0.926297
R13105 VDD.n2046 VDD.n2029 0.926297
R13106 VDD.n4473 VDD.n4472 0.926297
R13107 VDD.n4469 VDD.n2047 0.926297
R13108 VDD.n2090 VDD.n2089 0.926297
R13109 VDD.n4463 VDD.n2057 0.926297
R13110 VDD.n2068 VDD.n2058 0.926297
R13111 VDD.n4454 VDD.n2069 0.926297
R13112 VDD.n2074 VDD.n2070 0.926297
R13113 VDD.n4448 VDD.n2075 0.926297
R13114 VDD.n4439 VDD.n4438 0.926297
R13115 VDD.n4435 VDD.n2100 0.926297
R13116 VDD.n2111 VDD.n2106 0.926297
R13117 VDD.n4429 VDD.n2112 0.926297
R13118 VDD.n2130 VDD.n2113 0.926297
R13119 VDD.n4420 VDD.n4419 0.926297
R13120 VDD.n4416 VDD.n2136 0.926297
R13121 VDD.n2142 VDD.n2137 0.926297
R13122 VDD.n4410 VDD.n2143 0.926297
R13123 VDD.n2161 VDD.n2144 0.926297
R13124 VDD.n4401 VDD.n4400 0.926297
R13125 VDD.n4397 VDD.n2162 0.926297
R13126 VDD.n2173 VDD.n2168 0.926297
R13127 VDD.n4391 VDD.n2174 0.926297
R13128 VDD.n2183 VDD.n2175 0.926297
R13129 VDD.n4385 VDD.n4384 0.926297
R13130 VDD.n2200 VDD.n2184 0.926297
R13131 VDD.n4376 VDD.n4375 0.926297
R13132 VDD.n4372 VDD.n2201 0.926297
R13133 VDD.n2215 VDD.n2207 0.926297
R13134 VDD.n4366 VDD.n2216 0.926297
R13135 VDD.n2234 VDD.n2217 0.926297
R13136 VDD.n8769 VDD.n8767 0.906695
R13137 VDD.n8772 VDD.n8771 0.906695
R13138 VDD.n8775 VDD.n8755 0.906695
R13139 VDD.n8778 VDD.n8777 0.906695
R13140 VDD.n8781 VDD.n8753 0.906695
R13141 VDD.n8787 VDD.n8783 0.906695
R13142 VDD.n7914 VDD.n7912 0.906695
R13143 VDD.n7917 VDD.n7916 0.906695
R13144 VDD.n7920 VDD.n7900 0.906695
R13145 VDD.n7923 VDD.n7922 0.906695
R13146 VDD.n7926 VDD.n7898 0.906695
R13147 VDD.n7932 VDD.n7928 0.906695
R13148 VDD.n7060 VDD.n7058 0.906695
R13149 VDD.n7063 VDD.n7062 0.906695
R13150 VDD.n7066 VDD.n7046 0.906695
R13151 VDD.n7069 VDD.n7068 0.906695
R13152 VDD.n7072 VDD.n7044 0.906695
R13153 VDD.n7078 VDD.n7074 0.906695
R13154 VDD.n6205 VDD.n6203 0.906695
R13155 VDD.n6208 VDD.n6207 0.906695
R13156 VDD.n6211 VDD.n6191 0.906695
R13157 VDD.n6214 VDD.n6213 0.906695
R13158 VDD.n6217 VDD.n6189 0.906695
R13159 VDD.n6223 VDD.n6219 0.906695
R13160 VDD.n3701 VDD.n3700 0.903353
R13161 VDD.n3770 VDD.n3643 0.903353
R13162 VDD.n4329 VDD.n4328 0.902912
R13163 VDD.n1865 VDD.n1057 0.899959
R13164 VDD.n2395 VDD.n2391 0.899497
R13165 VDD.n4205 VDD.n2434 0.899497
R13166 VDD.n4131 VDD.n4064 0.899497
R13167 VDD.n4190 VDD.n4029 0.899497
R13168 VDD.n2903 VDD.n2901 0.884222
R13169 VDD.n2903 VDD.n2902 0.883499
R13170 VDD.n1437 VDD.n1412 0.880923
R13171 VDD.n4539 VDD.n4538 0.880923
R13172 VDD.n2051 VDD.n2050 0.880923
R13173 VDD.n4404 VDD.n4403 0.880923
R13174 VDD.n5159 VDD.n5158 0.880923
R13175 VDD.n1849 VDD.n1848 0.878931
R13176 VDD.n1828 VDD.n1079 0.878931
R13177 VDD.n5656 VDD.n5654 0.8405
R13178 VDD.n5654 VDD 0.8405
R13179 VDD.n7365 VDD.n7363 0.8405
R13180 VDD.n7363 VDD 0.8405
R13181 VDD.n3976 VDD.n3975 0.825441
R13182 VDD.n1704 VDD.n1703 0.824262
R13183 VDD.n3962 VDD.n3626 0.82077
R13184 VDD.n2378 VDD.n2377 0.813878
R13185 VDD.n4227 VDD.n4226 0.813878
R13186 VDD.n4078 VDD.n4073 0.813878
R13187 VDD.n4163 VDD.n4043 0.813878
R13188 VDD.n4573 VDD.n1006 0.813198
R13189 VDD.n2005 VDD.n1985 0.813198
R13190 VDD.n2103 VDD.n2083 0.813198
R13191 VDD.n2226 VDD.n2206 0.813198
R13192 VDD.n2360 VDD.n2224 0.813198
R13193 VDD.n1249 VDD.n1104 0.808921
R13194 VDD.n1230 VDD.n1114 0.808921
R13195 VDD.n1197 VDD.n1139 0.808921
R13196 VDD.n1178 VDD.n1149 0.808921
R13197 VDD.n4595 VDD.n990 0.808921
R13198 VDD.n983 VDD.n978 0.808921
R13199 VDD.n4649 VDD.n962 0.808921
R13200 VDD.n4667 VDD.n947 0.808921
R13201 VDD.n4706 VDD.n927 0.808921
R13202 VDD.n5452 VDD.n278 0.79598
R13203 VDD.n5394 VDD.n5393 0.79598
R13204 VDD.n5343 VDD.n344 0.79598
R13205 VDD.n388 VDD.n387 0.79598
R13206 VDD.n495 VDD.n434 0.79598
R13207 VDD.n554 VDD.n412 0.79598
R13208 VDD.n601 VDD.n600 0.79598
R13209 VDD.n5212 VDD.n637 0.79598
R13210 VDD.n5166 VDD.n675 0.79598
R13211 VDD.n4491 VDD.n2015 0.79404
R13212 VDD.n3354 VDD.n3353 0.775778
R13213 VDD.n3074 VDD.n3073 0.775778
R13214 VDD.n5649 VDD.n5648 0.761777
R13215 VDD.n6511 VDD.n6510 0.761777
R13216 VDD.n7358 VDD.n7357 0.761777
R13217 VDD.n8220 VDD.n8219 0.761777
R13218 VDD.n1866 VDD.n1055 0.761581
R13219 VDD.n3494 VDD.n3492 0.753441
R13220 VDD.n3501 VDD.n3492 0.753441
R13221 VDD.n3516 VDD.n3515 0.753441
R13222 VDD.n3515 VDD.n3507 0.753441
R13223 VDD.n3196 VDD.n3194 0.753441
R13224 VDD.n3203 VDD.n3194 0.753441
R13225 VDD.n3218 VDD.n3217 0.753441
R13226 VDD.n3217 VDD.n3209 0.753441
R13227 VDD.n3793 VDD.n3648 0.753441
R13228 VDD.n3744 VDD.n3742 0.753441
R13229 VDD.n3751 VDD.n3742 0.753441
R13230 VDD.n3836 VDD.n3835 0.753441
R13231 VDD.n3837 VDD.n3836 0.753441
R13232 VDD.n3841 VDD.n3735 0.753441
R13233 VDD.n3849 VDD.n3735 0.753441
R13234 VDD.n3886 VDD.n3885 0.753441
R13235 VDD.n3885 VDD.n3877 0.753441
R13236 VDD.n3859 VDD.n3858 0.753441
R13237 VDD.n3860 VDD.n3859 0.753441
R13238 VDD.n3863 VDD.n3707 0.753441
R13239 VDD.n3871 VDD.n3707 0.753441
R13240 VDD.n3917 VDD.n3916 0.753441
R13241 VDD.n3692 VDD.n3688 0.753441
R13242 VDD.n3779 VDD.n3778 0.753441
R13243 VDD.n2855 VDD.n2854 0.753441
R13244 VDD.n2824 VDD.n2822 0.753441
R13245 VDD.n2831 VDD.n2822 0.753441
R13246 VDD.n2879 VDD.n2878 0.753441
R13247 VDD.n2932 VDD.n2896 0.753441
R13248 VDD.n2966 VDD.n2964 0.753441
R13249 VDD.n2973 VDD.n2964 0.753441
R13250 VDD.n100 VDD.n43 0.753441
R13251 VDD.n51 VDD.n35 0.753441
R13252 VDD.n118 VDD.n111 0.753441
R13253 VDD.n130 VDD.n129 0.753441
R13254 VDD.n5546 VDD.n5543 0.753441
R13255 VDD.n5535 VDD.n5534 0.753441
R13256 VDD.n199 VDD.n188 0.753441
R13257 VDD.n227 VDD.n226 0.753441
R13258 VDD.n2527 VDD.n2515 0.753441
R13259 VDD.n2548 VDD.n2544 0.753441
R13260 VDD.n9001 VDD.n9000 0.750919
R13261 VDD.n8362 VDD.n8289 0.750919
R13262 VDD.n8146 VDD.n8145 0.750919
R13263 VDD.n7507 VDD.n7434 0.750919
R13264 VDD.n7292 VDD.n7291 0.750919
R13265 VDD.n6653 VDD.n6580 0.750919
R13266 VDD.n6437 VDD.n6436 0.750919
R13267 VDD.n5798 VDD.n5725 0.750919
R13268 VDD.n3919 VDD.n3657 0.743006
R13269 VDD.n2814 VDD.n2794 0.743006
R13270 VDD.n3806 VDD.n3762 0.742904
R13271 VDD.n4250 VDD.n2396 0.728259
R13272 VDD.n4204 VDD.n2435 0.728259
R13273 VDD.n4138 VDD.n4060 0.728259
R13274 VDD.n4194 VDD.n4193 0.728259
R13275 VDD.n2594 VDD.n2590 0.724685
R13276 VDD.n2593 VDD.n2590 0.724297
R13277 VDD.n4331 VDD.n4329 0.71293
R13278 VDD.n9001 VDD.n8271 0.708038
R13279 VDD.n8146 VDD.n7416 0.708038
R13280 VDD.n7292 VDD.n6562 0.708038
R13281 VDD.n6437 VDD.n5707 0.708038
R13282 VDD.n8403 VDD.n8282 0.700804
R13283 VDD.n7548 VDD.n7427 0.700804
R13284 VDD.n6694 VDD.n6573 0.700804
R13285 VDD.n5839 VDD.n5718 0.700804
R13286 VDD.n2357 VDD.n17 0.699924
R13287 VDD.n1506 VDD.n1504 0.69753
R13288 VDD.n1554 VDD.n1553 0.69753
R13289 VDD.n1306 VDD.n1305 0.69753
R13290 VDD.n1798 VDD.n1630 0.69753
R13291 VDD.n1663 VDD.n1660 0.69753
R13292 VDD.n1734 VDD.n1733 0.69753
R13293 VDD.n3975 VDD.n2507 0.692441
R13294 VDD.n3962 VDD.n3629 0.689368
R13295 VDD.n2454 VDD.n2442 0.687554
R13296 VDD.n5657 VDD 0.682932
R13297 VDD.n5657 VDD 0.682932
R13298 VDD.n7366 VDD 0.682932
R13299 VDD.n7366 VDD 0.682932
R13300 VDD.n138 VDD.n105 0.682531
R13301 VDD.n3454 VDD.n3453 0.682531
R13302 VDD.n3433 VDD.n3432 0.682531
R13303 VDD.n3424 VDD.n3423 0.682531
R13304 VDD.n3421 VDD.n3399 0.682531
R13305 VDD.n3316 VDD.n2767 0.6825
R13306 VDD.n3325 VDD.n2754 0.6825
R13307 VDD.n2870 VDD.n2775 0.6825
R13308 VDD.n8784 VDD.n8466 0.680146
R13309 VDD.n7929 VDD.n7611 0.680146
R13310 VDD.n7075 VDD.n6757 0.680146
R13311 VDD.n6220 VDD.n5902 0.680146
R13312 VDD.n4741 VDD.n909 0.677749
R13313 VDD.n4761 VDD.n4759 0.677749
R13314 VDD.n4799 VDD.n874 0.677749
R13315 VDD.n4817 VDD.n4816 0.677749
R13316 VDD.n4855 VDD.n847 0.677749
R13317 VDD.n4875 VDD.n4873 0.677749
R13318 VDD.n4913 VDD.n812 0.677749
R13319 VDD.n4931 VDD.n4930 0.677749
R13320 VDD.n4969 VDD.n785 0.677749
R13321 VDD.n4989 VDD.n4987 0.677749
R13322 VDD.n5027 VDD.n750 0.677749
R13323 VDD.n5045 VDD.n5044 0.677749
R13324 VDD.n5083 VDD.n723 0.677749
R13325 VDD.n5103 VDD.n5101 0.677749
R13326 VDD.n5141 VDD.n688 0.677749
R13327 VDD.t100 VDD.n1963 0.661784
R13328 VDD.t103 VDD.n2076 0.661784
R13329 VDD.n5406 VDD.n5405 0.651347
R13330 VDD.n5358 VDD.n334 0.651347
R13331 VDD.n375 VDD.n371 0.651347
R13332 VDD.n479 VDD.n440 0.651347
R13333 VDD.n539 VDD.n418 0.651347
R13334 VDD.n588 VDD.n584 0.651347
R13335 VDD.n5227 VDD.n628 0.651347
R13336 VDD.n5179 VDD.n5178 0.651347
R13337 VDD.n5456 VDD.n274 0.647691
R13338 VDD.n4278 VDD.n2373 0.64264
R13339 VDD.n2416 VDD.n2415 0.64264
R13340 VDD.n4105 VDD.n4104 0.64264
R13341 VDD.n4164 VDD.n4162 0.64264
R13342 VDD.n2451 VDD.n239 0.629701
R13343 VDD.n1844 VDD.n1066 0.627951
R13344 VDD.n1829 VDD.n1077 0.627951
R13345 VDD.n3111 VDD.n3108 0.614024
R13346 VDD.n8756 VDD.n8694 0.612674
R13347 VDD.n8834 VDD.n8833 0.612674
R13348 VDD.n8832 VDD.n8831 0.612674
R13349 VDD.n8711 VDD.n8699 0.612674
R13350 VDD.n7901 VDD.n7839 0.612674
R13351 VDD.n7979 VDD.n7978 0.612674
R13352 VDD.n7977 VDD.n7976 0.612674
R13353 VDD.n7856 VDD.n7844 0.612674
R13354 VDD.n7047 VDD.n6985 0.612674
R13355 VDD.n7125 VDD.n7124 0.612674
R13356 VDD.n7123 VDD.n7122 0.612674
R13357 VDD.n7002 VDD.n6990 0.612674
R13358 VDD.n6192 VDD.n6130 0.612674
R13359 VDD.n6270 VDD.n6269 0.612674
R13360 VDD.n6268 VDD.n6267 0.612674
R13361 VDD.n6147 VDD.n6135 0.612674
R13362 VDD.n1434 VDD.n1433 0.610024
R13363 VDD.n1946 VDD.n1945 0.610024
R13364 VDD.n2088 VDD.n2085 0.610024
R13365 VDD.n2166 VDD.n2165 0.610024
R13366 VDD.n8856 VDD.n8680 0.60463
R13367 VDD.n8691 VDD.n8689 0.60463
R13368 VDD.n8850 VDD.n8849 0.60463
R13369 VDD.n8847 VDD.n8846 0.60463
R13370 VDD.n8844 VDD.n8842 0.60463
R13371 VDD.n8840 VDD.n8692 0.60463
R13372 VDD.n8001 VDD.n7825 0.60463
R13373 VDD.n7836 VDD.n7834 0.60463
R13374 VDD.n7995 VDD.n7994 0.60463
R13375 VDD.n7992 VDD.n7991 0.60463
R13376 VDD.n7989 VDD.n7987 0.60463
R13377 VDD.n7985 VDD.n7837 0.60463
R13378 VDD.n7147 VDD.n6971 0.60463
R13379 VDD.n6982 VDD.n6980 0.60463
R13380 VDD.n7141 VDD.n7140 0.60463
R13381 VDD.n7138 VDD.n7137 0.60463
R13382 VDD.n7135 VDD.n7133 0.60463
R13383 VDD.n7131 VDD.n6983 0.60463
R13384 VDD.n6292 VDD.n6116 0.60463
R13385 VDD.n6127 VDD.n6125 0.60463
R13386 VDD.n6286 VDD.n6285 0.60463
R13387 VDD.n6283 VDD.n6282 0.60463
R13388 VDD.n6280 VDD.n6278 0.60463
R13389 VDD.n6276 VDD.n6128 0.60463
R13390 VDD.n2948 VDD.n2947 0.604026
R13391 VDD.n3021 VDD.n2890 0.603703
R13392 VDD.n2890 VDD.n2888 0.576974
R13393 VDD.n1471 VDD.n1469 0.570797
R13394 VDD.n1881 VDD.n1046 0.570797
R13395 VDD.n5600 VDD.n5599 0.568833
R13396 VDD.n5607 VDD.n0 0.55916
R13397 VDD.n4249 VDD.n2397 0.557022
R13398 VDD.n4201 VDD.n4200 0.557022
R13399 VDD.n4139 VDD.n4058 0.557022
R13400 VDD.n5457 VDD.n273 0.557022
R13401 VDD.n5655 VDD.n5612 0.544383
R13402 VDD.n6528 VDD.n6527 0.544383
R13403 VDD.n7364 VDD.n7321 0.544383
R13404 VDD.n8237 VDD.n8236 0.544383
R13405 VDD.n1895 VDD.n1005 0.542299
R13406 VDD.n1983 VDD.n1977 0.542299
R13407 VDD.n4442 VDD.n2082 0.542299
R13408 VDD.n2204 VDD.n2198 0.542299
R13409 VDD.n1246 VDD.n1245 0.539447
R13410 VDD.n1234 VDD.n1233 0.539447
R13411 VDD.n1194 VDD.n1193 0.539447
R13412 VDD.n1182 VDD.n1181 0.539447
R13413 VDD.n4600 VDD.n4598 0.539447
R13414 VDD.n4611 VDD.n4610 0.539447
R13415 VDD.n4656 VDD.n957 0.539447
R13416 VDD.n4668 VDD.n4666 0.539447
R13417 VDD.n4712 VDD.n4709 0.539447
R13418 VDD.n6526 VDD 0.530391
R13419 VDD.n8235 VDD 0.530391
R13420 VDD.n4356 VDD.n2235 0.529527
R13421 VDD.n2340 VDD.n2339 0.522949
R13422 VDD.n8364 VDD.n8363 0.515073
R13423 VDD.n7509 VDD.n7508 0.515073
R13424 VDD.n6655 VDD.n6654 0.515073
R13425 VDD.n5800 VDD.n5799 0.515073
R13426 VDD.n5453 VDD.n277 0.506715
R13427 VDD.n5397 VDD.n316 0.506715
R13428 VDD.n5344 VDD.n342 0.506715
R13429 VDD.n5299 VDD.n381 0.506715
R13430 VDD.n494 VDD.n436 0.506715
R13431 VDD.n551 VDD.n550 0.506715
R13432 VDD.n5266 VDD.n594 0.506715
R13433 VDD.n5216 VDD.n5215 0.506715
R13434 VDD.n5167 VDD.n672 0.506715
R13435 VDD.n1858 VDD.n1057 0.502461
R13436 VDD.n6525 VDD 0.497949
R13437 VDD.n8234 VDD 0.497949
R13438 VDD.n2629 VDD.n2628 0.491125
R13439 VDD.n3966 VDD.n3965 0.488891
R13440 VDD.n2630 VDD.n2629 0.488
R13441 VDD.n1870 VDD.n1869 0.484824
R13442 VDD.n3918 VDD.n3665 0.48381
R13443 VDD.n2809 VDD.n2808 0.483797
R13444 VDD.n123 VDD.n108 0.476817
R13445 VDD.n1404 VDD.n1401 0.474574
R13446 VDD.n1462 VDD.n1405 0.474574
R13447 VDD.n1459 VDD.n1458 0.474574
R13448 VDD.n1409 VDD.n1407 0.474574
R13449 VDD.n1451 VDD.n1448 0.474574
R13450 VDD.n1444 VDD.n1410 0.474574
R13451 VDD.n1441 VDD.n1440 0.474574
R13452 VDD.n1415 VDD.n1412 0.474574
R13453 VDD.n1433 VDD.n1430 0.474574
R13454 VDD.n1426 VDD.n1417 0.474574
R13455 VDD.n1423 VDD.n1422 0.474574
R13456 VDD.n1476 VDD.n1388 0.474574
R13457 VDD.n1894 VDD.n1028 0.474574
R13458 VDD.n1896 VDD.n1895 0.474574
R13459 VDD.n4574 VDD.n4573 0.474574
R13460 VDD.n1010 VDD.n1009 0.474574
R13461 VDD.n1905 VDD.n1904 0.474574
R13462 VDD.n4562 VDD.n1021 0.474574
R13463 VDD.n1025 VDD.n1022 0.474574
R13464 VDD.n4557 VDD.n1026 0.474574
R13465 VDD.n1916 VDD.n1915 0.474574
R13466 VDD.n1936 VDD.n1935 0.474574
R13467 VDD.n4543 VDD.n1926 0.474574
R13468 VDD.n1930 VDD.n1927 0.474574
R13469 VDD.n4538 VDD.n1931 0.474574
R13470 VDD.n1947 VDD.n1946 0.474574
R13471 VDD.n1971 VDD.n1970 0.474574
R13472 VDD.n4524 VDD.n1956 0.474574
R13473 VDD.n4517 VDD.n1961 0.474574
R13474 VDD.n1976 VDD.n1966 0.474574
R13475 VDD.n4513 VDD.n1977 0.474574
R13476 VDD.n1985 VDD.n1984 0.474574
R13477 VDD.n2008 VDD.n2007 0.474574
R13478 VDD.n4499 VDD.n1998 0.474574
R13479 VDD.n2002 VDD.n1999 0.474574
R13480 VDD.n4494 VDD.n2003 0.474574
R13481 VDD.n2020 VDD.n2019 0.474574
R13482 VDD.n2041 VDD.n2040 0.474574
R13483 VDD.n4480 VDD.n2031 0.474574
R13484 VDD.n2035 VDD.n2032 0.474574
R13485 VDD.n4475 VDD.n2036 0.474574
R13486 VDD.n2052 VDD.n2051 0.474574
R13487 VDD.n2088 VDD.n2087 0.474574
R13488 VDD.n4461 VDD.n2060 0.474574
R13489 VDD.n2064 VDD.n2061 0.474574
R13490 VDD.n2078 VDD.n2066 0.474574
R13491 VDD.n4446 VDD.n2079 0.474574
R13492 VDD.n2082 VDD.n2080 0.474574
R13493 VDD.n4441 VDD.n2083 0.474574
R13494 VDD.n2105 VDD.n2104 0.474574
R13495 VDD.n2125 VDD.n2124 0.474574
R13496 VDD.n4427 VDD.n2115 0.474574
R13497 VDD.n2119 VDD.n2116 0.474574
R13498 VDD.n4422 VDD.n2120 0.474574
R13499 VDD.n2135 VDD.n2134 0.474574
R13500 VDD.n2156 VDD.n2155 0.474574
R13501 VDD.n4408 VDD.n2146 0.474574
R13502 VDD.n2150 VDD.n2147 0.474574
R13503 VDD.n4403 VDD.n2151 0.474574
R13504 VDD.n2167 VDD.n2166 0.474574
R13505 VDD.n2192 VDD.n2191 0.474574
R13506 VDD.n4389 VDD.n2177 0.474574
R13507 VDD.n4382 VDD.n2182 0.474574
R13508 VDD.n2197 VDD.n2187 0.474574
R13509 VDD.n4378 VDD.n2198 0.474574
R13510 VDD.n2206 VDD.n2205 0.474574
R13511 VDD.n2229 VDD.n2228 0.474574
R13512 VDD.n4364 VDD.n2219 0.474574
R13513 VDD.n2223 VDD.n2220 0.474574
R13514 VDD.n3023 VDD.n3022 0.473002
R13515 VDD.n4279 VDD.n2371 0.471403
R13516 VDD.n4233 VDD.n2408 0.471403
R13517 VDD.n4099 VDD.n4077 0.471403
R13518 VDD.n4051 VDD.n4046 0.471403
R13519 VDD.n3680 VDD.n3671 0.469257
R13520 VDD.n3809 VDD.n3807 0.469245
R13521 VDD.n5491 VDD.n5489 0.461585
R13522 VDD.n5495 VDD.n252 0.452151
R13523 VDD.n2977 VDD.n2976 0.444775
R13524 VDD.n1367 VDD.n1366 0.444064
R13525 VDD.n1328 VDD.n1327 0.444064
R13526 VDD.n1584 VDD.n1309 0.444064
R13527 VDD.n1796 VDD.n1631 0.444064
R13528 VDD.n1658 VDD.n1651 0.444064
R13529 VDD.n1705 VDD.n1046 0.444064
R13530 VDD.n8239 VDD 0.435138
R13531 VDD.n5446 VDD.n5445 0.431961
R13532 VDD.n1465 VDD.n1372 0.428211
R13533 VDD.n6530 VDD 0.427658
R13534 VDD.n4122 VDD.t52 0.42104
R13535 VDD.n268 VDD.n245 0.42104
R13536 VDD.n5473 VDD.n248 0.42104
R13537 VDD.n5459 VDD.n247 0.42104
R13538 VDD.n4748 VDD.n904 0.406849
R13539 VDD.n902 VDD.n897 0.406849
R13540 VDD.n4804 VDD.n4802 0.406849
R13541 VDD.n4811 VDD.n867 0.406849
R13542 VDD.n4862 VDD.n842 0.406849
R13543 VDD.n840 VDD.n835 0.406849
R13544 VDD.n4918 VDD.n4916 0.406849
R13545 VDD.n4925 VDD.n805 0.406849
R13546 VDD.n4976 VDD.n780 0.406849
R13547 VDD.n778 VDD.n773 0.406849
R13548 VDD.n5032 VDD.n5030 0.406849
R13549 VDD.n5039 VDD.n743 0.406849
R13550 VDD.n5090 VDD.n718 0.406849
R13551 VDD.n716 VDD.n711 0.406849
R13552 VDD.n5146 VDD.n5144 0.406849
R13553 VDD.n5157 VDD.n681 0.406849
R13554 VDD.n3455 VDD.n2694 0.400769
R13555 VDD.n3445 VDD.n3444 0.400769
R13556 VDD.n3391 VDD.n3390 0.400769
R13557 VDD.n2721 VDD.n2714 0.400768
R13558 VDD.n3417 VDD.n3416 0.400768
R13559 VDD.n3361 VDD.n3360 0.400768
R13560 VDD.n3289 VDD.n3288 0.400768
R13561 VDD.n4564 VDD.n1019 0.39727
R13562 VDD.n4246 VDD.n4245 0.385784
R13563 VDD.n4086 VDD.n4085 0.385784
R13564 VDD.n4144 VDD.n4142 0.385784
R13565 VDD.n1494 VDD.n1371 0.380698
R13566 VDD.n1368 VDD.n1367 0.380698
R13567 VDD.n1504 VDD.n1362 0.380698
R13568 VDD.n1505 VDD.n1360 0.380698
R13569 VDD.n1510 VDD.n1357 0.380698
R13570 VDD.n1355 VDD.n1351 0.380698
R13571 VDD.n1520 VDD.n1349 0.380698
R13572 VDD.n1526 VDD.n1525 0.380698
R13573 VDD.n1533 VDD.n1532 0.380698
R13574 VDD.n1538 VDD.n1343 0.380698
R13575 VDD.n1340 VDD.n1339 0.380698
R13576 VDD.n1548 VDD.n1334 0.380698
R13577 VDD.n1549 VDD.n1332 0.380698
R13578 VDD.n1554 VDD.n1329 0.380698
R13579 VDD.n1327 VDD.n1322 0.380698
R13580 VDD.n1564 VDD.n1323 0.380698
R13581 VDD.n1579 VDD.n1311 0.380698
R13582 VDD.n1580 VDD.n1309 0.380698
R13583 VDD.n1585 VDD.n1306 0.380698
R13584 VDD.n1304 VDD.n1300 0.380698
R13585 VDD.n1595 VDD.n1298 0.380698
R13586 VDD.n1601 VDD.n1600 0.380698
R13587 VDD.n1608 VDD.n1607 0.380698
R13588 VDD.n1613 VDD.n1292 0.380698
R13589 VDD.n1289 VDD.n1288 0.380698
R13590 VDD.n1812 VDD.n1280 0.380698
R13591 VDD.n1284 VDD.n1281 0.380698
R13592 VDD.n1807 VDD.n1285 0.380698
R13593 VDD.n1627 VDD.n1626 0.380698
R13594 VDD.n1798 VDD.n1797 0.380698
R13595 VDD.n1634 VDD.n1631 0.380698
R13596 VDD.n1792 VDD.n1635 0.380698
R13597 VDD.n1650 VDD.n1649 0.380698
R13598 VDD.n1778 VDD.n1651 0.380698
R13599 VDD.n1660 VDD.n1659 0.380698
R13600 VDD.n1769 VDD.n1768 0.380698
R13601 VDD.n1667 VDD.n1664 0.380698
R13602 VDD.n1763 VDD.n1668 0.380698
R13603 VDD.n1677 VDD.n1676 0.380698
R13604 VDD.n1754 VDD.n1753 0.380698
R13605 VDD.n1684 VDD.n1681 0.380698
R13606 VDD.n1748 VDD.n1685 0.380698
R13607 VDD.n1694 VDD.n1693 0.380698
R13608 VDD.n1739 VDD.n1738 0.380698
R13609 VDD.n1701 VDD.n1698 0.380698
R13610 VDD.n1733 VDD.n1702 0.380698
R13611 VDD.n5455 VDD.n5454 0.378512
R13612 VDD.n3584 VDD.n2664 0.376971
R13613 VDD.n3584 VDD.n2665 0.376971
R13614 VDD.n3554 VDD.n3553 0.376971
R13615 VDD.n3550 VDD.n3549 0.376971
R13616 VDD.n3256 VDD.n3255 0.376971
R13617 VDD.n3252 VDD.n3251 0.376971
R13618 VDD.n3140 VDD.n3133 0.376971
R13619 VDD.n3140 VDD.n3134 0.376971
R13620 VDD.n3790 VDD.n3789 0.376971
R13621 VDD.n3789 VDD.n3766 0.376971
R13622 VDD.n3785 VDD.n3784 0.376971
R13623 VDD.n3640 VDD.n3637 0.376971
R13624 VDD.n2927 VDD.n2922 0.376971
R13625 VDD.n2927 VDD.n2919 0.376971
R13626 VDD.n2937 VDD.n2920 0.376971
R13627 VDD.n2912 VDD.n2910 0.376971
R13628 VDD.n2996 VDD.n2917 0.376971
R13629 VDD.n99 VDD.n45 0.376971
R13630 VDD.n96 VDD.n48 0.376971
R13631 VDD.n87 VDD.n49 0.376971
R13632 VDD.n79 VDD.n78 0.376971
R13633 VDD.n70 VDD.n69 0.376971
R13634 VDD.n69 VDD.n61 0.376971
R13635 VDD.n133 VDD.n113 0.376971
R13636 VDD.n5557 VDD.n5545 0.376971
R13637 VDD.n5554 VDD.n5549 0.376971
R13638 VDD.n5595 VDD.n5594 0.376971
R13639 VDD.n5562 VDD.n5533 0.376971
R13640 VDD.n5574 VDD.n5568 0.376971
R13641 VDD.n5574 VDD.n5573 0.376971
R13642 VDD.n198 VDD.n190 0.376971
R13643 VDD.n195 VDD.n193 0.376971
R13644 VDD.n236 VDD.n235 0.376971
R13645 VDD.n225 VDD.n224 0.376971
R13646 VDD.n216 VDD.n215 0.376971
R13647 VDD.n215 VDD.n207 0.376971
R13648 VDD.n1843 VDD.n1070 0.376971
R13649 VDD.n1833 VDD.n1832 0.376971
R13650 VDD.n5402 VDD.n309 0.362082
R13651 VDD.n5355 VDD.n5354 0.362082
R13652 VDD.n5304 VDD.n376 0.362082
R13653 VDD.n484 VDD.n482 0.362082
R13654 VDD.n540 VDD.n416 0.362082
R13655 VDD.n5271 VDD.n589 0.362082
R13656 VDD.n5226 VDD.n629 0.362082
R13657 VDD.n670 VDD.n666 0.362082
R13658 VDD.n2577 VDD.n2516 0.357498
R13659 VDD.n1880 VDD.n1047 0.346446
R13660 VDD.n8385 VDD.n8384 0.343549
R13661 VDD.n8380 VDD.n8297 0.343549
R13662 VDD.n8379 VDD.n8377 0.343549
R13663 VDD.n8376 VDD.n8374 0.343549
R13664 VDD.n8371 VDD.n8301 0.343549
R13665 VDD.n8370 VDD.n8369 0.343549
R13666 VDD.n7530 VDD.n7529 0.343549
R13667 VDD.n7525 VDD.n7442 0.343549
R13668 VDD.n7524 VDD.n7522 0.343549
R13669 VDD.n7521 VDD.n7519 0.343549
R13670 VDD.n7516 VDD.n7446 0.343549
R13671 VDD.n7515 VDD.n7514 0.343549
R13672 VDD.n6676 VDD.n6675 0.343549
R13673 VDD.n6671 VDD.n6588 0.343549
R13674 VDD.n6670 VDD.n6668 0.343549
R13675 VDD.n6667 VDD.n6665 0.343549
R13676 VDD.n6662 VDD.n6592 0.343549
R13677 VDD.n6661 VDD.n6660 0.343549
R13678 VDD.n5821 VDD.n5820 0.343549
R13679 VDD.n5816 VDD.n5733 0.343549
R13680 VDD.n5815 VDD.n5813 0.343549
R13681 VDD.n5812 VDD.n5810 0.343549
R13682 VDD.n5807 VDD.n5737 0.343549
R13683 VDD.n5806 VDD.n5805 0.343549
R13684 VDD.n2835 VDD.n2834 0.34084
R13685 VDD.n1427 VDD.n1426 0.339124
R13686 VDD.n1970 VDD.n1968 0.339124
R13687 VDD.n2086 VDD.n2060 0.339124
R13688 VDD.n2191 VDD.n2189 0.339124
R13689 VDD.n4722 VDD.n4721 0.337342
R13690 VDD.n2488 VDD.n2479 0.33059
R13691 VDD.n4008 VDD.n2480 0.33059
R13692 VDD.n2482 VDD.n394 0.33059
R13693 VDD.n6523 VDD 0.329892
R13694 VDD.n8232 VDD 0.329892
R13695 VDD.n3934 VDD.n3933 0.324719
R13696 VDD.n3931 VDD.n3930 0.324719
R13697 VDD.n3689 VDD.n3656 0.324719
R13698 VDD.n2688 VDD.n2687 0.324719
R13699 VDD.n3473 VDD.n3472 0.324719
R13700 VDD.n3300 VDD.n3068 0.324719
R13701 VDD.n3175 VDD.n3174 0.324719
R13702 VDD.n1377 VDD.n1373 0.317332
R13703 VDD.n1490 VDD.n1488 0.317332
R13704 VDD.n1569 VDD.n1568 0.317332
R13705 VDD.n1317 VDD.n1316 0.317332
R13706 VDD.n1644 VDD.n1643 0.317332
R13707 VDD.n1783 VDD.n1782 0.317332
R13708 VDD.n1867 VDD.n1056 0.313753
R13709 VDD.n4293 VDD.n2360 0.30922
R13710 VDD.n4283 VDD.n4282 0.300166
R13711 VDD.n4234 VDD.n2405 0.300166
R13712 VDD.n4100 VDD.n4098 0.300166
R13713 VDD.n4156 VDD.n4155 0.300166
R13714 VDD.n6527 VDD 0.299413
R13715 VDD.n8236 VDD 0.299413
R13716 VDD.n6529 VDD.n6466 0.292759
R13717 VDD.n8238 VDD.n8175 0.292759
R13718 VDD.n5674 VDD.n5673 0.292507
R13719 VDD.n7383 VDD.n7382 0.292507
R13720 VDD.n3381 VDD.n3380 0.278729
R13721 VDD.n3435 VDD.n3434 0.278729
R13722 VDD.n3471 VDD.n2691 0.278729
R13723 VDD.n3404 VDD.n2731 0.278729
R13724 VDD.n3177 VDD.n3086 0.278729
R13725 VDD.n3431 VDD.n2711 0.278729
R13726 VDD.n3475 VDD.n2680 0.278729
R13727 VDD.n5675 VDD 0.278033
R13728 VDD.n7384 VDD 0.278033
R13729 VDD.n4725 VDD.n917 0.27309
R13730 VDD.n1477 VDD.n1387 0.271399
R13731 VDD.n1897 VDD.n1894 0.271399
R13732 VDD.n1960 VDD.n1957 0.271399
R13733 VDD.n4514 VDD.n1976 0.271399
R13734 VDD.n4457 VDD.n4456 0.271399
R13735 VDD.n4446 VDD.n4445 0.271399
R13736 VDD.n2181 VDD.n2178 0.271399
R13737 VDD.n4379 VDD.n2197 0.271399
R13738 VDD.n1241 VDD.n1106 0.269974
R13739 VDD.n1113 VDD.n1110 0.269974
R13740 VDD.n1189 VDD.n1141 0.269974
R13741 VDD.n1148 VDD.n1145 0.269974
R13742 VDD.n4599 VDD.n985 0.269974
R13743 VDD.n986 VDD.n982 0.269974
R13744 VDD.n4657 VDD.n954 0.269974
R13745 VDD.n955 VDD.n950 0.269974
R13746 VDD.n4711 VDD.n4710 0.269974
R13747 VDD.n2866 VDD.n2864 0.26925
R13748 VDD.n9023 VDD.n9022 0.267107
R13749 VDD.n8168 VDD.n8167 0.267107
R13750 VDD.n7314 VDD.n7313 0.267107
R13751 VDD.n6459 VDD.n6458 0.267107
R13752 VDD.n1979 VDD.t100 0.265013
R13753 VDD.n2099 VDD.t103 0.265013
R13754 VDD.n5661 VDD.n5649 0.26137
R13755 VDD.n5661 VDD.n5660 0.26137
R13756 VDD.n5660 VDD.n5659 0.26137
R13757 VDD.n6512 VDD.n6511 0.26137
R13758 VDD.n6512 VDD.n6467 0.26137
R13759 VDD.n6520 VDD.n6467 0.26137
R13760 VDD.n7370 VDD.n7358 0.26137
R13761 VDD.n7370 VDD.n7369 0.26137
R13762 VDD.n7369 VDD.n7368 0.26137
R13763 VDD.n8221 VDD.n8220 0.26137
R13764 VDD.n8221 VDD.n8176 0.26137
R13765 VDD.n8229 VDD.n8176 0.26137
R13766 VDD.n2346 VDD 0.260619
R13767 VDD.n2355 VDD.n2354 0.25512
R13768 VDD.n5156 VDD.n674 0.236946
R13769 VDD.n5666 VDD.n5643 0.231925
R13770 VDD.n6517 VDD.n6506 0.231925
R13771 VDD.n7375 VDD.n7352 0.231925
R13772 VDD.n8226 VDD.n8215 0.231925
R13773 VDD.n5666 VDD.n5665 0.231891
R13774 VDD.n5666 VDD.n5644 0.231891
R13775 VDD.n6517 VDD.n6516 0.231891
R13776 VDD.n6518 VDD.n6517 0.231891
R13777 VDD.n7375 VDD.n7374 0.231891
R13778 VDD.n7375 VDD.n7353 0.231891
R13779 VDD.n8226 VDD.n8225 0.231891
R13780 VDD.n8227 VDD.n8226 0.231891
R13781 VDD.n3520 VDD.n3504 0.229427
R13782 VDD.n3520 VDD.n3519 0.229427
R13783 VDD.n3222 VDD.n3206 0.229427
R13784 VDD.n3222 VDD.n3221 0.229427
R13785 VDD.n3830 VDD.n3754 0.229427
R13786 VDD.n3832 VDD.n3830 0.229427
R13787 VDD.n3853 VDD.n3852 0.229427
R13788 VDD.n3855 VDD.n3853 0.229427
R13789 VDD.n3890 VDD.n3874 0.229427
R13790 VDD.n3890 VDD.n3889 0.229427
R13791 VDD.n6530 VDD.n6529 0.223437
R13792 VDD.n8239 VDD.n8238 0.22328
R13793 VDD.n5675 VDD.n5674 0.222418
R13794 VDD.n7384 VDD.n7383 0.222418
R13795 VDD.n5398 VDD.n315 0.217449
R13796 VDD.n5348 VDD.n5347 0.217449
R13797 VDD.n5300 VDD.n380 0.217449
R13798 VDD.n491 VDD.n490 0.217449
R13799 VDD.n545 VDD.n414 0.217449
R13800 VDD.n5267 VDD.n593 0.217449
R13801 VDD.n636 VDD.n632 0.217449
R13802 VDD.n5171 VDD.n5170 0.217449
R13803 VDD.n4292 VDD.n4291 0.216346
R13804 VDD.n3521 VDD.n3520 0.215848
R13805 VDD.n3223 VDD.n3222 0.215848
R13806 VDD.n3853 VDD.n3732 0.215848
R13807 VDD.n3891 VDD.n3890 0.215848
R13808 VDD.n3830 VDD.n3829 0.215848
R13809 VDD.n8245 VDD 0.215174
R13810 VDD.n7390 VDD 0.215174
R13811 VDD.n6536 VDD 0.215174
R13812 VDD.n5681 VDD 0.215174
R13813 VDD.n2403 VDD.n2400 0.214547
R13814 VDD.n4087 VDD.n4084 0.214547
R13815 VDD.n4143 VDD.n4053 0.214547
R13816 VDD.n1272 VDD.n1271 0.214355
R13817 VDD.n4292 VDD.n2359 0.211367
R13818 VDD.n2604 VDD.n1019 0.211364
R13819 VDD.n3983 VDD.n2499 0.211364
R13820 VDD.n143 VDD.n140 0.210656
R13821 VDD.n3612 VDD.n2635 0.210461
R13822 VDD.n3171 VDD.n3093 0.210461
R13823 VDD.n1054 VDD.n1050 0.208068
R13824 VDD.n5606 VDD.n2 0.204334
R13825 VDD.n1421 VDD.n1387 0.203675
R13826 VDD.n4523 VDD.n1957 0.203675
R13827 VDD.n4457 VDD.n2065 0.203675
R13828 VDD.n4388 VDD.n2178 0.203675
R13829 VDD.n3379 VDD.n3378 0.202844
R13830 VDD.n8363 VDD.n8362 0.193465
R13831 VDD.n7508 VDD.n7507 0.193465
R13832 VDD.n6654 VDD.n6653 0.193465
R13833 VDD.n5799 VDD.n5798 0.193465
R13834 VDD.n3552 VDD.n3551 0.190717
R13835 VDD.n3254 VDD.n3253 0.190717
R13836 VDD.n3846 VDD.n3736 0.190717
R13837 VDD.n3847 VDD.n3846 0.190717
R13838 VDD.n3868 VDD.n3708 0.190717
R13839 VDD.n3869 VDD.n3868 0.190717
R13840 VDD.n1494 VDD.n1493 0.190599
R13841 VDD.n1565 VDD.n1564 0.190599
R13842 VDD.n1581 VDD.n1579 0.190599
R13843 VDD.n1793 VDD.n1792 0.190599
R13844 VDD.n1779 VDD.n1650 0.190599
R13845 VDD.n2558 VDD.n2517 0.189124
R13846 VDD.n5492 VDD.n249 0.186007
R13847 VDD.n2576 VDD.n2519 0.178063
R13848 VDD.n5673 VDD 0.174685
R13849 VDD.n7382 VDD 0.174685
R13850 VDD VDD.n6466 0.174507
R13851 VDD VDD.n8175 0.174507
R13852 VDD.n5656 VDD 0.167831
R13853 VDD.n7365 VDD 0.167831
R13854 VDD.n8716 VDD.n8713 0.167457
R13855 VDD.n7861 VDD.n7858 0.167457
R13856 VDD.n7007 VDD.n7004 0.167457
R13857 VDD.n6152 VDD.n6149 0.167457
R13858 VDD.n2578 VDD.n2515 0.166946
R13859 VDD.n3522 VDD.n3521 0.164777
R13860 VDD.n3224 VDD.n3223 0.164777
R13861 VDD.n3732 VDD.n3731 0.164777
R13862 VDD.n3892 VDD.n3891 0.164777
R13863 VDD.n3829 VDD.n3828 0.164777
R13864 VDD.n2979 VDD.n2977 0.164777
R13865 VDD.n3580 VDD.n2681 0.161367
R13866 VDD.n3525 VDD.n2670 0.161367
R13867 VDD.n3469 VDD.n3468 0.161367
R13868 VDD.n3447 VDD.n3446 0.161367
R13869 VDD.n3429 VDD.n3428 0.161367
R13870 VDD.n3415 VDD.n3413 0.161367
R13871 VDD.n3393 VDD.n3392 0.161367
R13872 VDD.n3359 VDD.n3358 0.161367
R13873 VDD.n3287 VDD.n3286 0.161367
R13874 VDD.n3282 VDD.n3087 0.161367
R13875 VDD.n3227 VDD.n3076 0.161367
R13876 VDD.n3825 VDD.n3757 0.161367
R13877 VDD.n3728 VDD.n3666 0.161367
R13878 VDD.n3895 VDD.n3673 0.161367
R13879 VDD.n2839 VDD.n2810 0.161367
R13880 VDD.n3504 VDD.n3490 0.15935
R13881 VDD.n3519 VDD.n3518 0.15935
R13882 VDD.n3206 VDD.n3192 0.15935
R13883 VDD.n3221 VDD.n3220 0.15935
R13884 VDD.n3754 VDD.n3740 0.15935
R13885 VDD.n3833 VDD.n3832 0.15935
R13886 VDD.n3852 VDD.n3733 0.15935
R13887 VDD.n3856 VDD.n3855 0.15935
R13888 VDD.n3874 VDD.n3705 0.15935
R13889 VDD.n3889 VDD.n3888 0.15935
R13890 VDD.n2834 VDD.n2820 0.15935
R13891 VDD.n2976 VDD.n2962 0.15935
R13892 VDD.n4296 VDD.n4294 0.157987
R13893 VDD.n3574 VDD.n2679 0.150167
R13894 VDD.n3530 VDD.n2671 0.150167
R13895 VDD.n3464 VDD.n2695 0.150167
R13896 VDD.n3438 VDD.n3437 0.150167
R13897 VDD.n2720 VDD.n2719 0.150167
R13898 VDD.n3405 VDD.n3403 0.150167
R13899 VDD.n3384 VDD.n3383 0.150167
R13900 VDD.n3370 VDD.n3352 0.150167
R13901 VDD.n3297 VDD.n3295 0.150167
R13902 VDD.n3276 VDD.n3085 0.150167
R13903 VDD.n3232 VDD.n3077 0.150167
R13904 VDD.n3820 VDD.n3759 0.150167
R13905 VDD.n3723 VDD.n3661 0.150167
R13906 VDD.n3900 VDD.n3675 0.150167
R13907 VDD.n2848 VDD.n2812 0.150167
R13908 VDD.n9028 VDD 0.145785
R13909 VDD.n8173 VDD 0.145785
R13910 VDD.n7319 VDD 0.145785
R13911 VDD.n6464 VDD 0.145785
R13912 VDD.n3592 VDD.n2648 0.144522
R13913 VDD.n3590 VDD.n2660 0.144522
R13914 VDD.n3562 VDD.n3561 0.144522
R13915 VDD.n3557 VDD.n3556 0.144522
R13916 VDD.n3547 VDD.n3546 0.144522
R13917 VDD.n3542 VDD.n3541 0.144522
R13918 VDD.n3537 VDD.n3536 0.144522
R13919 VDD.n3532 VDD.n3531 0.144522
R13920 VDD.n3527 VDD.n3526 0.144522
R13921 VDD.n3264 VDD.n3263 0.144522
R13922 VDD.n3259 VDD.n3258 0.144522
R13923 VDD.n3249 VDD.n3248 0.144522
R13924 VDD.n3244 VDD.n3243 0.144522
R13925 VDD.n3239 VDD.n3238 0.144522
R13926 VDD.n3234 VDD.n3233 0.144522
R13927 VDD.n3229 VDD.n3228 0.144522
R13928 VDD.n3148 VDD.n3121 0.144522
R13929 VDD.n3146 VDD.n3129 0.144522
R13930 VDD.n3722 VDD.n3721 0.144522
R13931 VDD.n3727 VDD.n3726 0.144522
R13932 VDD.n3902 VDD.n3901 0.144522
R13933 VDD.n3897 VDD.n3896 0.144522
R13934 VDD.n3819 VDD.n3818 0.144522
R13935 VDD.n3824 VDD.n3823 0.144522
R13936 VDD.n2846 VDD.n2845 0.144522
R13937 VDD.n2841 VDD.n2840 0.144522
R13938 VDD.n2955 VDD.n2954 0.144522
R13939 VDD.n2961 VDD.n2960 0.144522
R13940 VDD.n73 VDD.n72 0.144522
R13941 VDD.n5577 VDD.n5565 0.144522
R13942 VDD.n219 VDD.n218 0.144522
R13943 VDD.n2836 VDD.n2835 0.141804
R13944 VDD.n3479 VDD.n2669 0.138912
R13945 VDD.n3535 VDD.n2672 0.138912
R13946 VDD.n3181 VDD.n3075 0.138912
R13947 VDD.n3237 VDD.n3078 0.138912
R13948 VDD.n4749 VDD.n901 0.13595
R13949 VDD.n4753 VDD.n4752 0.13595
R13950 VDD.n4803 VDD.n870 0.13595
R13951 VDD.n4812 VDD.n4810 0.13595
R13952 VDD.n4863 VDD.n839 0.13595
R13953 VDD.n4867 VDD.n4866 0.13595
R13954 VDD.n4917 VDD.n808 0.13595
R13955 VDD.n4926 VDD.n4924 0.13595
R13956 VDD.n4977 VDD.n777 0.13595
R13957 VDD.n4981 VDD.n4980 0.13595
R13958 VDD.n5031 VDD.n746 0.13595
R13959 VDD.n5040 VDD.n5038 0.13595
R13960 VDD.n5091 VDD.n715 0.13595
R13961 VDD.n5095 VDD.n5094 0.13595
R13962 VDD.n5145 VDD.n683 0.13595
R13963 VDD.n5154 VDD.n5153 0.13595
R13964 VDD.n8246 VDD.n8245 0.134558
R13965 VDD.n7391 VDD.n7390 0.134558
R13966 VDD.n6537 VDD.n6536 0.134558
R13967 VDD.n5682 VDD.n5681 0.134558
R13968 VDD.n3983 VDD.n2015 0.132757
R13969 VDD.n2370 VDD.n2364 0.128928
R13970 VDD.n4238 VDD.n4237 0.128928
R13971 VDD.n4091 VDD.n4080 0.128928
R13972 VDD.n4054 VDD.n4050 0.128928
R13973 VDD.n3563 VDD.n2677 0.127599
R13974 VDD.n3540 VDD.n2673 0.127599
R13975 VDD.n3265 VDD.n3083 0.127599
R13976 VDD.n3242 VDD.n3079 0.127599
R13977 VDD.n5605 VDD.n5604 0.1274
R13978 VDD.n1840 VDD.n1839 0.12599
R13979 VDD.n1076 VDD.n1072 0.12599
R13980 VDD.n5606 VDD.n5605 0.122353
R13981 VDD.n5607 VDD.n5606 0.119879
R13982 VDD.n5602 VDD.n17 0.117099
R13983 VDD.n3558 VDD.n2676 0.116231
R13984 VDD.n3545 VDD.n2674 0.116231
R13985 VDD.n3260 VDD.n3082 0.116231
R13986 VDD.n3247 VDD.n3080 0.116231
R13987 VDD.n2342 VDD 0.116103
R13988 VDD.n2343 VDD 0.116103
R13989 VDD.n3043 VDD.n2761 0.110519
R13990 VDD.n2901 VDD.n2490 0.110215
R13991 VDD.n3616 VDD.n3615 0.109875
R13992 VDD.n3943 VDD.n3942 0.109094
R13993 VDD.n1491 VDD.n1372 0.108934
R13994 VDD.n1492 VDD.n1491 0.108934
R13995 VDD.n1492 VDD.n1361 0.108934
R13996 VDD.n1507 VDD.n1361 0.108934
R13997 VDD.n1508 VDD.n1507 0.108934
R13998 VDD.n1508 VDD.n1350 0.108934
R13999 VDD.n1522 VDD.n1350 0.108934
R14000 VDD.n1523 VDD.n1522 0.108934
R14001 VDD.n1523 VDD.n1344 0.108934
R14002 VDD.n1535 VDD.n1344 0.108934
R14003 VDD.n1536 VDD.n1535 0.108934
R14004 VDD.n1536 VDD.n1333 0.108934
R14005 VDD.n1551 VDD.n1333 0.108934
R14006 VDD.n1552 VDD.n1551 0.108934
R14007 VDD.n1552 VDD.n1321 0.108934
R14008 VDD.n1566 VDD.n1321 0.108934
R14009 VDD.n1567 VDD.n1566 0.108934
R14010 VDD.n1567 VDD.n1310 0.108934
R14011 VDD.n1582 VDD.n1310 0.108934
R14012 VDD.n1583 VDD.n1582 0.108934
R14013 VDD.n1583 VDD.n1299 0.108934
R14014 VDD.n1597 VDD.n1299 0.108934
R14015 VDD.n1598 VDD.n1597 0.108934
R14016 VDD.n1598 VDD.n1293 0.108934
R14017 VDD.n1610 VDD.n1293 0.108934
R14018 VDD.n1611 VDD.n1610 0.108934
R14019 VDD.n1611 VDD.n1282 0.108934
R14020 VDD.n1810 VDD.n1282 0.108934
R14021 VDD.n1810 VDD.n1809 0.108934
R14022 VDD.n1809 VDD.n1283 0.108934
R14023 VDD.n1632 VDD.n1283 0.108934
R14024 VDD.n1795 VDD.n1632 0.108934
R14025 VDD.n1795 VDD.n1794 0.108934
R14026 VDD.n1794 VDD.n1633 0.108934
R14027 VDD.n1781 VDD.n1633 0.108934
R14028 VDD.n1781 VDD.n1780 0.108934
R14029 VDD.n1780 VDD.n1648 0.108934
R14030 VDD.n1665 VDD.n1648 0.108934
R14031 VDD.n1766 VDD.n1665 0.108934
R14032 VDD.n1766 VDD.n1765 0.108934
R14033 VDD.n1765 VDD.n1666 0.108934
R14034 VDD.n1682 VDD.n1666 0.108934
R14035 VDD.n1751 VDD.n1682 0.108934
R14036 VDD.n1751 VDD.n1750 0.108934
R14037 VDD.n1750 VDD.n1683 0.108934
R14038 VDD.n1699 VDD.n1683 0.108934
R14039 VDD.n1736 VDD.n1699 0.108934
R14040 VDD.n1736 VDD.n1735 0.108934
R14041 VDD.n1735 VDD.n1700 0.108934
R14042 VDD.n1700 VDD.n1048 0.108934
R14043 VDD.n1879 VDD.n1048 0.108934
R14044 VDD.n1879 VDD.n1878 0.108934
R14045 VDD.n1878 VDD.n1049 0.108934
R14046 VDD.n1868 VDD.n1049 0.108934
R14047 VDD.n1868 VDD.n1867 0.108934
R14048 VDD.n1851 VDD.n1056 0.108934
R14049 VDD.n1851 VDD.n1850 0.108934
R14050 VDD.n1850 VDD.n1065 0.108934
R14051 VDD.n1842 VDD.n1065 0.108934
R14052 VDD.n1842 VDD.n1841 0.108934
R14053 VDD.n1841 VDD.n1071 0.108934
R14054 VDD.n1831 VDD.n1071 0.108934
R14055 VDD.n1831 VDD.n1830 0.108934
R14056 VDD.n1830 VDD.n1078 0.108934
R14057 VDD.n1822 VDD.n1078 0.108934
R14058 VDD.n1822 VDD.n1821 0.108934
R14059 VDD.n1821 VDD.n1084 0.108934
R14060 VDD.n1273 VDD.n1084 0.108934
R14061 VDD.n1273 VDD.n1272 0.108934
R14062 VDD.n1271 VDD.n1090 0.108934
R14063 VDD.n1266 VDD.n1090 0.108934
R14064 VDD.n1266 VDD.n1265 0.108934
R14065 VDD.n1265 VDD.n1092 0.108934
R14066 VDD.n1257 VDD.n1092 0.108934
R14067 VDD.n1257 VDD.n1256 0.108934
R14068 VDD.n1256 VDD.n1099 0.108934
R14069 VDD.n1248 VDD.n1099 0.108934
R14070 VDD.n1248 VDD.n1247 0.108934
R14071 VDD.n1247 VDD.n1105 0.108934
R14072 VDD.n1111 VDD.n1105 0.108934
R14073 VDD.n1115 VDD.n1111 0.108934
R14074 VDD.n1232 VDD.n1115 0.108934
R14075 VDD.n1232 VDD.n1231 0.108934
R14076 VDD.n1231 VDD.n1116 0.108934
R14077 VDD.n1223 VDD.n1116 0.108934
R14078 VDD.n1223 VDD.n1222 0.108934
R14079 VDD.n1222 VDD.n1122 0.108934
R14080 VDD.n1214 VDD.n1122 0.108934
R14081 VDD.n1214 VDD.n1213 0.108934
R14082 VDD.n1213 VDD.n1128 0.108934
R14083 VDD.n1205 VDD.n1128 0.108934
R14084 VDD.n1205 VDD.n1204 0.108934
R14085 VDD.n1204 VDD.n1134 0.108934
R14086 VDD.n1196 VDD.n1134 0.108934
R14087 VDD.n1196 VDD.n1195 0.108934
R14088 VDD.n1195 VDD.n1140 0.108934
R14089 VDD.n1146 VDD.n1140 0.108934
R14090 VDD.n1150 VDD.n1146 0.108934
R14091 VDD.n1180 VDD.n1150 0.108934
R14092 VDD.n1180 VDD.n1179 0.108934
R14093 VDD.n1179 VDD.n1151 0.108934
R14094 VDD.n1171 VDD.n1151 0.108934
R14095 VDD.n1171 VDD.n1170 0.108934
R14096 VDD.n1170 VDD.n1157 0.108934
R14097 VDD.n1162 VDD.n1157 0.108934
R14098 VDD.n1162 VDD.n998 0.108934
R14099 VDD.n4584 VDD.n998 0.108934
R14100 VDD.n4585 VDD.n4584 0.108934
R14101 VDD.n4586 VDD.n4585 0.108934
R14102 VDD.n4586 VDD.n991 0.108934
R14103 VDD.n4596 VDD.n991 0.108934
R14104 VDD.n4597 VDD.n4596 0.108934
R14105 VDD.n4597 VDD.n984 0.108934
R14106 VDD.n4607 VDD.n984 0.108934
R14107 VDD.n4608 VDD.n4607 0.108934
R14108 VDD.n4609 VDD.n4608 0.108934
R14109 VDD.n4609 VDD.n977 0.108934
R14110 VDD.n4620 VDD.n977 0.108934
R14111 VDD.n4621 VDD.n4620 0.108934
R14112 VDD.n4622 VDD.n4621 0.108934
R14113 VDD.n4622 VDD.n970 0.108934
R14114 VDD.n4633 VDD.n970 0.108934
R14115 VDD.n4634 VDD.n4633 0.108934
R14116 VDD.n4635 VDD.n4634 0.108934
R14117 VDD.n4635 VDD.n963 0.108934
R14118 VDD.n4646 VDD.n963 0.108934
R14119 VDD.n4647 VDD.n4646 0.108934
R14120 VDD.n4648 VDD.n4647 0.108934
R14121 VDD.n4648 VDD.n956 0.108934
R14122 VDD.n4658 VDD.n956 0.108934
R14123 VDD.n4659 VDD.n4658 0.108934
R14124 VDD.n4659 VDD.n949 0.108934
R14125 VDD.n4669 VDD.n949 0.108934
R14126 VDD.n4670 VDD.n4669 0.108934
R14127 VDD.n4671 VDD.n4670 0.108934
R14128 VDD.n4671 VDD.n942 0.108934
R14129 VDD.n4682 VDD.n942 0.108934
R14130 VDD.n4683 VDD.n4682 0.108934
R14131 VDD.n4684 VDD.n4683 0.108934
R14132 VDD.n4684 VDD.n935 0.108934
R14133 VDD.n4695 VDD.n935 0.108934
R14134 VDD.n4696 VDD.n4695 0.108934
R14135 VDD.n4697 VDD.n4696 0.108934
R14136 VDD.n4697 VDD.n928 0.108934
R14137 VDD.n4707 VDD.n928 0.108934
R14138 VDD.n4708 VDD.n4707 0.108934
R14139 VDD.n4708 VDD.n917 0.108934
R14140 VDD.n4726 VDD.n4725 0.108934
R14141 VDD.n4727 VDD.n4726 0.108934
R14142 VDD.n4727 VDD.n910 0.108934
R14143 VDD.n4738 VDD.n910 0.108934
R14144 VDD.n4739 VDD.n4738 0.108934
R14145 VDD.n4740 VDD.n4739 0.108934
R14146 VDD.n4740 VDD.n903 0.108934
R14147 VDD.n4750 VDD.n903 0.108934
R14148 VDD.n4751 VDD.n4750 0.108934
R14149 VDD.n4751 VDD.n896 0.108934
R14150 VDD.n4762 VDD.n896 0.108934
R14151 VDD.n4763 VDD.n4762 0.108934
R14152 VDD.n4764 VDD.n4763 0.108934
R14153 VDD.n4764 VDD.n889 0.108934
R14154 VDD.n4775 VDD.n889 0.108934
R14155 VDD.n4776 VDD.n4775 0.108934
R14156 VDD.n4777 VDD.n4776 0.108934
R14157 VDD.n4777 VDD.n882 0.108934
R14158 VDD.n4788 VDD.n882 0.108934
R14159 VDD.n4789 VDD.n4788 0.108934
R14160 VDD.n4790 VDD.n4789 0.108934
R14161 VDD.n4790 VDD.n875 0.108934
R14162 VDD.n4800 VDD.n875 0.108934
R14163 VDD.n4801 VDD.n4800 0.108934
R14164 VDD.n4801 VDD.n869 0.108934
R14165 VDD.n4813 VDD.n869 0.108934
R14166 VDD.n4814 VDD.n4813 0.108934
R14167 VDD.n4815 VDD.n4814 0.108934
R14168 VDD.n4815 VDD.n862 0.108934
R14169 VDD.n4826 VDD.n862 0.108934
R14170 VDD.n4827 VDD.n4826 0.108934
R14171 VDD.n4828 VDD.n4827 0.108934
R14172 VDD.n4828 VDD.n855 0.108934
R14173 VDD.n4839 VDD.n855 0.108934
R14174 VDD.n4840 VDD.n4839 0.108934
R14175 VDD.n4841 VDD.n4840 0.108934
R14176 VDD.n4841 VDD.n848 0.108934
R14177 VDD.n4852 VDD.n848 0.108934
R14178 VDD.n4853 VDD.n4852 0.108934
R14179 VDD.n4854 VDD.n4853 0.108934
R14180 VDD.n4854 VDD.n841 0.108934
R14181 VDD.n4864 VDD.n841 0.108934
R14182 VDD.n4865 VDD.n4864 0.108934
R14183 VDD.n4865 VDD.n834 0.108934
R14184 VDD.n4876 VDD.n834 0.108934
R14185 VDD.n4877 VDD.n4876 0.108934
R14186 VDD.n4878 VDD.n4877 0.108934
R14187 VDD.n4878 VDD.n827 0.108934
R14188 VDD.n4889 VDD.n827 0.108934
R14189 VDD.n4890 VDD.n4889 0.108934
R14190 VDD.n4891 VDD.n4890 0.108934
R14191 VDD.n4891 VDD.n820 0.108934
R14192 VDD.n4902 VDD.n820 0.108934
R14193 VDD.n4903 VDD.n4902 0.108934
R14194 VDD.n4904 VDD.n4903 0.108934
R14195 VDD.n4904 VDD.n813 0.108934
R14196 VDD.n4914 VDD.n813 0.108934
R14197 VDD.n4915 VDD.n4914 0.108934
R14198 VDD.n4915 VDD.n807 0.108934
R14199 VDD.n4927 VDD.n807 0.108934
R14200 VDD.n4928 VDD.n4927 0.108934
R14201 VDD.n4929 VDD.n4928 0.108934
R14202 VDD.n4929 VDD.n800 0.108934
R14203 VDD.n4940 VDD.n800 0.108934
R14204 VDD.n4941 VDD.n4940 0.108934
R14205 VDD.n4942 VDD.n4941 0.108934
R14206 VDD.n4942 VDD.n793 0.108934
R14207 VDD.n4953 VDD.n793 0.108934
R14208 VDD.n4954 VDD.n4953 0.108934
R14209 VDD.n4955 VDD.n4954 0.108934
R14210 VDD.n4955 VDD.n786 0.108934
R14211 VDD.n4966 VDD.n786 0.108934
R14212 VDD.n4967 VDD.n4966 0.108934
R14213 VDD.n4968 VDD.n4967 0.108934
R14214 VDD.n4968 VDD.n779 0.108934
R14215 VDD.n4978 VDD.n779 0.108934
R14216 VDD.n4979 VDD.n4978 0.108934
R14217 VDD.n4979 VDD.n772 0.108934
R14218 VDD.n4990 VDD.n772 0.108934
R14219 VDD.n4991 VDD.n4990 0.108934
R14220 VDD.n4992 VDD.n4991 0.108934
R14221 VDD.n4992 VDD.n765 0.108934
R14222 VDD.n5003 VDD.n765 0.108934
R14223 VDD.n5004 VDD.n5003 0.108934
R14224 VDD.n5005 VDD.n5004 0.108934
R14225 VDD.n5005 VDD.n758 0.108934
R14226 VDD.n5016 VDD.n758 0.108934
R14227 VDD.n5017 VDD.n5016 0.108934
R14228 VDD.n5018 VDD.n5017 0.108934
R14229 VDD.n5018 VDD.n751 0.108934
R14230 VDD.n5028 VDD.n751 0.108934
R14231 VDD.n5029 VDD.n5028 0.108934
R14232 VDD.n5029 VDD.n745 0.108934
R14233 VDD.n5041 VDD.n745 0.108934
R14234 VDD.n5042 VDD.n5041 0.108934
R14235 VDD.n5043 VDD.n5042 0.108934
R14236 VDD.n5043 VDD.n738 0.108934
R14237 VDD.n5054 VDD.n738 0.108934
R14238 VDD.n5055 VDD.n5054 0.108934
R14239 VDD.n5056 VDD.n5055 0.108934
R14240 VDD.n5056 VDD.n731 0.108934
R14241 VDD.n5067 VDD.n731 0.108934
R14242 VDD.n5068 VDD.n5067 0.108934
R14243 VDD.n5069 VDD.n5068 0.108934
R14244 VDD.n5069 VDD.n724 0.108934
R14245 VDD.n5080 VDD.n724 0.108934
R14246 VDD.n5081 VDD.n5080 0.108934
R14247 VDD.n5082 VDD.n5081 0.108934
R14248 VDD.n5082 VDD.n717 0.108934
R14249 VDD.n5092 VDD.n717 0.108934
R14250 VDD.n5093 VDD.n5092 0.108934
R14251 VDD.n5093 VDD.n710 0.108934
R14252 VDD.n5104 VDD.n710 0.108934
R14253 VDD.n5105 VDD.n5104 0.108934
R14254 VDD.n5106 VDD.n5105 0.108934
R14255 VDD.n5106 VDD.n703 0.108934
R14256 VDD.n5117 VDD.n703 0.108934
R14257 VDD.n5118 VDD.n5117 0.108934
R14258 VDD.n5119 VDD.n5118 0.108934
R14259 VDD.n5119 VDD.n696 0.108934
R14260 VDD.n5130 VDD.n696 0.108934
R14261 VDD.n5131 VDD.n5130 0.108934
R14262 VDD.n5132 VDD.n5131 0.108934
R14263 VDD.n5132 VDD.n689 0.108934
R14264 VDD.n5142 VDD.n689 0.108934
R14265 VDD.n5143 VDD.n5142 0.108934
R14266 VDD.n5143 VDD.n682 0.108934
R14267 VDD.n5155 VDD.n682 0.108934
R14268 VDD.n5156 VDD.n5155 0.108934
R14269 VDD.n5454 VDD.n276 0.108934
R14270 VDD.n299 VDD.n276 0.108934
R14271 VDD.n5435 VDD.n299 0.108934
R14272 VDD.n5435 VDD.n5434 0.108934
R14273 VDD.n5434 VDD.n300 0.108934
R14274 VDD.n303 VDD.n300 0.108934
R14275 VDD.n5424 VDD.n303 0.108934
R14276 VDD.n5424 VDD.n5423 0.108934
R14277 VDD.n5423 VDD.n304 0.108934
R14278 VDD.n307 VDD.n304 0.108934
R14279 VDD.n5412 VDD.n307 0.108934
R14280 VDD.n5412 VDD.n5411 0.108934
R14281 VDD.n5411 VDD.n308 0.108934
R14282 VDD.n311 VDD.n308 0.108934
R14283 VDD.n5400 VDD.n311 0.108934
R14284 VDD.n5400 VDD.n5399 0.108934
R14285 VDD.n5399 VDD.n312 0.108934
R14286 VDD.n5392 VDD.n312 0.108934
R14287 VDD.n5392 VDD.n5391 0.108934
R14288 VDD.n5391 VDD.n318 0.108934
R14289 VDD.n321 VDD.n318 0.108934
R14290 VDD.n5380 VDD.n321 0.108934
R14291 VDD.n5380 VDD.n5379 0.108934
R14292 VDD.n5379 VDD.n322 0.108934
R14293 VDD.n325 VDD.n322 0.108934
R14294 VDD.n5368 VDD.n325 0.108934
R14295 VDD.n5368 VDD.n5367 0.108934
R14296 VDD.n5367 VDD.n326 0.108934
R14297 VDD.n335 VDD.n326 0.108934
R14298 VDD.n5357 VDD.n335 0.108934
R14299 VDD.n5357 VDD.n5356 0.108934
R14300 VDD.n5356 VDD.n336 0.108934
R14301 VDD.n5346 VDD.n336 0.108934
R14302 VDD.n5346 VDD.n5345 0.108934
R14303 VDD.n5345 VDD.n343 0.108934
R14304 VDD.n351 VDD.n343 0.108934
R14305 VDD.n5335 VDD.n351 0.108934
R14306 VDD.n5335 VDD.n5334 0.108934
R14307 VDD.n5334 VDD.n352 0.108934
R14308 VDD.n360 VDD.n352 0.108934
R14309 VDD.n5324 VDD.n360 0.108934
R14310 VDD.n5324 VDD.n5323 0.108934
R14311 VDD.n5323 VDD.n361 0.108934
R14312 VDD.n369 VDD.n361 0.108934
R14313 VDD.n5313 VDD.n369 0.108934
R14314 VDD.n5313 VDD.n5312 0.108934
R14315 VDD.n5312 VDD.n370 0.108934
R14316 VDD.n378 VDD.n370 0.108934
R14317 VDD.n5302 VDD.n378 0.108934
R14318 VDD.n5302 VDD.n5301 0.108934
R14319 VDD.n5301 VDD.n379 0.108934
R14320 VDD.n390 VDD.n379 0.108934
R14321 VDD.n5291 VDD.n390 0.108934
R14322 VDD.n5291 VDD.n5290 0.108934
R14323 VDD.n5290 VDD.n391 0.108934
R14324 VDD.n453 VDD.n391 0.108934
R14325 VDD.n453 VDD.n449 0.108934
R14326 VDD.n461 VDD.n449 0.108934
R14327 VDD.n462 VDD.n461 0.108934
R14328 VDD.n462 VDD.n445 0.108934
R14329 VDD.n471 VDD.n445 0.108934
R14330 VDD.n472 VDD.n471 0.108934
R14331 VDD.n472 VDD.n441 0.108934
R14332 VDD.n480 VDD.n441 0.108934
R14333 VDD.n481 VDD.n480 0.108934
R14334 VDD.n481 VDD.n437 0.108934
R14335 VDD.n492 VDD.n437 0.108934
R14336 VDD.n493 VDD.n492 0.108934
R14337 VDD.n493 VDD.n433 0.108934
R14338 VDD.n502 VDD.n433 0.108934
R14339 VDD.n503 VDD.n502 0.108934
R14340 VDD.n503 VDD.n429 0.108934
R14341 VDD.n511 VDD.n429 0.108934
R14342 VDD.n512 VDD.n511 0.108934
R14343 VDD.n512 VDD.n425 0.108934
R14344 VDD.n521 VDD.n425 0.108934
R14345 VDD.n522 VDD.n521 0.108934
R14346 VDD.n522 VDD.n421 0.108934
R14347 VDD.n530 VDD.n421 0.108934
R14348 VDD.n531 VDD.n530 0.108934
R14349 VDD.n531 VDD.n417 0.108934
R14350 VDD.n541 VDD.n417 0.108934
R14351 VDD.n542 VDD.n541 0.108934
R14352 VDD.n542 VDD.n413 0.108934
R14353 VDD.n552 VDD.n413 0.108934
R14354 VDD.n553 VDD.n552 0.108934
R14355 VDD.n553 VDD.n409 0.108934
R14356 VDD.n561 VDD.n409 0.108934
R14357 VDD.n562 VDD.n561 0.108934
R14358 VDD.n562 VDD.n405 0.108934
R14359 VDD.n571 VDD.n405 0.108934
R14360 VDD.n572 VDD.n571 0.108934
R14361 VDD.n572 VDD.n401 0.108934
R14362 VDD.n581 VDD.n401 0.108934
R14363 VDD.n582 VDD.n581 0.108934
R14364 VDD.n5280 VDD.n582 0.108934
R14365 VDD.n5280 VDD.n5279 0.108934
R14366 VDD.n5279 VDD.n583 0.108934
R14367 VDD.n591 VDD.n583 0.108934
R14368 VDD.n5269 VDD.n591 0.108934
R14369 VDD.n5269 VDD.n5268 0.108934
R14370 VDD.n5268 VDD.n592 0.108934
R14371 VDD.n603 VDD.n592 0.108934
R14372 VDD.n5258 VDD.n603 0.108934
R14373 VDD.n5258 VDD.n5257 0.108934
R14374 VDD.n5257 VDD.n604 0.108934
R14375 VDD.n612 VDD.n604 0.108934
R14376 VDD.n5247 VDD.n612 0.108934
R14377 VDD.n5247 VDD.n5246 0.108934
R14378 VDD.n5246 VDD.n613 0.108934
R14379 VDD.n621 VDD.n613 0.108934
R14380 VDD.n5236 VDD.n621 0.108934
R14381 VDD.n5236 VDD.n5235 0.108934
R14382 VDD.n5235 VDD.n622 0.108934
R14383 VDD.n630 VDD.n622 0.108934
R14384 VDD.n5225 VDD.n630 0.108934
R14385 VDD.n5225 VDD.n5224 0.108934
R14386 VDD.n5224 VDD.n631 0.108934
R14387 VDD.n5214 VDD.n631 0.108934
R14388 VDD.n5214 VDD.n5213 0.108934
R14389 VDD.n5213 VDD.n638 0.108934
R14390 VDD.n646 VDD.n638 0.108934
R14391 VDD.n5203 VDD.n646 0.108934
R14392 VDD.n5203 VDD.n5202 0.108934
R14393 VDD.n5202 VDD.n647 0.108934
R14394 VDD.n655 VDD.n647 0.108934
R14395 VDD.n5192 VDD.n655 0.108934
R14396 VDD.n5192 VDD.n5191 0.108934
R14397 VDD.n5191 VDD.n656 0.108934
R14398 VDD.n664 VDD.n656 0.108934
R14399 VDD.n5181 VDD.n664 0.108934
R14400 VDD.n5181 VDD.n5180 0.108934
R14401 VDD.n5180 VDD.n665 0.108934
R14402 VDD.n673 VDD.n665 0.108934
R14403 VDD.n5169 VDD.n673 0.108934
R14404 VDD.n5169 VDD.n5168 0.108934
R14405 VDD.n5168 VDD.n674 0.108934
R14406 VDD.n4291 VDD.n2363 0.108934
R14407 VDD.n4281 VDD.n2363 0.108934
R14408 VDD.n4281 VDD.n4280 0.108934
R14409 VDD.n4280 VDD.n2372 0.108934
R14410 VDD.n2380 VDD.n2372 0.108934
R14411 VDD.n4270 VDD.n2380 0.108934
R14412 VDD.n4270 VDD.n4269 0.108934
R14413 VDD.n4269 VDD.n2381 0.108934
R14414 VDD.n2389 VDD.n2381 0.108934
R14415 VDD.n4259 VDD.n2389 0.108934
R14416 VDD.n4259 VDD.n4258 0.108934
R14417 VDD.n4258 VDD.n2390 0.108934
R14418 VDD.n2398 VDD.n2390 0.108934
R14419 VDD.n4248 VDD.n2398 0.108934
R14420 VDD.n4248 VDD.n4247 0.108934
R14421 VDD.n4247 VDD.n2399 0.108934
R14422 VDD.n2406 VDD.n2399 0.108934
R14423 VDD.n4236 VDD.n2406 0.108934
R14424 VDD.n4236 VDD.n4235 0.108934
R14425 VDD.n4235 VDD.n2407 0.108934
R14426 VDD.n2418 VDD.n2407 0.108934
R14427 VDD.n4225 VDD.n2418 0.108934
R14428 VDD.n4225 VDD.n4224 0.108934
R14429 VDD.n4224 VDD.n2419 0.108934
R14430 VDD.n2427 VDD.n2419 0.108934
R14431 VDD.n4214 VDD.n2427 0.108934
R14432 VDD.n4214 VDD.n4213 0.108934
R14433 VDD.n4213 VDD.n2428 0.108934
R14434 VDD.n2436 VDD.n2428 0.108934
R14435 VDD.n4203 VDD.n2436 0.108934
R14436 VDD.n4203 VDD.n4202 0.108934
R14437 VDD.n4202 VDD.n2437 0.108934
R14438 VDD.n4088 VDD.n2437 0.108934
R14439 VDD.n4089 VDD.n4088 0.108934
R14440 VDD.n4089 VDD.n4079 0.108934
R14441 VDD.n4101 VDD.n4079 0.108934
R14442 VDD.n4102 VDD.n4101 0.108934
R14443 VDD.n4103 VDD.n4102 0.108934
R14444 VDD.n4103 VDD.n4072 0.108934
R14445 VDD.n4114 VDD.n4072 0.108934
R14446 VDD.n4115 VDD.n4114 0.108934
R14447 VDD.n4116 VDD.n4115 0.108934
R14448 VDD.n4116 VDD.n4065 0.108934
R14449 VDD.n4128 VDD.n4065 0.108934
R14450 VDD.n4129 VDD.n4128 0.108934
R14451 VDD.n4130 VDD.n4129 0.108934
R14452 VDD.n4130 VDD.n4059 0.108934
R14453 VDD.n4140 VDD.n4059 0.108934
R14454 VDD.n4141 VDD.n4140 0.108934
R14455 VDD.n4141 VDD.n4052 0.108934
R14456 VDD.n4152 VDD.n4052 0.108934
R14457 VDD.n4153 VDD.n4152 0.108934
R14458 VDD.n4154 VDD.n4153 0.108934
R14459 VDD.n4154 VDD.n4045 0.108934
R14460 VDD.n4165 VDD.n4045 0.108934
R14461 VDD.n4166 VDD.n4165 0.108934
R14462 VDD.n4167 VDD.n4166 0.108934
R14463 VDD.n4167 VDD.n4038 0.108934
R14464 VDD.n4178 VDD.n4038 0.108934
R14465 VDD.n4179 VDD.n4178 0.108934
R14466 VDD.n4180 VDD.n4179 0.108934
R14467 VDD.n4180 VDD.n4030 0.108934
R14468 VDD.n4191 VDD.n4030 0.108934
R14469 VDD.n4192 VDD.n4191 0.108934
R14470 VDD.n4192 VDD.n275 0.108934
R14471 VDD.n5455 VDD.n275 0.108934
R14472 VDD.n1465 VDD.n1464 0.108934
R14473 VDD.n1464 VDD.n1402 0.108934
R14474 VDD.n1454 VDD.n1402 0.108934
R14475 VDD.n1454 VDD.n1453 0.108934
R14476 VDD.n1453 VDD.n1408 0.108934
R14477 VDD.n1413 VDD.n1408 0.108934
R14478 VDD.n1436 VDD.n1413 0.108934
R14479 VDD.n1436 VDD.n1435 0.108934
R14480 VDD.n1435 VDD.n1414 0.108934
R14481 VDD.n1419 VDD.n1414 0.108934
R14482 VDD.n1419 VDD.n1418 0.108934
R14483 VDD.n1418 VDD.n1027 0.108934
R14484 VDD.n1898 VDD.n1027 0.108934
R14485 VDD.n1899 VDD.n1898 0.108934
R14486 VDD.n1900 VDD.n1899 0.108934
R14487 VDD.n1901 VDD.n1900 0.108934
R14488 VDD.n1901 VDD.n1023 0.108934
R14489 VDD.n4560 VDD.n1023 0.108934
R14490 VDD.n4560 VDD.n4559 0.108934
R14491 VDD.n4559 VDD.n1024 0.108934
R14492 VDD.n1932 VDD.n1024 0.108934
R14493 VDD.n1932 VDD.n1928 0.108934
R14494 VDD.n4541 VDD.n1928 0.108934
R14495 VDD.n4541 VDD.n4540 0.108934
R14496 VDD.n4540 VDD.n1929 0.108934
R14497 VDD.n1967 VDD.n1929 0.108934
R14498 VDD.n1973 VDD.n1967 0.108934
R14499 VDD.n1974 VDD.n1973 0.108934
R14500 VDD.n4516 VDD.n1974 0.108934
R14501 VDD.n4516 VDD.n4515 0.108934
R14502 VDD.n4515 VDD.n1975 0.108934
R14503 VDD.n2004 VDD.n1975 0.108934
R14504 VDD.n2004 VDD.n2000 0.108934
R14505 VDD.n4497 VDD.n2000 0.108934
R14506 VDD.n4497 VDD.n4496 0.108934
R14507 VDD.n4496 VDD.n2001 0.108934
R14508 VDD.n2037 VDD.n2001 0.108934
R14509 VDD.n2037 VDD.n2033 0.108934
R14510 VDD.n4478 VDD.n2033 0.108934
R14511 VDD.n4478 VDD.n4477 0.108934
R14512 VDD.n4477 VDD.n2034 0.108934
R14513 VDD.n2084 VDD.n2034 0.108934
R14514 VDD.n2084 VDD.n2062 0.108934
R14515 VDD.n4459 VDD.n2062 0.108934
R14516 VDD.n4459 VDD.n4458 0.108934
R14517 VDD.n4458 VDD.n2063 0.108934
R14518 VDD.n4444 VDD.n2063 0.108934
R14519 VDD.n4444 VDD.n4443 0.108934
R14520 VDD.n4443 VDD.n2081 0.108934
R14521 VDD.n2121 VDD.n2081 0.108934
R14522 VDD.n2121 VDD.n2117 0.108934
R14523 VDD.n4425 VDD.n2117 0.108934
R14524 VDD.n4425 VDD.n4424 0.108934
R14525 VDD.n4424 VDD.n2118 0.108934
R14526 VDD.n2152 VDD.n2118 0.108934
R14527 VDD.n2152 VDD.n2148 0.108934
R14528 VDD.n4406 VDD.n2148 0.108934
R14529 VDD.n4406 VDD.n4405 0.108934
R14530 VDD.n4405 VDD.n2149 0.108934
R14531 VDD.n2188 VDD.n2149 0.108934
R14532 VDD.n2194 VDD.n2188 0.108934
R14533 VDD.n2195 VDD.n2194 0.108934
R14534 VDD.n4381 VDD.n2195 0.108934
R14535 VDD.n4381 VDD.n4380 0.108934
R14536 VDD.n4380 VDD.n2196 0.108934
R14537 VDD.n2225 VDD.n2196 0.108934
R14538 VDD.n2225 VDD.n2221 0.108934
R14539 VDD.n4362 VDD.n2221 0.108934
R14540 VDD.n4362 VDD.n4361 0.108934
R14541 VDD.n4361 VDD.n2222 0.108934
R14542 VDD.n2362 VDD.n2222 0.108934
R14543 VDD.n2902 VDD.n2490 0.10877
R14544 VDD.n8398 VDD.n8290 0.107703
R14545 VDD.n7543 VDD.n7435 0.107703
R14546 VDD.n6689 VDD.n6581 0.107703
R14547 VDD.n5834 VDD.n5726 0.107703
R14548 VDD.n3602 VDD.n3601 0.0995999
R14549 VDD.n3567 VDD.n3566 0.0995999
R14550 VDD.n3269 VDD.n3268 0.0995999
R14551 VDD.n3158 VDD.n3157 0.0995999
R14552 VDD.n3977 VDD.n3976 0.0980399
R14553 VDD.n2454 VDD.n2453 0.0932536
R14554 VDD.n9027 VDD.n9026 0.0926226
R14555 VDD.n8172 VDD.n8171 0.0926226
R14556 VDD.n7318 VDD.n7317 0.0926226
R14557 VDD.n6463 VDD.n6462 0.0926226
R14558 VDD.n5654 VDD 0.0926053
R14559 VDD.n7363 VDD 0.0926053
R14560 VDD.n3617 VDD.n2507 0.0923441
R14561 VDD.n2627 VDD.n2594 0.0905941
R14562 VDD.n2627 VDD.n2593 0.0897616
R14563 VDD.n5511 VDD.n5510 0.0895625
R14564 VDD.n3115 VDD.n3107 0.0861908
R14565 VDD.n2908 VDD.n2907 0.0856562
R14566 VDD.n2561 VDD.n2535 0.0825312
R14567 VDD.n2551 VDD.n2550 0.0825312
R14568 VDD.n3115 VDD.n3108 0.0777426
R14569 VDD.n9028 VDD.n9027 0.0745132
R14570 VDD.n8173 VDD.n8172 0.0745132
R14571 VDD.n7319 VDD.n7318 0.0745132
R14572 VDD.n6464 VDD.n6463 0.0745132
R14573 VDD VDD.n3116 0.0739375
R14574 VDD.n3369 VDD.n3368 0.0736942
R14575 VDD.n3630 VDD.n3629 0.0736373
R14576 VDD.n5401 VDD.n310 0.0728164
R14577 VDD.n341 VDD.n337 0.0728164
R14578 VDD.n5303 VDD.n377 0.0728164
R14579 VDD.n483 VDD.n438 0.0728164
R14580 VDD.n544 VDD.n543 0.0728164
R14581 VDD.n5270 VDD.n590 0.0728164
R14582 VDD.n5223 VDD.n5222 0.0728164
R14583 VDD.n5172 VDD.n671 0.0728164
R14584 VDD.n3956 VDD.n3626 0.0717614
R14585 VDD.n4302 VDD.n2340 0.071743
R14586 VDD.n3626 VDD.n3623 0.0711193
R14587 VDD.n3701 VDD.n3677 0.0707228
R14588 VDD.n3935 VDD.n3643 0.0707228
R14589 VDD.n3956 VDD.n3629 0.0703248
R14590 VDD.n1877 VDD.n1876 0.0696892
R14591 VDD.n3772 VDD.n3771 0.0692474
R14592 VDD.n9022 VDD.n9021 0.0688877
R14593 VDD.n8167 VDD.n8166 0.0688877
R14594 VDD.n7313 VDD.n7312 0.0688877
R14595 VDD.n6458 VDD.n6457 0.0688877
R14596 VDD.n1423 VDD.n1420 0.0682249
R14597 VDD.n1972 VDD.n1956 0.0682249
R14598 VDD.n4460 VDD.n2061 0.0682249
R14599 VDD.n2193 VDD.n2177 0.0682249
R14600 VDD.n2943 VDD.n2942 0.0679494
R14601 VDD.n5508 VDD 0.0645625
R14602 VDD.n9021 VDD.n8246 0.0643587
R14603 VDD.n8166 VDD.n7391 0.0643587
R14604 VDD.n7312 VDD.n6537 0.0643587
R14605 VDD.n6457 VDD.n5682 0.0643587
R14606 VDD.n1378 VDD.n1377 0.0638663
R14607 VDD.n1490 VDD.n1489 0.0638663
R14608 VDD.n1568 VDD.n1320 0.0638663
R14609 VDD.n1316 VDD.n1315 0.0638663
R14610 VDD.n1643 VDD.n1642 0.0638663
R14611 VDD.n1782 VDD.n1647 0.0638663
R14612 VDD.n3108 VDD.n2486 0.0636644
R14613 VDD.n3466 VDD.n2693 0.0631347
R14614 VDD.n3411 VDD.n2732 0.0631347
R14615 VDD.n3097 VDD.n3094 0.0631347
R14616 VDD.n3280 VDD.n3089 0.0631347
R14617 VDD.n3426 VDD.n2713 0.0631347
R14618 VDD.n2685 VDD.n2637 0.0631347
R14619 VDD.n3578 VDD.n2683 0.0631347
R14620 VDD.n3449 VDD.n2702 0.0627929
R14621 VDD.n3395 VDD.n2738 0.0627929
R14622 VDD.n104 VDD.n34 0.0608156
R14623 VDD.n5655 VDD 0.060807
R14624 VDD.n7364 VDD 0.060807
R14625 VDD.n3923 VDD.n3920 0.0604712
R14626 VDD.n3651 VDD.n3649 0.0604712
R14627 VDD.n3941 VDD.n3636 0.0604712
R14628 VDD.n2863 VDD.n2798 0.0604712
R14629 VDD.n3762 VDD.n3646 0.0595872
R14630 VDD.n237 VDD.n174 0.0595049
R14631 VDD.n107 VDD.n106 0.0591683
R14632 VDD.n3929 VDD.n3657 0.0591603
R14633 VDD.n2814 VDD.n2796 0.0591603
R14634 VDD.n2451 VDD.n238 0.0589865
R14635 VDD.n3002 VDD.n2897 0.0586853
R14636 VDD.n3356 VDD.n3328 0.0581563
R14637 VDD.n5635 VDD.n5634 0.056838
R14638 VDD.n5636 VDD.n5635 0.056838
R14639 VDD.n5636 VDD.n5613 0.056838
R14640 VDD.n5672 VDD.n5613 0.056838
R14641 VDD.n6483 VDD.n6475 0.056838
R14642 VDD.n6494 VDD.n6475 0.056838
R14643 VDD.n6496 VDD.n6494 0.056838
R14644 VDD.n6496 VDD.n6495 0.056838
R14645 VDD.n7344 VDD.n7343 0.056838
R14646 VDD.n7345 VDD.n7344 0.056838
R14647 VDD.n7345 VDD.n7322 0.056838
R14648 VDD.n7381 VDD.n7322 0.056838
R14649 VDD.n8192 VDD.n8184 0.056838
R14650 VDD.n8203 VDD.n8184 0.056838
R14651 VDD.n8205 VDD.n8203 0.056838
R14652 VDD.n8205 VDD.n8204 0.056838
R14653 VDD VDD.n5507 0.05675
R14654 VDD.n3112 VDD.n3107 0.0566413
R14655 VDD.n3606 VDD.n3605 0.0565323
R14656 VDD.n3575 VDD.n3573 0.0565323
R14657 VDD.n3463 VDD.n3462 0.0565323
R14658 VDD.n2707 VDD.n2705 0.0565323
R14659 VDD.n2727 VDD.n2716 0.0565323
R14660 VDD.n3409 VDD.n3406 0.0565323
R14661 VDD.n2743 VDD.n2741 0.0565323
R14662 VDD.n3296 VDD.n3065 0.0565323
R14663 VDD.n3277 VDD.n3275 0.0565323
R14664 VDD.n3165 VDD.n3164 0.0565323
R14665 VDD.n2890 VDD.n2869 0.0561943
R14666 VDD.n2948 VDD.n2894 0.0558794
R14667 VDD.n57 VDD.n38 0.0547109
R14668 VDD.n5587 VDD.n5586 0.0547109
R14669 VDD.n203 VDD.n202 0.0547109
R14670 VDD VDD.n9029 0.0526991
R14671 VDD.n3979 VDD.n2507 0.0521995
R14672 VDD.n2593 VDD.n2592 0.0521189
R14673 VDD VDD.n7320 0.0517913
R14674 VDD.n2362 VDD.n2359 0.0517048
R14675 VDD.n2594 VDD.n2591 0.0513458
R14676 VDD.n2542 VDD.n2538 0.0493281
R14677 VDD.n3605 VDD.n2643 0.0487198
R14678 VDD.n3573 VDD.n3572 0.0487198
R14679 VDD.n3462 VDD.n3461 0.0487198
R14680 VDD.n3439 VDD.n2707 0.0487198
R14681 VDD.n2727 VDD.n2726 0.0487198
R14682 VDD.n3409 VDD.n3408 0.0487198
R14683 VDD.n3385 VDD.n2743 0.0487198
R14684 VDD.n3275 VDD.n3274 0.0487198
R14685 VDD.n3164 VDD.n3163 0.0487198
R14686 VDD VDD.n6465 0.0482611
R14687 VDD VDD.n8174 0.0482611
R14688 VDD.n3357 VDD.n3356 0.0479088
R14689 VDD.n3047 VDD.n3046 0.0472468
R14690 VDD.n5527 VDD.n161 0.0462851
R14691 VDD.n5631 VDD.n5626 0.0461081
R14692 VDD.n6484 VDD.n6480 0.0461081
R14693 VDD.n7340 VDD.n7335 0.0461081
R14694 VDD.n8193 VDD.n8189 0.0461081
R14695 VDD.n3699 VDD.n3686 0.0459877
R14696 VDD.n39 VDD.n32 0.0459833
R14697 VDD.n5509 VDD.n169 0.0459833
R14698 VDD.n3027 VDD.n2872 0.0457021
R14699 VDD.n3976 VDD.n3617 0.0456313
R14700 VDD.n139 VDD.n27 0.0456006
R14701 VDD.n5538 VDD.n160 0.0455549
R14702 VDD.n5538 VDD.n163 0.0454465
R14703 VDD.n2514 VDD.n2513 0.0454219
R14704 VDD.n2573 VDD.n2531 0.0454219
R14705 VDD.n2563 VDD.n2532 0.0454219
R14706 VDD.n27 VDD.n26 0.0454042
R14707 VDD.n2872 VDD.n2868 0.0453096
R14708 VDD.n3699 VDD.n3698 0.045025
R14709 VDD.n39 VDD.n33 0.0450203
R14710 VDD.n169 VDD.n165 0.0450203
R14711 VDD.n3071 VDD.n3070 0.0448136
R14712 VDD.n5596 VDD.n5527 0.0447244
R14713 VDD.n5505 VDD.n241 0.044241
R14714 VDD.n2666 VDD.n2660 0.0439783
R14715 VDD.n3556 VDD.n3483 0.0439783
R14716 VDD.n3547 VDD.n3484 0.0439783
R14717 VDD.n3258 VDD.n3185 0.0439783
R14718 VDD.n3249 VDD.n3186 0.0439783
R14719 VDD.n3135 VDD.n3129 0.0439783
R14720 VDD.n3772 VDD.n3769 0.0439783
R14721 VDD.n2942 VDD.n2918 0.0439783
R14722 VDD.n72 VDD.n59 0.0439783
R14723 VDD.n5577 VDD.n5576 0.0439783
R14724 VDD.n218 VDD.n205 0.0439783
R14725 VDD.n241 VDD.n238 0.0439172
R14726 VDD.n5632 VDD.n5621 0.0435743
R14727 VDD.n6481 VDD.n6476 0.0435743
R14728 VDD.n7341 VDD.n7330 0.0435743
R14729 VDD.n8190 VDD.n8185 0.0435743
R14730 VDD.n3041 VDD.n2867 0.0434688
R14731 VDD.n3041 VDD.n3040 0.0434688
R14732 VDD.n3040 VDD.n3039 0.0434688
R14733 VDD.n3035 VDD.n3034 0.0434688
R14734 VDD.n3034 VDD.n3033 0.0434688
R14735 VDD.n3033 VDD.n3031 0.0434688
R14736 VDD.n3031 VDD.n3030 0.0434688
R14737 VDD.n3018 VDD.n3017 0.0434688
R14738 VDD.n3017 VDD.n3016 0.0434688
R14739 VDD.n3016 VDD.n3014 0.0434688
R14740 VDD.n3010 VDD.n3009 0.0434688
R14741 VDD.n3009 VDD.n3008 0.0434688
R14742 VDD.n3008 VDD.n3006 0.0434688
R14743 VDD.n146 VDD.n144 0.0434688
R14744 VDD.n146 VDD.n145 0.0434688
R14745 VDD.n145 VDD.n9 0.0434688
R14746 VDD.n152 VDD.n9 0.0434688
R14747 VDD.n157 VDD.n155 0.0434688
R14748 VDD.n158 VDD.n157 0.0434688
R14749 VDD.n159 VDD.n158 0.0434688
R14750 VDD.n5599 VDD.n159 0.0434688
R14751 VDD.n5599 VDD.n5598 0.0434688
R14752 VDD.n5525 VDD.n5523 0.0434688
R14753 VDD.n5523 VDD.n5522 0.0434688
R14754 VDD.n5522 VDD.n5520 0.0434688
R14755 VDD.n5516 VDD.n5515 0.0434688
R14756 VDD.n5515 VDD.n5514 0.0434688
R14757 VDD.n2570 VDD.n2569 0.0434688
R14758 VDD.n2571 VDD.n2532 0.0434688
R14759 VDD.n3329 VDD.n2745 0.0434688
R14760 VDD.n3333 VDD.n3329 0.0434688
R14761 VDD.n3334 VDD.n3333 0.0434688
R14762 VDD.n3335 VDD.n3334 0.0434688
R14763 VDD.n3341 VDD.n3339 0.0434688
R14764 VDD.n3342 VDD.n3341 0.0434688
R14765 VDD.n3344 VDD.n3342 0.0434688
R14766 VDD.n3345 VDD.n3344 0.0434688
R14767 VDD.n3347 VDD.n3345 0.0434688
R14768 VDD.n3326 VDD.n3325 0.0434688
R14769 VDD.n3325 VDD.n3324 0.0434688
R14770 VDD.n3324 VDD.n3322 0.0434688
R14771 VDD.n3322 VDD.n3321 0.0434688
R14772 VDD.n3321 VDD.n3319 0.0434688
R14773 VDD.n3319 VDD.n3318 0.0434688
R14774 VDD.n3318 VDD.n2767 0.0434688
R14775 VDD.n3314 VDD.n2767 0.0434688
R14776 VDD.n3314 VDD.n3313 0.0434688
R14777 VDD.n3313 VDD.n3312 0.0434688
R14778 VDD.n3312 VDD.n2771 0.0434688
R14779 VDD.n3052 VDD.n2771 0.0434688
R14780 VDD.n3053 VDD.n3052 0.0434688
R14781 VDD.n3059 VDD.n3053 0.0434688
R14782 VDD.n4290 VDD.n4289 0.0433094
R14783 VDD.n4239 VDD.n2404 0.0433094
R14784 VDD.n4092 VDD.n4090 0.0433094
R14785 VDD.n4151 VDD.n4150 0.0433094
R14786 VDD.n3449 VDD.n3448 0.0430273
R14787 VDD.n3395 VDD.n3394 0.0430273
R14788 VDD.n3696 VDD.n3680 0.0429751
R14789 VDD.n3807 VDD.n3645 0.0429751
R14790 VDD.n81 VDD.n38 0.042958
R14791 VDD.n108 VDD.n25 0.042958
R14792 VDD.n5588 VDD.n5587 0.042958
R14793 VDD.n202 VDD.n166 0.042958
R14794 VDD.n3302 VDD.n3065 0.0428604
R14795 VDD.n3613 VDD.n2637 0.0426869
R14796 VDD.n3474 VDD.n2683 0.0426869
R14797 VDD.n3470 VDD.n2693 0.0426869
R14798 VDD.n3430 VDD.n2713 0.0426869
R14799 VDD.n3412 VDD.n3411 0.0426869
R14800 VDD.n3176 VDD.n3089 0.0426869
R14801 VDD.n3172 VDD.n3094 0.0426869
R14802 VDD.n3815 VDD.n3761 0.0420568
R14803 VDD.n3718 VDD.n3660 0.0420568
R14804 VDD.n3905 VDD.n3668 0.0420568
R14805 VDD.n2816 VDD.n2806 0.0420568
R14806 VDD.n2574 VDD.n2522 0.0415156
R14807 VDD.n2560 VDD.n2559 0.0415156
R14808 VDD.n2573 VDD.n2572 0.0415156
R14809 VDD VDD.n6526 0.0412609
R14810 VDD VDD.n8235 0.0412609
R14811 VDD.n3500 VDD.n3490 0.0412609
R14812 VDD.n3518 VDD.n3506 0.0412609
R14813 VDD.n3202 VDD.n3192 0.0412609
R14814 VDD.n3220 VDD.n3208 0.0412609
R14815 VDD.n3750 VDD.n3740 0.0412609
R14816 VDD.n3834 VDD.n3833 0.0412609
R14817 VDD.n3848 VDD.n3733 0.0412609
R14818 VDD.n3857 VDD.n3856 0.0412609
R14819 VDD.n3870 VDD.n3705 0.0412609
R14820 VDD.n3888 VDD.n3876 0.0412609
R14821 VDD.n2830 VDD.n2820 0.0412609
R14822 VDD.n2972 VDD.n2962 0.0412609
R14823 VDD.n3039 VDD.n3038 0.041125
R14824 VDD.n5519 VDD.n5516 0.041125
R14825 VDD.n3117 VDD 0.041125
R14826 VDD.n3030 VDD.n3028 0.0403437
R14827 VDD.n5526 VDD.n5525 0.0403437
R14828 VDD.n3373 VDD.n3326 0.0403437
R14829 VDD.n3022 VDD.n2871 0.0398734
R14830 VDD.n2531 VDD.n2524 0.0395625
R14831 VDD.n3592 VDD.n3591 0.0385435
R14832 VDD.n3561 VDD.n3482 0.0385435
R14833 VDD.n3542 VDD.n3485 0.0385435
R14834 VDD.n3263 VDD.n3184 0.0385435
R14835 VDD.n3244 VDD.n3187 0.0385435
R14836 VDD.n3148 VDD.n3147 0.0385435
R14837 VDD.n58 VDD.n57 0.0385435
R14838 VDD.n5586 VDD.n5561 0.0385435
R14839 VDD.n204 VDD.n203 0.0385435
R14840 VDD.n5638 VDD.n5621 0.0385068
R14841 VDD.n5671 VDD 0.0385068
R14842 VDD.n5615 VDD 0.0385068
R14843 VDD.n6492 VDD.n6476 0.0385068
R14844 VDD VDD.n6473 0.0385068
R14845 VDD.n6501 VDD 0.0385068
R14846 VDD.n7347 VDD.n7330 0.0385068
R14847 VDD.n7380 VDD 0.0385068
R14848 VDD.n7324 VDD 0.0385068
R14849 VDD.n8201 VDD.n8185 0.0385068
R14850 VDD VDD.n8182 0.0385068
R14851 VDD.n8210 VDD 0.0385068
R14852 VDD.n5505 VDD.n240 0.0380981
R14853 VDD.n41 VDD.n40 0.0380882
R14854 VDD.n110 VDD.n109 0.0380882
R14855 VDD.n5542 VDD.n5541 0.0380882
R14856 VDD.n186 VDD.n185 0.0380882
R14857 VDD.n3378 VDD.n2745 0.038
R14858 VDD.n3060 VDD.n3059 0.038
R14859 VDD.n2580 VDD.n2512 0.0376094
R14860 VDD.n2523 VDD.n2514 0.0376094
R14861 VDD.n8240 VDD.n5608 0.0364779
R14862 VDD.n6531 VDD.n5610 0.0358522
R14863 VDD.n2526 VDD.n2525 0.0356562
R14864 VDD.n2902 VDD.n2899 0.035222
R14865 VDD.n2995 VDD.n2948 0.0351381
R14866 VDD.n253 VDD.n240 0.0345604
R14867 VDD.n5657 VDD.n5656 0.0343645
R14868 VDD.n7366 VDD.n7365 0.0343645
R14869 VDD.n5605 VDD.n0 0.034112
R14870 VDD.n2906 VDD.n2901 0.0338623
R14871 VDD.n2564 VDD.n2534 0.0337031
R14872 VDD.n2563 VDD.n2562 0.0337031
R14873 VDD.n5676 VDD.n5611 0.033419
R14874 VDD.n7385 VDD.n5609 0.033419
R14875 VDD.n3601 VDD.n2645 0.0331087
R14876 VDD.n3566 VDD.n3481 0.0331087
R14877 VDD.n3537 VDD.n3486 0.0331087
R14878 VDD.n3268 VDD.n3183 0.0331087
R14879 VDD.n3239 VDD.n3188 0.0331087
R14880 VDD.n3157 VDD.n3118 0.0331087
R14881 VDD.n3070 VDD.n3063 0.0330948
R14882 VDD.n3368 VDD.n3367 0.0322427
R14883 VDD.n3004 VDD.n2897 0.0319008
R14884 VDD.n2513 VDD.n2508 0.03175
R14885 VDD.n107 VDD.n24 0.0314198
R14886 VDD.n3716 VDD.n3657 0.0312849
R14887 VDD.n2815 VDD.n2814 0.0312849
R14888 VDD.n2943 VDD.n2892 0.0311134
R14889 VDD.n174 VDD.n168 0.0310804
R14890 VDD.n3813 VDD.n3762 0.0308558
R14891 VDD.n3526 VDD.n3489 0.0303913
R14892 VDD.n3228 VDD.n3191 0.0303913
R14893 VDD.n3727 VDD.n3713 0.0303913
R14894 VDD.n3896 VDD.n3704 0.0303913
R14895 VDD.n3824 VDD.n3756 0.0303913
R14896 VDD.n2840 VDD.n2819 0.0303913
R14897 VDD.n2978 VDD.n2961 0.0303913
R14898 VDD.n3803 VDD.n3802 0.0303633
R14899 VDD.n3921 VDD.n3662 0.0303633
R14900 VDD.n3683 VDD.n3669 0.0303633
R14901 VDD.n2861 VDD.n2803 0.0303633
R14902 VDD.n3025 VDD.n2876 0.0303633
R14903 VDD.n2867 VDD.n2866 0.0301875
R14904 VDD.n144 VDD.n143 0.0301875
R14905 VDD.n5514 VDD.n5511 0.0301875
R14906 VDD.n3932 VDD.n3649 0.0301368
R14907 VDD.n3636 VDD.n3633 0.0301368
R14908 VDD.n3920 VDD.n3652 0.0301368
R14909 VDD.n2798 VDD.n2797 0.0301368
R14910 VDD.n5463 VDD.n259 0.0299811
R14911 VDD.n5462 VDD.n264 0.0299811
R14912 VDD.n101 VDD.n42 0.0297969
R14913 VDD.n135 VDD.n134 0.0297969
R14914 VDD.n5559 VDD.n5558 0.0297969
R14915 VDD.n200 VDD.n187 0.0297969
R14916 VDD.n2542 VDD.n2540 0.0297969
R14917 VDD.n34 VDD.n31 0.0297952
R14918 VDD.n3918 VDD.n3654 0.0291557
R14919 VDD.n3771 VDD.n3634 0.0291557
R14920 VDD.n2808 VDD.n2795 0.0291557
R14921 VDD.n5482 VDD.n256 0.0288019
R14922 VDD.n5466 VDD.n5465 0.0288019
R14923 VDD.n5484 VDD.n5483 0.0288019
R14924 VDD.n9029 VDD.n5608 0.0285752
R14925 VDD.n2452 VDD.n2451 0.0282045
R14926 VDD VDD.n5612 0.0281786
R14927 VDD.n6528 VDD 0.0281786
R14928 VDD VDD.n7321 0.0281786
R14929 VDD.n8237 VDD 0.0281786
R14930 VDD.n7320 VDD.n5610 0.028087
R14931 VDD.n4296 VDD.n4295 0.0280588
R14932 VDD.n3602 VDD.n2644 0.0278438
R14933 VDD.n3568 VDD.n3567 0.0278438
R14934 VDD.n3457 VDD.n3456 0.0278438
R14935 VDD.n3442 VDD.n2706 0.0278438
R14936 VDD.n2722 VDD.n2717 0.0278438
R14937 VDD.n3419 VDD.n3402 0.0278438
R14938 VDD.n3388 VDD.n2742 0.0278438
R14939 VDD.n3285 VDD.n3063 0.0278438
R14940 VDD.n3270 VDD.n3269 0.0278438
R14941 VDD.n3159 VDD.n3158 0.0278438
R14942 VDD.n3532 VDD.n3487 0.0276739
R14943 VDD.n3234 VDD.n3189 0.0276739
R14944 VDD.n5469 VDD.n257 0.0276226
R14945 VDD.n5637 VDD.n5625 0.027527
R14946 VDD.n5625 VDD.n5624 0.027527
R14947 VDD.n6493 VDD.n6474 0.027527
R14948 VDD.n6497 VDD.n6474 0.027527
R14949 VDD.n7346 VDD.n7334 0.027527
R14950 VDD.n7334 VDD.n7333 0.027527
R14951 VDD.n8202 VDD.n8183 0.027527
R14952 VDD.n8206 VDD.n8183 0.027527
R14953 VDD.n4295 VDD.n2341 0.0273817
R14954 VDD.n4297 VDD.n2358 0.0273817
R14955 VDD.n4299 VDD.n2358 0.0273817
R14956 VDD.n154 VDD.n152 0.0270625
R14957 VDD.n5468 VDD.n258 0.0264434
R14958 VDD.n5470 VDD.n5469 0.0264434
R14959 VDD.n6465 VDD.n5611 0.0261883
R14960 VDD.n8174 VDD.n5609 0.0261883
R14961 VDD.n2582 VDD.n2510 0.0258906
R14962 VDD.n2555 VDD.n2536 0.0258906
R14963 VDD.n2554 VDD.n2553 0.0258906
R14964 VDD.n2553 VDD.n2538 0.0258906
R14965 VDD.n2552 VDD.n2535 0.0258906
R14966 VDD.n2552 VDD.n2551 0.0258906
R14967 VDD.n5468 VDD.n5467 0.0252642
R14968 VDD.n5470 VDD.n5466 0.0252642
R14969 VDD.n3531 VDD.n3488 0.0249565
R14970 VDD.n3233 VDD.n3190 0.0249565
R14971 VDD.n3717 VDD.n3715 0.0249565
R14972 VDD.n3722 VDD.n3714 0.0249565
R14973 VDD.n3906 VDD.n3702 0.0249565
R14974 VDD.n3901 VDD.n3703 0.0249565
R14975 VDD.n3814 VDD.n3760 0.0249565
R14976 VDD.n3819 VDD.n3758 0.0249565
R14977 VDD.n2818 VDD.n2817 0.0249565
R14978 VDD.n2845 VDD.n2844 0.0249565
R14979 VDD.n2994 VDD.n2949 0.0249565
R14980 VDD.n2959 VDD.n2955 0.0249565
R14981 VDD.n3339 VDD.n3338 0.0247187
R14982 VDD.n5671 VDD.n5614 0.024466
R14983 VDD.n6499 VDD.n6473 0.024466
R14984 VDD.n7380 VDD.n7323 0.024466
R14985 VDD.n8208 VDD.n8182 0.024466
R14986 VDD.n3929 VDD.n3655 0.0239375
R14987 VDD.n3681 VDD.n3677 0.0239375
R14988 VDD.n3800 VDD.n3646 0.0239375
R14989 VDD.n3935 VDD.n3639 0.0239375
R14990 VDD.n2802 VDD.n2796 0.0239375
R14991 VDD.n2885 VDD.n2869 0.0239375
R14992 VDD.n2911 VDD.n2894 0.0239375
R14993 VDD.n92 VDD.n32 0.0239375
R14994 VDD.n139 VDD.n29 0.0239375
R14995 VDD.n5550 VDD.n160 0.0239375
R14996 VDD.n5509 VDD.n171 0.0239375
R14997 VDD.n2587 VDD.n2586 0.0239375
R14998 VDD.n2530 VDD.n2529 0.0239375
R14999 VDD VDD.n5654 0.0235263
R15000 VDD VDD.n7363 0.0235263
R15001 VDD.n3013 VDD.n3010 0.0231563
R15002 VDD.n3003 VDD.n2909 0.022375
R15003 VDD.n3527 VDD.n3488 0.0222391
R15004 VDD.n3229 VDD.n3190 0.0222391
R15005 VDD.n3721 VDD.n3715 0.0222391
R15006 VDD.n3726 VDD.n3714 0.0222391
R15007 VDD.n3902 VDD.n3702 0.0222391
R15008 VDD.n3897 VDD.n3703 0.0222391
R15009 VDD.n3818 VDD.n3760 0.0222391
R15010 VDD.n3823 VDD.n3758 0.0222391
R15011 VDD.n2846 VDD.n2818 0.0222391
R15012 VDD.n2844 VDD.n2841 0.0222391
R15013 VDD.n2954 VDD.n2949 0.0222391
R15014 VDD.n2960 VDD.n2959 0.0222391
R15015 VDD.n3914 VDD.n3913 0.0219844
R15016 VDD.n3695 VDD.n3691 0.0219844
R15017 VDD.n3796 VDD.n3795 0.0219844
R15018 VDD.n3776 VDD.n3775 0.0219844
R15019 VDD.n2852 VDD.n2851 0.0219844
R15020 VDD.n2882 VDD.n2881 0.0219844
R15021 VDD.n2935 VDD.n2934 0.0219844
R15022 VDD.n82 VDD.n80 0.0219844
R15023 VDD.n127 VDD.n126 0.0219844
R15024 VDD.n5589 VDD.n5537 0.0219844
R15025 VDD.n230 VDD.n229 0.0219844
R15026 VDD.n2546 VDD.n2545 0.0219844
R15027 VDD.n5464 VDD.n262 0.0217264
R15028 VDD.n5481 VDD.n5480 0.0217264
R15029 VDD.n5485 VDD.n252 0.0217264
R15030 VDD.n5623 VDD.n5614 0.0215953
R15031 VDD.n6499 VDD.n6498 0.0215953
R15032 VDD.n7332 VDD.n7323 0.0215953
R15033 VDD.n8208 VDD.n8207 0.0215953
R15034 VDD.n5607 VDD.n1 0.0211408
R15035 VDD.n3306 VDD.n17 0.0210308
R15036 VDD.n3014 VDD.n3013 0.0208125
R15037 VDD.n3363 VDD.n3362 0.0205059
R15038 VDD.n3291 VDD.n3290 0.0205059
R15039 VDD.n8240 VDD.n8239 0.0202566
R15040 VDD.n3367 VDD.n3327 0.0200312
R15041 VDD.n3069 VDD.n3066 0.0200312
R15042 VDD.n2588 VDD.n2587 0.0200312
R15043 VDD.n2589 VDD.n2508 0.0200312
R15044 VDD.n6531 VDD.n6530 0.019913
R15045 VDD.n3632 VDD.n3628 0.0198977
R15046 VDD.n3974 VDD.n3973 0.0197278
R15047 VDD.n3907 VDD.n3701 0.0196275
R15048 VDD.n3536 VDD.n3487 0.0195217
R15049 VDD.n3238 VDD.n3189 0.0195217
R15050 VDD.n5490 VDD.n239 0.0193679
R15051 VDD.n3338 VDD.n3335 0.01925
R15052 VDD.n3798 VDD.n3797 0.0186403
R15053 VDD.n3912 VDD.n3663 0.0186403
R15054 VDD.n3694 VDD.n3670 0.0186403
R15055 VDD.n2850 VDD.n2805 0.0186403
R15056 VDD.n2884 VDD.n2883 0.0186403
R15057 VDD.n3603 VDD.n2643 0.0185773
R15058 VDD.n3439 VDD.n2708 0.0185773
R15059 VDD.n2726 VDD.n2718 0.0185773
R15060 VDD.n3385 VDD.n2744 0.0185773
R15061 VDD.n5676 VDD.n5675 0.0185769
R15062 VDD.n7385 VDD.n7384 0.0185769
R15063 VDD.n5495 VDD.n5494 0.0181887
R15064 VDD.n2568 VDD.n2533 0.0180781
R15065 VDD.n2560 VDD.n2534 0.0180781
R15066 VDD.n2549 VDD.n2541 0.0180781
R15067 VDD.n2562 VDD.n2561 0.0180781
R15068 VDD.n2550 VDD.n2539 0.0180781
R15069 VDD.n3919 VDD.n3656 0.0176875
R15070 VDD.n2864 VDD.n2794 0.0176875
R15071 VDD.n242 VDD.n239 0.0176875
R15072 VDD.n2628 VDD.n2590 0.0176875
R15073 VDD.n3961 VDD.n3631 0.0169062
R15074 VDD.n155 VDD.n154 0.0169062
R15075 VDD.n2595 VDD.n2590 0.0169062
R15076 VDD.n3975 VDD.n2630 0.0169062
R15077 VDD.n3717 VDD.n3716 0.0168893
R15078 VDD.n3907 VDD.n3906 0.0168893
R15079 VDD.n3814 VDD.n3813 0.0168893
R15080 VDD.n2817 VDD.n2815 0.0168893
R15081 VDD.n2995 VDD.n2994 0.0168893
R15082 VDD.n3522 VDD.n3489 0.0168043
R15083 VDD.n3224 VDD.n3191 0.0168043
R15084 VDD.n3731 VDD.n3713 0.0168043
R15085 VDD.n3892 VDD.n3704 0.0168043
R15086 VDD.n3828 VDD.n3756 0.0168043
R15087 VDD.n2836 VDD.n2819 0.0168043
R15088 VDD.n2979 VDD.n2978 0.0168043
R15089 VDD.n5638 VDD.n5637 0.0165473
R15090 VDD.n6493 VDD.n6492 0.0165473
R15091 VDD.n7347 VDD.n7346 0.0165473
R15092 VDD.n8202 VDD.n8201 0.0165473
R15093 VDD.n3614 VDD.n3613 0.016125
R15094 VDD.n2686 VDD.n2685 0.016125
R15095 VDD.n3475 VDD.n3474 0.016125
R15096 VDD.n3578 VDD.n3577 0.016125
R15097 VDD.n3572 VDD.n3478 0.016125
R15098 VDD.n3471 VDD.n3470 0.016125
R15099 VDD.n3466 VDD.n2689 0.016125
R15100 VDD.n3461 VDD.n2698 0.016125
R15101 VDD.n3448 VDD.n3434 0.016125
R15102 VDD.n3452 VDD.n2702 0.016125
R15103 VDD.n3431 VDD.n3430 0.016125
R15104 VDD.n3426 VDD.n3425 0.016125
R15105 VDD.n3412 VDD.n2731 0.016125
R15106 VDD.n3422 VDD.n2732 0.016125
R15107 VDD.n3408 VDD.n3400 0.016125
R15108 VDD.n3394 VDD.n3380 0.016125
R15109 VDD.n3398 VDD.n2738 0.016125
R15110 VDD.n3357 VDD.n2766 0.016125
R15111 VDD.n3372 VDD.n3328 0.016125
R15112 VDD.n3285 VDD.n3067 0.016125
R15113 VDD.n3299 VDD.n3071 0.016125
R15114 VDD.n3177 VDD.n3176 0.016125
R15115 VDD.n3280 VDD.n3279 0.016125
R15116 VDD.n3274 VDD.n3180 0.016125
R15117 VDD.n3173 VDD.n3172 0.016125
R15118 VDD.n3097 VDD.n3090 0.016125
R15119 VDD.n3163 VDD.n3103 0.016125
R15120 VDD.n2947 VDD.n2898 0.016125
R15121 VDD.n2574 VDD.n2521 0.016125
R15122 VDD.n2569 VDD.n2568 0.016125
R15123 VDD.n2629 VDD.n2589 0.016125
R15124 VDD.n3978 VDD.n2632 0.016125
R15125 VDD.n5629 VDD.n5626 0.0157415
R15126 VDD.n6485 VDD.n6484 0.0157415
R15127 VDD.n7338 VDD.n7335 0.0157415
R15128 VDD.n8194 VDD.n8193 0.0157415
R15129 VDD.n5560 VDD.n5539 0.0145625
R15130 VDD.n3374 VDD.n2765 0.0145625
R15131 VDD.n3042 VDD.n2787 0.0143978
R15132 VDD.n3042 VDD.n2790 0.0143978
R15133 VDD.n2790 VDD.n2779 0.0143978
R15134 VDD.n3036 VDD.n2776 0.0143978
R15135 VDD.n3032 VDD.n2776 0.0143978
R15136 VDD.n3032 VDD.n2780 0.0143978
R15137 VDD.n3029 VDD.n2780 0.0143978
R15138 VDD.n3029 VDD.n2775 0.0143978
R15139 VDD.n3019 VDD.n2781 0.0143978
R15140 VDD.n3015 VDD.n2781 0.0143978
R15141 VDD.n3015 VDD.n2774 0.0143978
R15142 VDD.n3011 VDD.n2782 0.0143978
R15143 VDD.n3007 VDD.n2782 0.0143978
R15144 VDD.n3007 VDD.n2773 0.0143978
R15145 VDD.n147 VDD.n22 0.0143978
R15146 VDD.n147 VDD.n3 0.0143978
R15147 VDD.n5603 VDD.n7 0.0143978
R15148 VDD.n156 VDD.n148 0.0143978
R15149 VDD.n156 VDD.n10 0.0143978
R15150 VDD.n149 VDD.n10 0.0143978
R15151 VDD.n5600 VDD.n149 0.0143978
R15152 VDD.n5600 VDD.n151 0.0143978
R15153 VDD.n5524 VDD.n18 0.0143978
R15154 VDD.n5524 VDD.n19 0.0143978
R15155 VDD.n5521 VDD.n19 0.0143978
R15156 VDD.n5521 VDD.n13 0.0143978
R15157 VDD.n5517 VDD.n21 0.0143978
R15158 VDD.n5513 VDD.n21 0.0143978
R15159 VDD.n3331 VDD.n2748 0.0143978
R15160 VDD.n3332 VDD.n3331 0.0143978
R15161 VDD.n3332 VDD.n2757 0.0143978
R15162 VDD.n3336 VDD.n2757 0.0143978
R15163 VDD.n3340 VDD.n2750 0.0143978
R15164 VDD.n3340 VDD.n2758 0.0143978
R15165 VDD.n3343 VDD.n2758 0.0143978
R15166 VDD.n3343 VDD.n2749 0.0143978
R15167 VDD.n3346 VDD.n2749 0.0143978
R15168 VDD.n3375 VDD.n2763 0.0143978
R15169 VDD.n2763 VDD.n2754 0.0143978
R15170 VDD.n3323 VDD.n2754 0.0143978
R15171 VDD.n3323 VDD.n2755 0.0143978
R15172 VDD.n3320 VDD.n2755 0.0143978
R15173 VDD.n3320 VDD.n2753 0.0143978
R15174 VDD.n3317 VDD.n2753 0.0143978
R15175 VDD.n3317 VDD.n3316 0.0143978
R15176 VDD.n3316 VDD.n3315 0.0143978
R15177 VDD.n3315 VDD.n2770 0.0143978
R15178 VDD.n3311 VDD.n2770 0.0143978
R15179 VDD.n3311 VDD.n3310 0.0143978
R15180 VDD.n3310 VDD.n3049 0.0143978
R15181 VDD.n3307 VDD.n3049 0.0143978
R15182 VDD.n3307 VDD.n3055 0.0143978
R15183 VDD.n2644 VDD.n2634 0.0141719
R15184 VDD.n3569 VDD.n3568 0.0141719
R15185 VDD.n3458 VDD.n3457 0.0141719
R15186 VDD.n3442 VDD.n2700 0.0141719
R15187 VDD.n2722 VDD.n2710 0.0141719
R15188 VDD.n3420 VDD.n3419 0.0141719
R15189 VDD.n3388 VDD.n2736 0.0141719
R15190 VDD.n3363 VDD.n3327 0.0141719
R15191 VDD.n3291 VDD.n3069 0.0141719
R15192 VDD.n3271 VDD.n3270 0.0141719
R15193 VDD.n3160 VDD.n3159 0.0141719
R15194 VDD.n44 VDD.n33 0.0141719
R15195 VDD.n112 VDD.n26 0.0141719
R15196 VDD.n5544 VDD.n163 0.0141719
R15197 VDD.n189 VDD.n165 0.0141719
R15198 VDD.n2581 VDD.n2580 0.0141719
R15199 VDD.n2648 VDD.n2645 0.014087
R15200 VDD.n3562 VDD.n3481 0.014087
R15201 VDD.n3541 VDD.n3486 0.014087
R15202 VDD.n3264 VDD.n3183 0.014087
R15203 VDD.n3243 VDD.n3188 0.014087
R15204 VDD.n3121 VDD.n3118 0.014087
R15205 VDD.n5604 VDD.n3 0.0138925
R15206 VDD.n3021 VDD.n2870 0.0137813
R15207 VDD.n3037 VDD.n2779 0.0136398
R15208 VDD.n5518 VDD.n5517 0.0136398
R15209 VDD.n3018 VDD.n2873 0.013
R15210 VDD.n5598 VDD.n5597 0.013
R15211 VDD.n3348 VDD.n3347 0.013
R15212 VDD.n3970 VDD.n3968 0.0128788
R15213 VDD.n3944 VDD.n3627 0.0128788
R15214 VDD.n3959 VDD.n3627 0.0128788
R15215 VDD.n3971 VDD.n3970 0.0128788
R15216 VDD.n3576 VDD.n3575 0.0127111
R15217 VDD.n3463 VDD.n2696 0.0127111
R15218 VDD.n3406 VDD.n2734 0.0127111
R15219 VDD.n3278 VDD.n3277 0.0127111
R15220 VDD.n3165 VDD.n3101 0.0127111
R15221 VDD.n3377 VDD.n2748 0.012629
R15222 VDD.n3056 VDD.n3055 0.012629
R15223 VDD.n5487 VDD.n254 0.0122925
R15224 VDD.n5491 VDD.n5490 0.0122925
R15225 VDD.n5493 VDD.n253 0.0122925
R15226 VDD.n2686 VDD.n2642 0.0122188
R15227 VDD.n3452 VDD.n3451 0.0122188
R15228 VDD.n3425 VDD.n2729 0.0122188
R15229 VDD.n3398 VDD.n3397 0.0122188
R15230 VDD.n3372 VDD.n3350 0.0122188
R15231 VDD.n3299 VDD.n3062 0.0122188
R15232 VDD.n3915 VDD.n3914 0.0122188
R15233 VDD.n3923 VDD.n3922 0.0122188
R15234 VDD.n3691 VDD.n3687 0.0122188
R15235 VDD.n3686 VDD.n3684 0.0122188
R15236 VDD.n3795 VDD.n3647 0.0122188
R15237 VDD.n3801 VDD.n3651 0.0122188
R15238 VDD.n3777 VDD.n3776 0.0122188
R15239 VDD.n3941 VDD.n3940 0.0122188
R15240 VDD.n2853 VDD.n2852 0.0122188
R15241 VDD.n2863 VDD.n2862 0.0122188
R15242 VDD.n2881 VDD.n2880 0.0122188
R15243 VDD.n3027 VDD.n2874 0.0122188
R15244 VDD.n2934 VDD.n2895 0.0122188
R15245 VDD.n3002 VDD.n3001 0.0122188
R15246 VDD.n91 VDD.n31 0.0122188
R15247 VDD.n80 VDD.n36 0.0122188
R15248 VDD.n115 VDD.n106 0.0122188
R15249 VDD.n128 VDD.n127 0.0122188
R15250 VDD.n5596 VDD.n164 0.0122188
R15251 VDD.n5537 VDD.n5536 0.0122188
R15252 VDD.n237 VDD.n173 0.0122188
R15253 VDD.n229 VDD.n228 0.0122188
R15254 VDD.n2525 VDD.n2512 0.0122188
R15255 VDD.n2564 VDD.n2533 0.0122188
R15256 VDD.n2546 VDD.n2541 0.0122188
R15257 VDD.n2524 VDD.n2523 0.0122188
R15258 VDD.n5633 VDD.n5632 0.0114797
R15259 VDD.n5624 VDD.n5623 0.0114797
R15260 VDD.n6482 VDD.n6481 0.0114797
R15261 VDD.n6498 VDD.n6497 0.0114797
R15262 VDD.n7342 VDD.n7341 0.0114797
R15263 VDD.n7333 VDD.n7332 0.0114797
R15264 VDD.n8191 VDD.n8190 0.0114797
R15265 VDD.n8207 VDD.n8206 0.0114797
R15266 VDD.n3006 VDD.n3005 0.0114375
R15267 VDD.n9024 VDD.n8241 0.0111838
R15268 VDD.n8169 VDD.n7386 0.0111838
R15269 VDD.n7315 VDD.n6532 0.0111838
R15270 VDD.n6460 VDD.n5677 0.0111838
R15271 VDD.n5478 VDD.n263 0.0111132
R15272 VDD.n5489 VDD.n254 0.0111132
R15273 VDD.n3303 VDD.n3064 0.0106562
R15274 VDD.n3301 VDD.n3064 0.0106562
R15275 VDD.n3922 VDD.n3655 0.0102656
R15276 VDD.n3684 VDD.n3681 0.0102656
R15277 VDD.n3801 VDD.n3800 0.0102656
R15278 VDD.n3940 VDD.n3639 0.0102656
R15279 VDD.n2862 VDD.n2802 0.0102656
R15280 VDD.n2885 VDD.n2874 0.0102656
R15281 VDD.n3001 VDD.n2911 0.0102656
R15282 VDD.n92 VDD.n91 0.0102656
R15283 VDD.n115 VDD.n29 0.0102656
R15284 VDD.n5550 VDD.n164 0.0102656
R15285 VDD.n173 VDD.n171 0.0102656
R15286 VDD.n2865 VDD.n2787 0.0101021
R15287 VDD.n3020 VDD.n3019 0.0101021
R15288 VDD.n142 VDD.n22 0.0101021
R15289 VDD.n5513 VDD.n5512 0.0101021
R15290 VDD.n9026 VDD.n9025 0.0100583
R15291 VDD.n8171 VDD.n8170 0.0100583
R15292 VDD.n7317 VDD.n7316 0.0100583
R15293 VDD.n6462 VDD.n6461 0.0100583
R15294 VDD.n9030 VDD 0.00994196
R15295 VDD.n5478 VDD.n5477 0.00993396
R15296 VDD.n5487 VDD.n5486 0.00993396
R15297 VDD.n5540 VDD.n151 0.00984946
R15298 VDD.n3346 VDD.n2759 0.00984946
R15299 VDD.n3770 VDD.n3638 0.00957737
R15300 VDD.n3931 VDD.n3650 0.00957737
R15301 VDD.n3697 VDD.n3679 0.00957737
R15302 VDD.n3934 VDD.n3638 0.00957737
R15303 VDD.n3806 VDD.n3650 0.00957737
R15304 VDD.n3700 VDD.n3679 0.00957737
R15305 VDD.n2891 VDD.n2873 0.00957737
R15306 VDD.n2905 VDD.n2904 0.00957737
R15307 VDD.n3021 VDD.n2891 0.00957737
R15308 VDD.n2904 VDD.n2903 0.00957737
R15309 VDD.n105 VDD.n30 0.00957737
R15310 VDD.n140 VDD.n23 0.00957737
R15311 VDD.n5508 VDD.n172 0.00957737
R15312 VDD.n102 VDD.n30 0.00957737
R15313 VDD.n136 VDD.n23 0.00957737
R15314 VDD.n201 VDD.n172 0.00957737
R15315 VDD.n3604 VDD.n2636 0.00957737
R15316 VDD.n3480 VDD.n3477 0.00957737
R15317 VDD.n3454 VDD.n2692 0.00957737
R15318 VDD.n3433 VDD.n2703 0.00957737
R15319 VDD.n2728 VDD.n2712 0.00957737
R15320 VDD.n3421 VDD.n2735 0.00957737
R15321 VDD.n3379 VDD.n2739 0.00957737
R15322 VDD.n3182 VDD.n3179 0.00957737
R15323 VDD.n3117 VDD.n3092 0.00957737
R15324 VDD.n3114 VDD.n3113 0.00957737
R15325 VDD.n3102 VDD.n3092 0.00957737
R15326 VDD.n3396 VDD.n2739 0.00957737
R15327 VDD.n3410 VDD.n2735 0.00957737
R15328 VDD.n3450 VDD.n2703 0.00957737
R15329 VDD.n3424 VDD.n2712 0.00957737
R15330 VDD.n2697 VDD.n2692 0.00957737
R15331 VDD.n2687 VDD.n2636 0.00957737
R15332 VDD.n3480 VDD.n3473 0.00957737
R15333 VDD.n3182 VDD.n3175 0.00957737
R15334 VDD.n3113 VDD.n3111 0.00957737
R15335 VDD.n3962 VDD.n3624 0.00955797
R15336 VDD.n3969 VDD.n2631 0.00955797
R15337 VDD.n2946 VDD.n2773 0.00934409
R15338 VDD.n5656 VDD.n5655 0.00927193
R15339 VDD.n7365 VDD.n7364 0.00927193
R15340 VDD.n3111 VDD.n3106 0.00923422
R15341 VDD.n3962 VDD.n3625 0.0091882
R15342 VDD.n3942 VDD.n3635 0.0091882
R15343 VDD.n3806 VDD.n3644 0.0091882
R15344 VDD.n3919 VDD.n3653 0.0091882
R15345 VDD.n3700 VDD.n3678 0.0091882
R15346 VDD.n3770 VDD.n3635 0.0091882
R15347 VDD.n3689 VDD.n3678 0.0091882
R15348 VDD.n3930 VDD.n3653 0.0091882
R15349 VDD.n3933 VDD.n3644 0.0091882
R15350 VDD.n3957 VDD.n3625 0.0091882
R15351 VDD.n2801 VDD.n2794 0.0091882
R15352 VDD.n2947 VDD.n2893 0.0091882
R15353 VDD.n2907 VDD.n2900 0.0091882
R15354 VDD.n3005 VDD.n2893 0.0091882
R15355 VDD.n2903 VDD.n2900 0.0091882
R15356 VDD.n2801 VDD.n2800 0.0091882
R15357 VDD.n103 VDD.n37 0.0091882
R15358 VDD.n138 VDD.n137 0.0091882
R15359 VDD.n5597 VDD.n162 0.0091882
R15360 VDD.n5510 VDD.n167 0.0091882
R15361 VDD.n5507 VDD.n5506 0.0091882
R15362 VDD.n5560 VDD.n162 0.0091882
R15363 VDD.n103 VDD.n102 0.0091882
R15364 VDD.n201 VDD.n167 0.0091882
R15365 VDD.n137 VDD.n136 0.0091882
R15366 VDD.n5506 VDD.n239 0.0091882
R15367 VDD.n3604 VDD.n2633 0.0091882
R15368 VDD.n3477 VDD.n3476 0.0091882
R15369 VDD.n3472 VDD.n2690 0.0091882
R15370 VDD.n3453 VDD.n2701 0.0091882
R15371 VDD.n2728 VDD.n2709 0.0091882
R15372 VDD.n3410 VDD.n2730 0.0091882
R15373 VDD.n3399 VDD.n2737 0.0091882
R15374 VDD.n3349 VDD.n3348 0.0091882
R15375 VDD.n3179 VDD.n3178 0.0091882
R15376 VDD.n3174 VDD.n3091 0.0091882
R15377 VDD.n3396 VDD.n2737 0.0091882
R15378 VDD.n3178 VDD.n3068 0.0091882
R15379 VDD.n3102 VDD.n3091 0.0091882
R15380 VDD.n3349 VDD.n2765 0.0091882
R15381 VDD.n3423 VDD.n2730 0.0091882
R15382 VDD.n3432 VDD.n2709 0.0091882
R15383 VDD.n3450 VDD.n2701 0.0091882
R15384 VDD.n3615 VDD.n2633 0.0091882
R15385 VDD.n3476 VDD.n2688 0.0091882
R15386 VDD.n2697 VDD.n2690 0.0091882
R15387 VDD.n3116 VDD.n3106 0.00914234
R15388 VDD.n153 VDD.n7 0.0090914
R15389 VDD.n5633 VDD.n5631 0.00894595
R15390 VDD.n6482 VDD.n6480 0.00894595
R15391 VDD.n7342 VDD.n7340 0.00894595
R15392 VDD.n8191 VDD.n8189 0.00894595
R15393 VDD.n6526 VDD.n6523 0.00887321
R15394 VDD.n6526 VDD.n6525 0.00887321
R15395 VDD.n8235 VDD.n8232 0.00887321
R15396 VDD.n8235 VDD.n8234 0.00887321
R15397 VDD.n3967 VDD.n3966 0.00867391
R15398 VDD.n3591 VDD.n3590 0.00865217
R15399 VDD.n3557 VDD.n3482 0.00865217
R15400 VDD.n3546 VDD.n3485 0.00865217
R15401 VDD.n3259 VDD.n3184 0.00865217
R15402 VDD.n3248 VDD.n3187 0.00865217
R15403 VDD.n3147 VDD.n3146 0.00865217
R15404 VDD.n73 VDD.n58 0.00865217
R15405 VDD.n5565 VDD.n5561 0.00865217
R15406 VDD.n219 VDD.n204 0.00865217
R15407 VDD.n3972 VDD.n3969 0.00865217
R15408 VDD.n3337 VDD.n2750 0.00833333
R15409 VDD.n3913 VDD.n3654 0.0083125
R15410 VDD.n3696 VDD.n3695 0.0083125
R15411 VDD.n3796 VDD.n3645 0.0083125
R15412 VDD.n3775 VDD.n3634 0.0083125
R15413 VDD.n2851 VDD.n2795 0.0083125
R15414 VDD.n2882 VDD.n2871 0.0083125
R15415 VDD.n2935 VDD.n2892 0.0083125
R15416 VDD.n82 VDD.n81 0.0083125
R15417 VDD.n126 VDD.n25 0.0083125
R15418 VDD.n5589 VDD.n5588 0.0083125
R15419 VDD.n230 VDD.n166 0.0083125
R15420 VDD.n2586 VDD.n2510 0.0083125
R15421 VDD.n2559 VDD.n2536 0.0083125
R15422 VDD.n2555 VDD.n2554 0.0083125
R15423 VDD.n255 VDD.n2 0.0081375
R15424 VDD.n2945 VDD.n2944 0.00808064
R15425 VDD.n9024 VDD.n9023 0.00794532
R15426 VDD.n8169 VDD.n8168 0.00794532
R15427 VDD.n7315 VDD.n7314 0.00794532
R15428 VDD.n6460 VDD.n6459 0.00794532
R15429 VDD.n3012 VDD.n3011 0.00782796
R15430 VDD.n3962 VDD.n3622 0.00774638
R15431 VDD.n5467 VDD.n262 0.00757547
R15432 VDD.n3301 VDD.n3300 0.00753125
R15433 VDD.n3012 VDD.n2774 0.00706989
R15434 VDD.n261 VDD.n260 0.00694587
R15435 VDD.n3101 VDD.n3090 0.00685176
R15436 VDD.n3279 VDD.n3278 0.00685176
R15437 VDD.n3422 VDD.n2734 0.00685176
R15438 VDD.n2696 VDD.n2689 0.00685176
R15439 VDD.n3577 VDD.n3576 0.00685176
R15440 VDD.n2752 VDD.n2746 0.0068172
R15441 VDD.n3973 VDD.n3971 0.00678574
R15442 VDD.n2909 VDD.n2908 0.00675
R15443 VDD.n3303 VDD.n3061 0.00675
R15444 VDD.n3944 VDD.n3632 0.00661507
R15445 VDD.n3337 VDD.n3336 0.00656452
R15446 VDD.n5480 VDD.n258 0.00639623
R15447 VDD.n9025 VDD.n8242 0.00638768
R15448 VDD.n8170 VDD.n7387 0.00638768
R15449 VDD.n7316 VDD.n6533 0.00638768
R15450 VDD.n6461 VDD.n5678 0.00638768
R15451 VDD.n3606 VDD.n2642 0.00635938
R15452 VDD.n3451 VDD.n2705 0.00635938
R15453 VDD.n2729 VDD.n2716 0.00635938
R15454 VDD.n3397 VDD.n2741 0.00635938
R15455 VDD.n3369 VDD.n3350 0.00635938
R15456 VDD.n3296 VDD.n3062 0.00635938
R15457 VDD.n3302 VDD.n3066 0.00635938
R15458 VDD.n3963 VDD.n3623 0.00635938
R15459 VDD.n2582 VDD.n2581 0.00635938
R15460 VDD.n2529 VDD.n2521 0.00635938
R15461 VDD VDD.n9030 0.0061055
R15462 VDD.n3500 VDD.n3499 0.00593478
R15463 VDD.n3508 VDD.n3506 0.00593478
R15464 VDD.n3202 VDD.n3201 0.00593478
R15465 VDD.n3210 VDD.n3208 0.00593478
R15466 VDD.n3750 VDD.n3749 0.00593478
R15467 VDD.n3834 VDD.n3736 0.00593478
R15468 VDD.n3848 VDD.n3847 0.00593478
R15469 VDD.n3857 VDD.n3708 0.00593478
R15470 VDD.n3870 VDD.n3869 0.00593478
R15471 VDD.n3878 VDD.n3876 0.00593478
R15472 VDD.n2830 VDD.n2829 0.00593478
R15473 VDD.n2972 VDD.n2971 0.00593478
R15474 VDD.n153 VDD.n148 0.00580645
R15475 VDD.n3965 VDD.n3621 0.0056087
R15476 VDD.n2946 VDD.n2945 0.00555376
R15477 VDD.n3943 VDD.n3631 0.0051875
R15478 VDD.n3978 VDD.n3616 0.0051875
R15479 VDD.n5540 VDD.n18 0.00504839
R15480 VDD.n3375 VDD.n2759 0.00504839
R15481 VDD.n3628 VDD.n3621 0.00492754
R15482 VDD.n3073 VDD.n3067 0.00490286
R15483 VDD.n3353 VDD.n2766 0.00490286
R15484 VDD.n2865 VDD.n2778 0.0047957
R15485 VDD.n3020 VDD.n2775 0.0047957
R15486 VDD.n3045 VDD.n2783 0.0047957
R15487 VDD.n142 VDD.n12 0.0047957
R15488 VDD.n5512 VDD.n16 0.0047957
R15489 VDD.n5488 VDD.n255 0.00449057
R15490 VDD.n3569 VDD.n3478 0.00440625
R15491 VDD.n3458 VDD.n2698 0.00440625
R15492 VDD.n3420 VDD.n3400 0.00440625
R15493 VDD.n3271 VDD.n3180 0.00440625
R15494 VDD.n3160 VDD.n3103 0.00440625
R15495 VDD.n3915 VDD.n3652 0.00440625
R15496 VDD.n3698 VDD.n3687 0.00440625
R15497 VDD.n3932 VDD.n3647 0.00440625
R15498 VDD.n3777 VDD.n3633 0.00440625
R15499 VDD.n3958 VDD.n3957 0.00440625
R15500 VDD.n2853 VDD.n2797 0.00440625
R15501 VDD.n2880 VDD.n2868 0.00440625
R15502 VDD.n3004 VDD.n2895 0.00440625
R15503 VDD.n101 VDD.n41 0.00440625
R15504 VDD.n104 VDD.n36 0.00440625
R15505 VDD.n135 VDD.n110 0.00440625
R15506 VDD.n128 VDD.n24 0.00440625
R15507 VDD.n5559 VDD.n5542 0.00440625
R15508 VDD.n5536 VDD.n161 0.00440625
R15509 VDD.n200 VDD.n186 0.00440625
R15510 VDD.n228 VDD.n168 0.00440625
R15511 VDD.n2530 VDD.n2526 0.00440625
R15512 VDD.n2570 VDD.n2522 0.00440625
R15513 VDD.n2549 VDD.n2540 0.00440625
R15514 VDD.n2572 VDD.n2571 0.00440625
R15515 VDD.n3977 VDD.n3618 0.00433093
R15516 VDD.n3045 VDD.n2785 0.00429032
R15517 VDD.n12 VDD.n11 0.00429032
R15518 VDD.n16 VDD.n15 0.00429032
R15519 VDD.n5479 VDD.n261 0.00397228
R15520 VDD.n3028 VDD.n2870 0.003625
R15521 VDD.n5539 VDD.n5526 0.003625
R15522 VDD.n3374 VDD.n3373 0.003625
R15523 VDD.n3061 VDD.n3060 0.003625
R15524 VDD.n3583 VDD.n2666 0.00321739
R15525 VDD.n3552 VDD.n3483 0.00321739
R15526 VDD.n3551 VDD.n3484 0.00321739
R15527 VDD.n3254 VDD.n3185 0.00321739
R15528 VDD.n3253 VDD.n3186 0.00321739
R15529 VDD.n3139 VDD.n3135 0.00321739
R15530 VDD.n3769 VDD.n3767 0.00321739
R15531 VDD.n2926 VDD.n2918 0.00321739
R15532 VDD.n62 VDD.n59 0.00321739
R15533 VDD.n5576 VDD.n5575 0.00321739
R15534 VDD.n208 VDD.n205 0.00321739
R15535 VDD VDD.n5615 0.00303378
R15536 VDD VDD.n6501 0.00303378
R15537 VDD VDD.n7324 0.00303378
R15538 VDD VDD.n8210 0.00303378
R15539 VDD VDD.n5607 0.0029675
R15540 VDD.n3603 VDD.n2634 0.00295228
R15541 VDD.n2708 VDD.n2700 0.00295228
R15542 VDD.n2718 VDD.n2710 0.00295228
R15543 VDD.n2744 VDD.n2736 0.00295228
R15544 VDD.n5482 VDD.n5481 0.00285849
R15545 VDD.n5483 VDD.n257 0.00285849
R15546 VDD.n5494 VDD.n5493 0.00285849
R15547 VDD.n3038 VDD.n3035 0.00284375
R15548 VDD.n5520 VDD.n5519 0.00284375
R15549 VDD.n141 VDD.n6 0.00278115
R15550 VDD.n141 VDD.n8 0.00278115
R15551 VDD.n2756 VDD.n2747 0.00262546
R15552 VDD.n3376 VDD.n2756 0.00262546
R15553 VDD.n2944 VDD.n2783 0.00252151
R15554 VDD.n4294 VDD.n2359 0.00251613
R15555 VDD.n44 VDD.n42 0.00245312
R15556 VDD.n134 VDD.n112 0.00245312
R15557 VDD.n5558 VDD.n5544 0.00245312
R15558 VDD.n189 VDD.n187 0.00245312
R15559 VDD.n2448 VDD.n2447 0.00244542
R15560 VDD.n3058 VDD.n3050 0.00243946
R15561 VDD.n2793 VDD.n2791 0.00243946
R15562 VDD.n2791 VDD.n2789 0.00243946
R15563 VDD.n3058 VDD.n2772 0.00243946
R15564 VDD.n3377 VDD.n2746 0.00226882
R15565 VDD.n3305 VDD.n3056 0.00226882
R15566 VDD.n3960 VDD.n3959 0.0022029
R15567 VDD.n5502 VDD.n5501 0.00207156
R15568 VDD.n2445 VDD.n246 0.00207156
R15569 VDD.n2624 VDD.n2623 0.00207156
R15570 VDD.n2606 VDD.n2605 0.00207156
R15571 VDD.n4000 VDD.n3999 0.00207156
R15572 VDD.n3995 VDD.n3994 0.00207156
R15573 VDD.n3953 VDD.n2500 0.00207156
R15574 VDD.n3003 VDD.n2898 0.0020625
R15575 VDD.n269 VDD.n266 0.00194557
R15576 VDD.n269 VDD.n248 0.00194557
R15577 VDD.n5461 VDD.n5460 0.00194557
R15578 VDD.n5460 VDD.n248 0.00194557
R15579 VDD.n5501 VDD.n243 0.00194557
R15580 VDD.n246 VDD.n244 0.00194557
R15581 VDD.n2449 VDD.n2448 0.00194557
R15582 VDD.n2625 VDD.n2624 0.00194557
R15583 VDD.n2606 VDD.n2596 0.00194557
R15584 VDD.n3999 VDD.n3998 0.00194557
R15585 VDD.n3996 VDD.n3995 0.00194557
R15586 VDD.n2485 VDD.n2483 0.00194557
R15587 VDD.n2483 VDD.n2480 0.00194557
R15588 VDD.n3109 VDD.n2478 0.00194557
R15589 VDD.n2480 VDD.n2478 0.00194557
R15590 VDD.n3954 VDD.n3953 0.00194557
R15591 VDD.n3949 VDD.n2501 0.00194557
R15592 VDD.n3983 VDD.n2501 0.00194557
R15593 VDD.n3982 VDD.n3981 0.00194557
R15594 VDD.n3983 VDD.n3982 0.00194557
R15595 VDD.n3619 VDD.n2497 0.00194557
R15596 VDD.n3983 VDD.n2497 0.00194557
R15597 VDD.n3968 VDD.n3967 0.00186232
R15598 VDD.n3305 VDD.n3304 0.00176344
R15599 VDD.n4026 VDD.n2288 0.00175186
R15600 VDD.n5477 VDD.n259 0.00167925
R15601 VDD.n5464 VDD.n5463 0.00167925
R15602 VDD.n5486 VDD.n256 0.00167925
R15603 VDD.n5476 VDD.n264 0.00167925
R15604 VDD.n5465 VDD.n5462 0.00167925
R15605 VDD.n5485 VDD.n5484 0.00167925
R15606 VDD.n5601 VDD.n4 0.00145036
R15607 VDD.n5602 VDD.n5601 0.00145036
R15608 VDD.n14 VDD.n1 0.00143078
R15609 VDD.n14 VDD.n5 0.00143078
R15610 VDD.n2769 VDD.n2761 0.00141098
R15611 VDD.n2769 VDD.n2764 0.00141098
R15612 VDD.n3964 VDD.n3622 0.0014058
R15613 VDD.n2768 VDD.n2760 0.00139311
R15614 VDD.n2768 VDD.n2762 0.00139311
R15615 VDD.n5502 VDD.n248 0.00137395
R15616 VDD.n2445 VDD.n248 0.00137395
R15617 VDD.n2623 VDD.n1019 0.00137395
R15618 VDD.n2605 VDD.n1019 0.00137395
R15619 VDD.n3994 VDD.n2480 0.00137395
R15620 VDD.n4000 VDD.n2480 0.00137395
R15621 VDD.n3983 VDD.n2500 0.00137395
R15622 VDD.n3051 VDD.n3047 0.00136393
R15623 VDD.n3044 VDD.n2786 0.00136393
R15624 VDD.n3308 VDD.n3051 0.00136393
R15625 VDD.n3044 VDD.n3043 0.00136393
R15626 VDD.n3057 VDD.n3048 0.00134811
R15627 VDD.n2784 VDD.n2777 0.00134811
R15628 VDD.n3046 VDD.n2777 0.00134811
R15629 VDD.n3306 VDD.n3048 0.00134811
R15630 VDD.n3962 VDD.n3961 0.00128125
R15631 VDD.n3975 VDD.n3969 0.00128125
R15632 VDD.n3969 VDD.n2632 0.00128125
R15633 VDD.n3037 VDD.n3036 0.00125806
R15634 VDD.n5518 VDD.n13 0.00125806
R15635 VDD.n150 VDD.n5 0.00119582
R15636 VDD.n150 VDD.n8 0.00119582
R15637 VDD.n3330 VDD.n2747 0.0011787
R15638 VDD.n3330 VDD.n2762 0.0011787
R15639 VDD.n4297 VDD.n4296 0.00117707
R15640 VDD.n20 VDD.n6 0.00117624
R15641 VDD.n20 VDD.n4 0.00117624
R15642 VDD.n2764 VDD.n2751 0.00116083
R15643 VDD.n3376 VDD.n2751 0.00116083
R15644 VDD.n3057 VDD.n3054 0.00115824
R15645 VDD.n2789 VDD.n2788 0.00115824
R15646 VDD.n2788 VDD.n2784 0.00115824
R15647 VDD.n3054 VDD.n2772 0.00115824
R15648 VDD.n3309 VDD.n3308 0.00114242
R15649 VDD.n2793 VDD.n2792 0.00114242
R15650 VDD.n2792 VDD.n2786 0.00114242
R15651 VDD.n3309 VDD.n3050 0.00114242
R15652 VDD.n4010 VDD.n2477 0.00105433
R15653 VDD.n3984 VDD.n2494 0.00104275
R15654 VDD.n4027 VDD.n4026 0.00104275
R15655 VDD.n2477 VDD.n2474 0.00104275
R15656 VDD.n4028 VDD.n248 0.00103737
R15657 VDD.n4026 VDD.n4025 0.00103651
R15658 VDD.n3985 VDD.n3984 0.00101611
R15659 VDD.n5499 VDD.n5498 0.00101576
R15660 VDD.n3992 VDD.n3991 0.00101522
R15661 VDD.n2457 VDD.n2456 0.00100772
R15662 VDD.n4196 VDD.n4028 0.00100538
R15663 VDD.n5604 VDD.n5603 0.00100538
R15664 VDD.n2505 VDD.n2498 0.00100409
R15665 VDD.n4002 VDD.n2484 0.00100409
R15666 VDD.n2447 VDD.n2443 0.00100372
R15667 VDD.n2609 VDD.n2608 0.00100292
R15668 VDD.n2608 VDD.n2601 0.00100251
R15669 VDD.n4003 VDD.n4002 0.00100251
R15670 VDD.n3946 VDD.n2498 0.00100251
R15671 VDD.n5499 VDD.n248 0.00100095
R15672 VDD.n3992 VDD.n2480 0.00100089
R15673 VDD.n2456 VDD.n248 0.00100024
R15674 VDD.n4301 VDD.n4300 0.00100002
R15675 VDD.n9023 VDD.n8242 0.00100001
R15676 VDD.n8168 VDD.n7387 0.00100001
R15677 VDD.n7314 VDD.n6533 0.00100001
R15678 VDD.n6459 VDD.n5678 0.00100001
R15679 VDD.n6462 VDD.n5677 0.001
R15680 VDD.n7317 VDD.n6532 0.001
R15681 VDD.n8171 VDD.n7386 0.001
R15682 VDD.n9026 VDD.n8241 0.001
R15683 VDD.n2447 VDD.n248 0.001
R15684 VDD.n2608 VDD.n1019 0.001
R15685 VDD.n4002 VDD.n2480 0.001
R15686 VDD.n2480 VDD.n2477 0.001
R15687 VDD.n3984 VDD.n3983 0.001
R15688 VDD.n3983 VDD.n2498 0.001
R15689 VDD.n4299 VDD.n4298 0.000855023
R15690 VDD.n4298 VDD.n4297 0.000855023
R15691 VDD.n4299 VDD.n2341 0.000855004
R15692 VDD.n5479 VDD.n255 0.00079375
R15693 VDD.n4011 VDD.n4010 0.000554326
R15694 VDD.n2459 VDD.n2441 0.000542748
R15695 VDD.n2441 VDD.n248 0.000542748
R15696 VDD.n4196 VDD.n4195 0.000542748
R15697 VDD.n4027 VDD.n2287 0.000542748
R15698 VDD.n4024 VDD.n2340 0.000542748
R15699 VDD.n4025 VDD.n4024 0.000542748
R15700 VDD.n4012 VDD.n2474 0.000542748
R15701 VDD.n3989 VDD.n2492 0.000542748
R15702 VDD.n2492 VDD.n2480 0.000542748
R15703 VDD.n3987 VDD.n2494 0.000542748
R15704 VDD.n2613 VDD.n2612 0.000542748
R15705 VDD.n2613 VDD.n1019 0.000542748
R15706 VDD.n2603 VDD.n1019 0.000523923
R15707 VDD.n3983 VDD.n2473 0.000523923
R15708 VDD.n2475 VDD.n2473 0.000523923
R15709 VDD.n2618 VDD.n2603 0.000523923
R15710 VDD.n5498 VDD.n5497 0.000516711
R15711 VDD.n3991 VDD.n3990 0.000516107
R15712 VDD.n3986 VDD.n3985 0.000516107
R15713 VDD.n2458 VDD.n2457 0.000507966
R15714 VDD.n4005 VDD.n2484 0.000504095
R15715 VDD.n2506 VDD.n2505 0.000504095
R15716 VDD.n2450 VDD.n2443 0.000503718
R15717 VDD.n2611 VDD.n2609 0.000502918
R15718 VDD.n2615 VDD.n2614 0.000502851
R15719 VDD.n2614 VDD.n2493 0.000502851
R15720 VDD.n2610 VDD.n2601 0.000502515
R15721 VDD.n4004 VDD.n4003 0.000502515
R15722 VDD.n3946 VDD.n3945 0.000502515
R15723 VDD.n4329 VDD.n2288 0.000501859
R15724 VDD.n2617 VDD.n2616 0.000501425
R15725 VDD.n2616 VDD.n2615 0.000501425
R15726 VDD.n8363 VDD.n8242 0.000500887
R15727 VDD.n7508 VDD.n7387 0.000500887
R15728 VDD.n6654 VDD.n6533 0.000500887
R15729 VDD.n5799 VDD.n5678 0.000500887
R15730 VDD.n9025 VDD.n9024 0.000500755
R15731 VDD.n8170 VDD.n8169 0.000500755
R15732 VDD.n7316 VDD.n7315 0.000500755
R15733 VDD.n6461 VDD.n6460 0.000500755
R15734 VDD.n2461 VDD.n2460 0.000500648
R15735 VDD.t54 VDD.n2461 0.000500648
R15736 VDD.n4197 VDD.n2438 0.000500648
R15737 VDD.t54 VDD.n4197 0.000500648
R15738 VDD.n6465 VDD.n6464 0.0005006
R15739 VDD.n7320 VDD.n7319 0.0005006
R15740 VDD.n8174 VDD.n8173 0.0005006
R15741 VDD.n9029 VDD.n9028 0.0005006
R15742 VDD.n4014 VDD.n4013 0.000500389
R15743 VDD.n4015 VDD.n4014 0.000500389
R15744 VDD.n3988 VDD.n2472 0.000500389
R15745 VDD.n4015 VDD.n2472 0.000500389
R15746 VDD.n8716 VDD.n8246 0.000500314
R15747 VDD.n7861 VDD.n7391 0.000500314
R15748 VDD.n7007 VDD.n6537 0.000500314
R15749 VDD.n6152 VDD.n5682 0.000500314
R15750 VDD.n5677 VDD.n5676 0.000500314
R15751 VDD.n6532 VDD.n6531 0.000500314
R15752 VDD.n7386 VDD.n7385 0.000500314
R15753 VDD.n8241 VDD.n8240 0.000500314
R15754 VDD.n6463 VDD.n5611 0.000500311
R15755 VDD.n7318 VDD.n5610 0.000500311
R15756 VDD.n8172 VDD.n5609 0.000500311
R15757 VDD.n9027 VDD.n5608 0.000500311
R15758 VDD.n9021 VDD.n9020 0.000500201
R15759 VDD.n8166 VDD.n8165 0.000500201
R15760 VDD.n7312 VDD.n7311 0.000500201
R15761 VDD.n6457 VDD.n6456 0.000500201
R15762 VDD.n4302 VDD.n4301 0.000500031
R15763 VSS.n1272 VSS.n196 5581.17
R15764 VSS.n1279 VSS.n192 4777.48
R15765 VSS.n1264 VSS.n192 4777.48
R15766 VSS.n1272 VSS.n195 3889.41
R15767 VSS.n1883 VSS.n1706 1956.7
R15768 VSS.n1878 VSS.n1706 1956.7
R15769 VSS.n1886 VSS.n1703 1892.49
R15770 VSS.n1709 VSS.n1703 1892.49
R15771 VSS.n1875 VSS.t60 1049.46
R15772 VSS.t38 VSS.n1704 1045.16
R15773 VSS.t60 VSS.t14 984.947
R15774 VSS.t14 VSS.t12 984.947
R15775 VSS.t41 VSS.t10 984.947
R15776 VSS.t10 VSS.t38 984.947
R15777 VSS.n1034 VSS.n204 927.715
R15778 VSS.n588 VSS.n191 803.688
R15779 VSS.n1279 VSS.n191 803.688
R15780 VSS.t53 VSS.t50 671.51
R15781 VSS.t50 VSS.t8 671.51
R15782 VSS.t8 VSS.t35 671.51
R15783 VSS.t35 VSS.t0 671.51
R15784 VSS.t0 VSS.t27 671.51
R15785 VSS.t27 VSS.t68 671.51
R15786 VSS.t4 VSS.t20 671.51
R15787 VSS.t2 VSS.t4 671.51
R15788 VSS.t29 VSS.t2 671.51
R15789 VSS.t24 VSS.t29 671.51
R15790 VSS.t18 VSS.t24 671.51
R15791 VSS.t16 VSS.t18 671.51
R15792 VSS.t46 VSS.t16 671.51
R15793 VSS.n590 VSS.t6 617.261
R15794 VSS.n1273 VSS.t22 614.33
R15795 VSS.n1034 VSS.n1033 585
R15796 VSS.n1033 VSS.n199 585
R15797 VSS.n1033 VSS.n1032 585
R15798 VSS.n1259 VSS.n1258 585
R15799 VSS.n1259 VSS.n214 585
R15800 VSS.n1260 VSS.n211 585
R15801 VSS.n1258 VSS.n211 585
R15802 VSS.n214 VSS.n211 585
R15803 VSS.n1260 VSS.n1259 585
R15804 VSS.n1275 VSS.n1274 585
R15805 VSS.n1274 VSS.n182 585
R15806 VSS.n1274 VSS.n184 585
R15807 VSS.n598 VSS.n184 585
R15808 VSS.n598 VSS.n182 585
R15809 VSS.n1274 VSS.t53 561.547
R15810 VSS.n1259 VSS.t46 561.547
R15811 VSS.t12 VSS.n1874 492.474
R15812 VSS.n1874 VSS.t41 492.474
R15813 VSS.n1271 VSS.n1270 417.392
R15814 VSS.n1278 VSS.n194 357.288
R15815 VSS.n1263 VSS.n194 357.288
R15816 VSS.n599 VSS.n597 340.154
R15817 VSS.t30 VSS.n596 338.688
R15818 VSS.n212 VSS.t22 335.755
R15819 VSS.t20 VSS.n212 335.755
R15820 VSS.n1271 VSS.n197 291.457
R15821 VSS.n1275 VSS.n190 260.455
R15822 VSS.n1260 VSS.n208 260.455
R15823 VSS.n596 VSS.n583 236.055
R15824 VSS.n597 VSS.t30 197.935
R15825 VSS.n1749 VSS.n1748 185
R15826 VSS.n1745 VSS.n1744 185
R15827 VSS.n1741 VSS.n1740 185
R15828 VSS.n1737 VSS.n1736 185
R15829 VSS.n1733 VSS.n1732 185
R15830 VSS.n1810 VSS.n1731 185
R15831 VSS.n1726 VSS.n1725 185
R15832 VSS.n1820 VSS.n1819 185
R15833 VSS.n1828 VSS.n1720 185
R15834 VSS.n1839 VSS.n1838 185
R15835 VSS.n1858 VSS.n1716 185
R15836 VSS.n1845 VSS.n1844 185
R15837 VSS.n1777 VSS.n1776 185
R15838 VSS.n1784 VSS.n1783 185
R15839 VSS.n1791 VSS.n1790 185
R15840 VSS.n1798 VSS.n1797 185
R15841 VSS.n1805 VSS.n1804 185
R15842 VSS.n1809 VSS.n1808 185
R15843 VSS.n1807 VSS.n1806 185
R15844 VSS.n1818 VSS.n1724 185
R15845 VSS.n1827 VSS.n1826 185
R15846 VSS.n1837 VSS.n1717 185
R15847 VSS.n1842 VSS.n1841 185
R15848 VSS.n1860 VSS.n1859 185
R15849 VSS.n1585 VSS.n1584 185
R15850 VSS.n1581 VSS.n1580 185
R15851 VSS.n1577 VSS.n1576 185
R15852 VSS.n1573 VSS.n1572 185
R15853 VSS.n1569 VSS.n1568 185
R15854 VSS.n1646 VSS.n1567 185
R15855 VSS.n1562 VSS.n1561 185
R15856 VSS.n1656 VSS.n1655 185
R15857 VSS.n1664 VSS.n1556 185
R15858 VSS.n1675 VSS.n1674 185
R15859 VSS.n1694 VSS.n1552 185
R15860 VSS.n1681 VSS.n1680 185
R15861 VSS.n1613 VSS.n1612 185
R15862 VSS.n1620 VSS.n1619 185
R15863 VSS.n1627 VSS.n1626 185
R15864 VSS.n1634 VSS.n1633 185
R15865 VSS.n1641 VSS.n1640 185
R15866 VSS.n1645 VSS.n1644 185
R15867 VSS.n1643 VSS.n1642 185
R15868 VSS.n1654 VSS.n1560 185
R15869 VSS.n1663 VSS.n1662 185
R15870 VSS.n1673 VSS.n1553 185
R15871 VSS.n1696 VSS.n1695 185
R15872 VSS.n1678 VSS.n1677 185
R15873 VSS.n1364 VSS.n1363 185
R15874 VSS.n1363 VSS.n1362 185
R15875 VSS.n1495 VSS.n1494 185
R15876 VSS.n1495 VSS.n61 185
R15877 VSS.n1496 VSS.n52 185
R15878 VSS.n1496 VSS.n44 185
R15879 VSS.n1305 VSS.n1304 185
R15880 VSS.n176 VSS.n172 185
R15881 VSS.n174 VSS.n158 185
R15882 VSS.n166 VSS.n165 185
R15883 VSS.n164 VSS.n163 185
R15884 VSS.n1306 VSS.n156 185
R15885 VSS.n1119 VSS.n1118 185
R15886 VSS.n1119 VSS.n1107 185
R15887 VSS.n1139 VSS.n1136 185
R15888 VSS.n1240 VSS.n1239 185
R15889 VSS.n1241 VSS.n1157 185
R15890 VSS.n1230 VSS.n1229 185
R15891 VSS.n1232 VSS.n1231 185
R15892 VSS.n1220 VSS.n1219 185
R15893 VSS.n1222 VSS.n1221 185
R15894 VSS.n1159 VSS.n1158 185
R15895 VSS.n1163 VSS.n1162 185
R15896 VSS.n1167 VSS.n1166 185
R15897 VSS.n1211 VSS.n1210 185
R15898 VSS.n1202 VSS.n1201 185
R15899 VSS.n1195 VSS.n1194 185
R15900 VSS.n366 VSS.n259 185
R15901 VSS.n995 VSS.n994 185
R15902 VSS.n965 VSS.n964 185
R15903 VSS.n969 VSS.n968 185
R15904 VSS.n973 VSS.n972 185
R15905 VSS.n975 VSS.n974 185
R15906 VSS.n981 VSS.n980 185
R15907 VSS.n988 VSS.n987 185
R15908 VSS.n1017 VSS.n1016 185
R15909 VSS.n1006 VSS.n1005 185
R15910 VSS.n1015 VSS.n229 185
R15911 VSS.n1004 VSS.n959 185
R15912 VSS.n961 VSS.n960 185
R15913 VSS.n644 VSS.n643 185
R15914 VSS.n614 VSS.n613 185
R15915 VSS.n618 VSS.n617 185
R15916 VSS.n622 VSS.n621 185
R15917 VSS.n624 VSS.n623 185
R15918 VSS.n630 VSS.n629 185
R15919 VSS.n637 VSS.n636 185
R15920 VSS.n657 VSS.n608 185
R15921 VSS.n506 VSS.n505 185
R15922 VSS.n659 VSS.n658 185
R15923 VSS.n652 VSS.n651 185
R15924 VSS.n610 VSS.n609 185
R15925 VSS.n786 VSS.n493 185
R15926 VSS.n535 VSS.n512 185
R15927 VSS.n526 VSS.n512 185
R15928 VSS.n1759 VSS.n1758 152
R15929 VSS.n1760 VSS.n1754 152
R15930 VSS.n1927 VSS.n1926 152
R15931 VSS.n1925 VSS.n1924 152
R15932 VSS.n1595 VSS.n1594 152
R15933 VSS.n1593 VSS.n1592 152
R15934 VSS.n124 VSS.n121 152
R15935 VSS.n123 VSS.n122 152
R15936 VSS.n1433 VSS.n1427 152
R15937 VSS.n1432 VSS.n1431 152
R15938 VSS.n1410 VSS.n75 152
R15939 VSS.n1418 VSS.n69 152
R15940 VSS.n1409 VSS.n72 152
R15941 VSS.n1417 VSS.n1416 152
R15942 VSS.n1389 VSS.n117 152
R15943 VSS.n1397 VSS.n111 152
R15944 VSS.n1388 VSS.n114 152
R15945 VSS.n1396 VSS.n1395 152
R15946 VSS.n1080 VSS.n1074 152
R15947 VSS.n1079 VSS.n1078 152
R15948 VSS.n1178 VSS.n1172 152
R15949 VSS.n1177 VSS.n1176 152
R15950 VSS.n268 VSS.n265 152
R15951 VSS.n267 VSS.n266 152
R15952 VSS.n285 VSS.n279 152
R15953 VSS.n284 VSS.n283 152
R15954 VSS.n689 VSS.n686 152
R15955 VSS.n688 VSS.n687 152
R15956 VSS.n706 VSS.n700 152
R15957 VSS.n705 VSS.n704 152
R15958 VSS.n1037 VSS.n204 151.312
R15959 VSS.n1882 VSS.n1880 146.495
R15960 VSS.n1880 VSS.n1879 146.495
R15961 VSS.n1870 VSS.n1701 142.119
R15962 VSS.n1887 VSS.n1701 142.119
R15963 VSS.n1298 VSS.n1297 136.728
R15964 VSS.n1771 VSS.n1770 133.951
R15965 VSS.n1607 VSS.n1606 133.951
R15966 VSS.n1189 VSS.n1188 133.951
R15967 VSS.n1019 VSS.n1018 133.951
R15968 VSS.n668 VSS.n667 133.951
R15969 VSS.n587 VSS.n585 113.809
R15970 VSS.n1268 VSS.n199 109.144
R15971 VSS.n1778 VSS.n1777 104.172
R15972 VSS.n1785 VSS.n1784 104.172
R15973 VSS.n1792 VSS.n1791 104.172
R15974 VSS.n1799 VSS.n1798 104.172
R15975 VSS.n1811 VSS.n1805 104.172
R15976 VSS.n1818 VSS.n1817 104.172
R15977 VSS.n1827 VSS.n1721 104.172
R15978 VSS.n1829 VSS.n1717 104.172
R15979 VSS.n1859 VSS.n1840 104.172
R15980 VSS.n1857 VSS.n1841 104.172
R15981 VSS.n1614 VSS.n1613 104.172
R15982 VSS.n1621 VSS.n1620 104.172
R15983 VSS.n1628 VSS.n1627 104.172
R15984 VSS.n1635 VSS.n1634 104.172
R15985 VSS.n1647 VSS.n1641 104.172
R15986 VSS.n1654 VSS.n1653 104.172
R15987 VSS.n1663 VSS.n1557 104.172
R15988 VSS.n1665 VSS.n1553 104.172
R15989 VSS.n1695 VSS.n1676 104.172
R15990 VSS.n1693 VSS.n1677 104.172
R15991 VSS.n1307 VSS.n158 104.172
R15992 VSS.n1305 VSS.n159 104.172
R15993 VSS.n1196 VSS.n1195 104.172
R15994 VSS.n1203 VSS.n1202 104.172
R15995 VSS.n1242 VSS.n1211 104.172
R15996 VSS.n1240 VSS.n1212 104.172
R15997 VSS.n1230 VSS.n1216 104.172
R15998 VSS.n980 VSS.n979 104.172
R15999 VSS.n987 VSS.n986 104.172
R16000 VSS.n994 VSS.n993 104.172
R16001 VSS.n1005 VSS.n1001 104.172
R16002 VSS.n1003 VSS.n229 104.172
R16003 VSS.n629 VSS.n628 104.172
R16004 VSS.n636 VSS.n635 104.172
R16005 VSS.n643 VSS.n642 104.172
R16006 VSS.n658 VSS.n650 104.172
R16007 VSS.n656 VSS.n651 104.172
R16008 VSS.t6 VSS.n583 96.7682
R16009 VSS.n541 VSS.n512 91.5693
R16010 VSS.n579 VSS.n188 83.0979
R16011 VSS.n591 VSS.n586 83.0979
R16012 VSS.n591 VSS.n584 71.2233
R16013 VSS.n1036 VSS.n1035 69.3802
R16014 VSS.n162 VSS.t66 68.2323
R16015 VSS.n976 VSS.t64 68.2323
R16016 VSS.n625 VSS.t54 68.2323
R16017 VSS.t48 VSS.n1218 68.2319
R16018 VSS.n1705 VSS.n1702 64.0037
R16019 VSS.n1873 VSS.n1708 64.0037
R16020 VSS.n1756 VSS.t59 60.2505
R16021 VSS.n1923 VSS.t40 60.2505
R16022 VSS.n1591 VSS.t37 60.2505
R16023 VSS.n113 VSS.t57 60.2505
R16024 VSS.n125 VSS.t65 60.2505
R16025 VSS.n71 VSS.t43 60.2505
R16026 VSS.n1429 VSS.t34 60.2505
R16027 VSS.n1076 VSS.t55 60.2505
R16028 VSS.n1174 VSS.t45 60.2505
R16029 VSS.n281 VSS.t62 60.2505
R16030 VSS.n269 VSS.t32 60.2505
R16031 VSS.n702 VSS.t49 60.2505
R16032 VSS.n690 VSS.t52 60.2505
R16033 VSS.n587 VSS.n193 60.1048
R16034 VSS.n1278 VSS.n193 60.1048
R16035 VSS.n1257 VSS.n1038 58.0643
R16036 VSS.n580 VSS.n183 58.0643
R16037 VSS.n1886 VSS.n1702 57.9466
R16038 VSS.n1873 VSS.n1709 57.9466
R16039 VSS.t68 VSS.n1273 57.1814
R16040 VSS.n595 VSS.n582 53.5273
R16041 VSS.n1274 VSS.n187 48.3844
R16042 VSS.n1266 VSS.n200 48.3844
R16043 VSS.n211 VSS.n206 48.3844
R16044 VSS.n598 VSS.n185 45.2735
R16045 VSS.n1275 VSS.n189 44.6499
R16046 VSS.n189 VSS.n182 44.6499
R16047 VSS.n1283 VSS.n184 44.6499
R16048 VSS.n214 VSS.n213 44.6499
R16049 VSS.n1258 VSS.n215 44.6499
R16050 VSS.n1034 VSS.n207 44.6499
R16051 VSS.n1032 VSS.n207 44.6499
R16052 VSS.n1032 VSS.n205 44.6499
R16053 VSS.n205 VSS.n199 44.6499
R16054 VSS.n1761 VSS.n1752 44.3237
R16055 VSS.n1933 VSS.n1921 44.3237
R16056 VSS.n1601 VSS.n1589 44.3237
R16057 VSS.n131 VSS.n119 44.3237
R16058 VSS.n1434 VSS.n1425 44.3237
R16059 VSS.n1411 VSS.n1408 44.3237
R16060 VSS.n1419 VSS.n67 44.3237
R16061 VSS.n1390 VSS.n1387 44.3237
R16062 VSS.n1398 VSS.n109 44.3237
R16063 VSS.n1081 VSS.n1072 44.3237
R16064 VSS.n1179 VSS.n1170 44.3237
R16065 VSS.n275 VSS.n263 44.3237
R16066 VSS.n286 VSS.n277 44.3237
R16067 VSS.n696 VSS.n684 44.3237
R16068 VSS.n707 VSS.n698 44.3237
R16069 VSS.n1809 VSS.t61 35.3798
R16070 VSS.n1806 VSS.t61 35.3798
R16071 VSS.n1645 VSS.t39 35.3798
R16072 VSS.n1642 VSS.t39 35.3798
R16073 VSS.n164 VSS.t66 35.3798
R16074 VSS.n1220 VSS.t48 35.3798
R16075 VSS.t64 VSS.n975 35.3798
R16076 VSS.n623 VSS.t54 35.3798
R16077 VSS.n600 VSS.n582 33.9301
R16078 VSS.n1810 VSS.n1809 31.4488
R16079 VSS.n1806 VSS.n1725 31.4488
R16080 VSS.n1646 VSS.n1645 31.4488
R16081 VSS.n1642 VSS.n1561 31.4488
R16082 VSS.n165 VSS.n164 31.4488
R16083 VSS.n1221 VSS.n1220 31.4488
R16084 VSS.n975 VSS.n972 31.4488
R16085 VSS.n623 VSS.n621 31.4488
R16086 VSS.n1846 VSS.n1845 30.0212
R16087 VSS.n1682 VSS.n1681 30.0212
R16088 VSS.n1759 VSS.n1756 29.03
R16089 VSS.n1926 VSS.n1923 29.03
R16090 VSS.n1594 VSS.n1591 29.03
R16091 VSS.n125 VSS.n124 29.03
R16092 VSS.n1432 VSS.n1429 29.03
R16093 VSS.n1409 VSS.n71 29.03
R16094 VSS.n1417 VSS.n71 29.03
R16095 VSS.n1388 VSS.n113 29.03
R16096 VSS.n1396 VSS.n113 29.03
R16097 VSS.n1079 VSS.n1076 29.03
R16098 VSS.n1177 VSS.n1174 29.03
R16099 VSS.n269 VSS.n268 29.03
R16100 VSS.n284 VSS.n281 29.03
R16101 VSS.n690 VSS.n689 29.03
R16102 VSS.n705 VSS.n702 29.03
R16103 VSS.n1805 VSS.n1732 27.5177
R16104 VSS.n1819 VSS.n1818 27.5177
R16105 VSS.n1641 VSS.n1568 27.5177
R16106 VSS.n1655 VSS.n1654 27.5177
R16107 VSS.n1306 VSS.n1305 27.5177
R16108 VSS.n1231 VSS.n1230 27.5177
R16109 VSS.n980 VSS.n968 27.5177
R16110 VSS.n629 VSS.n617 27.5177
R16111 VSS.n200 VSS.n199 26.5914
R16112 VSS.n1032 VSS.n200 26.5914
R16113 VSS.n1034 VSS.n200 26.5914
R16114 VSS.n1798 VSS.n1736 23.5867
R16115 VSS.n1828 VSS.n1827 23.5867
R16116 VSS.n1634 VSS.n1572 23.5867
R16117 VSS.n1664 VSS.n1663 23.5867
R16118 VSS.n172 VSS.n158 23.5867
R16119 VSS.n1241 VSS.n1240 23.5867
R16120 VSS.n987 VSS.n964 23.5867
R16121 VSS.n636 VSS.n613 23.5867
R16122 VSS.n595 VSS.n584 23.5464
R16123 VSS.n599 VSS.n598 23.4593
R16124 VSS.n1263 VSS.n1262 22.9106
R16125 VSS.n1278 VSS.n1277 22.9106
R16126 VSS.n1771 VSS.n1748 21.6212
R16127 VSS.n1607 VSS.n1584 21.6212
R16128 VSS.n1189 VSS.n1166 21.6212
R16129 VSS.n1018 VSS.n1017 21.6212
R16130 VSS.n667 VSS.n505 21.6212
R16131 VSS.n1498 VSS.n1497 20.6425
R16132 VSS.n1110 VSS.n1109 20.6425
R16133 VSS.n1138 VSS.n1137 20.6425
R16134 VSS.n1332 VSS.n144 20.6425
R16135 VSS.n1468 VSS.n60 20.6425
R16136 VSS.n126 VSS.n121 20.4805
R16137 VSS.n270 VSS.n265 20.4805
R16138 VSS.n691 VSS.n686 20.4805
R16139 VSS.n1078 VSS.n1077 20.4803
R16140 VSS.n1176 VSS.n1175 20.4803
R16141 VSS.n1758 VSS.n1757 20.4802
R16142 VSS.n1928 VSS.n1927 20.4802
R16143 VSS.n1596 VSS.n1595 20.4802
R16144 VSS.n1431 VSS.n1430 20.4802
R16145 VSS.n283 VSS.n282 20.4802
R16146 VSS.n704 VSS.n703 20.4802
R16147 VSS.n1415 VSS.n72 19.9534
R16148 VSS.n1416 VSS.n1415 19.9534
R16149 VSS.n1394 VSS.n114 19.9534
R16150 VSS.n1395 VSS.n1394 19.9534
R16151 VSS.n1791 VSS.n1740 19.6557
R16152 VSS.n1839 VSS.n1717 19.6557
R16153 VSS.n1627 VSS.n1576 19.6557
R16154 VSS.n1675 VSS.n1553 19.6557
R16155 VSS.n1211 VSS.n1158 19.6557
R16156 VSS.n994 VSS.n960 19.6557
R16157 VSS.n643 VSS.n609 19.6557
R16158 VSS.n1262 VSS.n1261 19.4788
R16159 VSS.n1277 VSS.n1276 19.4788
R16160 VSS.n1966 VSS.n1907 19.4149
R16161 VSS.n314 VSS.n257 19.4149
R16162 VSS.n748 VSS.n491 19.4149
R16163 VSS.n1959 VSS.n1905 19.4144
R16164 VSS.n321 VSS.n255 19.4144
R16165 VSS.n741 VSS.n489 19.4144
R16166 VSS.n1971 VSS.n1908 19.3738
R16167 VSS.n309 VSS.n258 19.3738
R16168 VSS.n753 VSS.n492 19.3738
R16169 VSS.n1954 VSS.n1904 19.3733
R16170 VSS.n326 VSS.n254 19.3733
R16171 VSS.n736 VSS.n488 19.3733
R16172 VSS.n1976 VSS.n1909 19.3278
R16173 VSS.n1534 VSS.n1533 19.3273
R16174 VSS.n1948 VSS.n1903 19.3273
R16175 VSS.n331 VSS.n253 19.3273
R16176 VSS.n731 VSS.n487 19.3273
R16177 VSS.n1981 VSS.n1910 19.277
R16178 VSS.n2012 VSS.n2011 19.2765
R16179 VSS.n1996 VSS.n1995 19.2765
R16180 VSS.n1370 VSS.n137 19.2765
R16181 VSS.n1453 VSS.n55 19.2765
R16182 VSS.n96 VSS.n41 19.2765
R16183 VSS.n1099 VSS.n1068 19.2765
R16184 VSS.n893 VSS.n447 19.2765
R16185 VSS.n422 VSS.n421 19.2765
R16186 VSS.n921 VSS.n920 19.2765
R16187 VSS.n928 VSS.n392 19.2765
R16188 VSS.n367 VSS.n246 19.2765
R16189 VSS.n336 VSS.n252 19.2765
R16190 VSS.n250 VSS.n249 19.2765
R16191 VSS.n726 VSS.n486 19.2765
R16192 VSS.n778 VSS.n484 19.2765
R16193 VSS.n801 VSS.n800 19.2765
R16194 VSS.n820 VSS.n819 19.2765
R16195 VSS.n553 VSS.n517 19.2765
R16196 VSS.n1986 VSS.n1911 19.2214
R16197 VSS.n1540 VSS.n1526 19.2209
R16198 VSS.n1914 VSS.n1902 19.2209
R16199 VSS.n1375 VSS.n135 19.2209
R16200 VSS.n1448 VSS.n54 19.2209
R16201 VSS.n101 VSS.n53 19.2209
R16202 VSS.n1094 VSS.n1066 19.2209
R16203 VSS.n445 VSS.n444 19.2209
R16204 VSS.n427 VSS.n420 19.2209
R16205 VSS.n404 VSS.n403 19.2209
R16206 VSS.n390 VSS.n389 19.2209
R16207 VSS.n372 VSS.n245 19.2209
R16208 VSS.n341 VSS.n251 19.2209
R16209 VSS.n356 VSS.n260 19.2209
R16210 VSS.n721 VSS.n485 19.2209
R16211 VSS.n773 VSS.n494 19.2209
R16212 VSS.n789 VSS.n787 19.2209
R16213 VSS.n833 VSS.n832 19.2209
R16214 VSS.n564 VSS.n563 19.2209
R16215 VSS.n349 VSS.n261 19.161
R16216 VSS.n716 VSS.n495 19.161
R16217 VSS.n1993 VSS.n1992 19.1605
R16218 VSS.n1380 VSS.n133 19.1605
R16219 VSS.n1443 VSS.n59 19.1605
R16220 VSS.n106 VSS.n43 19.1605
R16221 VSS.n1089 VSS.n1067 19.1605
R16222 VSS.n898 VSS.n896 19.1605
R16223 VSS.n912 VSS.n911 19.1605
R16224 VSS.n407 VSS.n405 19.1605
R16225 VSS.n933 VSS.n931 19.1605
R16226 VSS.n947 VSS.n946 19.1605
R16227 VSS.n365 VSS.n364 19.1605
R16228 VSS.n785 VSS.n784 19.1605
R16229 VSS.n798 VSS.n797 19.1605
R16230 VSS.n837 VSS.n836 19.1605
R16231 VSS.n574 VSS.n573 19.1605
R16232 VSS.n1764 VSS.n1752 18.9796
R16233 VSS.n1933 VSS.n1932 18.9796
R16234 VSS.n1601 VSS.n1600 18.9796
R16235 VSS.n131 VSS.n130 18.9796
R16236 VSS.n1437 VSS.n1425 18.9796
R16237 VSS.n1408 VSS.n1407 18.9796
R16238 VSS.n1422 VSS.n67 18.9796
R16239 VSS.n1387 VSS.n1386 18.9796
R16240 VSS.n1401 VSS.n109 18.9796
R16241 VSS.n1084 VSS.n1072 18.9796
R16242 VSS.n1182 VSS.n1170 18.9796
R16243 VSS.n275 VSS.n274 18.9796
R16244 VSS.n289 VSS.n277 18.9796
R16245 VSS.n696 VSS.n695 18.9796
R16246 VSS.n710 VSS.n698 18.9796
R16247 VSS.n163 VSS.n162 18.7663
R16248 VSS.n976 VSS.n974 18.7663
R16249 VSS.n625 VSS.n624 18.7663
R16250 VSS.n1219 VSS.n1218 18.7661
R16251 VSS.n1146 VSS.n1128 18.5279
R16252 VSS.n1770 VSS.n1769 18.0631
R16253 VSS.n1606 VSS.n1605 18.0631
R16254 VSS.n1188 VSS.n1187 18.0631
R16255 VSS.n1020 VSS.n1019 18.0631
R16256 VSS.n669 VSS.n668 18.0631
R16257 VSS.n1778 VSS.n1744 17.6902
R16258 VSS.n1858 VSS.n1857 17.6902
R16259 VSS.n1614 VSS.n1580 17.6902
R16260 VSS.n1694 VSS.n1693 17.6902
R16261 VSS.n1196 VSS.n1162 17.6902
R16262 VSS.n1004 VSS.n1003 17.6902
R16263 VSS.n657 VSS.n656 17.6902
R16264 VSS.n1298 VSS.n171 16.9684
R16265 VSS.n1784 VSS.n1744 15.7246
R16266 VSS.n1859 VSS.n1858 15.7246
R16267 VSS.n1620 VSS.n1580 15.7246
R16268 VSS.n1695 VSS.n1694 15.7246
R16269 VSS.n1202 VSS.n1162 15.7246
R16270 VSS.n1005 VSS.n1004 15.7246
R16271 VSS.n658 VSS.n657 15.7246
R16272 VSS.n542 VSS.n541 15.4173
R16273 VSS.n1785 VSS.n1740 13.7591
R16274 VSS.n1840 VSS.n1839 13.7591
R16275 VSS.n1621 VSS.n1576 13.7591
R16276 VSS.n1676 VSS.n1675 13.7591
R16277 VSS.n1203 VSS.n1158 13.7591
R16278 VSS.n1001 VSS.n960 13.7591
R16279 VSS.n650 VSS.n609 13.7591
R16280 VSS.n1776 VSS.n1775 13.5534
R16281 VSS.n1783 VSS.n1782 13.5534
R16282 VSS.n1790 VSS.n1789 13.5534
R16283 VSS.n1797 VSS.n1796 13.5534
R16284 VSS.n1804 VSS.n1803 13.5534
R16285 VSS.n1808 VSS.n1807 13.5534
R16286 VSS.n1727 VSS.n1724 13.5534
R16287 VSS.n1826 VSS.n1825 13.5534
R16288 VSS.n1837 VSS.n1836 13.5534
R16289 VSS.n1861 VSS.n1860 13.5534
R16290 VSS.n1851 VSS.n1842 13.5534
R16291 VSS.n1612 VSS.n1611 13.5534
R16292 VSS.n1619 VSS.n1618 13.5534
R16293 VSS.n1626 VSS.n1625 13.5534
R16294 VSS.n1633 VSS.n1632 13.5534
R16295 VSS.n1640 VSS.n1639 13.5534
R16296 VSS.n1644 VSS.n1643 13.5534
R16297 VSS.n1563 VSS.n1560 13.5534
R16298 VSS.n1662 VSS.n1661 13.5534
R16299 VSS.n1673 VSS.n1672 13.5534
R16300 VSS.n1697 VSS.n1696 13.5534
R16301 VSS.n1687 VSS.n1678 13.5534
R16302 VSS.n1364 VSS.n141 13.5534
R16303 VSS.n1494 VSS.n1493 13.5534
R16304 VSS.n89 VSS.n44 13.5534
R16305 VSS.n1304 VSS.n1303 13.5534
R16306 VSS.n1107 VSS.n1106 13.5534
R16307 VSS.n1194 VSS.n1193 13.5534
R16308 VSS.n1201 VSS.n1200 13.5534
R16309 VSS.n1210 VSS.n1209 13.5534
R16310 VSS.n1229 VSS.n1228 13.5534
R16311 VSS.n304 VSS.n259 13.5534
R16312 VSS.n982 VSS.n981 13.5534
R16313 VSS.n989 VSS.n988 13.5534
R16314 VSS.n996 VSS.n995 13.5534
R16315 VSS.n1007 VSS.n1006 13.5534
R16316 VSS.n1015 VSS.n1014 13.5534
R16317 VSS.n631 VSS.n630 13.5534
R16318 VSS.n638 VSS.n637 13.5534
R16319 VSS.n645 VSS.n644 13.5534
R16320 VSS.n660 VSS.n659 13.5534
R16321 VSS.n653 VSS.n652 13.5534
R16322 VSS.n758 VSS.n493 13.5534
R16323 VSS.n535 VSS.n534 13.5534
R16324 VSS.n1362 VSS.n1361 13.177
R16325 VSS.n1471 VSS.n61 13.177
R16326 VSS.n52 VSS.n51 13.177
R16327 VSS.n174 VSS.n153 13.177
R16328 VSS.n1118 VSS.n1117 13.177
R16329 VSS.n1136 VSS.n1051 13.177
R16330 VSS.n1239 VSS.n1238 13.177
R16331 VSS.n2014 VSS.n2013 12.0077
R16332 VSS.n1994 VSS.n1919 12.0077
R16333 VSS.n1777 VSS.n1748 11.7936
R16334 VSS.n1845 VSS.n1841 11.7936
R16335 VSS.n1613 VSS.n1584 11.7936
R16336 VSS.n1681 VSS.n1677 11.7936
R16337 VSS.n1195 VSS.n1166 11.7936
R16338 VSS.n1017 VSS.n229 11.7936
R16339 VSS.n651 VSS.n505 11.7936
R16340 VSS.n1270 VSS.n1269 11.5947
R16341 VSS.n1038 VSS.n1036 11.3164
R16342 VSS.n1792 VSS.n1736 9.82809
R16343 VSS.n1829 VSS.n1828 9.82809
R16344 VSS.n1628 VSS.n1572 9.82809
R16345 VSS.n1665 VSS.n1664 9.82809
R16346 VSS.n1297 VSS.n172 9.82809
R16347 VSS.n1242 VSS.n1241 9.82809
R16348 VSS.n993 VSS.n964 9.82809
R16349 VSS.n642 VSS.n613 9.82809
R16350 VSS.n1539 VSS.n1538 9.3005
R16351 VSS.n1536 VSS.n1535 9.3005
R16352 VSS.n1529 VSS.n1528 9.3005
R16353 VSS.n1533 VSS.n1532 9.3005
R16354 VSS.n1540 VSS.n1525 9.3005
R16355 VSS.n2016 VSS.n2015 9.3005
R16356 VSS.n2011 VSS.n2010 9.3005
R16357 VSS.n1763 VSS.n1753 9.3005
R16358 VSS.n1765 VSS.n1764 9.3005
R16359 VSS.n1762 VSS.n1755 9.3005
R16360 VSS.n1762 VSS.n1761 9.3005
R16361 VSS.n1823 VSS.n1722 9.3005
R16362 VSS.n1814 VSS.n1728 9.3005
R16363 VSS.n1730 VSS.n1729 9.3005
R16364 VSS.n1735 VSS.n1734 9.3005
R16365 VSS.n1739 VSS.n1738 9.3005
R16366 VSS.n1743 VSS.n1742 9.3005
R16367 VSS.n1747 VSS.n1746 9.3005
R16368 VSS.n1751 VSS.n1750 9.3005
R16369 VSS.n1769 VSS.n1768 9.3005
R16370 VSS.n1773 VSS.n1772 9.3005
R16371 VSS.n1772 VSS.n1771 9.3005
R16372 VSS.n1775 VSS.n1774 9.3005
R16373 VSS.n1780 VSS.n1779 9.3005
R16374 VSS.n1779 VSS.n1778 9.3005
R16375 VSS.n1782 VSS.n1781 9.3005
R16376 VSS.n1787 VSS.n1786 9.3005
R16377 VSS.n1786 VSS.n1785 9.3005
R16378 VSS.n1789 VSS.n1788 9.3005
R16379 VSS.n1794 VSS.n1793 9.3005
R16380 VSS.n1793 VSS.n1792 9.3005
R16381 VSS.n1796 VSS.n1795 9.3005
R16382 VSS.n1801 VSS.n1800 9.3005
R16383 VSS.n1800 VSS.n1799 9.3005
R16384 VSS.n1803 VSS.n1802 9.3005
R16385 VSS.n1813 VSS.n1812 9.3005
R16386 VSS.n1812 VSS.n1811 9.3005
R16387 VSS.n1816 VSS.n1815 9.3005
R16388 VSS.n1817 VSS.n1816 9.3005
R16389 VSS.n1727 VSS.n1723 9.3005
R16390 VSS.n1822 VSS.n1821 9.3005
R16391 VSS.n1821 VSS.n1721 9.3005
R16392 VSS.n1825 VSS.n1824 9.3005
R16393 VSS.n1831 VSS.n1830 9.3005
R16394 VSS.n1830 VSS.n1829 9.3005
R16395 VSS.n1836 VSS.n1835 9.3005
R16396 VSS.n1715 VSS.n1713 9.3005
R16397 VSS.n1840 VSS.n1715 9.3005
R16398 VSS.n1848 VSS.n1847 9.3005
R16399 VSS.n1851 VSS.n1850 9.3005
R16400 VSS.n1856 VSS.n1855 9.3005
R16401 VSS.n1857 VSS.n1856 9.3005
R16402 VSS.n1861 VSS.n1714 9.3005
R16403 VSS.n1931 VSS.n1930 9.3005
R16404 VSS.n1932 VSS.n1920 9.3005
R16405 VSS.n1929 VSS.n1922 9.3005
R16406 VSS.n1922 VSS.n1921 9.3005
R16407 VSS.n1955 VSS.n1943 9.3005
R16408 VSS.n1960 VSS.n1942 9.3005
R16409 VSS.n1965 VSS.n1941 9.3005
R16410 VSS.n1970 VSS.n1940 9.3005
R16411 VSS.n1975 VSS.n1939 9.3005
R16412 VSS.n1980 VSS.n1938 9.3005
R16413 VSS.n1985 VSS.n1937 9.3005
R16414 VSS.n1990 VSS.n1936 9.3005
R16415 VSS.n1992 VSS.n1991 9.3005
R16416 VSS.n1989 VSS.n1988 9.3005
R16417 VSS.n1987 VSS.n1986 9.3005
R16418 VSS.n1984 VSS.n1983 9.3005
R16419 VSS.n1982 VSS.n1981 9.3005
R16420 VSS.n1979 VSS.n1978 9.3005
R16421 VSS.n1977 VSS.n1976 9.3005
R16422 VSS.n1974 VSS.n1973 9.3005
R16423 VSS.n1972 VSS.n1971 9.3005
R16424 VSS.n1969 VSS.n1968 9.3005
R16425 VSS.n1967 VSS.n1966 9.3005
R16426 VSS.n1964 VSS.n1963 9.3005
R16427 VSS.n1962 VSS.n1961 9.3005
R16428 VSS.n1959 VSS.n1958 9.3005
R16429 VSS.n1957 VSS.n1956 9.3005
R16430 VSS.n1954 VSS.n1953 9.3005
R16431 VSS.n1951 VSS.n1950 9.3005
R16432 VSS.n1948 VSS.n1947 9.3005
R16433 VSS.n1897 VSS.n1546 9.3005
R16434 VSS.n1996 VSS.n1896 9.3005
R16435 VSS.n1901 VSS.n1900 9.3005
R16436 VSS.n1915 VSS.n1914 9.3005
R16437 VSS.n1918 VSS.n1917 9.3005
R16438 VSS.n1599 VSS.n1598 9.3005
R16439 VSS.n1600 VSS.n1588 9.3005
R16440 VSS.n1597 VSS.n1590 9.3005
R16441 VSS.n1590 VSS.n1589 9.3005
R16442 VSS.n1659 VSS.n1558 9.3005
R16443 VSS.n1650 VSS.n1564 9.3005
R16444 VSS.n1566 VSS.n1565 9.3005
R16445 VSS.n1571 VSS.n1570 9.3005
R16446 VSS.n1575 VSS.n1574 9.3005
R16447 VSS.n1579 VSS.n1578 9.3005
R16448 VSS.n1583 VSS.n1582 9.3005
R16449 VSS.n1587 VSS.n1586 9.3005
R16450 VSS.n1605 VSS.n1604 9.3005
R16451 VSS.n1609 VSS.n1608 9.3005
R16452 VSS.n1608 VSS.n1607 9.3005
R16453 VSS.n1611 VSS.n1610 9.3005
R16454 VSS.n1616 VSS.n1615 9.3005
R16455 VSS.n1615 VSS.n1614 9.3005
R16456 VSS.n1618 VSS.n1617 9.3005
R16457 VSS.n1623 VSS.n1622 9.3005
R16458 VSS.n1622 VSS.n1621 9.3005
R16459 VSS.n1625 VSS.n1624 9.3005
R16460 VSS.n1630 VSS.n1629 9.3005
R16461 VSS.n1629 VSS.n1628 9.3005
R16462 VSS.n1632 VSS.n1631 9.3005
R16463 VSS.n1637 VSS.n1636 9.3005
R16464 VSS.n1636 VSS.n1635 9.3005
R16465 VSS.n1639 VSS.n1638 9.3005
R16466 VSS.n1649 VSS.n1648 9.3005
R16467 VSS.n1648 VSS.n1647 9.3005
R16468 VSS.n1652 VSS.n1651 9.3005
R16469 VSS.n1653 VSS.n1652 9.3005
R16470 VSS.n1563 VSS.n1559 9.3005
R16471 VSS.n1658 VSS.n1657 9.3005
R16472 VSS.n1657 VSS.n1557 9.3005
R16473 VSS.n1661 VSS.n1660 9.3005
R16474 VSS.n1692 VSS.n1691 9.3005
R16475 VSS.n1693 VSS.n1692 9.3005
R16476 VSS.n1667 VSS.n1666 9.3005
R16477 VSS.n1666 VSS.n1665 9.3005
R16478 VSS.n1672 VSS.n1671 9.3005
R16479 VSS.n1551 VSS.n1549 9.3005
R16480 VSS.n1676 VSS.n1551 9.3005
R16481 VSS.n1697 VSS.n1550 9.3005
R16482 VSS.n1687 VSS.n1686 9.3005
R16483 VSS.n1684 VSS.n1683 9.3005
R16484 VSS.n1889 VSS.n1888 9.3005
R16485 VSS.n1462 VSS.n1460 9.3005
R16486 VSS.n1475 VSS.n1472 9.3005
R16487 VSS.n1493 VSS.n1492 9.3005
R16488 VSS.n1474 VSS.n1473 9.3005
R16489 VSS.n1477 VSS.n1476 9.3005
R16490 VSS.n1464 VSS.n1463 9.3005
R16491 VSS.n1444 VSS.n66 9.3005
R16492 VSS.n1449 VSS.n65 9.3005
R16493 VSS.n1454 VSS.n64 9.3005
R16494 VSS.n1456 VSS.n1455 9.3005
R16495 VSS.n1453 VSS.n1452 9.3005
R16496 VSS.n1451 VSS.n1450 9.3005
R16497 VSS.n1448 VSS.n1447 9.3005
R16498 VSS.n1446 VSS.n1445 9.3005
R16499 VSS.n1443 VSS.n1442 9.3005
R16500 VSS.n87 VSS.n86 9.3005
R16501 VSS.n48 VSS.n47 9.3005
R16502 VSS.n85 VSS.n84 9.3005
R16503 VSS.n90 VSS.n89 9.3005
R16504 VSS.n46 VSS.n36 9.3005
R16505 VSS.n50 VSS.n49 9.3005
R16506 VSS.n104 VSS.n103 9.3005
R16507 VSS.n100 VSS.n77 9.3005
R16508 VSS.n102 VSS.n101 9.3005
R16509 VSS.n99 VSS.n98 9.3005
R16510 VSS.n97 VSS.n96 9.3005
R16511 VSS.n94 VSS.n93 9.3005
R16512 VSS.n95 VSS.n78 9.3005
R16513 VSS.n105 VSS.n76 9.3005
R16514 VSS.n107 VSS.n106 9.3005
R16515 VSS.n74 VSS.n73 9.3005
R16516 VSS.n1421 VSS.n68 9.3005
R16517 VSS.n1436 VSS.n1426 9.3005
R16518 VSS.n1438 VSS.n1437 9.3005
R16519 VSS.n1435 VSS.n1428 9.3005
R16520 VSS.n1435 VSS.n1434 9.3005
R16521 VSS.n1407 VSS.n1406 9.3005
R16522 VSS.n1413 VSS.n1412 9.3005
R16523 VSS.n1412 VSS.n1411 9.3005
R16524 VSS.n1420 VSS.n70 9.3005
R16525 VSS.n1420 VSS.n1419 9.3005
R16526 VSS.n1423 VSS.n1422 9.3005
R16527 VSS.n130 VSS.n118 9.3005
R16528 VSS.n129 VSS.n128 9.3005
R16529 VSS.n127 VSS.n120 9.3005
R16530 VSS.n120 VSS.n119 9.3005
R16531 VSS.n1386 VSS.n1385 9.3005
R16532 VSS.n1392 VSS.n1391 9.3005
R16533 VSS.n1391 VSS.n1390 9.3005
R16534 VSS.n116 VSS.n115 9.3005
R16535 VSS.n1399 VSS.n112 9.3005
R16536 VSS.n1399 VSS.n1398 9.3005
R16537 VSS.n1402 VSS.n1401 9.3005
R16538 VSS.n1400 VSS.n110 9.3005
R16539 VSS.n1379 VSS.n134 9.3005
R16540 VSS.n1374 VSS.n136 9.3005
R16541 VSS.n1369 VSS.n138 9.3005
R16542 VSS.n1368 VSS.n1367 9.3005
R16543 VSS.n1371 VSS.n1370 9.3005
R16544 VSS.n1373 VSS.n1372 9.3005
R16545 VSS.n1376 VSS.n1375 9.3005
R16546 VSS.n1378 VSS.n1377 9.3005
R16547 VSS.n1381 VSS.n1380 9.3005
R16548 VSS.n1355 VSS.n1351 9.3005
R16549 VSS.n1329 VSS.n1328 9.3005
R16550 VSS.n1352 VSS.n141 9.3005
R16551 VSS.n1357 VSS.n1356 9.3005
R16552 VSS.n1331 VSS.n1330 9.3005
R16553 VSS.n148 VSS.n146 9.3005
R16554 VSS.n168 VSS.n167 9.3005
R16555 VSS.n167 VSS.n159 9.3005
R16556 VSS.n169 VSS.n161 9.3005
R16557 VSS.n1311 VSS.n1310 9.3005
R16558 VSS.n1294 VSS.n173 9.3005
R16559 VSS.n1296 VSS.n1295 9.3005
R16560 VSS.n1297 VSS.n1296 9.3005
R16561 VSS.n171 VSS.n170 9.3005
R16562 VSS.n1303 VSS.n1302 9.3005
R16563 VSS.n1308 VSS.n157 9.3005
R16564 VSS.n1308 VSS.n1307 9.3005
R16565 VSS.n1309 VSS.n155 9.3005
R16566 VSS.n1082 VSS.n1075 9.3005
R16567 VSS.n1082 VSS.n1081 9.3005
R16568 VSS.n1085 VSS.n1084 9.3005
R16569 VSS.n1083 VSS.n1073 9.3005
R16570 VSS.n1090 VSS.n1071 9.3005
R16571 VSS.n1095 VSS.n1070 9.3005
R16572 VSS.n1100 VSS.n1069 9.3005
R16573 VSS.n1099 VSS.n1098 9.3005
R16574 VSS.n1097 VSS.n1096 9.3005
R16575 VSS.n1094 VSS.n1093 9.3005
R16576 VSS.n1092 VSS.n1091 9.3005
R16577 VSS.n1089 VSS.n1088 9.3005
R16578 VSS.n1102 VSS.n1101 9.3005
R16579 VSS.n1123 VSS.n1122 9.3005
R16580 VSS.n1106 VSS.n1058 9.3005
R16581 VSS.n1114 VSS.n1111 9.3005
R16582 VSS.n1113 VSS.n1112 9.3005
R16583 VSS.n1116 VSS.n1115 9.3005
R16584 VSS.n1121 VSS.n1062 9.3005
R16585 VSS.n1130 VSS.n1052 9.3005
R16586 VSS.n1144 VSS.n1143 9.3005
R16587 VSS.n1142 VSS.n1141 9.3005
R16588 VSS.n1147 VSS.n1146 9.3005
R16589 VSS.n1134 VSS.n1133 9.3005
R16590 VSS.n1132 VSS.n1131 9.3005
R16591 VSS.n1225 VSS.n1217 9.3005
R16592 VSS.n1224 VSS.n1223 9.3005
R16593 VSS.n1223 VSS.n1216 9.3005
R16594 VSS.n1180 VSS.n1173 9.3005
R16595 VSS.n1180 VSS.n1179 9.3005
R16596 VSS.n1183 VSS.n1182 9.3005
R16597 VSS.n1181 VSS.n1171 9.3005
R16598 VSS.n1169 VSS.n1168 9.3005
R16599 VSS.n1165 VSS.n1164 9.3005
R16600 VSS.n1161 VSS.n1160 9.3005
R16601 VSS.n1205 VSS.n1204 9.3005
R16602 VSS.n1204 VSS.n1203 9.3005
R16603 VSS.n1200 VSS.n1199 9.3005
R16604 VSS.n1198 VSS.n1197 9.3005
R16605 VSS.n1197 VSS.n1196 9.3005
R16606 VSS.n1193 VSS.n1192 9.3005
R16607 VSS.n1191 VSS.n1190 9.3005
R16608 VSS.n1190 VSS.n1189 9.3005
R16609 VSS.n1187 VSS.n1186 9.3005
R16610 VSS.n1245 VSS.n1244 9.3005
R16611 VSS.n1209 VSS.n1045 9.3005
R16612 VSS.n1235 VSS.n1214 9.3005
R16613 VSS.n1228 VSS.n1227 9.3005
R16614 VSS.n1234 VSS.n1233 9.3005
R16615 VSS.n1233 VSS.n1212 9.3005
R16616 VSS.n1237 VSS.n1236 9.3005
R16617 VSS.n1243 VSS.n1156 9.3005
R16618 VSS.n1243 VSS.n1242 9.3005
R16619 VSS.n446 VSS.n437 9.3005
R16620 VSS.n901 VSS.n900 9.3005
R16621 VSS.n893 VSS.n892 9.3005
R16622 VSS.n898 VSS.n897 9.3005
R16623 VSS.n444 VSS.n440 9.3005
R16624 VSS.n434 VSS.n422 9.3005
R16625 VSS.n425 VSS.n423 9.3005
R16626 VSS.n913 VSS.n912 9.3005
R16627 VSS.n430 VSS.n429 9.3005
R16628 VSS.n428 VSS.n427 9.3005
R16629 VSS.n407 VSS.n406 9.3005
R16630 VSS.n410 VSS.n409 9.3005
R16631 VSS.n403 VSS.n400 9.3005
R16632 VSS.n919 VSS.n918 9.3005
R16633 VSS.n921 VSS.n396 9.3005
R16634 VSS.n928 VSS.n927 9.3005
R16635 VSS.n391 VSS.n382 9.3005
R16636 VSS.n389 VSS.n385 9.3005
R16637 VSS.n936 VSS.n935 9.3005
R16638 VSS.n933 VSS.n932 9.3005
R16639 VSS.n379 VSS.n367 9.3005
R16640 VSS.n370 VSS.n368 9.3005
R16641 VSS.n948 VSS.n947 9.3005
R16642 VSS.n375 VSS.n374 9.3005
R16643 VSS.n373 VSS.n372 9.3005
R16644 VSS.n274 VSS.n262 9.3005
R16645 VSS.n273 VSS.n272 9.3005
R16646 VSS.n271 VSS.n264 9.3005
R16647 VSS.n264 VSS.n263 9.3005
R16648 VSS.n290 VSS.n289 9.3005
R16649 VSS.n287 VSS.n280 9.3005
R16650 VSS.n287 VSS.n286 9.3005
R16651 VSS.n288 VSS.n278 9.3005
R16652 VSS.n346 VSS.n345 9.3005
R16653 VSS.n340 VSS.n293 9.3005
R16654 VSS.n335 VSS.n294 9.3005
R16655 VSS.n330 VSS.n295 9.3005
R16656 VSS.n325 VSS.n296 9.3005
R16657 VSS.n320 VSS.n297 9.3005
R16658 VSS.n315 VSS.n298 9.3005
R16659 VSS.n310 VSS.n299 9.3005
R16660 VSS.n305 VSS.n300 9.3005
R16661 VSS.n304 VSS.n303 9.3005
R16662 VSS.n307 VSS.n306 9.3005
R16663 VSS.n309 VSS.n308 9.3005
R16664 VSS.n312 VSS.n311 9.3005
R16665 VSS.n314 VSS.n313 9.3005
R16666 VSS.n317 VSS.n316 9.3005
R16667 VSS.n319 VSS.n318 9.3005
R16668 VSS.n322 VSS.n321 9.3005
R16669 VSS.n324 VSS.n323 9.3005
R16670 VSS.n327 VSS.n326 9.3005
R16671 VSS.n329 VSS.n328 9.3005
R16672 VSS.n332 VSS.n331 9.3005
R16673 VSS.n334 VSS.n333 9.3005
R16674 VSS.n337 VSS.n336 9.3005
R16675 VSS.n339 VSS.n338 9.3005
R16676 VSS.n342 VSS.n341 9.3005
R16677 VSS.n344 VSS.n343 9.3005
R16678 VSS.n347 VSS.n261 9.3005
R16679 VSS.n302 VSS.n301 9.3005
R16680 VSS.n364 VSS.n363 9.3005
R16681 VSS.n361 VSS.n360 9.3005
R16682 VSS.n357 VSS.n356 9.3005
R16683 VSS.n354 VSS.n353 9.3005
R16684 VSS.n249 VSS.n238 9.3005
R16685 VSS.n247 VSS.n236 9.3005
R16686 VSS.n971 VSS.n970 9.3005
R16687 VSS.n967 VSS.n966 9.3005
R16688 VSS.n978 VSS.n977 9.3005
R16689 VSS.n979 VSS.n978 9.3005
R16690 VSS.n983 VSS.n982 9.3005
R16691 VSS.n985 VSS.n984 9.3005
R16692 VSS.n986 VSS.n985 9.3005
R16693 VSS.n990 VSS.n989 9.3005
R16694 VSS.n992 VSS.n991 9.3005
R16695 VSS.n993 VSS.n992 9.3005
R16696 VSS.n997 VSS.n996 9.3005
R16697 VSS.n963 VSS.n962 9.3005
R16698 VSS.n1008 VSS.n1007 9.3005
R16699 VSS.n1020 VSS.n225 9.3005
R16700 VSS.n1011 VSS.n227 9.3005
R16701 VSS.n1018 VSS.n227 9.3005
R16702 VSS.n1014 VSS.n1013 9.3005
R16703 VSS.n1002 VSS.n232 9.3005
R16704 VSS.n1003 VSS.n1002 9.3005
R16705 VSS.n1000 VSS.n999 9.3005
R16706 VSS.n1001 VSS.n1000 9.3005
R16707 VSS.n998 VSS.n961 9.3005
R16708 VSS.n620 VSS.n619 9.3005
R16709 VSS.n616 VSS.n615 9.3005
R16710 VSS.n627 VSS.n626 9.3005
R16711 VSS.n628 VSS.n627 9.3005
R16712 VSS.n632 VSS.n631 9.3005
R16713 VSS.n634 VSS.n633 9.3005
R16714 VSS.n635 VSS.n634 9.3005
R16715 VSS.n639 VSS.n638 9.3005
R16716 VSS.n641 VSS.n640 9.3005
R16717 VSS.n642 VSS.n641 9.3005
R16718 VSS.n646 VSS.n645 9.3005
R16719 VSS.n612 VSS.n611 9.3005
R16720 VSS.n661 VSS.n660 9.3005
R16721 VSS.n655 VSS.n509 9.3005
R16722 VSS.n656 VSS.n655 9.3005
R16723 VSS.n670 VSS.n669 9.3005
R16724 VSS.n666 VSS.n665 9.3005
R16725 VSS.n667 VSS.n666 9.3005
R16726 VSS.n653 VSS.n507 9.3005
R16727 VSS.n649 VSS.n648 9.3005
R16728 VSS.n650 VSS.n649 9.3005
R16729 VSS.n647 VSS.n610 9.3005
R16730 VSS.n695 VSS.n683 9.3005
R16731 VSS.n694 VSS.n693 9.3005
R16732 VSS.n692 VSS.n685 9.3005
R16733 VSS.n685 VSS.n684 9.3005
R16734 VSS.n711 VSS.n710 9.3005
R16735 VSS.n708 VSS.n701 9.3005
R16736 VSS.n708 VSS.n707 9.3005
R16737 VSS.n709 VSS.n699 9.3005
R16738 VSS.n717 VSS.n682 9.3005
R16739 VSS.n722 VSS.n681 9.3005
R16740 VSS.n727 VSS.n680 9.3005
R16741 VSS.n732 VSS.n679 9.3005
R16742 VSS.n737 VSS.n678 9.3005
R16743 VSS.n742 VSS.n677 9.3005
R16744 VSS.n747 VSS.n676 9.3005
R16745 VSS.n752 VSS.n675 9.3005
R16746 VSS.n757 VSS.n674 9.3005
R16747 VSS.n759 VSS.n758 9.3005
R16748 VSS.n756 VSS.n755 9.3005
R16749 VSS.n754 VSS.n753 9.3005
R16750 VSS.n751 VSS.n750 9.3005
R16751 VSS.n749 VSS.n748 9.3005
R16752 VSS.n746 VSS.n745 9.3005
R16753 VSS.n744 VSS.n743 9.3005
R16754 VSS.n741 VSS.n740 9.3005
R16755 VSS.n739 VSS.n738 9.3005
R16756 VSS.n736 VSS.n735 9.3005
R16757 VSS.n734 VSS.n733 9.3005
R16758 VSS.n731 VSS.n730 9.3005
R16759 VSS.n729 VSS.n728 9.3005
R16760 VSS.n726 VSS.n725 9.3005
R16761 VSS.n724 VSS.n723 9.3005
R16762 VSS.n721 VSS.n720 9.3005
R16763 VSS.n719 VSS.n718 9.3005
R16764 VSS.n716 VSS.n715 9.3005
R16765 VSS.n761 VSS.n760 9.3005
R16766 VSS.n784 VSS.n783 9.3005
R16767 VSS.n770 VSS.n769 9.3005
R16768 VSS.n773 VSS.n772 9.3005
R16769 VSS.n776 VSS.n775 9.3005
R16770 VSS.n779 VSS.n778 9.3005
R16771 VSS.n763 VSS.n762 9.3005
R16772 VSS.n802 VSS.n801 9.3005
R16773 VSS.n482 VSS.n475 9.3005
R16774 VSS.n794 VSS.n793 9.3005
R16775 VSS.n797 VSS.n796 9.3005
R16776 VSS.n790 VSS.n789 9.3005
R16777 VSS.n838 VSS.n837 9.3005
R16778 VSS.n821 VSS.n816 9.3005
R16779 VSS.n832 VSS.n831 9.3005
R16780 VSS.n825 VSS.n824 9.3005
R16781 VSS.n819 VSS.n812 9.3005
R16782 VSS.n539 VSS.n538 9.3005
R16783 VSS.n542 VSS.n525 9.3005
R16784 VSS.n549 VSS.n521 9.3005
R16785 VSS.n573 VSS.n511 9.3005
R16786 VSS.n570 VSS.n513 9.3005
R16787 VSS.n565 VSS.n564 9.3005
R16788 VSS.n561 VSS.n560 9.3005
R16789 VSS.n554 VSS.n553 9.3005
R16790 VSS.n551 VSS.n550 9.3005
R16791 VSS.n551 VSS.n512 9.3005
R16792 VSS.n534 VSS.n533 9.3005
R16793 VSS.n540 VSS.n524 9.3005
R16794 VSS.n540 VSS.n512 9.3005
R16795 VSS.n206 VSS.n199 9.3005
R16796 VSS.n1032 VSS.n206 9.3005
R16797 VSS.n1034 VSS.n206 9.3005
R16798 VSS.n601 VSS.n600 9.3005
R16799 VSS.n600 VSS.n599 9.3005
R16800 VSS.n186 VSS.n184 9.19092
R16801 VSS.n1258 VSS.n203 9.19092
R16802 VSS.n1261 VSS.n1260 9.01392
R16803 VSS.n1258 VSS.n1257 9.01392
R16804 VSS.n1252 VSS.n214 9.01392
R16805 VSS.n184 VSS.n183 9.01392
R16806 VSS.n1285 VSS.n182 9.01392
R16807 VSS.n1276 VSS.n1275 9.01392
R16808 VSS.n1495 VSS.n58 8.80469
R16809 VSS.n1496 VSS.n39 8.80469
R16810 VSS.n1363 VSS.n142 8.80469
R16811 VSS.n1119 VSS.n1064 8.80469
R16812 VSS.n1139 VSS.n1135 8.80469
R16813 VSS.n1495 VSS.n57 8.7709
R16814 VSS.n1496 VSS.n42 8.7709
R16815 VSS.n1363 VSS.n143 8.7709
R16816 VSS.n1120 VSS.n1119 8.7709
R16817 VSS.n1140 VSS.n1139 8.7709
R16818 VSS.n1415 VSS.n71 8.76429
R16819 VSS.n1394 VSS.n113 8.76429
R16820 VSS.n1495 VSS.n56 8.73737
R16821 VSS.n1496 VSS.n40 8.73737
R16822 VSS.n1363 VSS.n139 8.73737
R16823 VSS.n1119 VSS.n1065 8.73737
R16824 VSS.n366 VSS.n248 8.73737
R16825 VSS.n786 VSS.n483 8.73737
R16826 VSS.n1885 VSS.n1704 8.50504
R16827 VSS.n1275 VSS.n185 8.44701
R16828 VSS.n1760 VSS.n1759 8.21641
R16829 VSS.n1926 VSS.n1925 8.21641
R16830 VSS.n1594 VSS.n1593 8.21641
R16831 VSS.n124 VSS.n123 8.21641
R16832 VSS.n1433 VSS.n1432 8.21641
R16833 VSS.n1410 VSS.n1409 8.21641
R16834 VSS.n1418 VSS.n1417 8.21641
R16835 VSS.n1389 VSS.n1388 8.21641
R16836 VSS.n1397 VSS.n1396 8.21641
R16837 VSS.n1080 VSS.n1079 8.21641
R16838 VSS.n1178 VSS.n1177 8.21641
R16839 VSS.n268 VSS.n267 8.21641
R16840 VSS.n285 VSS.n284 8.21641
R16841 VSS.n689 VSS.n688 8.21641
R16842 VSS.n706 VSS.n705 8.21641
R16843 VSS.n1269 VSS.n198 8.16282
R16844 VSS.n1994 VSS.n1905 8.139
R16845 VSS.n366 VSS.n255 8.139
R16846 VSS.n786 VSS.n489 8.139
R16847 VSS.n1994 VSS.n1907 8.13855
R16848 VSS.n366 VSS.n257 8.13855
R16849 VSS.n786 VSS.n491 8.13855
R16850 VSS.n1994 VSS.n1904 8.11104
R16851 VSS.n366 VSS.n254 8.11104
R16852 VSS.n786 VSS.n488 8.11104
R16853 VSS.n1994 VSS.n1908 8.11059
R16854 VSS.n366 VSS.n258 8.11059
R16855 VSS.n786 VSS.n492 8.11059
R16856 VSS.n2013 VSS.n1534 8.08351
R16857 VSS.n1994 VSS.n1903 8.08351
R16858 VSS.n366 VSS.n253 8.08351
R16859 VSS.n786 VSS.n487 8.08351
R16860 VSS.n1994 VSS.n1909 8.08305
R16861 VSS.n2013 VSS.n2012 8.05639
R16862 VSS.n1995 VSS.n1994 8.05639
R16863 VSS.n1495 VSS.n55 8.05639
R16864 VSS.n1496 VSS.n41 8.05639
R16865 VSS.n1363 VSS.n137 8.05639
R16866 VSS.n1119 VSS.n1068 8.05639
R16867 VSS.n895 VSS.n447 8.05639
R16868 VSS.n910 VSS.n421 8.05639
R16869 VSS.n920 VSS.n397 8.05639
R16870 VSS.n930 VSS.n392 8.05639
R16871 VSS.n945 VSS.n246 8.05639
R16872 VSS.n366 VSS.n252 8.05639
R16873 VSS.n366 VSS.n250 8.05639
R16874 VSS.n786 VSS.n486 8.05639
R16875 VSS.n786 VSS.n484 8.05639
R16876 VSS.n800 VSS.n799 8.05639
R16877 VSS.n835 VSS.n820 8.05639
R16878 VSS.n517 VSS.n512 8.05639
R16879 VSS.n1994 VSS.n1910 8.05594
R16880 VSS.n2013 VSS.n1526 8.02969
R16881 VSS.n1994 VSS.n1902 8.02969
R16882 VSS.n1495 VSS.n54 8.02969
R16883 VSS.n1496 VSS.n53 8.02969
R16884 VSS.n1363 VSS.n135 8.02969
R16885 VSS.n1119 VSS.n1066 8.02969
R16886 VSS.n895 VSS.n445 8.02969
R16887 VSS.n910 VSS.n420 8.02969
R16888 VSS.n404 VSS.n397 8.02969
R16889 VSS.n930 VSS.n390 8.02969
R16890 VSS.n945 VSS.n245 8.02969
R16891 VSS.n366 VSS.n260 8.02969
R16892 VSS.n366 VSS.n251 8.02969
R16893 VSS.n786 VSS.n494 8.02969
R16894 VSS.n786 VSS.n485 8.02969
R16895 VSS.n799 VSS.n787 8.02969
R16896 VSS.n835 VSS.n833 8.02969
R16897 VSS.n563 VSS.n512 8.02969
R16898 VSS.n1994 VSS.n1911 8.02924
R16899 VSS.n1994 VSS.n1993 8.00339
R16900 VSS.n1363 VSS.n133 8.00339
R16901 VSS.n1495 VSS.n59 8.00339
R16902 VSS.n1496 VSS.n43 8.00339
R16903 VSS.n1119 VSS.n1067 8.00339
R16904 VSS.n896 VSS.n895 8.00339
R16905 VSS.n911 VSS.n910 8.00339
R16906 VSS.n405 VSS.n397 8.00339
R16907 VSS.n931 VSS.n930 8.00339
R16908 VSS.n946 VSS.n945 8.00339
R16909 VSS.n366 VSS.n365 8.00339
R16910 VSS.n786 VSS.n785 8.00339
R16911 VSS.n799 VSS.n798 8.00339
R16912 VSS.n836 VSS.n835 8.00339
R16913 VSS.n574 VSS.n512 8.00339
R16914 VSS.n366 VSS.n349 8.00293
R16915 VSS.n786 VSS.n495 8.00293
R16916 VSS.n1282 VSS.n182 7.69718
R16917 VSS.n1260 VSS.n201 7.69718
R16918 VSS.n214 VSS.n202 7.69718
R16919 VSS.n600 VSS.n188 7.3129
R16920 VSS.n592 VSS.n585 6.95702
R16921 VSS.n581 VSS.n580 6.95702
R16922 VSS.n126 VSS.n125 6.92242
R16923 VSS.n270 VSS.n269 6.92242
R16924 VSS.n691 VSS.n690 6.92242
R16925 VSS.n1928 VSS.n1923 6.92012
R16926 VSS.n1596 VSS.n1591 6.92012
R16927 VSS.n1430 VSS.n1429 6.92012
R16928 VSS.n282 VSS.n281 6.92012
R16929 VSS.n703 VSS.n702 6.92012
R16930 VSS.n1757 VSS.n1756 6.92011
R16931 VSS.n1077 VSS.n1076 6.92007
R16932 VSS.n1175 VSS.n1174 6.92007
R16933 VSS.n199 VSS.n198 6.81049
R16934 VSS.n1032 VSS.n1031 6.81049
R16935 VSS.n1035 VSS.n1034 6.81049
R16936 VSS.n1019 VSS.n228 6.55106
R16937 VSS.n668 VSS.n504 6.55006
R16938 VSS.n1188 VSS.n1185 6.43466
R16939 VSS.n1770 VSS.n1767 6.43466
R16940 VSS.n1606 VSS.n1603 6.43466
R16941 VSS.n834 VSS.n814 6.4167
R16942 VSS.n1528 VSS.n1527 6.11953
R16943 VSS.n1803 VSS.n1730 6.02403
R16944 VSS.n1808 VSS.n1731 6.02403
R16945 VSS.n1807 VSS.n1726 6.02403
R16946 VSS.n1728 VSS.n1727 6.02403
R16947 VSS.n1966 VSS.n1965 6.02403
R16948 VSS.n1960 VSS.n1959 6.02403
R16949 VSS.n1639 VSS.n1566 6.02403
R16950 VSS.n1644 VSS.n1567 6.02403
R16951 VSS.n1643 VSS.n1562 6.02403
R16952 VSS.n1564 VSS.n1563 6.02403
R16953 VSS.n1303 VSS.n161 6.02403
R16954 VSS.n166 VSS.n163 6.02403
R16955 VSS.n1228 VSS.n1217 6.02403
R16956 VSS.n1222 VSS.n1219 6.02403
R16957 VSS.n321 VSS.n320 6.02403
R16958 VSS.n315 VSS.n314 6.02403
R16959 VSS.n974 VSS.n973 6.02403
R16960 VSS.n982 VSS.n971 6.02403
R16961 VSS.n624 VSS.n622 6.02403
R16962 VSS.n631 VSS.n620 6.02403
R16963 VSS.n742 VSS.n741 6.02403
R16964 VSS.n748 VSS.n747 6.02403
R16965 VSS.n1799 VSS.n1732 5.89705
R16966 VSS.n1819 VSS.n1721 5.89705
R16967 VSS.n1635 VSS.n1568 5.89705
R16968 VSS.n1655 VSS.n1557 5.89705
R16969 VSS.n1307 VSS.n1306 5.89705
R16970 VSS.n1231 VSS.n1212 5.89705
R16971 VSS.n986 VSS.n968 5.89705
R16972 VSS.n635 VSS.n617 5.89705
R16973 VSS.n1764 VSS.n1763 5.64756
R16974 VSS.n1758 VSS.n1754 5.64756
R16975 VSS.n1927 VSS.n1924 5.64756
R16976 VSS.n1932 VSS.n1931 5.64756
R16977 VSS.n1595 VSS.n1592 5.64756
R16978 VSS.n1600 VSS.n1599 5.64756
R16979 VSS.n122 VSS.n121 5.64756
R16980 VSS.n130 VSS.n129 5.64756
R16981 VSS.n1437 VSS.n1436 5.64756
R16982 VSS.n1431 VSS.n1427 5.64756
R16983 VSS.n1407 VSS.n74 5.64756
R16984 VSS.n75 VSS.n72 5.64756
R16985 VSS.n1416 VSS.n69 5.64756
R16986 VSS.n1422 VSS.n1421 5.64756
R16987 VSS.n1386 VSS.n116 5.64756
R16988 VSS.n117 VSS.n114 5.64756
R16989 VSS.n1395 VSS.n111 5.64756
R16990 VSS.n1401 VSS.n1400 5.64756
R16991 VSS.n1078 VSS.n1074 5.64756
R16992 VSS.n1084 VSS.n1083 5.64756
R16993 VSS.n1176 VSS.n1172 5.64756
R16994 VSS.n1182 VSS.n1181 5.64756
R16995 VSS.n266 VSS.n265 5.64756
R16996 VSS.n274 VSS.n273 5.64756
R16997 VSS.n289 VSS.n288 5.64756
R16998 VSS.n283 VSS.n279 5.64756
R16999 VSS.n687 VSS.n686 5.64756
R17000 VSS.n695 VSS.n694 5.64756
R17001 VSS.n710 VSS.n709 5.64756
R17002 VSS.n704 VSS.n700 5.64756
R17003 VSS.n2015 VSS.n2014 5.61038
R17004 VSS.n1919 VSS.n1918 5.61038
R17005 VSS.n836 VSS.n818 5.39982
R17006 VSS.n405 VSS.n401 5.39151
R17007 VSS.n365 VSS.n350 5.39151
R17008 VSS.n785 VSS.n496 5.39151
R17009 VSS.n896 VSS.n441 5.39051
R17010 VSS.n911 VSS.n419 5.39051
R17011 VSS.n931 VSS.n386 5.39051
R17012 VSS.n946 VSS.n244 5.39051
R17013 VSS.n798 VSS.n788 5.39051
R17014 VSS.n575 VSS.n574 5.38802
R17015 VSS.n1846 VSS.n1843 5.3711
R17016 VSS.n1682 VSS.n1679 5.3711
R17017 VSS.n1087 VSS.n1067 5.28653
R17018 VSS.n1993 VSS.n1935 5.28613
R17019 VSS.n1382 VSS.n133 5.2751
R17020 VSS.n1441 VSS.n59 5.2751
R17021 VSS.n108 VSS.n43 5.2751
R17022 VSS.n349 VSS.n348 5.27461
R17023 VSS.n714 VSS.n495 5.27461
R17024 VSS.n1796 VSS.n1735 5.27109
R17025 VSS.n1804 VSS.n1733 5.27109
R17026 VSS.n1820 VSS.n1724 5.27109
R17027 VSS.n1825 VSS.n1722 5.27109
R17028 VSS.n1971 VSS.n1970 5.27109
R17029 VSS.n1955 VSS.n1954 5.27109
R17030 VSS.n1632 VSS.n1571 5.27109
R17031 VSS.n1640 VSS.n1569 5.27109
R17032 VSS.n1656 VSS.n1560 5.27109
R17033 VSS.n1661 VSS.n1558 5.27109
R17034 VSS.n326 VSS.n325 5.27109
R17035 VSS.n310 VSS.n309 5.27109
R17036 VSS.n981 VSS.n969 5.27109
R17037 VSS.n989 VSS.n967 5.27109
R17038 VSS.n630 VSS.n618 5.27109
R17039 VSS.n638 VSS.n616 5.27109
R17040 VSS.n737 VSS.n736 5.27109
R17041 VSS.n753 VSS.n752 5.27109
R17042 VSS.n316 VSS.n256 5.26828
R17043 VSS.n746 VSS.n490 5.26828
R17044 VSS.n1964 VSS.n1906 5.26828
R17045 VSS.n319 VSS.n256 5.26748
R17046 VSS.n743 VSS.n490 5.26748
R17047 VSS.n1961 VSS.n1906 5.26748
R17048 VSS.n894 VSS.n893 5.13412
R17049 VSS.n909 VSS.n422 5.13412
R17050 VSS.n922 VSS.n921 5.13412
R17051 VSS.n929 VSS.n928 5.13412
R17052 VSS.n944 VSS.n367 5.13412
R17053 VSS.n801 VSS.n480 5.13412
R17054 VSS.n543 VSS.n540 4.89462
R17055 VSS.n593 VSS.n592 4.83275
R17056 VSS.n1766 VSS.n1752 4.76425
R17057 VSS.n1934 VSS.n1933 4.76425
R17058 VSS.n1602 VSS.n1601 4.76425
R17059 VSS.n132 VSS.n131 4.76425
R17060 VSS.n1439 VSS.n1425 4.76425
R17061 VSS.n1408 VSS.n1405 4.76425
R17062 VSS.n1424 VSS.n67 4.76425
R17063 VSS.n1387 VSS.n1384 4.76425
R17064 VSS.n1403 VSS.n109 4.76425
R17065 VSS.n1086 VSS.n1072 4.76425
R17066 VSS.n1184 VSS.n1170 4.76425
R17067 VSS.n276 VSS.n275 4.76425
R17068 VSS.n291 VSS.n277 4.76425
R17069 VSS.n697 VSS.n696 4.76425
R17070 VSS.n712 VSS.n698 4.76425
R17071 VSS.n1224 VSS.n1218 4.68469
R17072 VSS.n168 VSS.n162 4.68392
R17073 VSS.n977 VSS.n976 4.68392
R17074 VSS.n626 VSS.n625 4.68392
R17075 VSS.n1415 VSS.n1414 4.6505
R17076 VSS.n1394 VSS.n1393 4.6505
R17077 VSS.n1533 VSS.n1531 4.51815
R17078 VSS.n1789 VSS.n1739 4.51815
R17079 VSS.n1797 VSS.n1737 4.51815
R17080 VSS.n1826 VSS.n1720 4.51815
R17081 VSS.n1836 VSS.n1718 4.51815
R17082 VSS.n1976 VSS.n1975 4.51815
R17083 VSS.n1949 VSS.n1948 4.51815
R17084 VSS.n1625 VSS.n1575 4.51815
R17085 VSS.n1633 VSS.n1573 4.51815
R17086 VSS.n1662 VSS.n1556 4.51815
R17087 VSS.n1672 VSS.n1554 4.51815
R17088 VSS.n1304 VSS.n160 4.51815
R17089 VSS.n1229 VSS.n1215 4.51815
R17090 VSS.n331 VSS.n330 4.51815
R17091 VSS.n305 VSS.n304 4.51815
R17092 VSS.n988 VSS.n965 4.51815
R17093 VSS.n996 VSS.n963 4.51815
R17094 VSS.n637 VSS.n614 4.51815
R17095 VSS.n645 VSS.n612 4.51815
R17096 VSS.n732 VSS.n731 4.51815
R17097 VSS.n758 VSS.n757 4.51815
R17098 VSS.n903 VSS.n441 4.51417
R17099 VSS.n432 VSS.n419 4.51417
R17100 VSS.n412 VSS.n401 4.51417
R17101 VSS.n938 VSS.n386 4.51417
R17102 VSS.n377 VSS.n244 4.51417
R17103 VSS.n350 VSS.n235 4.51417
R17104 VSS.n1010 VSS.n228 4.51417
R17105 VSS.n663 VSS.n504 4.51417
R17106 VSS.n766 VSS.n496 4.51417
R17107 VSS.n788 VSS.n478 4.51417
R17108 VSS.n2018 VSS.n1518 4.5005
R17109 VSS.n1531 VSS.n1530 4.5005
R17110 VSS.n1832 VSS.n1718 4.5005
R17111 VSS.n1719 VSS.n1712 4.5005
R17112 VSS.n1949 VSS.n1944 4.5005
R17113 VSS.n1952 VSS.n1545 4.5005
R17114 VSS.n1668 VSS.n1554 4.5005
R17115 VSS.n1555 VSS.n1548 4.5005
R17116 VSS.n1890 VSS.n1547 4.5005
R17117 VSS.n1893 VSS.n1547 4.5005
R17118 VSS.n1999 VSS.n1544 4.5005
R17119 VSS.n1913 VSS.n1544 4.5005
R17120 VSS.n1894 VSS.n1544 4.5005
R17121 VSS.n1999 VSS.n1998 4.5005
R17122 VSS.n1998 VSS.n1997 4.5005
R17123 VSS.n1893 VSS.n1892 4.5005
R17124 VSS.n1892 VSS.n1698 4.5005
R17125 VSS.n1868 VSS.n1711 4.5005
R17126 VSS.n1852 VSS.n1711 4.5005
R17127 VSS.n1864 VSS.n1711 4.5005
R17128 VSS.n1866 VSS.n1862 4.5005
R17129 VSS.n1542 VSS.n1516 4.5005
R17130 VSS.n1542 VSS.n1541 4.5005
R17131 VSS.n2008 VSS.n1542 4.5005
R17132 VSS.n2009 VSS.n1537 4.5005
R17133 VSS.n2009 VSS.n2008 4.5005
R17134 VSS.n1688 VSS.n1547 4.5005
R17135 VSS.n1457 VSS.n62 4.5005
R17136 VSS.n92 VSS.n79 4.5005
R17137 VSS.n1366 VSS.n1365 4.5005
R17138 VSS.n1105 VSS.n1104 4.5005
R17139 VSS.n1208 VSS.n1207 4.5005
R17140 VSS.n1254 VSS.n209 4.5005
R17141 VSS.n1247 VSS.n1043 4.5005
R17142 VSS.n1154 VSS.n1043 4.5005
R17143 VSS.n1154 VSS.n1041 4.5005
R17144 VSS.n1247 VSS.n1044 4.5005
R17145 VSS.n1154 VSS.n1044 4.5005
R17146 VSS.n1256 VSS.n1248 4.5005
R17147 VSS.n1253 VSS.n1248 4.5005
R17148 VSS.n1254 VSS.n1253 4.5005
R17149 VSS.n1151 VSS.n1126 4.5005
R17150 VSS.n1137 VSS.n1126 4.5005
R17151 VSS.n1152 VSS.n1151 4.5005
R17152 VSS.n1152 VSS.n1051 4.5005
R17153 VSS.n1129 VSS.n1048 4.5005
R17154 VSS.n1153 VSS.n1049 4.5005
R17155 VSS.n1145 VSS.n1049 4.5005
R17156 VSS.n1125 VSS.n1056 4.5005
R17157 VSS.n1060 VSS.n1056 4.5005
R17158 VSS.n1060 VSS.n1054 4.5005
R17159 VSS.n1125 VSS.n1057 4.5005
R17160 VSS.n1060 VSS.n1057 4.5005
R17161 VSS.n1109 VSS.n1057 4.5005
R17162 VSS.n1117 VSS.n1054 4.5005
R17163 VSS.n1125 VSS.n1054 4.5005
R17164 VSS.n1063 VSS.n1056 4.5005
R17165 VSS.n1124 VSS.n1059 4.5005
R17166 VSS.n1125 VSS.n1124 4.5005
R17167 VSS.n1153 VSS.n1048 4.5005
R17168 VSS.n1153 VSS.n1152 4.5005
R17169 VSS.n1151 VSS.n1048 4.5005
R17170 VSS.n1215 VSS.n1044 4.5005
R17171 VSS.n1238 VSS.n1041 4.5005
R17172 VSS.n1247 VSS.n1041 4.5005
R17173 VSS.n1213 VSS.n1043 4.5005
R17174 VSS.n1246 VSS.n1046 4.5005
R17175 VSS.n1247 VSS.n1246 4.5005
R17176 VSS.n566 VSS.n565 4.5005
R17177 VSS.n556 VSS.n555 4.5005
R17178 VSS.n546 VSS.n522 4.5005
R17179 VSS.n530 VSS.n527 4.5005
R17180 VSS.n548 VSS.n547 4.5005
R17181 VSS.n557 VSS.n518 4.5005
R17182 VSS.n559 VSS.n558 4.5005
R17183 VSS.n567 VSS.n514 4.5005
R17184 VSS.n569 VSS.n568 4.5005
R17185 VSS.n576 VSS.n575 4.5005
R17186 VSS.n572 VSS.n571 4.5005
R17187 VSS.n562 VSS.n516 4.5005
R17188 VSS.n552 VSS.n520 4.5005
R17189 VSS.n544 VSS.n543 4.5005
R17190 VSS.n537 VSS.n536 4.5005
R17191 VSS.n532 VSS.n531 4.5005
R17192 VSS.n868 VSS.n811 4.5005
R17193 VSS.n822 VSS.n811 4.5005
R17194 VSS.n866 VSS.n811 4.5005
R17195 VSS.n867 VSS.n814 4.5005
R17196 VSS.n804 VSS.n803 4.5005
R17197 VSS.n781 VSS.n780 4.5005
R17198 VSS.n782 VSS.n781 4.5005
R17199 VSS.n782 VSS.n479 4.5005
R17200 VSS.n782 VSS.n497 4.5005
R17201 VSS.n767 VSS.n479 4.5005
R17202 VSS.n774 VSS.n767 4.5005
R17203 VSS.n606 VSS.n605 4.5005
R17204 VSS.n607 VSS.n606 4.5005
R17205 VSS.n671 VSS.n502 4.5005
R17206 VSS.n1029 VSS.n217 4.5005
R17207 VSS.n957 VSS.n956 4.5005
R17208 VSS.n958 VSS.n957 4.5005
R17209 VSS.n953 VSS.n952 4.5005
R17210 VSS.n952 VSS.n234 4.5005
R17211 VSS.n955 VSS.n234 4.5005
R17212 VSS.n362 VSS.n234 4.5005
R17213 VSS.n955 VSS.n233 4.5005
R17214 VSS.n355 VSS.n233 4.5005
R17215 VSS.n943 VSS.n942 4.5005
R17216 VSS.n949 VSS.n242 4.5005
R17217 VSS.n925 VSS.n381 4.5005
R17218 VSS.n934 VSS.n381 4.5005
R17219 VSS.n941 VSS.n381 4.5005
R17220 VSS.n940 VSS.n383 4.5005
R17221 VSS.n956 VSS.n223 4.5005
R17222 VSS.n230 VSS.n223 4.5005
R17223 VSS.n1023 VSS.n223 4.5005
R17224 VSS.n1023 VSS.n1022 4.5005
R17225 VSS.n1027 VSS.n1024 4.5005
R17226 VSS.n1030 VSS.n1024 4.5005
R17227 VSS.n1030 VSS.n1029 4.5005
R17228 VSS.n1010 VSS.n224 4.5005
R17229 VSS.n1022 VSS.n1021 4.5005
R17230 VSS.n351 VSS.n235 4.5005
R17231 VSS.n942 VSS.n240 4.5005
R17232 VSS.n371 VSS.n240 4.5005
R17233 VSS.n950 VSS.n240 4.5005
R17234 VSS.n917 VSS.n916 4.5005
R17235 VSS.n917 VSS.n398 4.5005
R17236 VSS.n926 VSS.n925 4.5005
R17237 VSS.n908 VSS.n907 4.5005
R17238 VSS.n914 VSS.n417 4.5005
R17239 VSS.n916 VSS.n394 4.5005
R17240 VSS.n408 VSS.n394 4.5005
R17241 VSS.n924 VSS.n394 4.5005
R17242 VSS.n804 VSS.n474 4.5005
R17243 VSS.n795 VSS.n474 4.5005
R17244 VSS.n807 VSS.n474 4.5005
R17245 VSS.n806 VSS.n476 4.5005
R17246 VSS.n605 VSS.n500 4.5005
R17247 VSS.n654 VSS.n500 4.5005
R17248 VSS.n672 VSS.n500 4.5005
R17249 VSS.n768 VSS.n766 4.5005
R17250 VSS.n478 VSS.n477 4.5005
R17251 VSS.n807 VSS.n806 4.5005
R17252 VSS.n839 VSS.n817 4.5005
R17253 VSS.n866 VSS.n839 4.5005
R17254 VSS.n868 VSS.n867 4.5005
R17255 VSS.n890 VSS.n436 4.5005
R17256 VSS.n899 VSS.n436 4.5005
R17257 VSS.n906 VSS.n436 4.5005
R17258 VSS.n891 VSS.n890 4.5005
R17259 VSS.n905 VSS.n438 4.5005
R17260 VSS.n907 VSS.n415 4.5005
R17261 VSS.n426 VSS.n415 4.5005
R17262 VSS.n915 VSS.n415 4.5005
R17263 VSS.n904 VSS.n903 4.5005
R17264 VSS.n906 VSS.n905 4.5005
R17265 VSS.n432 VSS.n416 4.5005
R17266 VSS.n915 VSS.n914 4.5005
R17267 VSS.n924 VSS.n923 4.5005
R17268 VSS.n413 VSS.n412 4.5005
R17269 VSS.n939 VSS.n938 4.5005
R17270 VSS.n941 VSS.n940 4.5005
R17271 VSS.n377 VSS.n241 4.5005
R17272 VSS.n950 VSS.n949 4.5005
R17273 VSS.n953 VSS.n237 4.5005
R17274 VSS.n663 VSS.n501 4.5005
R17275 VSS.n672 VSS.n671 4.5005
R17276 VSS.n780 VSS.n764 4.5005
R17277 VSS.n867 VSS.n866 4.5005
R17278 VSS.n1290 VSS.n179 4.5005
R17279 VSS.n1291 VSS.n150 4.5005
R17280 VSS.n160 VSS.n150 4.5005
R17281 VSS.n1313 VSS.n150 4.5005
R17282 VSS.n1312 VSS.n153 4.5005
R17283 VSS.n1293 VSS.n1291 4.5005
R17284 VSS.n175 VSS.n151 4.5005
R17285 VSS.n1313 VSS.n151 4.5005
R17286 VSS.n1293 VSS.n1292 4.5005
R17287 VSS.n1313 VSS.n1312 4.5005
R17288 VSS.n1291 VSS.n151 4.5005
R17289 VSS.n88 VSS.n33 4.5005
R17290 VSS.n1500 VSS.n33 4.5005
R17291 VSS.n1500 VSS.n35 4.5005
R17292 VSS.n1500 VSS.n32 4.5005
R17293 VSS.n1500 VSS.n1499 4.5005
R17294 VSS.n1488 VSS.n1466 4.5005
R17295 VSS.n1489 VSS.n1488 4.5005
R17296 VSS.n1488 VSS.n1469 4.5005
R17297 VSS.n1490 VSS.n1469 4.5005
R17298 VSS.n1469 VSS.n1468 4.5005
R17299 VSS.n1489 VSS.n1471 4.5005
R17300 VSS.n1490 VSS.n1489 4.5005
R17301 VSS.n1490 VSS.n1466 4.5005
R17302 VSS.n1466 VSS.n1465 4.5005
R17303 VSS.n1491 VSS.n63 4.5005
R17304 VSS.n1491 VSS.n1490 4.5005
R17305 VSS.n1353 VSS.n1327 4.5005
R17306 VSS.n1358 VSS.n1327 4.5005
R17307 VSS.n1360 VSS.n1327 4.5005
R17308 VSS.n1333 VSS.n1327 4.5005
R17309 VSS.n1354 VSS.n1353 4.5005
R17310 VSS.n1359 VSS.n1358 4.5005
R17311 VSS.n1358 VSS.n145 4.5005
R17312 VSS.n1359 VSS.n1333 4.5005
R17313 VSS.n1333 VSS.n1332 4.5005
R17314 VSS.n1361 VSS.n1360 4.5005
R17315 VSS.n1360 VSS.n1359 4.5005
R17316 VSS.n37 VSS.n35 4.5005
R17317 VSS.n45 VSS.n35 4.5005
R17318 VSS.n1499 VSS.n37 4.5005
R17319 VSS.n1499 VSS.n1498 4.5005
R17320 VSS.n51 VSS.n32 4.5005
R17321 VSS.n37 VSS.n32 4.5005
R17322 VSS.n1288 VSS.n178 4.5005
R17323 VSS.n1290 VSS.n178 4.5005
R17324 VSS.n1289 VSS.n1288 4.5005
R17325 VSS.n1290 VSS.n1289 4.5005
R17326 VSS.n1871 VSS.n1869 4.28946
R17327 VSS.n1772 VSS.n1751 4.14168
R17328 VSS.n1772 VSS.n1749 4.14168
R17329 VSS.n1847 VSS.n1844 4.14168
R17330 VSS.n1988 VSS.n1936 4.14168
R17331 VSS.n1608 VSS.n1587 4.14168
R17332 VSS.n1608 VSS.n1585 4.14168
R17333 VSS.n1683 VSS.n1680 4.14168
R17334 VSS.n1379 VSS.n1378 4.14168
R17335 VSS.n1355 VSS.n1354 4.14168
R17336 VSS.n1330 VSS.n1329 4.14168
R17337 VSS.n1445 VSS.n1444 4.14168
R17338 VSS.n1462 VSS.n63 4.14168
R17339 VSS.n1475 VSS.n1474 4.14168
R17340 VSS.n105 VSS.n104 4.14168
R17341 VSS.n88 VSS.n87 4.14168
R17342 VSS.n47 VSS.n46 4.14168
R17343 VSS.n1292 VSS.n173 4.14168
R17344 VSS.n1309 VSS.n1308 4.14168
R17345 VSS.n1091 VSS.n1090 4.14168
R17346 VSS.n1122 VSS.n1059 4.14168
R17347 VSS.n1112 VSS.n1111 4.14168
R17348 VSS.n1145 VSS.n1144 4.14168
R17349 VSS.n1134 VSS.n1131 4.14168
R17350 VSS.n1190 VSS.n1169 4.14168
R17351 VSS.n1190 VSS.n1167 4.14168
R17352 VSS.n1244 VSS.n1046 4.14168
R17353 VSS.n1233 VSS.n1214 4.14168
R17354 VSS.n900 VSS.n899 4.14168
R17355 VSS.n429 VSS.n417 4.14168
R17356 VSS.n409 VSS.n408 4.14168
R17357 VSS.n935 VSS.n934 4.14168
R17358 VSS.n374 VSS.n242 4.14168
R17359 VSS.n345 VSS.n344 4.14168
R17360 VSS.n362 VSS.n361 4.14168
R17361 VSS.n1016 VSS.n227 4.14168
R17362 VSS.n1021 VSS.n227 4.14168
R17363 VSS.n666 VSS.n506 4.14168
R17364 VSS.n666 VSS.n502 4.14168
R17365 VSS.n718 VSS.n717 4.14168
R17366 VSS.n769 VSS.n497 4.14168
R17367 VSS.n795 VSS.n794 4.14168
R17368 VSS.n821 VSS.n817 4.14168
R17369 VSS.n552 VSS.n551 4.14168
R17370 VSS.n572 VSS.n513 4.14168
R17371 VSS.n1710 VSS.n1707 4.1033
R17372 VSS.n1881 VSS.n1699 4.10304
R17373 VSS.n1882 VSS.n1881 3.93684
R17374 VSS.n1879 VSS.n1707 3.93684
R17375 VSS.n2011 VSS.n1537 3.76521
R17376 VSS.n1782 VSS.n1743 3.76521
R17377 VSS.n1790 VSS.n1741 3.76521
R17378 VSS.n1838 VSS.n1837 3.76521
R17379 VSS.n1862 VSS.n1861 3.76521
R17380 VSS.n1981 VSS.n1980 3.76521
R17381 VSS.n1997 VSS.n1996 3.76521
R17382 VSS.n1618 VSS.n1579 3.76521
R17383 VSS.n1626 VSS.n1577 3.76521
R17384 VSS.n1674 VSS.n1673 3.76521
R17385 VSS.n1698 VSS.n1697 3.76521
R17386 VSS.n1362 VSS.n145 3.76521
R17387 VSS.n1465 VSS.n61 3.76521
R17388 VSS.n52 VSS.n45 3.76521
R17389 VSS.n175 VSS.n174 3.76521
R17390 VSS.n1118 VSS.n1063 3.76521
R17391 VSS.n1136 VSS.n1129 3.76521
R17392 VSS.n1239 VSS.n1213 3.76521
R17393 VSS.n336 VSS.n335 3.76521
R17394 VSS.n301 VSS.n259 3.76521
R17395 VSS.n247 VSS.n237 3.76521
R17396 VSS.n995 VSS.n961 3.76521
R17397 VSS.n1000 VSS.n958 3.76521
R17398 VSS.n644 VSS.n610 3.76521
R17399 VSS.n649 VSS.n607 3.76521
R17400 VSS.n727 VSS.n726 3.76521
R17401 VSS.n760 VSS.n493 3.76521
R17402 VSS.n764 VSS.n763 3.76521
R17403 VSS.n534 VSS.n528 3.49117
R17404 VSS.n1077 VSS.n1075 3.47842
R17405 VSS.n1175 VSS.n1173 3.47842
R17406 VSS.n1430 VSS.n1428 3.47756
R17407 VSS.n1929 VSS.n1928 3.47756
R17408 VSS.n1597 VSS.n1596 3.47756
R17409 VSS.n282 VSS.n280 3.47756
R17410 VSS.n703 VSS.n701 3.47756
R17411 VSS.n1757 VSS.n1755 3.47753
R17412 VSS.n127 VSS.n126 3.4767
R17413 VSS.n271 VSS.n270 3.4767
R17414 VSS.n692 VSS.n691 3.4767
R17415 VSS.n594 VSS.n577 3.41629
R17416 VSS.n22 VSS.n11 3.4105
R17417 VSS.n1502 VSS.n22 3.4105
R17418 VSS.n22 VSS.n12 3.4105
R17419 VSS.n22 VSS.n19 3.4105
R17420 VSS.n22 VSS.n13 3.4105
R17421 VSS.n22 VSS.n15 3.4105
R17422 VSS.n22 VSS.n17 3.4105
R17423 VSS.n22 VSS.n18 3.4105
R17424 VSS.n24 VSS.n11 3.4105
R17425 VSS.n1502 VSS.n24 3.4105
R17426 VSS.n24 VSS.n12 3.4105
R17427 VSS.n24 VSS.n19 3.4105
R17428 VSS.n24 VSS.n13 3.4105
R17429 VSS.n24 VSS.n15 3.4105
R17430 VSS.n24 VSS.n17 3.4105
R17431 VSS.n24 VSS.n18 3.4105
R17432 VSS.n842 VSS.n451 3.4105
R17433 VSS.n845 VSS.n842 3.4105
R17434 VSS.n842 VSS.n461 3.4105
R17435 VSS.n842 VSS.n458 3.4105
R17436 VSS.n842 VSS.n462 3.4105
R17437 VSS.n842 VSS.n457 3.4105
R17438 VSS.n842 VSS.n463 3.4105
R17439 VSS.n842 VSS.n456 3.4105
R17440 VSS.n842 VSS.n464 3.4105
R17441 VSS.n842 VSS.n455 3.4105
R17442 VSS.n842 VSS.n465 3.4105
R17443 VSS.n842 VSS.n466 3.4105
R17444 VSS.n843 VSS.n842 3.4105
R17445 VSS.n472 VSS.n461 3.4105
R17446 VSS.n472 VSS.n458 3.4105
R17447 VSS.n472 VSS.n462 3.4105
R17448 VSS.n472 VSS.n457 3.4105
R17449 VSS.n472 VSS.n463 3.4105
R17450 VSS.n472 VSS.n456 3.4105
R17451 VSS.n472 VSS.n464 3.4105
R17452 VSS.n472 VSS.n455 3.4105
R17453 VSS.n472 VSS.n465 3.4105
R17454 VSS.n472 VSS.n454 3.4105
R17455 VSS.n472 VSS.n466 3.4105
R17456 VSS.n886 VSS.n472 3.4105
R17457 VSS.n887 VSS.n459 3.4105
R17458 VSS.n459 VSS.n450 3.4105
R17459 VSS.n886 VSS.n450 3.4105
R17460 VSS.n466 VSS.n450 3.4105
R17461 VSS.n465 VSS.n450 3.4105
R17462 VSS.n455 VSS.n450 3.4105
R17463 VSS.n464 VSS.n450 3.4105
R17464 VSS.n456 VSS.n450 3.4105
R17465 VSS.n463 VSS.n450 3.4105
R17466 VSS.n457 VSS.n450 3.4105
R17467 VSS.n462 VSS.n450 3.4105
R17468 VSS.n458 VSS.n450 3.4105
R17469 VSS.n461 VSS.n450 3.4105
R17470 VSS.n845 VSS.n450 3.4105
R17471 VSS.n888 VSS.n450 3.4105
R17472 VSS.n453 VSS.n450 3.4105
R17473 VSS.n844 VSS.n843 3.4105
R17474 VSS.n844 VSS.n466 3.4105
R17475 VSS.n844 VSS.n454 3.4105
R17476 VSS.n844 VSS.n465 3.4105
R17477 VSS.n844 VSS.n455 3.4105
R17478 VSS.n844 VSS.n464 3.4105
R17479 VSS.n844 VSS.n456 3.4105
R17480 VSS.n844 VSS.n463 3.4105
R17481 VSS.n844 VSS.n457 3.4105
R17482 VSS.n844 VSS.n462 3.4105
R17483 VSS.n844 VSS.n458 3.4105
R17484 VSS.n844 VSS.n461 3.4105
R17485 VSS.n845 VSS.n844 3.4105
R17486 VSS.n844 VSS.n451 3.4105
R17487 VSS.n888 VSS.n887 3.4105
R17488 VSS.n887 VSS.n461 3.4105
R17489 VSS.n887 VSS.n458 3.4105
R17490 VSS.n887 VSS.n462 3.4105
R17491 VSS.n887 VSS.n457 3.4105
R17492 VSS.n887 VSS.n463 3.4105
R17493 VSS.n887 VSS.n456 3.4105
R17494 VSS.n887 VSS.n464 3.4105
R17495 VSS.n887 VSS.n455 3.4105
R17496 VSS.n887 VSS.n465 3.4105
R17497 VSS.n887 VSS.n454 3.4105
R17498 VSS.n887 VSS.n466 3.4105
R17499 VSS.n887 VSS.n453 3.4105
R17500 VSS.n845 VSS.n468 3.4105
R17501 VSS.n468 VSS.n461 3.4105
R17502 VSS.n468 VSS.n458 3.4105
R17503 VSS.n468 VSS.n462 3.4105
R17504 VSS.n468 VSS.n457 3.4105
R17505 VSS.n468 VSS.n463 3.4105
R17506 VSS.n468 VSS.n456 3.4105
R17507 VSS.n468 VSS.n464 3.4105
R17508 VSS.n468 VSS.n455 3.4105
R17509 VSS.n468 VSS.n465 3.4105
R17510 VSS.n468 VSS.n454 3.4105
R17511 VSS.n468 VSS.n466 3.4105
R17512 VSS.n886 VSS.n468 3.4105
R17513 VSS.n887 VSS.n886 3.4105
R17514 VSS.n1503 VSS.n15 3.4105
R17515 VSS.n21 VSS.n13 3.4105
R17516 VSS.n21 VSS.n15 3.4105
R17517 VSS.n21 VSS.n17 3.4105
R17518 VSS.n21 VSS.n14 3.4105
R17519 VSS.n21 VSS.n18 3.4105
R17520 VSS.n21 VSS.n19 3.4105
R17521 VSS.n21 VSS.n12 3.4105
R17522 VSS.n1502 VSS.n21 3.4105
R17523 VSS.n21 VSS.n11 3.4105
R17524 VSS.n1484 VSS.n26 3.4105
R17525 VSS.n1503 VSS.n17 3.4105
R17526 VSS.n1503 VSS.n14 3.4105
R17527 VSS.n1503 VSS.n18 3.4105
R17528 VSS.n26 VSS.n17 3.4105
R17529 VSS.n1315 VSS.n26 3.4105
R17530 VSS.n28 VSS.n26 3.4105
R17531 VSS.n1486 VSS.n26 3.4105
R17532 VSS.n26 VSS.n11 3.4105
R17533 VSS.n1502 VSS.n26 3.4105
R17534 VSS.n26 VSS.n12 3.4105
R17535 VSS.n26 VSS.n13 3.4105
R17536 VSS.n1503 VSS.n13 3.4105
R17537 VSS.n1503 VSS.n19 3.4105
R17538 VSS.n1503 VSS.n12 3.4105
R17539 VSS.n1503 VSS.n1502 3.4105
R17540 VSS.n1503 VSS.n11 3.4105
R17541 VSS.n30 VSS.n12 3.4105
R17542 VSS.n1502 VSS.n30 3.4105
R17543 VSS.n30 VSS.n11 3.4105
R17544 VSS.n1486 VSS.n30 3.4105
R17545 VSS.n1484 VSS.n30 3.4105
R17546 VSS.n30 VSS.n28 3.4105
R17547 VSS.n1315 VSS.n30 3.4105
R17548 VSS.n30 VSS.n17 3.4105
R17549 VSS.n30 VSS.n15 3.4105
R17550 VSS.n30 VSS.n13 3.4105
R17551 VSS.n26 VSS.n15 3.4105
R17552 VSS.n843 VSS.n468 3.4105
R17553 VSS.n843 VSS.n472 3.4105
R17554 VSS.n2042 VSS.n1513 3.4105
R17555 VSS.n1513 VSS.n9 3.4105
R17556 VSS.n1513 VSS.n1 3.4105
R17557 VSS.n1513 VSS.n8 3.4105
R17558 VSS.n1513 VSS.n2 3.4105
R17559 VSS.n1513 VSS.n7 3.4105
R17560 VSS.n1513 VSS.n3 3.4105
R17561 VSS.n1513 VSS.n6 3.4105
R17562 VSS.n2001 VSS.n1513 3.4105
R17563 VSS.n2001 VSS.n1508 3.4105
R17564 VSS.n1508 VSS.n4 3.4105
R17565 VSS.n1508 VSS.n6 3.4105
R17566 VSS.n1508 VSS.n3 3.4105
R17567 VSS.n1508 VSS.n7 3.4105
R17568 VSS.n1508 VSS.n2 3.4105
R17569 VSS.n1508 VSS.n8 3.4105
R17570 VSS.n1508 VSS.n1 3.4105
R17571 VSS.n1508 VSS.n9 3.4105
R17572 VSS.n1513 VSS.n10 3.4105
R17573 VSS.n1508 VSS.n10 3.4105
R17574 VSS.n2045 VSS.n1504 3.4105
R17575 VSS.n2042 VSS.n1504 3.4105
R17576 VSS.n1504 VSS.n9 3.4105
R17577 VSS.n1504 VSS.n1 3.4105
R17578 VSS.n1504 VSS.n8 3.4105
R17579 VSS.n1504 VSS.n2 3.4105
R17580 VSS.n1504 VSS.n7 3.4105
R17581 VSS.n1504 VSS.n3 3.4105
R17582 VSS.n1504 VSS.n6 3.4105
R17583 VSS.n1504 VSS.n5 3.4105
R17584 VSS.n2045 VSS.n1506 3.4105
R17585 VSS.n1506 VSS.n9 3.4105
R17586 VSS.n1506 VSS.n1 3.4105
R17587 VSS.n1506 VSS.n8 3.4105
R17588 VSS.n1506 VSS.n2 3.4105
R17589 VSS.n1506 VSS.n7 3.4105
R17590 VSS.n1506 VSS.n3 3.4105
R17591 VSS.n1506 VSS.n6 3.4105
R17592 VSS.n2046 VSS.n5 3.4105
R17593 VSS.n2046 VSS.n4 3.4105
R17594 VSS.n2046 VSS.n6 3.4105
R17595 VSS.n2046 VSS.n3 3.4105
R17596 VSS.n2046 VSS.n7 3.4105
R17597 VSS.n2046 VSS.n2 3.4105
R17598 VSS.n2046 VSS.n8 3.4105
R17599 VSS.n2046 VSS.n1 3.4105
R17600 VSS.n2046 VSS.n9 3.4105
R17601 VSS.n2046 VSS.n2045 3.4105
R17602 VSS.n1513 VSS.n1512 3.4105
R17603 VSS.n1506 VSS.n5 3.4105
R17604 VSS.n2045 VSS.n2044 3.4105
R17605 VSS.n2044 VSS.n9 3.4105
R17606 VSS.n2044 VSS.n1 3.4105
R17607 VSS.n2044 VSS.n8 3.4105
R17608 VSS.n2044 VSS.n2 3.4105
R17609 VSS.n2044 VSS.n7 3.4105
R17610 VSS.n2044 VSS.n3 3.4105
R17611 VSS.n2044 VSS.n6 3.4105
R17612 VSS.n2044 VSS.n5 3.4105
R17613 VSS.n1512 VSS.n1508 3.4105
R17614 VSS.n1541 VSS.n1536 3.38874
R17615 VSS.n1779 VSS.n1747 3.38874
R17616 VSS.n1779 VSS.n1745 3.38874
R17617 VSS.n1856 VSS.n1716 3.38874
R17618 VSS.n1856 VSS.n1852 3.38874
R17619 VSS.n1985 VSS.n1984 3.38874
R17620 VSS.n1913 VSS.n1901 3.38874
R17621 VSS.n1615 VSS.n1583 3.38874
R17622 VSS.n1615 VSS.n1581 3.38874
R17623 VSS.n1692 VSS.n1552 3.38874
R17624 VSS.n1692 VSS.n1688 3.38874
R17625 VSS.n1374 VSS.n1373 3.38874
R17626 VSS.n1370 VSS.n1369 3.38874
R17627 VSS.n1450 VSS.n1449 3.38874
R17628 VSS.n1454 VSS.n1453 3.38874
R17629 VSS.n100 VSS.n99 3.38874
R17630 VSS.n96 VSS.n95 3.38874
R17631 VSS.n1096 VSS.n1095 3.38874
R17632 VSS.n1100 VSS.n1099 3.38874
R17633 VSS.n1197 VSS.n1165 3.38874
R17634 VSS.n1197 VSS.n1163 3.38874
R17635 VSS.n1200 VSS.n1161 3.38874
R17636 VSS.n446 VSS.n438 3.38874
R17637 VSS.n426 VSS.n425 3.38874
R17638 VSS.n919 VSS.n398 3.38874
R17639 VSS.n391 VSS.n383 3.38874
R17640 VSS.n371 VSS.n370 3.38874
R17641 VSS.n340 VSS.n339 3.38874
R17642 VSS.n355 VSS.n354 3.38874
R17643 VSS.n1002 VSS.n959 3.38874
R17644 VSS.n1002 VSS.n230 3.38874
R17645 VSS.n655 VSS.n608 3.38874
R17646 VSS.n655 VSS.n654 3.38874
R17647 VSS.n723 VSS.n722 3.38874
R17648 VSS.n775 VSS.n774 3.38874
R17649 VSS.n482 VSS.n476 3.38874
R17650 VSS.n824 VSS.n822 3.38874
R17651 VSS.n562 VSS.n561 3.38874
R17652 VSS.n1261 VSS.n210 3.33963
R17653 VSS.n1252 VSS.n210 3.33963
R17654 VSS.n1252 VSS.n216 3.33963
R17655 VSS.n1257 VSS.n216 3.33963
R17656 VSS.n1035 VSS.n218 3.33963
R17657 VSS.n1031 VSS.n218 3.33963
R17658 VSS.n1031 VSS.n219 3.33963
R17659 VSS.n219 VSS.n198 3.33963
R17660 VSS.n1276 VSS.n181 3.33963
R17661 VSS.n1285 VSS.n181 3.33963
R17662 VSS.n1285 VSS.n1284 3.33963
R17663 VSS.n1284 VSS.n183 3.33963
R17664 VSS.n2013 VSS.t15 3.3065
R17665 VSS.n2013 VSS.t13 3.3065
R17666 VSS.n1994 VSS.t42 3.3065
R17667 VSS.n1994 VSS.t11 3.3065
R17668 VSS.n1363 VSS.t66 3.3065
R17669 VSS.n1363 VSS.t58 3.3065
R17670 VSS.t44 VSS.n1495 3.3065
R17671 VSS.n1495 VSS.t36 3.3065
R17672 VSS.n1496 VSS.t58 3.3065
R17673 VSS.n1496 VSS.t44 3.3065
R17674 VSS.n1119 VSS.t56 3.3065
R17675 VSS.n1119 VSS.t19 3.3065
R17676 VSS.n1139 VSS.t17 3.3065
R17677 VSS.n1139 VSS.t47 3.3065
R17678 VSS.n895 VSS.t28 3.3065
R17679 VSS.n895 VSS.t69 3.3065
R17680 VSS.n910 VSS.t23 3.3065
R17681 VSS.n910 VSS.t21 3.3065
R17682 VSS.n397 VSS.t5 3.3065
R17683 VSS.n397 VSS.t3 3.3065
R17684 VSS.n930 VSS.t70 3.3065
R17685 VSS.n930 VSS.t25 3.3065
R17686 VSS.n945 VSS.t26 3.3065
R17687 VSS.n945 VSS.t33 3.3065
R17688 VSS.t33 VSS.n366 3.3065
R17689 VSS.n366 VSS.t63 3.3065
R17690 VSS.n786 VSS.t54 3.3065
R17691 VSS.t51 VSS.n786 3.3065
R17692 VSS.n799 VSS.t51 3.3065
R17693 VSS.n799 VSS.t9 3.3065
R17694 VSS.n835 VSS.t67 3.3065
R17695 VSS.n835 VSS.t1 3.3065
R17696 VSS.n512 VSS.t7 3.3065
R17697 VSS.n512 VSS.t31 3.3065
R17698 VSS.n1365 VSS.n139 3.22952
R17699 VSS.n62 VSS.n56 3.22952
R17700 VSS.n79 VSS.n40 3.22952
R17701 VSS.n1105 VSS.n1065 3.22952
R17702 VSS.n1035 VSS.n217 3.03311
R17703 VSS.n1261 VSS.n209 3.03311
R17704 VSS.n1027 VSS.n198 3.03311
R17705 VSS.n1031 VSS.n1030 3.03311
R17706 VSS.n1257 VSS.n1256 3.03311
R17707 VSS.n1253 VSS.n1252 3.03311
R17708 VSS.n183 VSS.n178 3.03311
R17709 VSS.n1276 VSS.n179 3.03311
R17710 VSS.n1289 VSS.n1285 3.03311
R17711 VSS.n1871 VSS.n1870 3.02152
R17712 VSS.n1541 VSS.n1540 3.01226
R17713 VSS.n1775 VSS.n1747 3.01226
R17714 VSS.n1783 VSS.n1745 3.01226
R17715 VSS.n1860 VSS.n1716 3.01226
R17716 VSS.n1852 VSS.n1851 3.01226
R17717 VSS.n1986 VSS.n1985 3.01226
R17718 VSS.n1914 VSS.n1913 3.01226
R17719 VSS.n1611 VSS.n1583 3.01226
R17720 VSS.n1619 VSS.n1581 3.01226
R17721 VSS.n1696 VSS.n1552 3.01226
R17722 VSS.n1688 VSS.n1687 3.01226
R17723 VSS.n1375 VSS.n1374 3.01226
R17724 VSS.n1369 VSS.n1368 3.01226
R17725 VSS.n1365 VSS.n1364 3.01226
R17726 VSS.n1449 VSS.n1448 3.01226
R17727 VSS.n1455 VSS.n1454 3.01226
R17728 VSS.n1494 VSS.n62 3.01226
R17729 VSS.n101 VSS.n100 3.01226
R17730 VSS.n95 VSS.n94 3.01226
R17731 VSS.n79 VSS.n44 3.01226
R17732 VSS.n1095 VSS.n1094 3.01226
R17733 VSS.n1101 VSS.n1100 3.01226
R17734 VSS.n1107 VSS.n1105 3.01226
R17735 VSS.n1193 VSS.n1165 3.01226
R17736 VSS.n1201 VSS.n1163 3.01226
R17737 VSS.n1204 VSS.n1161 3.01226
R17738 VSS.n1210 VSS.n1208 3.01226
R17739 VSS.n444 VSS.n438 3.01226
R17740 VSS.n427 VSS.n426 3.01226
R17741 VSS.n403 VSS.n398 3.01226
R17742 VSS.n389 VSS.n383 3.01226
R17743 VSS.n372 VSS.n371 3.01226
R17744 VSS.n341 VSS.n340 3.01226
R17745 VSS.n356 VSS.n355 3.01226
R17746 VSS.n1006 VSS.n959 3.01226
R17747 VSS.n1014 VSS.n230 3.01226
R17748 VSS.n659 VSS.n608 3.01226
R17749 VSS.n654 VSS.n653 3.01226
R17750 VSS.n722 VSS.n721 3.01226
R17751 VSS.n774 VSS.n773 3.01226
R17752 VSS.n789 VSS.n476 3.01226
R17753 VSS.n832 VSS.n822 3.01226
R17754 VSS.n564 VSS.n562 3.01226
R17755 VSS.n1139 VSS.n1128 2.66358
R17756 VSS.n1538 VSS.n1537 2.63579
R17757 VSS.n1786 VSS.n1743 2.63579
R17758 VSS.n1786 VSS.n1741 2.63579
R17759 VSS.n1838 VSS.n1715 2.63579
R17760 VSS.n1862 VSS.n1715 2.63579
R17761 VSS.n1980 VSS.n1979 2.63579
R17762 VSS.n1997 VSS.n1897 2.63579
R17763 VSS.n1622 VSS.n1579 2.63579
R17764 VSS.n1622 VSS.n1577 2.63579
R17765 VSS.n1674 VSS.n1551 2.63579
R17766 VSS.n1698 VSS.n1551 2.63579
R17767 VSS.n1204 VSS.n1159 2.63579
R17768 VSS.n335 VSS.n334 2.63579
R17769 VSS.n249 VSS.n237 2.63579
R17770 VSS.n1000 VSS.n961 2.63579
R17771 VSS.n1007 VSS.n958 2.63579
R17772 VSS.n649 VSS.n610 2.63579
R17773 VSS.n660 VSS.n607 2.63579
R17774 VSS.n728 VSS.n727 2.63579
R17775 VSS.n778 VSS.n764 2.63579
R17776 VSS.n819 VSS.n814 2.63579
R17777 VSS.n536 VSS.n535 2.63579
R17778 VSS.n145 VSS.n143 2.529
R17779 VSS.n1465 VSS.n57 2.529
R17780 VSS.n45 VSS.n42 2.529
R17781 VSS.n1120 VSS.n1063 2.529
R17782 VSS.n1140 VSS.n1129 2.529
R17783 VSS.n301 VSS.n248 2.47658
R17784 VSS.n760 VSS.n483 2.47658
R17785 VSS.n1299 VSS.n1298 2.35698
R17786 VSS.n1256 VSS.n1255 2.2603
R17787 VSS.n1028 VSS.n1027 2.2603
R17788 VSS.n1769 VSS.n1751 2.25932
R17789 VSS.n1776 VSS.n1749 2.25932
R17790 VSS.n1844 VSS.n1842 2.25932
R17791 VSS.n1992 VSS.n1936 2.25932
R17792 VSS.n1605 VSS.n1587 2.25932
R17793 VSS.n1612 VSS.n1585 2.25932
R17794 VSS.n1680 VSS.n1678 2.25932
R17795 VSS.n1380 VSS.n1379 2.25932
R17796 VSS.n1329 VSS.n146 2.25932
R17797 VSS.n1444 VSS.n1443 2.25932
R17798 VSS.n1476 VSS.n1475 2.25932
R17799 VSS.n106 VSS.n105 2.25932
R17800 VSS.n50 VSS.n47 2.25932
R17801 VSS.n1310 VSS.n1309 2.25932
R17802 VSS.n1090 VSS.n1089 2.25932
R17803 VSS.n1116 VSS.n1111 2.25932
R17804 VSS.n1131 VSS.n1130 2.25932
R17805 VSS.n1187 VSS.n1169 2.25932
R17806 VSS.n1194 VSS.n1167 2.25932
R17807 VSS.n1237 VSS.n1214 2.25932
R17808 VSS.n899 VSS.n898 2.25932
R17809 VSS.n912 VSS.n417 2.25932
R17810 VSS.n408 VSS.n407 2.25932
R17811 VSS.n934 VSS.n933 2.25932
R17812 VSS.n947 VSS.n242 2.25932
R17813 VSS.n345 VSS.n261 2.25932
R17814 VSS.n364 VSS.n362 2.25932
R17815 VSS.n1016 VSS.n1015 2.25932
R17816 VSS.n1021 VSS.n1020 2.25932
R17817 VSS.n652 VSS.n506 2.25932
R17818 VSS.n669 VSS.n502 2.25932
R17819 VSS.n717 VSS.n716 2.25932
R17820 VSS.n784 VSS.n497 2.25932
R17821 VSS.n797 VSS.n795 2.25932
R17822 VSS.n837 VSS.n817 2.25932
R17823 VSS.n551 VSS.n521 2.25932
R17824 VSS.n553 VSS.n552 2.25932
R17825 VSS.n573 VSS.n572 2.25932
R17826 VSS.n829 VSS.n818 2.25051
R17827 VSS.n766 VSS.n498 2.25002
R17828 VSS.n359 VSS.n235 2.25002
R17829 VSS.n938 VSS.n388 2.25002
R17830 VSS.n412 VSS.n411 2.25002
R17831 VSS.n792 VSS.n478 2.25002
R17832 VSS.n903 VSS.n443 2.25002
R17833 VSS.n829 VSS.n813 2.24905
R17834 VSS.n1010 VSS.n231 2.24807
R17835 VSS.n377 VSS.n369 2.24807
R17836 VSS.n663 VSS.n508 2.24807
R17837 VSS.n432 VSS.n424 2.24807
R17838 VSS.n1854 VSS.n1712 2.2471
R17839 VSS.n1899 VSS.n1545 2.2471
R17840 VSS.n1690 VSS.n1548 2.2471
R17841 VSS.n1867 VSS.n1866 2.24691
R17842 VSS.n1150 VSS.n1049 2.24691
R17843 VSS.n1124 VSS.n1061 2.24691
R17844 VSS.n1246 VSS.n1155 2.24691
R17845 VSS.n767 VSS.n673 2.24691
R17846 VSS.n671 VSS.n503 2.24691
R17847 VSS.n951 VSS.n233 2.24691
R17848 VSS.n949 VSS.n243 2.24691
R17849 VSS.n940 VSS.n384 2.24691
R17850 VSS.n1022 VSS.n226 2.24691
R17851 VSS.n914 VSS.n418 2.24691
R17852 VSS.n923 VSS.n395 2.24691
R17853 VSS.n806 VSS.n805 2.24691
R17854 VSS.n839 VSS.n810 2.24691
R17855 VSS.n905 VSS.n439 2.24691
R17856 VSS.n1312 VSS.n154 2.24691
R17857 VSS.n1491 VSS.n1459 2.24691
R17858 VSS.n1866 VSS.n1865 2.24671
R17859 VSS.n1126 VSS.n1047 2.24671
R17860 VSS.n803 VSS.n473 2.24671
R17861 VSS.n606 VSS.n499 2.24671
R17862 VSS.n957 VSS.n222 2.24671
R17863 VSS.n943 VSS.n239 2.24671
R17864 VSS.n917 VSS.n393 2.24671
R17865 VSS.n926 VSS.n380 2.24671
R17866 VSS.n908 VSS.n414 2.24671
R17867 VSS.n891 VSS.n435 2.24671
R17868 VSS.n954 VSS.n953 2.24671
R17869 VSS.n780 VSS.n765 2.24671
R17870 VSS.n1293 VSS.n149 2.24671
R17871 VSS.n81 VSS.n33 2.24671
R17872 VSS.n1353 VSS.n1339 2.24671
R17873 VSS.n1149 VSS.n1127 2.24613
R17874 VSS.n1888 VSS.n1887 2.24394
R17875 VSS.n541 VSS.n521 2.24086
R17876 VSS.n1689 VSS.n1548 2.23886
R17877 VSS.n1853 VSS.n1712 2.23886
R17878 VSS.n1834 VSS.n1712 2.23886
R17879 VSS.n2018 VSS.n1523 2.23886
R17880 VSS.n2018 VSS.n1521 2.23886
R17881 VSS.n1946 VSS.n1545 2.23886
R17882 VSS.n1898 VSS.n1545 2.23886
R17883 VSS.n1670 VSS.n1548 2.23886
R17884 VSS.n771 VSS.n766 2.23886
R17885 VSS.n664 VSS.n663 2.23886
R17886 VSS.n358 VSS.n235 2.23886
R17887 VSS.n377 VSS.n376 2.23886
R17888 VSS.n938 VSS.n937 2.23886
R17889 VSS.n1012 VSS.n1010 2.23886
R17890 VSS.n432 VSS.n431 2.23886
R17891 VSS.n412 VSS.n402 2.23886
R17892 VSS.n791 VSS.n478 2.23886
R17893 VSS.n903 VSS.n902 2.23886
R17894 VSS.n1811 VSS.n1810 1.96602
R17895 VSS.n1817 VSS.n1725 1.96602
R17896 VSS.n1647 VSS.n1646 1.96602
R17897 VSS.n1653 VSS.n1561 1.96602
R17898 VSS.n165 VSS.n159 1.96602
R17899 VSS.n1221 VSS.n1216 1.96602
R17900 VSS.n979 VSS.n972 1.96602
R17901 VSS.n628 VSS.n621 1.96602
R17902 VSS.n829 VSS.n823 1.93808
R17903 VSS.n2018 VSS.n1520 1.93713
R17904 VSS.n1531 VSS.n1528 1.88285
R17905 VSS.n1793 VSS.n1739 1.88285
R17906 VSS.n1793 VSS.n1737 1.88285
R17907 VSS.n1830 VSS.n1720 1.88285
R17908 VSS.n1830 VSS.n1718 1.88285
R17909 VSS.n1975 VSS.n1974 1.88285
R17910 VSS.n1950 VSS.n1949 1.88285
R17911 VSS.n1629 VSS.n1575 1.88285
R17912 VSS.n1629 VSS.n1573 1.88285
R17913 VSS.n1666 VSS.n1556 1.88285
R17914 VSS.n1666 VSS.n1554 1.88285
R17915 VSS.n1356 VSS.n1355 1.88285
R17916 VSS.n1463 VSS.n1462 1.88285
R17917 VSS.n87 VSS.n84 1.88285
R17918 VSS.n1296 VSS.n173 1.88285
R17919 VSS.n1296 VSS.n176 1.88285
R17920 VSS.n1122 VSS.n1121 1.88285
R17921 VSS.n1144 VSS.n1141 1.88285
R17922 VSS.n1244 VSS.n1243 1.88285
R17923 VSS.n1243 VSS.n1157 1.88285
R17924 VSS.n330 VSS.n329 1.88285
R17925 VSS.n306 VSS.n305 1.88285
R17926 VSS.n992 VSS.n965 1.88285
R17927 VSS.n992 VSS.n963 1.88285
R17928 VSS.n641 VSS.n614 1.88285
R17929 VSS.n641 VSS.n612 1.88285
R17930 VSS.n733 VSS.n732 1.88285
R17931 VSS.n757 VSS.n756 1.88285
R17932 VSS.n536 VSS.n526 1.88285
R17933 VSS.n1332 VSS.n142 1.82308
R17934 VSS.n1468 VSS.n58 1.82308
R17935 VSS.n1498 VSS.n39 1.82308
R17936 VSS.n1109 VSS.n1064 1.82308
R17937 VSS.n1137 VSS.n1135 1.82308
R17938 VSS.n843 VSS.n452 1.71198
R17939 VSS.n1888 VSS.n1700 1.70717
R17940 VSS.n27 VSS.n14 1.70597
R17941 VSS.n845 VSS.n460 1.70597
R17942 VSS.n841 VSS.n454 1.70596
R17943 VSS.n25 VSS.n14 1.70596
R17944 VSS.n886 VSS.n469 1.70592
R17945 VSS.n1485 VSS.n16 1.70592
R17946 VSS.n471 VSS.n451 1.70592
R17947 VSS.n1485 VSS.n1483 1.70592
R17948 VSS.n2043 VSS.n2042 1.70591
R17949 VSS.n1510 VSS.n4 1.7059
R17950 VSS.n2042 VSS.n0 1.70578
R17951 VSS.n1507 VSS.n4 1.70577
R17952 VSS.n29 VSS.n19 1.70567
R17953 VSS.n2019 VSS.n2018 1.7055
R17954 VSS.n2002 VSS.n1543 1.7055
R17955 VSS.n2007 VSS.n2006 1.7055
R17956 VSS.n2021 VSS.n2020 1.7055
R17957 VSS.n2024 VSS.n2023 1.7055
R17958 VSS.n2027 VSS.n2026 1.7055
R17959 VSS.n2030 VSS.n2029 1.7055
R17960 VSS.n2035 VSS.n2034 1.7055
R17961 VSS.n2038 VSS.n2037 1.7055
R17962 VSS.n2040 VSS.n1514 1.7055
R17963 VSS.n1515 VSS.n1509 1.7055
R17964 VSS.n2033 VSS.n2032 1.7055
R17965 VSS.n2004 VSS.n2003 1.7055
R17966 VSS.n809 VSS.n467 1.7055
R17967 VSS.n449 VSS.n448 1.7055
R17968 VSS.n847 VSS.n846 1.7055
R17969 VSS.n850 VSS.n849 1.7055
R17970 VSS.n853 VSS.n852 1.7055
R17971 VSS.n858 VSS.n857 1.7055
R17972 VSS.n861 VSS.n860 1.7055
R17973 VSS.n864 VSS.n863 1.7055
R17974 VSS.n827 VSS.n815 1.7055
R17975 VSS.n871 VSS.n870 1.7055
R17976 VSS.n874 VSS.n873 1.7055
R17977 VSS.n877 VSS.n876 1.7055
R17978 VSS.n882 VSS.n881 1.7055
R17979 VSS.n884 VSS.n470 1.7055
R17980 VSS.n1349 VSS.n1348 1.7055
R17981 VSS.n1344 VSS.n1343 1.7055
R17982 VSS.n31 VSS.n20 1.7055
R17983 VSS.n34 VSS.n23 1.7055
R17984 VSS.n1481 VSS.n1480 1.7055
R17985 VSS.n1317 VSS.n1316 1.7055
R17986 VSS.n1320 VSS.n1319 1.7055
R17987 VSS.n1325 VSS.n1324 1.7055
R17988 VSS.n1336 VSS.n1334 1.7055
R17989 VSS.n808 VSS.n459 1.7055
R17990 VSS.n889 VSS.n888 1.7055
R17991 VSS.n845 VSS.n840 1.7055
R17992 VSS.n848 VSS.n461 1.7055
R17993 VSS.n851 VSS.n458 1.7055
R17994 VSS.n856 VSS.n462 1.7055
R17995 VSS.n859 VSS.n457 1.7055
R17996 VSS.n862 VSS.n463 1.7055
R17997 VSS.n869 VSS.n464 1.7055
R17998 VSS.n872 VSS.n455 1.7055
R17999 VSS.n875 VSS.n465 1.7055
R18000 VSS.n878 VSS.n454 1.7055
R18001 VSS.n883 VSS.n466 1.7055
R18002 VSS.n886 VSS.n885 1.7055
R18003 VSS.n1345 VSS.n19 1.7055
R18004 VSS.n1340 VSS.n12 1.7055
R18005 VSS.n1502 VSS.n1501 1.7055
R18006 VSS.n1479 VSS.n11 1.7055
R18007 VSS.n1487 VSS.n1486 1.7055
R18008 VSS.n1315 VSS.n1314 1.7055
R18009 VSS.n1318 VSS.n14 1.7055
R18010 VSS.n1323 VSS.n17 1.7055
R18011 VSS.n1350 VSS.n13 1.7055
R18012 VSS.n1326 VSS.n15 1.7055
R18013 VSS.n1863 VSS.n1505 1.7055
R18014 VSS.n2001 VSS.n2000 1.7055
R18015 VSS.n2005 VSS.n4 1.7055
R18016 VSS.n1522 VSS.n6 1.7055
R18017 VSS.n2022 VSS.n3 1.7055
R18018 VSS.n2025 VSS.n7 1.7055
R18019 VSS.n2031 VSS.n8 1.7055
R18020 VSS.n2036 VSS.n1 1.7055
R18021 VSS.n2039 VSS.n9 1.7055
R18022 VSS.n2042 VSS.n2041 1.7055
R18023 VSS.n1511 VSS.n1505 1.70511
R18024 VSS.n604 VSS.n576 1.6655
R18025 VSS.n528 VSS.n512 1.60574
R18026 VSS.n366 VSS.n256 1.60111
R18027 VSS.n786 VSS.n490 1.60111
R18028 VSS.n1994 VSS.n1906 1.60111
R18029 VSS.n594 VSS.n593 1.59802
R18030 VSS.n531 VSS.n529 1.5255
R18031 VSS.n1527 VSS.n1518 1.52198
R18032 VSS.n2018 VSS.n1519 1.51434
R18033 VSS.n1912 VSS.n1545 1.51434
R18034 VSS.n1679 VSS.n1548 1.51434
R18035 VSS.n1843 VSS.n1712 1.51289
R18036 VSS.n543 VSS.n542 1.50638
R18037 VSS.n1025 VSS.n217 1.50296
R18038 VSS.n1249 VSS.n209 1.50296
R18039 VSS.n1287 VSS.n179 1.50296
R18040 VSS.n516 VSS.n515 1.5005
R18041 VSS.n520 VSS.n519 1.5005
R18042 VSS.n545 VSS.n544 1.5005
R18043 VSS.n537 VSS.n523 1.5005
R18044 VSS.n1892 VSS.n1891 1.49719
R18045 VSS.n1998 VSS.n1895 1.49719
R18046 VSS.n1300 VSS.n152 1.49076
R18047 VSS.n1301 VSS.n1300 1.4899
R18048 VSS.n1467 VSS.n1461 1.4899
R18049 VSS.n1108 VSS.n1053 1.4899
R18050 VSS.n1226 VSS.n1040 1.4899
R18051 VSS.n2018 VSS.n2017 1.48477
R18052 VSS.n1916 VSS.n1545 1.48477
R18053 VSS.n1685 VSS.n1548 1.48477
R18054 VSS.n1849 VSS.n1712 1.48477
R18055 VSS.n1010 VSS.n1009 1.48392
R18056 VSS.n378 VSS.n377 1.48392
R18057 VSS.n938 VSS.n387 1.48392
R18058 VSS.n481 VSS.n478 1.48392
R18059 VSS.n663 VSS.n662 1.48392
R18060 VSS.n903 VSS.n442 1.48392
R18061 VSS.n433 VSS.n432 1.48392
R18062 VSS.n777 VSS.n766 1.48392
R18063 VSS.n352 VSS.n235 1.48392
R18064 VSS.n412 VSS.n399 1.48392
R18065 VSS.n1251 VSS.n1250 1.48264
R18066 VSS.n1026 VSS.n220 1.48264
R18067 VSS.n180 VSS.n177 1.48264
R18068 VSS.n1497 VSS.n1496 1.46886
R18069 VSS.n1119 VSS.n1110 1.46886
R18070 VSS.n1363 VSS.n144 1.46879
R18071 VSS.n1495 VSS.n60 1.46879
R18072 VSS.n1139 VSS.n1138 1.46878
R18073 VSS.n1281 VSS.n187 1.46668
R18074 VSS.n1259 VSS.n200 1.46668
R18075 VSS.n1266 VSS.n206 1.46668
R18076 VSS.n1033 VSS.n211 1.46668
R18077 VSS.n895 VSS.n894 1.41292
R18078 VSS.n910 VSS.n909 1.41292
R18079 VSS.n922 VSS.n397 1.41292
R18080 VSS.n930 VSS.n929 1.41292
R18081 VSS.n945 VSS.n944 1.41292
R18082 VSS.n799 VSS.n480 1.41292
R18083 VSS.n2009 VSS.n1524 1.35312
R18084 VSS.n829 VSS.n826 1.34465
R18085 VSS.n830 VSS.n829 1.34235
R18086 VSS.n880 VSS.n879 1.13717
R18087 VSS.n829 VSS.n828 1.13717
R18088 VSS.n855 VSS.n854 1.13717
R18089 VSS.n1347 VSS.n1346 1.13717
R18090 VSS.n1342 VSS.n1341 1.13717
R18091 VSS.n1482 VSS.n1478 1.13717
R18092 VSS.n83 VSS.n82 1.13717
R18093 VSS.n1338 VSS.n1337 1.13717
R18094 VSS.n1322 VSS.n1321 1.13717
R18095 VSS.n2018 VSS.n1517 1.13083
R18096 VSS.n1945 VSS.n1545 1.13027
R18097 VSS.n1669 VSS.n1548 1.13027
R18098 VSS.n1833 VSS.n1712 1.13002
R18099 VSS.n1800 VSS.n1735 1.12991
R18100 VSS.n1800 VSS.n1733 1.12991
R18101 VSS.n1821 VSS.n1820 1.12991
R18102 VSS.n1821 VSS.n1722 1.12991
R18103 VSS.n1970 VSS.n1969 1.12991
R18104 VSS.n1956 VSS.n1955 1.12991
R18105 VSS.n1636 VSS.n1571 1.12991
R18106 VSS.n1636 VSS.n1569 1.12991
R18107 VSS.n1657 VSS.n1656 1.12991
R18108 VSS.n1657 VSS.n1558 1.12991
R18109 VSS.n1308 VSS.n156 1.12991
R18110 VSS.n1233 VSS.n1232 1.12991
R18111 VSS.n325 VSS.n324 1.12991
R18112 VSS.n311 VSS.n310 1.12991
R18113 VSS.n985 VSS.n969 1.12991
R18114 VSS.n985 VSS.n967 1.12991
R18115 VSS.n634 VSS.n618 1.12991
R18116 VSS.n634 VSS.n616 1.12991
R18117 VSS.n738 VSS.n737 1.12991
R18118 VSS.n752 VSS.n751 1.12991
R18119 VSS.n540 VSS.n539 1.12991
R18120 VSS.n571 VSS.n510 1.1255
R18121 VSS.n1470 VSS.n1461 1.10942
R18122 VSS.n1149 VSS.n1050 1.10935
R18123 VSS.n1055 VSS.n1053 1.10935
R18124 VSS.n1042 VSS.n1040 1.10935
R18125 VSS.n1761 VSS.n1760 1.09595
R18126 VSS.n1925 VSS.n1921 1.09595
R18127 VSS.n1593 VSS.n1589 1.09595
R18128 VSS.n123 VSS.n119 1.09595
R18129 VSS.n1434 VSS.n1433 1.09595
R18130 VSS.n1411 VSS.n1410 1.09595
R18131 VSS.n1419 VSS.n1418 1.09595
R18132 VSS.n1390 VSS.n1389 1.09595
R18133 VSS.n1398 VSS.n1397 1.09595
R18134 VSS.n1081 VSS.n1080 1.09595
R18135 VSS.n1179 VSS.n1178 1.09595
R18136 VSS.n267 VSS.n263 1.09595
R18137 VSS.n286 VSS.n285 1.09595
R18138 VSS.n688 VSS.n684 1.09595
R18139 VSS.n707 VSS.n706 1.09595
R18140 VSS.n835 VSS.n834 1.0555
R18141 VSS.n1338 VSS.n1335 1.02924
R18142 VSS.n83 VSS.n38 1.02924
R18143 VSS.n1338 VSS.n147 1.02693
R18144 VSS.n83 VSS.n80 1.02693
R18145 VSS.n1149 VSS.n1148 0.903813
R18146 VSS.n1461 VSS.n1458 0.903813
R18147 VSS.n1300 VSS.n1299 0.903541
R18148 VSS.n1103 VSS.n1053 0.90354
R18149 VSS.n1206 VSS.n1040 0.90354
R18150 VSS.n1872 VSS.n1871 0.787987
R18151 VSS.n1763 VSS.n1762 0.753441
R18152 VSS.n1762 VSS.n1754 0.753441
R18153 VSS.n1924 VSS.n1922 0.753441
R18154 VSS.n1931 VSS.n1922 0.753441
R18155 VSS.n1592 VSS.n1590 0.753441
R18156 VSS.n1599 VSS.n1590 0.753441
R18157 VSS.n122 VSS.n120 0.753441
R18158 VSS.n129 VSS.n120 0.753441
R18159 VSS.n1436 VSS.n1435 0.753441
R18160 VSS.n1435 VSS.n1427 0.753441
R18161 VSS.n1412 VSS.n74 0.753441
R18162 VSS.n1412 VSS.n75 0.753441
R18163 VSS.n1420 VSS.n69 0.753441
R18164 VSS.n1421 VSS.n1420 0.753441
R18165 VSS.n1391 VSS.n116 0.753441
R18166 VSS.n1391 VSS.n117 0.753441
R18167 VSS.n1399 VSS.n111 0.753441
R18168 VSS.n1400 VSS.n1399 0.753441
R18169 VSS.n176 VSS.n175 0.753441
R18170 VSS.n160 VSS.n156 0.753441
R18171 VSS.n1082 VSS.n1074 0.753441
R18172 VSS.n1083 VSS.n1082 0.753441
R18173 VSS.n1208 VSS.n1159 0.753441
R18174 VSS.n1213 VSS.n1157 0.753441
R18175 VSS.n1232 VSS.n1215 0.753441
R18176 VSS.n1180 VSS.n1172 0.753441
R18177 VSS.n1181 VSS.n1180 0.753441
R18178 VSS.n266 VSS.n264 0.753441
R18179 VSS.n273 VSS.n264 0.753441
R18180 VSS.n288 VSS.n287 0.753441
R18181 VSS.n287 VSS.n279 0.753441
R18182 VSS.n687 VSS.n685 0.753441
R18183 VSS.n694 VSS.n685 0.753441
R18184 VSS.n709 VSS.n708 0.753441
R18185 VSS.n708 VSS.n700 0.753441
R18186 VSS.n539 VSS.n526 0.753441
R18187 VSS.n1026 VSS.n221 0.720975
R18188 VSS.n1250 VSS.n1039 0.720975
R18189 VSS.n1281 VSS.n185 0.720717
R18190 VSS.n91 VSS.n83 0.707257
R18191 VSS.n1338 VSS.n140 0.707257
R18192 VSS.n1894 VSS.n1893 0.682531
R18193 VSS.n1151 VSS.n1125 0.682531
R18194 VSS.n907 VSS.n906 0.682531
R18195 VSS.n916 VSS.n915 0.682531
R18196 VSS.n925 VSS.n924 0.682531
R18197 VSS.n942 VSS.n941 0.682531
R18198 VSS.n865 VSS.n456 0.6825
R18199 VSS.n834 VSS.n813 0.640088
R18200 VSS.n1286 VSS.n177 0.614024
R18201 VSS.n1148 VSS.n1128 0.594417
R18202 VSS.n1110 VSS.n1108 0.575661
R18203 VSS.n1467 VSS.n60 0.575335
R18204 VSS.n1335 VSS.n144 0.574421
R18205 VSS.n1497 VSS.n38 0.574409
R18206 VSS.n2028 VSS.n2 0.568833
R18207 VSS.n1138 VSS.n1127 0.561441
R18208 VSS.n2000 VSS.n1999 0.534875
R18209 VSS.n2047 VSS 0.524115
R18210 VSS.n601 VSS.n581 0.496624
R18211 VSS.n2015 VSS.n1526 0.461175
R18212 VSS.n1918 VSS.n1902 0.461175
R18213 VSS.n1378 VSS.n135 0.461175
R18214 VSS.n1445 VSS.n54 0.461175
R18215 VSS.n104 VSS.n53 0.461175
R18216 VSS.n1091 VSS.n1066 0.461175
R18217 VSS.n900 VSS.n445 0.461175
R18218 VSS.n429 VSS.n420 0.461175
R18219 VSS.n409 VSS.n404 0.461175
R18220 VSS.n935 VSS.n390 0.461175
R18221 VSS.n374 VSS.n245 0.461175
R18222 VSS.n344 VSS.n251 0.461175
R18223 VSS.n361 VSS.n260 0.461175
R18224 VSS.n718 VSS.n485 0.461175
R18225 VSS.n769 VSS.n494 0.461175
R18226 VSS.n794 VSS.n787 0.461175
R18227 VSS.n833 VSS.n821 0.461175
R18228 VSS.n563 VSS.n513 0.461175
R18229 VSS.n1988 VSS.n1911 0.460679
R18230 VSS.n602 VSS.n601 0.430441
R18231 VSS.n2012 VSS.n1536 0.430121
R18232 VSS.n1995 VSS.n1901 0.430121
R18233 VSS.n1373 VSS.n137 0.430121
R18234 VSS.n1450 VSS.n55 0.430121
R18235 VSS.n99 VSS.n41 0.430121
R18236 VSS.n1096 VSS.n1068 0.430121
R18237 VSS.n447 VSS.n446 0.430121
R18238 VSS.n425 VSS.n421 0.430121
R18239 VSS.n920 VSS.n919 0.430121
R18240 VSS.n392 VSS.n391 0.430121
R18241 VSS.n370 VSS.n246 0.430121
R18242 VSS.n339 VSS.n252 0.430121
R18243 VSS.n354 VSS.n250 0.430121
R18244 VSS.n723 VSS.n486 0.430121
R18245 VSS.n775 VSS.n484 0.430121
R18246 VSS.n800 VSS.n482 0.430121
R18247 VSS.n824 VSS.n820 0.430121
R18248 VSS.n561 VSS.n517 0.430121
R18249 VSS.n1984 VSS.n1910 0.429625
R18250 VSS.n1767 VSS.n1766 0.420318
R18251 VSS.n1603 VSS.n1602 0.420318
R18252 VSS.n1185 VSS.n1184 0.420318
R18253 VSS.n1538 VSS.n1534 0.398603
R18254 VSS.n1903 VSS.n1897 0.398603
R18255 VSS.n334 VSS.n253 0.398603
R18256 VSS.n728 VSS.n487 0.398603
R18257 VSS.n1979 VSS.n1909 0.398108
R18258 VSS.n1869 VSS.n1868 0.382531
R18259 VSS.n2013 VSS.n1527 0.378264
R18260 VSS.n1812 VSS.n1730 0.376971
R18261 VSS.n1812 VSS.n1731 0.376971
R18262 VSS.n1816 VSS.n1726 0.376971
R18263 VSS.n1816 VSS.n1728 0.376971
R18264 VSS.n1965 VSS.n1964 0.376971
R18265 VSS.n1961 VSS.n1960 0.376971
R18266 VSS.n1648 VSS.n1566 0.376971
R18267 VSS.n1648 VSS.n1567 0.376971
R18268 VSS.n1652 VSS.n1562 0.376971
R18269 VSS.n1652 VSS.n1564 0.376971
R18270 VSS.n1354 VSS.n141 0.376971
R18271 VSS.n1361 VSS.n146 0.376971
R18272 VSS.n1493 VSS.n63 0.376971
R18273 VSS.n1476 VSS.n1471 0.376971
R18274 VSS.n89 VSS.n88 0.376971
R18275 VSS.n51 VSS.n50 0.376971
R18276 VSS.n1292 VSS.n171 0.376971
R18277 VSS.n1310 VSS.n153 0.376971
R18278 VSS.n167 VSS.n161 0.376971
R18279 VSS.n167 VSS.n166 0.376971
R18280 VSS.n1106 VSS.n1059 0.376971
R18281 VSS.n1117 VSS.n1116 0.376971
R18282 VSS.n1146 VSS.n1145 0.376971
R18283 VSS.n1130 VSS.n1051 0.376971
R18284 VSS.n1209 VSS.n1046 0.376971
R18285 VSS.n1238 VSS.n1237 0.376971
R18286 VSS.n1223 VSS.n1217 0.376971
R18287 VSS.n1223 VSS.n1222 0.376971
R18288 VSS.n320 VSS.n319 0.376971
R18289 VSS.n316 VSS.n315 0.376971
R18290 VSS.n978 VSS.n973 0.376971
R18291 VSS.n978 VSS.n971 0.376971
R18292 VSS.n627 VSS.n622 0.376971
R18293 VSS.n627 VSS.n620 0.376971
R18294 VSS.n743 VSS.n742 0.376971
R18295 VSS.n747 VSS.n746 0.376971
R18296 VSS.n1950 VSS.n1904 0.366615
R18297 VSS.n329 VSS.n254 0.366615
R18298 VSS.n733 VSS.n488 0.366615
R18299 VSS.n1974 VSS.n1908 0.366119
R18300 VSS.n306 VSS.n258 0.366119
R18301 VSS.n756 VSS.n492 0.366119
R18302 VSS.n602 VSS.n578 0.35821
R18303 VSS.n1847 VSS.n1846 0.337513
R18304 VSS.n1683 VSS.n1682 0.337513
R18305 VSS.n1956 VSS.n1905 0.334147
R18306 VSS.n324 VSS.n255 0.334147
R18307 VSS.n738 VSS.n489 0.334147
R18308 VSS.n1969 VSS.n1907 0.333652
R18309 VSS.n311 VSS.n257 0.333652
R18310 VSS.n751 VSS.n491 0.333652
R18311 VSS.n1154 VSS.n1153 0.324719
R18312 VSS.n781 VSS.n672 0.324719
R18313 VSS.n804 VSS.n479 0.324719
R18314 VSS.n952 VSS.n950 0.324719
R18315 VSS.n956 VSS.n955 0.324719
R18316 VSS.n1935 VSS.n1934 0.316384
R18317 VSS.n1087 VSS.n1086 0.316384
R18318 VSS VSS.n1889 0.313
R18319 VSS.n605 VSS.n604 0.298156
R18320 VSS.n2014 VSS.n1519 0.297854
R18321 VSS.n1919 VSS.n1912 0.297854
R18322 VSS.n909 VSS.n908 0.251319
R18323 VSS.n944 VSS.n943 0.251319
R18324 VSS.n803 VSS.n480 0.251319
R18325 VSS.n923 VSS.n922 0.251319
R18326 VSS.n929 VSS.n926 0.251319
R18327 VSS.n894 VSS.n891 0.251319
R18328 VSS.n1488 VSS.n1487 0.234094
R18329 VSS.n529 VSS.n528 0.23152
R18330 VSS.n1383 VSS.n132 0.229427
R18331 VSS.n1384 VSS.n1383 0.229427
R18332 VSS.n1404 VSS.n1403 0.229427
R18333 VSS.n1405 VSS.n1404 0.229427
R18334 VSS.n1440 VSS.n1424 0.229427
R18335 VSS.n1440 VSS.n1439 0.229427
R18336 VSS.n292 VSS.n276 0.229427
R18337 VSS.n292 VSS.n291 0.229427
R18338 VSS.n713 VSS.n697 0.229427
R18339 VSS.n713 VSS.n712 0.229427
R18340 VSS.n1441 VSS.n1440 0.191391
R18341 VSS.n1404 VSS.n108 0.191391
R18342 VSS.n1383 VSS.n1382 0.191391
R18343 VSS.n348 VSS.n292 0.191391
R18344 VSS.n714 VSS.n713 0.191391
R18345 VSS.n1815 VSS.n1813 0.190717
R18346 VSS.n1963 VSS.n1962 0.190717
R18347 VSS.n1651 VSS.n1649 0.190717
R18348 VSS.n1393 VSS.n1392 0.190717
R18349 VSS.n1393 VSS.n112 0.190717
R18350 VSS.n1414 VSS.n1413 0.190717
R18351 VSS.n1414 VSS.n70 0.190717
R18352 VSS.n318 VSS.n317 0.190717
R18353 VSS.n745 VSS.n744 0.190717
R18354 VSS.n1768 VSS.n1767 0.164777
R18355 VSS.n1604 VSS.n1603 0.164777
R18356 VSS.n1442 VSS.n1441 0.164777
R18357 VSS.n108 VSS.n107 0.164777
R18358 VSS.n1382 VSS.n1381 0.164777
R18359 VSS.n1186 VSS.n1185 0.164777
R18360 VSS.n348 VSS.n347 0.164777
R18361 VSS.n715 VSS.n714 0.164777
R18362 VSS.n1766 VSS.n1765 0.15935
R18363 VSS.n1934 VSS.n1920 0.15935
R18364 VSS.n1602 VSS.n1588 0.15935
R18365 VSS.n132 VSS.n118 0.15935
R18366 VSS.n1385 VSS.n1384 0.15935
R18367 VSS.n1403 VSS.n1402 0.15935
R18368 VSS.n1406 VSS.n1405 0.15935
R18369 VSS.n1424 VSS.n1423 0.15935
R18370 VSS.n1439 VSS.n1438 0.15935
R18371 VSS.n1086 VSS.n1085 0.15935
R18372 VSS.n1184 VSS.n1183 0.15935
R18373 VSS.n276 VSS.n262 0.15935
R18374 VSS.n291 VSS.n290 0.15935
R18375 VSS.n697 VSS.n683 0.15935
R18376 VSS.n712 VSS.n711 0.15935
R18377 VSS.n808 VSS.n807 0.15675
R18378 VSS.n1504 VSS.n1503 0.149462
R18379 VSS.n195 VSS.n188 0.146748
R18380 VSS.n1774 VSS.n1773 0.144522
R18381 VSS.n1781 VSS.n1780 0.144522
R18382 VSS.n1788 VSS.n1787 0.144522
R18383 VSS.n1795 VSS.n1794 0.144522
R18384 VSS.n1802 VSS.n1801 0.144522
R18385 VSS.n1822 VSS.n1723 0.144522
R18386 VSS.n1989 VSS.n1987 0.144522
R18387 VSS.n1983 VSS.n1982 0.144522
R18388 VSS.n1978 VSS.n1977 0.144522
R18389 VSS.n1973 VSS.n1972 0.144522
R18390 VSS.n1968 VSS.n1967 0.144522
R18391 VSS.n1958 VSS.n1957 0.144522
R18392 VSS.n1610 VSS.n1609 0.144522
R18393 VSS.n1617 VSS.n1616 0.144522
R18394 VSS.n1624 VSS.n1623 0.144522
R18395 VSS.n1631 VSS.n1630 0.144522
R18396 VSS.n1638 VSS.n1637 0.144522
R18397 VSS.n1658 VSS.n1559 0.144522
R18398 VSS.n1447 VSS.n1446 0.144522
R18399 VSS.n1452 VSS.n1451 0.144522
R18400 VSS.n103 VSS.n102 0.144522
R18401 VSS.n98 VSS.n97 0.144522
R18402 VSS.n1377 VSS.n1376 0.144522
R18403 VSS.n1372 VSS.n1371 0.144522
R18404 VSS.n1093 VSS.n1092 0.144522
R18405 VSS.n1098 VSS.n1097 0.144522
R18406 VSS.n1192 VSS.n1191 0.144522
R18407 VSS.n1199 VSS.n1198 0.144522
R18408 VSS.n343 VSS.n342 0.144522
R18409 VSS.n338 VSS.n337 0.144522
R18410 VSS.n333 VSS.n332 0.144522
R18411 VSS.n328 VSS.n327 0.144522
R18412 VSS.n323 VSS.n322 0.144522
R18413 VSS.n313 VSS.n312 0.144522
R18414 VSS.n308 VSS.n307 0.144522
R18415 VSS.n984 VSS.n983 0.144522
R18416 VSS.n991 VSS.n990 0.144522
R18417 VSS.n633 VSS.n632 0.144522
R18418 VSS.n640 VSS.n639 0.144522
R18419 VSS.n720 VSS.n719 0.144522
R18420 VSS.n725 VSS.n724 0.144522
R18421 VSS.n730 VSS.n729 0.144522
R18422 VSS.n735 VSS.n734 0.144522
R18423 VSS.n740 VSS.n739 0.144522
R18424 VSS.n750 VSS.n749 0.144522
R18425 VSS.n755 VSS.n754 0.144522
R18426 VSS.n1991 VSS.n1935 0.141804
R18427 VSS.n1088 VSS.n1087 0.141804
R18428 VSS.n1368 VSS.n139 0.125448
R18429 VSS.n1455 VSS.n56 0.125448
R18430 VSS.n94 VSS.n40 0.125448
R18431 VSS.n1101 VSS.n1065 0.125448
R18432 VSS.n248 VSS.n247 0.125448
R18433 VSS.n763 VSS.n483 0.125448
R18434 VSS.n303 VSS.n302 0.122443
R18435 VSS.n998 VSS.n997 0.122443
R18436 VSS.n647 VSS.n646 0.122443
R18437 VSS.n761 VSS.n759 0.122443
R18438 VSS VSS.n2046 0.11659
R18439 VSS.n1248 VSS.n1247 0.113781
R18440 VSS.n1291 VSS.n1290 0.113781
R18441 VSS.n1824 VSS.n1719 0.106563
R18442 VSS.n1953 VSS.n1952 0.106563
R18443 VSS.n1660 VSS.n1555 0.106563
R18444 VSS.n1356 VSS.n143 0.0902327
R18445 VSS.n1463 VSS.n57 0.0902327
R18446 VSS.n84 VSS.n42 0.0902327
R18447 VSS.n1121 VSS.n1120 0.0902327
R18448 VSS.n1141 VSS.n1140 0.0902327
R18449 VSS.n1253 VSS.n1251 0.0861908
R18450 VSS.n1030 VSS.n220 0.0861908
R18451 VSS.n1289 VSS.n180 0.0861908
R18452 VSS.n1289 VSS.n1286 0.0777426
R18453 VSS.n831 VSS.n830 0.07529
R18454 VSS.n1027 VSS.n221 0.0740544
R18455 VSS.n1256 VSS.n1039 0.0740544
R18456 VSS.n1103 VSS.n1058 0.0699908
R18457 VSS.n1206 VSS.n1045 0.0699908
R18458 VSS.n1299 VSS.n170 0.0699908
R18459 VSS.n1492 VSS.n1458 0.0695895
R18460 VSS.n1148 VSS.n1147 0.0695894
R18461 VSS.n1253 VSS.n1039 0.0683603
R18462 VSS.n1030 VSS.n221 0.0683603
R18463 VSS.n1227 VSS.n1226 0.0679423
R18464 VSS.n1302 VSS.n1301 0.0676044
R18465 VSS.n1890 VSS 0.066125
R18466 VSS.n1024 VSS 0.066125
R18467 VSS.n91 VSS.n90 0.0638939
R18468 VSS.n1352 VSS.n140 0.0638939
R18469 VSS.n1286 VSS.n178 0.0636644
R18470 VSS.n2017 VSS.n1525 0.0618569
R18471 VSS.n1916 VSS.n1915 0.0618569
R18472 VSS.n1686 VSS.n1685 0.0618569
R18473 VSS.n1850 VSS.n1849 0.0615154
R18474 VSS.n433 VSS.n423 0.0611815
R18475 VSS.n378 VSS.n368 0.0611815
R18476 VSS.n1009 VSS.n232 0.0611815
R18477 VSS.n662 VSS.n509 0.0611815
R18478 VSS.n481 VSS.n475 0.0611815
R18479 VSS.n387 VSS.n382 0.0611815
R18480 VSS.n442 VSS.n437 0.0611815
R18481 VSS.n918 VSS.n399 0.0608398
R18482 VSS.n353 VSS.n352 0.0608398
R18483 VSS.n777 VSS.n776 0.0608398
R18484 VSS.n1312 VSS.n152 0.0604712
R18485 VSS.n902 VSS.n440 0.0584854
R18486 VSS.n431 VSS.n428 0.0584854
R18487 VSS.n402 VSS.n400 0.0584854
R18488 VSS.n937 VSS.n385 0.0584854
R18489 VSS.n376 VSS.n373 0.0584854
R18490 VSS.n358 VSS.n357 0.0584854
R18491 VSS.n1013 VSS.n1012 0.0584854
R18492 VSS.n664 VSS.n507 0.0584854
R18493 VSS.n772 VSS.n771 0.0584854
R18494 VSS.n791 VSS.n790 0.0584854
R18495 VSS.n1251 VSS.n209 0.0566413
R18496 VSS.n220 VSS.n217 0.0566413
R18497 VSS.n180 VSS.n179 0.0566413
R18498 VSS.n1535 VSS.n1523 0.0565323
R18499 VSS.n1855 VSS.n1853 0.0565323
R18500 VSS.n1900 VSS.n1898 0.0565323
R18501 VSS.n1691 VSS.n1689 0.0565323
R18502 VSS.n826 VSS.n825 0.0558464
R18503 VSS.n1330 VSS.n142 0.0547459
R18504 VSS.n1474 VSS.n58 0.0547459
R18505 VSS.n46 VSS.n39 0.0547459
R18506 VSS.n1112 VSS.n1064 0.0547459
R18507 VSS.n1135 VSS.n1134 0.0547459
R18508 VSS.n547 VSS.n519 0.053
R18509 VSS.n1532 VSS.n1521 0.0526261
R18510 VSS.n1539 VSS.n1521 0.0526261
R18511 VSS.n1835 VSS.n1834 0.0526261
R18512 VSS.n1834 VSS.n1713 0.0526261
R18513 VSS.n1947 VSS.n1946 0.0526261
R18514 VSS.n1946 VSS.n1546 0.0526261
R18515 VSS.n1671 VSS.n1670 0.0526261
R18516 VSS.n1670 VSS.n1549 0.0526261
R18517 VSS.n826 VSS.n812 0.0502162
R18518 VSS.n890 VSS.n889 0.0497188
R18519 VSS.n549 VSS.n548 0.0493281
R18520 VSS.n559 VSS.n518 0.0493281
R18521 VSS.n569 VSS.n514 0.0493281
R18522 VSS VSS.n1023 0.0489375
R18523 VSS.n2010 VSS.n1523 0.0487198
R18524 VSS.n1853 VSS.n1714 0.0487198
R18525 VSS.n1898 VSS.n1896 0.0487198
R18526 VSS.n1689 VSS.n1550 0.0487198
R18527 VSS.n1314 VSS.n1313 0.0481562
R18528 VSS.n902 VSS.n901 0.0467667
R18529 VSS.n431 VSS.n430 0.0467667
R18530 VSS.n410 VSS.n402 0.0467667
R18531 VSS.n937 VSS.n936 0.0467667
R18532 VSS.n376 VSS.n375 0.0467667
R18533 VSS.n360 VSS.n358 0.0467667
R18534 VSS.n1012 VSS.n1011 0.0467667
R18535 VSS.n665 VSS.n664 0.0467667
R18536 VSS.n771 VSS.n770 0.0467667
R18537 VSS.n793 VSS.n791 0.0467667
R18538 VSS.n1360 VSS.n147 0.0464244
R18539 VSS.n80 VSS.n32 0.0464244
R18540 VSS.n1152 VSS.n1050 0.0461141
R18541 VSS.n1055 VSS.n1054 0.0461141
R18542 VSS.n1042 VSS.n1041 0.0461141
R18543 VSS.n1489 VSS.n1470 0.045605
R18544 VSS.n1470 VSS.n1466 0.0454086
R18545 VSS.n399 VSS.n396 0.0449804
R18546 VSS.n352 VSS.n238 0.0449804
R18547 VSS.n779 VSS.n777 0.0449804
R18548 VSS.n1056 VSS.n1055 0.0448907
R18549 VSS.n1050 VSS.n1048 0.0448907
R18550 VSS.n1043 VSS.n1042 0.0448907
R18551 VSS.n892 VSS.n442 0.04464
R18552 VSS.n434 VSS.n433 0.04464
R18553 VSS.n927 VSS.n387 0.04464
R18554 VSS.n379 VSS.n378 0.04464
R18555 VSS.n1009 VSS.n1008 0.04464
R18556 VSS.n662 VSS.n661 0.04464
R18557 VSS.n802 VSS.n481 0.04464
R18558 VSS.n80 VSS.n35 0.0445792
R18559 VSS.n1358 VSS.n147 0.0445792
R18560 VSS.n1849 VSS.n1848 0.0443642
R18561 VSS.n2017 VSS.n2016 0.0440244
R18562 VSS.n1917 VSS.n1916 0.0440244
R18563 VSS.n1685 VSS.n1684 0.0440244
R18564 VSS.n1802 VSS.n1729 0.0439783
R18565 VSS.n1814 VSS.n1723 0.0439783
R18566 VSS.n1967 VSS.n1941 0.0439783
R18567 VSS.n1958 VSS.n1942 0.0439783
R18568 VSS.n1638 VSS.n1565 0.0439783
R18569 VSS.n1650 VSS.n1559 0.0439783
R18570 VSS.n1302 VSS.n169 0.0439783
R18571 VSS.n1227 VSS.n1225 0.0439783
R18572 VSS.n322 VSS.n297 0.0439783
R18573 VSS.n313 VSS.n298 0.0439783
R18574 VSS.n983 VSS.n970 0.0439783
R18575 VSS.n632 VSS.n619 0.0439783
R18576 VSS.n740 VSS.n677 0.0439783
R18577 VSS.n749 VSS.n676 0.0439783
R18578 VSS.n2041 VSS.n1515 0.0434688
R18579 VSS.n2041 VSS.n2040 0.0434688
R18580 VSS.n2040 VSS.n2039 0.0434688
R18581 VSS.n2039 VSS.n2038 0.0434688
R18582 VSS.n2038 VSS.n2036 0.0434688
R18583 VSS.n2036 VSS.n2035 0.0434688
R18584 VSS.n2031 VSS.n2030 0.0434688
R18585 VSS.n2030 VSS.n2028 0.0434688
R18586 VSS.n2028 VSS.n2027 0.0434688
R18587 VSS.n2027 VSS.n2025 0.0434688
R18588 VSS.n2025 VSS.n2024 0.0434688
R18589 VSS.n2024 VSS.n2022 0.0434688
R18590 VSS.n2022 VSS.n2021 0.0434688
R18591 VSS.n2007 VSS.n2005 0.0434688
R18592 VSS.n885 VSS.n809 0.0434688
R18593 VSS.n885 VSS.n884 0.0434688
R18594 VSS.n884 VSS.n883 0.0434688
R18595 VSS.n883 VSS.n882 0.0434688
R18596 VSS.n878 VSS.n877 0.0434688
R18597 VSS.n877 VSS.n875 0.0434688
R18598 VSS.n875 VSS.n874 0.0434688
R18599 VSS.n874 VSS.n872 0.0434688
R18600 VSS.n872 VSS.n871 0.0434688
R18601 VSS.n871 VSS.n869 0.0434688
R18602 VSS.n865 VSS.n864 0.0434688
R18603 VSS.n864 VSS.n862 0.0434688
R18604 VSS.n862 VSS.n861 0.0434688
R18605 VSS.n861 VSS.n859 0.0434688
R18606 VSS.n859 VSS.n858 0.0434688
R18607 VSS.n858 VSS.n856 0.0434688
R18608 VSS.n852 VSS.n851 0.0434688
R18609 VSS.n851 VSS.n850 0.0434688
R18610 VSS.n850 VSS.n848 0.0434688
R18611 VSS.n848 VSS.n847 0.0434688
R18612 VSS.n847 VSS.n840 0.0434688
R18613 VSS.n840 VSS.n448 0.0434688
R18614 VSS.n1318 VSS.n1317 0.0434688
R18615 VSS.n1319 VSS.n1318 0.0434688
R18616 VSS.n1325 VSS.n1323 0.0434688
R18617 VSS.n1326 VSS.n1325 0.0434688
R18618 VSS.n1350 VSS.n1349 0.0434688
R18619 VSS.n1345 VSS.n1344 0.0434688
R18620 VSS.n1340 VSS.n31 0.0434688
R18621 VSS.n1501 VSS.n31 0.0434688
R18622 VSS.n1480 VSS.n1479 0.0434688
R18623 VSS.n882 VSS.n879 0.0426875
R18624 VSS.n1127 VSS.n1126 0.0419945
R18625 VSS.n1501 VSS.n1500 0.0419063
R18626 VSS.n537 VSS.n527 0.0415156
R18627 VSS.n1765 VSS.n1753 0.0412609
R18628 VSS.n1930 VSS.n1920 0.0412609
R18629 VSS.n1598 VSS.n1588 0.0412609
R18630 VSS.n128 VSS.n118 0.0412609
R18631 VSS.n1385 VSS.n115 0.0412609
R18632 VSS.n1402 VSS.n110 0.0412609
R18633 VSS.n1406 VSS.n73 0.0412609
R18634 VSS.n1423 VSS.n68 0.0412609
R18635 VSS.n1438 VSS.n1426 0.0412609
R18636 VSS.n1085 VSS.n1073 0.0412609
R18637 VSS.n1183 VSS.n1171 0.0412609
R18638 VSS.n272 VSS.n262 0.0412609
R18639 VSS.n290 VSS.n278 0.0412609
R18640 VSS.n693 VSS.n683 0.0412609
R18641 VSS.n711 VSS.n699 0.0412609
R18642 VSS.n1346 VSS.n1345 0.041125
R18643 VSS.n1795 VSS.n1734 0.0385435
R18644 VSS.n1824 VSS.n1823 0.0385435
R18645 VSS.n1972 VSS.n1940 0.0385435
R18646 VSS.n1953 VSS.n1943 0.0385435
R18647 VSS.n1631 VSS.n1570 0.0385435
R18648 VSS.n1660 VSS.n1659 0.0385435
R18649 VSS.n327 VSS.n296 0.0385435
R18650 VSS.n308 VSS.n299 0.0385435
R18651 VSS.n990 VSS.n966 0.0385435
R18652 VSS.n639 VSS.n615 0.0385435
R18653 VSS.n735 VSS.n678 0.0385435
R18654 VSS.n754 VSS.n675 0.0385435
R18655 VSS.n809 VSS.n808 0.038
R18656 VSS.n889 VSS.n448 0.038
R18657 VSS.n2004 VSS.n1543 0.0372187
R18658 VSS.n866 VSS.n865 0.0372187
R18659 VSS.n533 VSS.n532 0.0356562
R18660 VSS.n565 VSS.n514 0.0356562
R18661 VSS.n1323 VSS.n1322 0.0356562
R18662 VSS.n1341 VSS.n1340 0.0356562
R18663 VSS.n1317 VSS.n1314 0.034875
R18664 VSS.n1487 VSS.n1478 0.034875
R18665 VSS.n856 VSS.n855 0.0340938
R18666 VSS.n1788 VSS.n1738 0.0331087
R18667 VSS.n1977 VSS.n1939 0.0331087
R18668 VSS.n1624 VSS.n1574 0.0331087
R18669 VSS.n332 VSS.n295 0.0331087
R18670 VSS.n303 VSS.n300 0.0331087
R18671 VSS.n997 VSS.n962 0.0331087
R18672 VSS.n646 VSS.n611 0.0331087
R18673 VSS.n730 VSS.n679 0.0331087
R18674 VSS.n759 VSS.n674 0.0331087
R18675 VSS.n2008 VSS.n2007 0.0325312
R18676 VSS.n575 VSS.n511 0.03175
R18677 VSS.n558 VSS.n557 0.03175
R18678 VSS.n568 VSS.n567 0.03175
R18679 VSS.n1864 VSS.n1863 0.0309688
R18680 VSS.n2035 VSS.n2032 0.0309688
R18681 VSS.n830 VSS.n816 0.0306452
R18682 VSS.n1335 VSS.n1333 0.0304205
R18683 VSS.n1499 VSS.n38 0.0304205
R18684 VSS.n1773 VSS.n1750 0.0303913
R18685 VSS.n1990 VSS.n1989 0.0303913
R18686 VSS.n1609 VSS.n1586 0.0303913
R18687 VSS.n1446 VSS.n66 0.0303913
R18688 VSS.n103 VSS.n76 0.0303913
R18689 VSS.n1377 VSS.n134 0.0303913
R18690 VSS.n1092 VSS.n1071 0.0303913
R18691 VSS.n1191 VSS.n1168 0.0303913
R18692 VSS.n346 VSS.n343 0.0303913
R18693 VSS.n719 VSS.n682 0.0303913
R18694 VSS.n1863 VSS.n1515 0.0301875
R18695 VSS.n2000 VSS.n1543 0.0301875
R18696 VSS.n152 VSS.n151 0.0301368
R18697 VSS.n897 VSS.n441 0.0297969
R18698 VSS.n913 VSS.n419 0.0297969
R18699 VSS.n406 VSS.n401 0.0297969
R18700 VSS.n932 VSS.n386 0.0297969
R18701 VSS.n948 VSS.n244 0.0297969
R18702 VSS.n363 VSS.n350 0.0297969
R18703 VSS.n228 VSS.n225 0.0297969
R18704 VSS.n670 VSS.n504 0.0297969
R18705 VSS.n783 VSS.n496 0.0297969
R18706 VSS.n796 VSS.n788 0.0297969
R18707 VSS.n545 VSS.n523 0.02925
R18708 VSS.n1301 VSS.n150 0.0288505
R18709 VSS.n1469 VSS.n1467 0.0288505
R18710 VSS.n1108 VSS.n1057 0.0285117
R18711 VSS.n1226 VSS.n1044 0.0285117
R18712 VSS.n576 VSS.n510 0.028
R18713 VSS.n555 VSS.n518 0.0278438
R18714 VSS.n1327 VSS.n1326 0.0278438
R18715 VSS.n1781 VSS.n1742 0.0276739
R18716 VSS.n1982 VSS.n1938 0.0276739
R18717 VSS.n1617 VSS.n1578 0.0276739
R18718 VSS.n337 VSS.n294 0.0276739
R18719 VSS.n725 VSS.n680 0.0276739
R18720 VSS.n530 VSS.n523 0.02675
R18721 VSS.n568 VSS.n510 0.02675
R18722 VSS.n544 VSS.n524 0.0258906
R18723 VSS.n1359 VSS.n1350 0.0255
R18724 VSS.n92 VSS.n91 0.0250149
R18725 VSS.n1366 VSS.n140 0.0250149
R18726 VSS.n1780 VSS.n1746 0.0249565
R18727 VSS.n1983 VSS.n1937 0.0249565
R18728 VSS.n1616 VSS.n1582 0.0249565
R18729 VSS.n1451 VSS.n65 0.0249565
R18730 VSS.n1452 VSS.n64 0.0249565
R18731 VSS.n98 VSS.n77 0.0249565
R18732 VSS.n97 VSS.n78 0.0249565
R18733 VSS.n1372 VSS.n136 0.0249565
R18734 VSS.n1371 VSS.n138 0.0249565
R18735 VSS.n1097 VSS.n1070 0.0249565
R18736 VSS.n1098 VSS.n1069 0.0249565
R18737 VSS.n1198 VSS.n1164 0.0249565
R18738 VSS.n1199 VSS.n1160 0.0249565
R18739 VSS.n338 VSS.n293 0.0249565
R18740 VSS.n724 VSS.n681 0.0249565
R18741 VSS.n1529 VSS.n1518 0.0239375
R18742 VSS.n1831 VSS.n1719 0.0239375
R18743 VSS.n1952 VSS.n1951 0.0239375
R18744 VSS.n1667 VSS.n1555 0.0239375
R18745 VSS.n525 VSS.n522 0.0239375
R18746 VSS.n603 VSS.n577 0.0232776
R18747 VSS.n567 VSS.n566 0.023
R18748 VSS.n838 VSS.n818 0.022459
R18749 VSS.n844 VSS.n21 0.0223109
R18750 VSS.n1774 VSS.n1746 0.0222391
R18751 VSS.n1987 VSS.n1937 0.0222391
R18752 VSS.n1610 VSS.n1582 0.0222391
R18753 VSS.n1447 VSS.n65 0.0222391
R18754 VSS.n1456 VSS.n64 0.0222391
R18755 VSS.n102 VSS.n77 0.0222391
R18756 VSS.n93 VSS.n78 0.0222391
R18757 VSS.n1376 VSS.n136 0.0222391
R18758 VSS.n1367 VSS.n138 0.0222391
R18759 VSS.n1093 VSS.n1070 0.0222391
R18760 VSS.n1102 VSS.n1069 0.0222391
R18761 VSS.n1192 VSS.n1164 0.0222391
R18762 VSS.n1205 VSS.n1160 0.0222391
R18763 VSS.n342 VSS.n293 0.0222391
R18764 VSS.n720 VSS.n681 0.0222391
R18765 VSS.n1491 VSS.n1460 0.0219844
R18766 VSS.n1473 VSS.n1472 0.0219844
R18767 VSS.n86 VSS.n33 0.0219844
R18768 VSS.n48 VSS.n36 0.0219844
R18769 VSS.n1353 VSS.n1351 0.0219844
R18770 VSS.n1331 VSS.n1328 0.0219844
R18771 VSS.n1294 VSS.n1293 0.0219844
R18772 VSS.n157 VSS.n155 0.0219844
R18773 VSS.n1124 VSS.n1123 0.0219844
R18774 VSS.n1114 VSS.n1113 0.0219844
R18775 VSS.n1143 VSS.n1049 0.0219844
R18776 VSS.n1133 VSS.n1132 0.0219844
R18777 VSS.n1246 VSS.n1245 0.0219844
R18778 VSS.n1235 VSS.n1234 0.0219844
R18779 VSS.n839 VSS.n816 0.0219844
R18780 VSS.n550 VSS.n520 0.0219844
R18781 VSS.n571 VSS.n570 0.0219844
R18782 VSS.n558 VSS.n515 0.02175
R18783 VSS.n2021 VSS.n1516 0.0208125
R18784 VSS.n901 VSS.n443 0.0205304
R18785 VSS.n411 VSS.n410 0.0205304
R18786 VSS.n936 VSS.n388 0.0205304
R18787 VSS.n360 VSS.n359 0.0205304
R18788 VSS.n770 VSS.n498 0.0205304
R18789 VSS.n793 VSS.n792 0.0205304
R18790 VSS.n546 VSS.n545 0.0205
R18791 VSS.n1835 VSS.n1833 0.0204768
R18792 VSS.n1947 VSS.n1945 0.0204759
R18793 VSS.n1671 VSS.n1669 0.0204759
R18794 VSS.n1532 VSS.n1517 0.020474
R18795 VSS.n2010 VSS.n2009 0.0200312
R18796 VSS.n1866 VSS.n1714 0.0200312
R18797 VSS.n1998 VSS.n1896 0.0200312
R18798 VSS.n1892 VSS.n1550 0.0200312
R18799 VSS.n953 VSS.n236 0.0200312
R18800 VSS.n999 VSS.n957 0.0200312
R18801 VSS.n648 VSS.n606 0.0200312
R18802 VSS.n780 VSS.n762 0.0200312
R18803 VSS.n548 VSS.n522 0.0200312
R18804 VSS.n570 VSS.n569 0.0200312
R18805 VSS.n1787 VSS.n1742 0.0195217
R18806 VSS.n1978 VSS.n1938 0.0195217
R18807 VSS.n1623 VSS.n1578 0.0195217
R18808 VSS.n333 VSS.n294 0.0195217
R18809 VSS.n729 VSS.n680 0.0195217
R18810 VSS.n1458 VSS.n1457 0.0188525
R18811 VSS.n1457 VSS.n1456 0.0188424
R18812 VSS.n93 VSS.n92 0.0188424
R18813 VSS.n1367 VSS.n1366 0.0188424
R18814 VSS.n1104 VSS.n1102 0.0188424
R18815 VSS.n1207 VSS.n1205 0.0188424
R18816 VSS.n1104 VSS.n1103 0.0184465
R18817 VSS.n1207 VSS.n1206 0.0184465
R18818 VSS.n905 VSS.n437 0.0180781
R18819 VSS.n423 VSS.n415 0.0180781
R18820 VSS.n430 VSS.n416 0.0180781
R18821 VSS.n918 VSS.n917 0.0180781
R18822 VSS.n940 VSS.n382 0.0180781
R18823 VSS.n368 VSS.n240 0.0180781
R18824 VSS.n375 VSS.n241 0.0180781
R18825 VSS.n353 VSS.n233 0.0180781
R18826 VSS.n232 VSS.n223 0.0180781
R18827 VSS.n1011 VSS.n224 0.0180781
R18828 VSS.n509 VSS.n500 0.0180781
R18829 VSS.n665 VSS.n501 0.0180781
R18830 VSS.n776 VSS.n767 0.0180781
R18831 VSS.n806 VSS.n475 0.0180781
R18832 VSS.n825 VSS.n811 0.0180781
R18833 VSS.n560 VSS.n516 0.0180781
R18834 VSS.n557 VSS.n556 0.018
R18835 VSS.n1125 VSS.n1053 0.0176875
R18836 VSS.n1247 VSS.n1040 0.0176875
R18837 VSS.n1290 VSS.n177 0.0176875
R18838 VSS.n1490 VSS.n1461 0.0176875
R18839 VSS.n1999 VSS.n1545 0.0169062
R18840 VSS.n1893 VSS.n1548 0.0169062
R18841 VSS.n1768 VSS.n1750 0.0168043
R18842 VSS.n1991 VSS.n1990 0.0168043
R18843 VSS.n1604 VSS.n1586 0.0168043
R18844 VSS.n1442 VSS.n66 0.0168043
R18845 VSS.n107 VSS.n76 0.0168043
R18846 VSS.n1381 VSS.n134 0.0168043
R18847 VSS.n1088 VSS.n1071 0.0168043
R18848 VSS.n1186 VSS.n1168 0.0168043
R18849 VSS.n347 VSS.n346 0.0168043
R18850 VSS.n715 VSS.n682 0.0168043
R18851 VSS.n1542 VSS.n1525 0.016125
R18852 VSS.n2016 VSS.n1519 0.016125
R18853 VSS.n1850 VSS.n1711 0.016125
R18854 VSS.n1848 VSS.n1843 0.016125
R18855 VSS.n1915 VSS.n1544 0.016125
R18856 VSS.n1917 VSS.n1912 0.016125
R18857 VSS.n1686 VSS.n1547 0.016125
R18858 VSS.n1684 VSS.n1679 0.016125
R18859 VSS.n560 VSS.n559 0.016125
R18860 VSS.n565 VSS.n516 0.016125
R18861 VSS.n869 VSS.n868 0.016125
R18862 VSS.n1334 VSS.n1327 0.016125
R18863 VSS.n556 VSS.n519 0.0155
R18864 VSS.n83 VSS.n34 0.0153437
R18865 VSS.n2042 VSS.n1509 0.0143978
R18866 VSS.n2042 VSS.n1514 0.0143978
R18867 VSS.n1514 VSS.n9 0.0143978
R18868 VSS.n2037 VSS.n9 0.0143978
R18869 VSS.n2037 VSS.n1 0.0143978
R18870 VSS.n2034 VSS.n1 0.0143978
R18871 VSS.n2029 VSS.n8 0.0143978
R18872 VSS.n2029 VSS.n2 0.0143978
R18873 VSS.n2026 VSS.n2 0.0143978
R18874 VSS.n2026 VSS.n7 0.0143978
R18875 VSS.n2023 VSS.n7 0.0143978
R18876 VSS.n2023 VSS.n3 0.0143978
R18877 VSS.n2020 VSS.n3 0.0143978
R18878 VSS.n2006 VSS.n6 0.0143978
R18879 VSS.n2006 VSS.n4 0.0143978
R18880 VSS.n886 VSS.n467 0.0143978
R18881 VSS.n886 VSS.n470 0.0143978
R18882 VSS.n470 VSS.n466 0.0143978
R18883 VSS.n881 VSS.n466 0.0143978
R18884 VSS.n876 VSS.n454 0.0143978
R18885 VSS.n876 VSS.n465 0.0143978
R18886 VSS.n873 VSS.n465 0.0143978
R18887 VSS.n873 VSS.n455 0.0143978
R18888 VSS.n870 VSS.n455 0.0143978
R18889 VSS.n870 VSS.n464 0.0143978
R18890 VSS.n827 VSS.n456 0.0143978
R18891 VSS.n863 VSS.n456 0.0143978
R18892 VSS.n863 VSS.n463 0.0143978
R18893 VSS.n860 VSS.n463 0.0143978
R18894 VSS.n860 VSS.n457 0.0143978
R18895 VSS.n857 VSS.n457 0.0143978
R18896 VSS.n857 VSS.n462 0.0143978
R18897 VSS.n853 VSS.n458 0.0143978
R18898 VSS.n849 VSS.n458 0.0143978
R18899 VSS.n849 VSS.n461 0.0143978
R18900 VSS.n846 VSS.n461 0.0143978
R18901 VSS.n846 VSS.n845 0.0143978
R18902 VSS.n845 VSS.n449 0.0143978
R18903 VSS.n1316 VSS.n14 0.0143978
R18904 VSS.n1320 VSS.n14 0.0143978
R18905 VSS.n1324 VSS.n17 0.0143978
R18906 VSS.n1324 VSS.n15 0.0143978
R18907 VSS.n1336 VSS.n15 0.0143978
R18908 VSS.n1348 VSS.n13 0.0143978
R18909 VSS.n1343 VSS.n19 0.0143978
R18910 VSS.n20 VSS.n12 0.0143978
R18911 VSS.n1502 VSS.n20 0.0143978
R18912 VSS.n1502 VSS.n23 0.0143978
R18913 VSS.n1481 VSS.n11 0.0143978
R18914 VSS.n2009 VSS.n1539 0.0141719
R18915 VSS.n1866 VSS.n1713 0.0141719
R18916 VSS.n1998 VSS.n1546 0.0141719
R18917 VSS.n1892 VSS.n1549 0.0141719
R18918 VSS.n1466 VSS.n1464 0.0141719
R18919 VSS.n85 VSS.n35 0.0141719
R18920 VSS.n1358 VSS.n1357 0.0141719
R18921 VSS.n1295 VSS.n151 0.0141719
R18922 VSS.n1062 VSS.n1056 0.0141719
R18923 VSS.n1142 VSS.n1048 0.0141719
R18924 VSS.n1156 VSS.n1043 0.0141719
R18925 VSS.n892 VSS.n891 0.0141719
R18926 VSS.n908 VSS.n434 0.0141719
R18927 VSS.n923 VSS.n396 0.0141719
R18928 VSS.n927 VSS.n926 0.0141719
R18929 VSS.n943 VSS.n379 0.0141719
R18930 VSS.n302 VSS.n236 0.0141719
R18931 VSS.n953 VSS.n238 0.0141719
R18932 VSS.n999 VSS.n998 0.0141719
R18933 VSS.n1008 VSS.n957 0.0141719
R18934 VSS.n648 VSS.n647 0.0141719
R18935 VSS.n661 VSS.n606 0.0141719
R18936 VSS.n762 VSS.n761 0.0141719
R18937 VSS.n780 VSS.n779 0.0141719
R18938 VSS.n803 VSS.n802 0.0141719
R18939 VSS.n867 VSS.n812 0.0141719
R18940 VSS.n538 VSS.n537 0.0141719
R18941 VSS.n881 VSS.n880 0.0141452
R18942 VSS.n1337 VSS.n13 0.0141452
R18943 VSS.n1794 VSS.n1738 0.014087
R18944 VSS.n1973 VSS.n1939 0.014087
R18945 VSS.n1630 VSS.n1574 0.014087
R18946 VSS.n328 VSS.n295 0.014087
R18947 VSS.n307 VSS.n300 0.014087
R18948 VSS.n991 VSS.n962 0.014087
R18949 VSS.n640 VSS.n611 0.014087
R18950 VSS.n734 VSS.n679 0.014087
R18951 VSS.n755 VSS.n674 0.014087
R18952 VSS.n1347 VSS.n19 0.0136398
R18953 VSS.n2032 VSS.n2031 0.013
R18954 VSS.n547 VSS.n546 0.013
R18955 VSS.n467 VSS.n459 0.012629
R18956 VSS.n888 VSS.n449 0.012629
R18957 VSS.n1524 VSS.n1516 0.012435
R18958 VSS.n1891 VSS.n1890 0.0124292
R18959 VSS.n1895 VSS.n1894 0.0124292
R18960 VSS.n2020 VSS.n2019 0.0123763
R18961 VSS.n2003 VSS.n2002 0.0123763
R18962 VSS.n1477 VSS.n1472 0.0122188
R18963 VSS.n49 VSS.n48 0.0122188
R18964 VSS.n1328 VSS.n148 0.0122188
R18965 VSS.n1311 VSS.n155 0.0122188
R18966 VSS.n1115 VSS.n1114 0.0122188
R18967 VSS.n1132 VSS.n1052 0.0122188
R18968 VSS.n1236 VSS.n1235 0.0122188
R18969 VSS.n905 VSS.n904 0.0122188
R18970 VSS.n897 VSS.n436 0.0122188
R18971 VSS.n914 VSS.n913 0.0122188
R18972 VSS.n917 VSS.n413 0.0122188
R18973 VSS.n406 VSS.n394 0.0122188
R18974 VSS.n940 VSS.n939 0.0122188
R18975 VSS.n932 VSS.n381 0.0122188
R18976 VSS.n949 VSS.n948 0.0122188
R18977 VSS.n351 VSS.n233 0.0122188
R18978 VSS.n363 VSS.n234 0.0122188
R18979 VSS.n1022 VSS.n225 0.0122188
R18980 VSS.n671 VSS.n670 0.0122188
R18981 VSS.n768 VSS.n767 0.0122188
R18982 VSS.n783 VSS.n782 0.0122188
R18983 VSS.n806 VSS.n477 0.0122188
R18984 VSS.n796 VSS.n474 0.0122188
R18985 VSS.n839 VSS.n838 0.0122188
R18986 VSS.n550 VSS.n549 0.0122188
R18987 VSS.n554 VSS.n520 0.0122188
R18988 VSS.n555 VSS.n554 0.0122188
R18989 VSS.n571 VSS.n511 0.0122188
R18990 VSS.n1249 VSS.n1248 0.0118907
R18991 VSS.n1025 VSS.n1024 0.0118907
R18992 VSS.n1288 VSS.n1287 0.0118907
R18993 VSS.n1321 VSS.n17 0.011871
R18994 VSS.n1342 VSS.n12 0.011871
R18995 VSS.n1316 VSS.n1315 0.0116183
R18996 VSS.n1486 VSS.n1482 0.0116183
R18997 VSS.n2008 VSS.n1522 0.0114375
R18998 VSS.n829 VSS.n815 0.0114375
R18999 VSS.n1479 VSS.n37 0.0114375
R19000 VSS.n854 VSS.n462 0.0113656
R19001 VSS.n828 VSS.n464 0.0108602
R19002 VSS.n428 VSS.n424 0.010758
R19003 VSS.n373 VSS.n369 0.010758
R19004 VSS.n1013 VSS.n231 0.010758
R19005 VSS.n508 VSS.n507 0.010758
R19006 VSS.n1855 VSS.n1854 0.0107521
R19007 VSS.n1900 VSS.n1899 0.0107521
R19008 VSS.n1691 VSS.n1690 0.0107521
R19009 VSS.n566 VSS.n515 0.0105
R19010 VSS.n581 VSS.n197 0.0104225
R19011 VSS.n2034 VSS.n2033 0.0103548
R19012 VSS.n1530 VSS.n1529 0.0102656
R19013 VSS.n1832 VSS.n1831 0.0102656
R19014 VSS.n1951 VSS.n1944 0.0102656
R19015 VSS.n1668 VSS.n1667 0.0102656
R19016 VSS.n1464 VSS.n1460 0.0102656
R19017 VSS.n1473 VSS.n1469 0.0102656
R19018 VSS.n86 VSS.n85 0.0102656
R19019 VSS.n1499 VSS.n36 0.0102656
R19020 VSS.n1357 VSS.n1351 0.0102656
R19021 VSS.n1333 VSS.n1331 0.0102656
R19022 VSS.n1295 VSS.n1294 0.0102656
R19023 VSS.n157 VSS.n150 0.0102656
R19024 VSS.n1123 VSS.n1062 0.0102656
R19025 VSS.n1113 VSS.n1057 0.0102656
R19026 VSS.n1143 VSS.n1142 0.0102656
R19027 VSS.n1133 VSS.n1126 0.0102656
R19028 VSS.n1245 VSS.n1156 0.0102656
R19029 VSS.n1234 VSS.n1044 0.0102656
R19030 VSS.n1509 VSS.n1505 0.0101021
R19031 VSS.n2002 VSS.n2001 0.0101021
R19032 VSS.n831 VSS.n823 0.00995073
R19033 VSS.n855 VSS.n852 0.009875
R19034 VSS.n1542 VSS.n1520 0.00987154
R19035 VSS.n1535 VSS.n1520 0.00967578
R19036 VSS.n1255 VSS.n1250 0.00962927
R19037 VSS.n1028 VSS.n1026 0.00962927
R19038 VSS.n82 VSS.n11 0.00959677
R19039 VSS.n1865 VSS.n1864 0.00957737
R19040 VSS.n1865 VSS.n1712 0.00957737
R19041 VSS.n1153 VSS.n1047 0.00957737
R19042 VSS.n1149 VSS.n1047 0.00957737
R19043 VSS.n672 VSS.n499 0.00957737
R19044 VSS.n766 VSS.n765 0.00957737
R19045 VSS.n807 VSS.n473 0.00957737
R19046 VSS.n903 VSS.n435 0.00957737
R19047 VSS.n915 VSS.n414 0.00957737
R19048 VSS.n924 VSS.n393 0.00957737
R19049 VSS.n938 VSS.n380 0.00957737
R19050 VSS.n950 VSS.n239 0.00957737
R19051 VSS.n954 VSS.n235 0.00957737
R19052 VSS.n1023 VSS.n222 0.00957737
R19053 VSS.n478 VSS.n473 0.00957737
R19054 VSS.n765 VSS.n479 0.00957737
R19055 VSS.n663 VSS.n499 0.00957737
R19056 VSS.n1010 VSS.n222 0.00957737
R19057 VSS.n955 VSS.n954 0.00957737
R19058 VSS.n377 VSS.n239 0.00957737
R19059 VSS.n412 VSS.n393 0.00957737
R19060 VSS.n941 VSS.n380 0.00957737
R19061 VSS.n432 VSS.n414 0.00957737
R19062 VSS.n906 VSS.n435 0.00957737
R19063 VSS.n1313 VSS.n149 0.00957737
R19064 VSS.n1339 VSS.n1338 0.00957737
R19065 VSS.n83 VSS.n81 0.00957737
R19066 VSS.n1300 VSS.n149 0.00957737
R19067 VSS.n81 VSS.n37 0.00957737
R19068 VSS.n1359 VSS.n1339 0.00957737
R19069 VSS.n1255 VSS.n1254 0.00952566
R19070 VSS.n1029 VSS.n1028 0.00952566
R19071 VSS.n1868 VSS.n1867 0.0091882
R19072 VSS.n1867 VSS.n1712 0.0091882
R19073 VSS.n1061 VSS.n1053 0.0091882
R19074 VSS.n1151 VSS.n1150 0.0091882
R19075 VSS.n1155 VSS.n1040 0.0091882
R19076 VSS.n1155 VSS.n1154 0.0091882
R19077 VSS.n1150 VSS.n1149 0.0091882
R19078 VSS.n1061 VSS.n1060 0.0091882
R19079 VSS.n663 VSS.n503 0.0091882
R19080 VSS.n766 VSS.n673 0.0091882
R19081 VSS.n805 VSS.n804 0.0091882
R19082 VSS.n829 VSS.n810 0.0091882
R19083 VSS.n903 VSS.n439 0.0091882
R19084 VSS.n432 VSS.n418 0.0091882
R19085 VSS.n916 VSS.n395 0.0091882
R19086 VSS.n938 VSS.n384 0.0091882
R19087 VSS.n377 VSS.n243 0.0091882
R19088 VSS.n951 VSS.n235 0.0091882
R19089 VSS.n956 VSS.n226 0.0091882
R19090 VSS.n781 VSS.n673 0.0091882
R19091 VSS.n605 VSS.n503 0.0091882
R19092 VSS.n952 VSS.n951 0.0091882
R19093 VSS.n942 VSS.n243 0.0091882
R19094 VSS.n925 VSS.n384 0.0091882
R19095 VSS.n1010 VSS.n226 0.0091882
R19096 VSS.n412 VSS.n395 0.0091882
R19097 VSS.n907 VSS.n418 0.0091882
R19098 VSS.n805 VSS.n478 0.0091882
R19099 VSS.n868 VSS.n810 0.0091882
R19100 VSS.n890 VSS.n439 0.0091882
R19101 VSS.n1300 VSS.n154 0.0091882
R19102 VSS.n1461 VSS.n1459 0.0091882
R19103 VSS.n1291 VSS.n154 0.0091882
R19104 VSS.n1488 VSS.n1459 0.0091882
R19105 VSS.n1854 VSS.n1711 0.00879896
R19106 VSS.n1899 VSS.n1544 0.00879896
R19107 VSS.n1690 VSS.n1547 0.00879896
R19108 VSS.n1801 VSS.n1734 0.00865217
R19109 VSS.n1823 VSS.n1822 0.00865217
R19110 VSS.n1968 VSS.n1940 0.00865217
R19111 VSS.n1957 VSS.n1943 0.00865217
R19112 VSS.n1637 VSS.n1570 0.00865217
R19113 VSS.n1659 VSS.n1658 0.00865217
R19114 VSS.n323 VSS.n296 0.00865217
R19115 VSS.n312 VSS.n299 0.00865217
R19116 VSS.n984 VSS.n966 0.00865217
R19117 VSS.n633 VSS.n615 0.00865217
R19118 VSS.n739 VSS.n678 0.00865217
R19119 VSS.n750 VSS.n675 0.00865217
R19120 VSS.n532 VSS.n527 0.0083125
R19121 VSS.n544 VSS.n525 0.0083125
R19122 VSS.n1322 VSS.n1319 0.0083125
R19123 VSS.n1344 VSS.n1341 0.0083125
R19124 VSS.n823 VSS.n811 0.00765694
R19125 VSS.n231 VSS.n223 0.00685176
R19126 VSS.n369 VSS.n240 0.00685176
R19127 VSS.n508 VSS.n500 0.00685176
R19128 VSS.n424 VSS.n415 0.00685176
R19129 VSS.n453 VSS.n451 0.0068172
R19130 VSS.n2018 VSS.n1522 0.00675
R19131 VSS.n2005 VSS.n2004 0.00675
R19132 VSS.n866 VSS.n815 0.00675
R19133 VSS.n1895 VSS.n1545 0.00671462
R19134 VSS.n1891 VSS.n1548 0.00671462
R19135 VSS.n1485 VSS.n1484 0.00656452
R19136 VSS.n1250 VSS.n1249 0.00647588
R19137 VSS.n1026 VSS.n1025 0.00647588
R19138 VSS.n1287 VSS.n177 0.00647588
R19139 VSS.n538 VSS.n524 0.00635938
R19140 VSS.n2047 VSS 0.00595359
R19141 VSS.n1755 VSS.n1753 0.00593478
R19142 VSS.n1930 VSS.n1929 0.00593478
R19143 VSS.n1598 VSS.n1597 0.00593478
R19144 VSS.n128 VSS.n127 0.00593478
R19145 VSS.n1392 VSS.n115 0.00593478
R19146 VSS.n112 VSS.n110 0.00593478
R19147 VSS.n1413 VSS.n73 0.00593478
R19148 VSS.n70 VSS.n68 0.00593478
R19149 VSS.n1428 VSS.n1426 0.00593478
R19150 VSS.n1075 VSS.n1073 0.00593478
R19151 VSS.n1173 VSS.n1171 0.00593478
R19152 VSS.n272 VSS.n271 0.00593478
R19153 VSS.n280 VSS.n278 0.00593478
R19154 VSS.n693 VSS.n692 0.00593478
R19155 VSS.n701 VSS.n699 0.00593478
R19156 VSS.n2018 VSS.n1524 0.00592961
R19157 VSS.n28 VSS.n18 0.00580645
R19158 VSS.n531 VSS.n530 0.0055
R19159 VSS.n82 VSS.n23 0.00530108
R19160 VSS.n219 VSS.n205 0.00507113
R19161 VSS.n1266 VSS.n205 0.00507113
R19162 VSS.n218 VSS.n207 0.00507113
R19163 VSS.n1266 VSS.n207 0.00507113
R19164 VSS.n216 VSS.n215 0.00507113
R19165 VSS.n213 VSS.n210 0.00507113
R19166 VSS.n189 VSS.n181 0.00507113
R19167 VSS.n1281 VSS.n189 0.00507113
R19168 VSS.n1284 VSS.n1283 0.00507113
R19169 VSS.n1530 VSS.n1517 0.00492302
R19170 VSS.n1945 VSS.n1944 0.00492108
R19171 VSS.n1669 VSS.n1668 0.00492108
R19172 VSS.n1833 VSS.n1832 0.00492021
R19173 VSS.n867 VSS.n813 0.00490286
R19174 VSS.n2045 VSS.n1505 0.0047957
R19175 VSS.n2001 VSS.n5 0.0047957
R19176 VSS.n215 VSS.n202 0.00478282
R19177 VSS.n213 VSS.n201 0.00478282
R19178 VSS.n1283 VSS.n1282 0.00478282
R19179 VSS.n2033 VSS.n8 0.00454301
R19180 VSS.n904 VSS.n440 0.00440625
R19181 VSS.n914 VSS.n416 0.00440625
R19182 VSS.n413 VSS.n400 0.00440625
R19183 VSS.n939 VSS.n385 0.00440625
R19184 VSS.n949 VSS.n241 0.00440625
R19185 VSS.n357 VSS.n351 0.00440625
R19186 VSS.n1022 VSS.n224 0.00440625
R19187 VSS.n671 VSS.n501 0.00440625
R19188 VSS.n772 VSS.n768 0.00440625
R19189 VSS.n790 VSS.n477 0.00440625
R19190 VSS.n533 VSS.n529 0.00440625
R19191 VSS.n2045 VSS.n10 0.00429032
R19192 VSS.n1512 VSS.n5 0.00429032
R19193 VSS.n828 VSS.n827 0.00403763
R19194 VSS VSS.n2047 0.00379439
R19195 VSS.n854 VSS.n853 0.00353226
R19196 VSS.n1315 VSS.n18 0.00327957
R19197 VSS.n1813 VSS.n1729 0.00321739
R19198 VSS.n1815 VSS.n1814 0.00321739
R19199 VSS.n1963 VSS.n1941 0.00321739
R19200 VSS.n1962 VSS.n1942 0.00321739
R19201 VSS.n1649 VSS.n1565 0.00321739
R19202 VSS.n1651 VSS.n1650 0.00321739
R19203 VSS.n169 VSS.n168 0.00321739
R19204 VSS.n1225 VSS.n1224 0.00321739
R19205 VSS.n318 VSS.n297 0.00321739
R19206 VSS.n317 VSS.n298 0.00321739
R19207 VSS.n977 VSS.n970 0.00321739
R19208 VSS.n626 VSS.n619 0.00321739
R19209 VSS.n744 VSS.n677 0.00321739
R19210 VSS.n745 VSS.n676 0.00321739
R19211 VSS.n1321 VSS.n1320 0.00302688
R19212 VSS.n1343 VSS.n1342 0.00302688
R19213 VSS.n443 VSS.n436 0.00295228
R19214 VSS.n411 VSS.n394 0.00295228
R19215 VSS.n388 VSS.n381 0.00295228
R19216 VSS.n359 VSS.n234 0.00295228
R19217 VSS.n782 VSS.n498 0.00295228
R19218 VSS.n792 VSS.n474 0.00295228
R19219 VSS.n1349 VSS.n1346 0.00284375
R19220 VSS.n1480 VSS.n1478 0.00284375
R19221 VSS.n1511 VSS.n1508 0.00278115
R19222 VSS.n1513 VSS.n1511 0.00278115
R19223 VSS.n1889 VSS.n1699 0.00269167
R19224 VSS.n2019 VSS.n6 0.00252151
R19225 VSS.n2003 VSS.n4 0.00252151
R19226 VSS.n1486 VSS.n1485 0.00252151
R19227 VSS.n1492 VSS.n1491 0.00245312
R19228 VSS.n1489 VSS.n1477 0.00245312
R19229 VSS.n90 VSS.n33 0.00245312
R19230 VSS.n49 VSS.n32 0.00245312
R19231 VSS.n1353 VSS.n1352 0.00245312
R19232 VSS.n1360 VSS.n148 0.00245312
R19233 VSS.n1293 VSS.n170 0.00245312
R19234 VSS.n1312 VSS.n1311 0.00245312
R19235 VSS.n1124 VSS.n1058 0.00245312
R19236 VSS.n1115 VSS.n1054 0.00245312
R19237 VSS.n1147 VSS.n1049 0.00245312
R19238 VSS.n1152 VSS.n1052 0.00245312
R19239 VSS.n1246 VSS.n1045 0.00245312
R19240 VSS.n1236 VSS.n1041 0.00245312
R19241 VSS.n843 VSS.n459 0.00226882
R19242 VSS.n888 VSS.n451 0.00226882
R19243 VSS.n1500 VSS.n34 0.0020625
R19244 VSS.n1266 VSS.n202 0.00178792
R19245 VSS.n1266 VSS.n201 0.00178792
R19246 VSS.n1282 VSS.n1281 0.00178792
R19247 VSS.n29 VSS.n26 0.00166815
R19248 VSS.n887 VSS.n452 0.00166815
R19249 VSS.n452 VSS.n450 0.00166815
R19250 VSS.n30 VSS.n29 0.00166815
R19251 VSS.n1704 VSS.n1702 0.00149427
R19252 VSS.n1507 VSS.n1504 0.00145036
R19253 VSS.n2044 VSS.n1507 0.00145036
R19254 VSS.n1506 VSS.n0 0.00143078
R19255 VSS.n2046 VSS.n0 0.00143078
R19256 VSS.n1700 VSS.n1699 0.00130794
R19257 VSS.n879 VSS.n878 0.00128125
R19258 VSS.n1338 VSS.n1334 0.00128125
R19259 VSS.n1348 VSS.n1347 0.00125806
R19260 VSS.n1482 VSS.n1481 0.00125806
R19261 VSS.n1513 VSS.n1510 0.00119582
R19262 VSS.n1510 VSS.n1506 0.00119582
R19263 VSS.n2043 VSS.n1508 0.00117624
R19264 VSS.n2044 VSS.n2043 0.00117624
R19265 VSS.n1268 VSS.n1267 0.00117024
R19266 VSS.n1483 VSS.n21 0.0011689
R19267 VSS.n472 VSS.n471 0.0011689
R19268 VSS.n1483 VSS.n24 0.0011689
R19269 VSS.n471 VSS.n468 0.0011689
R19270 VSS.n1503 VSS.n16 0.00116156
R19271 VSS.n842 VSS.n469 0.00116156
R19272 VSS.n22 VSS.n16 0.00116156
R19273 VSS.n844 VSS.n469 0.00116156
R19274 VSS.n589 VSS.n588 0.00113518
R19275 VSS.n1280 VSS.n1279 0.00113518
R19276 VSS.n1265 VSS.n1264 0.00113518
R19277 VSS.n1267 VSS.n196 0.00113518
R19278 VSS.n26 VSS.n25 0.00107344
R19279 VSS.n841 VSS.n450 0.00107344
R19280 VSS.n25 VSS.n22 0.00107344
R19281 VSS.n842 VSS.n841 0.00107344
R19282 VSS.n27 VSS.n24 0.00106609
R19283 VSS.n887 VSS.n460 0.00106609
R19284 VSS.n472 VSS.n460 0.00106609
R19285 VSS.n30 VSS.n27 0.00106609
R19286 VSS.n1265 VSS.n208 0.00105224
R19287 VSS.n1280 VSS.n190 0.00105224
R19288 VSS.n1037 VSS.n203 0.00100786
R19289 VSS.n579 VSS.n186 0.00100786
R19290 VSS.n589 VSS.n586 0.00100398
R19291 VSS.n1884 VSS.n1883 0.00100166
R19292 VSS.n1878 VSS.n1877 0.00100166
R19293 VSS.n1884 VSS.n1705 0.00100102
R19294 VSS.n1877 VSS.n1708 0.00100102
R19295 VSS.n1876 VSS.n1875 0.00100018
R19296 VSS.n1266 VSS.n203 0.00100009
R19297 VSS.n1281 VSS.n186 0.00100009
R19298 VSS.n578 VSS.n577 0.00100007
R19299 VSS.n1869 VSS.n1710 0.00100006
R19300 VSS.n603 VSS.n602 0.00100002
R19301 VSS.n1872 VSS.n1710 0.00100001
R19302 VSS.n1267 VSS.n1266 0.001
R19303 VSS.n1885 VSS.n1884 0.001
R19304 VSS.n1875 VSS.n1873 0.001
R19305 VSS.n1877 VSS.n1876 0.001
R19306 VSS.n590 VSS.n589 0.001
R19307 VSS.n1281 VSS.n1280 0.001
R19308 VSS.n1266 VSS.n1265 0.001
R19309 VSS.n880 VSS.n454 0.000752688
R19310 VSS.n1337 VSS.n1336 0.000752688
R19311 VSS.n1269 VSS.n1268 0.000670243
R19312 VSS.n588 VSS.n587 0.000635176
R19313 VSS.n1279 VSS.n1278 0.000635176
R19314 VSS.n1264 VSS.n1263 0.000635176
R19315 VSS.n1270 VSS.n196 0.000635176
R19316 VSS.n591 VSS.n590 0.000635176
R19317 VSS.n592 VSS.n591 0.000635176
R19318 VSS.n197 VSS.n195 0.000631513
R19319 VSS.n195 VSS.n187 0.000631513
R19320 VSS.n1262 VSS.n208 0.000552238
R19321 VSS.n1277 VSS.n190 0.000552238
R19322 VSS.n1036 VSS.n204 0.000512877
R19323 VSS.n1266 VSS.n204 0.000512877
R19324 VSS.n593 VSS.n584 0.00051244
R19325 VSS.n584 VSS.n583 0.00051244
R19326 VSS.n581 VSS.n188 0.000511972
R19327 VSS.n1281 VSS.n188 0.000511972
R19328 VSS.n193 VSS.n191 0.000509014
R19329 VSS.n596 VSS.n191 0.000509014
R19330 VSS.n1038 VSS.n1037 0.000507954
R19331 VSS.n580 VSS.n579 0.000507954
R19332 VSS.n1887 VSS.n1886 0.000505303
R19333 VSS.n1886 VSS.n1885 0.000505303
R19334 VSS.n1870 VSS.n1709 0.000505303
R19335 VSS.n1876 VSS.n1709 0.000505303
R19336 VSS.n586 VSS.n585 0.000503977
R19337 VSS.n1703 VSS.n1701 0.000503145
R19338 VSS.n1874 VSS.n1703 0.000503145
R19339 VSS.n1874 VSS.n1706 0.000503145
R19340 VSS.n1880 VSS.n1706 0.000503145
R19341 VSS.n1883 VSS.n1882 0.000501661
R19342 VSS.n1879 VSS.n1878 0.000501661
R19343 VSS.n194 VSS.n192 0.000501229
R19344 VSS.n212 VSS.n192 0.000501229
R19345 VSS.n1272 VSS.n1271 0.000501048
R19346 VSS.n1273 VSS.n1272 0.000501048
R19347 VSS.n1881 VSS.n1705 0.000501025
R19348 VSS.n1708 VSS.n1707 0.000501025
R19349 VSS.n596 VSS.n595 0.000500725
R19350 VSS.n595 VSS.n594 0.000500725
R19351 VSS.n582 VSS.n578 0.000500479
R19352 VSS.n597 VSS.n582 0.000500479
R19353 VSS.n1702 VSS.n1700 0.000500181
R19354 VSS.n1873 VSS.n1872 0.000500181
R19355 VSS.n604 VSS.n603 0.000500106
R19356 a_2151_4783.n51 a_2151_4783.t8 60.2505
R19357 a_2151_4783.n72 a_2151_4783.t9 60.2505
R19358 a_2151_4783.n94 a_2151_4783.t6 60.2505
R19359 a_2151_4783.n39 a_2151_4783.t4 60.2505
R19360 a_2151_4783.n5 a_2151_4783.n60 9.3005
R19361 a_2151_4783.n7 a_2151_4783.n64 9.3005
R19362 a_2151_4783.n8 a_2151_4783.n82 9.3005
R19363 a_2151_4783.n10 a_2151_4783.n86 9.3005
R19364 a_2151_4783.n11 a_2151_4783.n104 9.3005
R19365 a_2151_4783.n12 a_2151_4783.n48 9.3005
R19366 a_2151_4783.n12 a_2151_4783.n47 9.3005
R19367 a_2151_4783.n12 a_2151_4783.n46 9.3005
R19368 a_2151_4783.n46 a_2151_4783.n45 9.3005
R19369 a_2151_4783.n11 a_2151_4783.n103 9.3005
R19370 a_2151_4783.n11 a_2151_4783.n102 9.3005
R19371 a_2151_4783.n102 a_2151_4783.n101 9.3005
R19372 a_2151_4783.n10 a_2151_4783.n87 9.3005
R19373 a_2151_4783.n10 a_2151_4783.n93 9.3005
R19374 a_2151_4783.n93 a_2151_4783.n92 9.3005
R19375 a_2151_4783.n8 a_2151_4783.n81 9.3005
R19376 a_2151_4783.n8 a_2151_4783.n80 9.3005
R19377 a_2151_4783.n80 a_2151_4783.n79 9.3005
R19378 a_2151_4783.n7 a_2151_4783.n65 9.3005
R19379 a_2151_4783.n7 a_2151_4783.n71 9.3005
R19380 a_2151_4783.n71 a_2151_4783.n70 9.3005
R19381 a_2151_4783.n5 a_2151_4783.n58 9.3005
R19382 a_2151_4783.n58 a_2151_4783.n57 9.3005
R19383 a_2151_4783.n5 a_2151_4783.n59 9.3005
R19384 a_2151_4783.n0 a_2151_4783.n109 9.3005
R19385 a_2151_4783.n95 a_2151_4783.n94 8.76429
R19386 a_2151_4783.n73 a_2151_4783.n72 8.76429
R19387 a_2151_4783.n44 a_2151_4783.n43 7.45411
R19388 a_2151_4783.n100 a_2151_4783.n99 7.45411
R19389 a_2151_4783.n91 a_2151_4783.n90 7.45411
R19390 a_2151_4783.n78 a_2151_4783.n77 7.45411
R19391 a_2151_4783.n69 a_2151_4783.n68 7.45411
R19392 a_2151_4783.n56 a_2151_4783.n55 7.45411
R19393 a_2151_4783.n40 a_2151_4783.n39 6.80334
R19394 a_2151_4783.n52 a_2151_4783.n51 6.80105
R19395 a_2151_4783.n111 a_2151_4783.n110 6.31679
R19396 a_2151_4783.n42 a_2151_4783.n41 5.64756
R19397 a_2151_4783.n98 a_2151_4783.n97 5.64756
R19398 a_2151_4783.n89 a_2151_4783.n88 5.64756
R19399 a_2151_4783.n76 a_2151_4783.n75 5.64756
R19400 a_2151_4783.n67 a_2151_4783.n66 5.64756
R19401 a_2151_4783.n54 a_2151_4783.n53 5.64756
R19402 a_2151_4783.n112 a_2151_4783.t5 5.5395
R19403 a_2151_4783.t7 a_2151_4783.n112 5.5395
R19404 a_2151_4783.n0 a_2151_4783.n108 4.95534
R19405 a_2151_4783.n50 a_2151_4783.n49 4.73575
R19406 a_2151_4783.n106 a_2151_4783.n105 4.73575
R19407 a_2151_4783.n9 a_2151_4783.n85 4.73575
R19408 a_2151_4783.n84 a_2151_4783.n83 4.73575
R19409 a_2151_4783.n6 a_2151_4783.n63 4.73575
R19410 a_2151_4783.n62 a_2151_4783.n61 4.73575
R19411 a_2151_4783.n1 a_2151_4783.n13 4.6673
R19412 a_2151_4783.n96 a_2151_4783.n95 4.6505
R19413 a_2151_4783.n74 a_2151_4783.n73 4.6505
R19414 a_2151_4783.n4 a_2151_4783.n31 4.5005
R19415 a_2151_4783.n4 a_2151_4783.n28 4.5005
R19416 a_2151_4783.n2 a_2151_4783.n20 4.5005
R19417 a_2151_4783.n2 a_2151_4783.n23 4.5005
R19418 a_2151_4783.n0 a_2151_4783.n38 4.5005
R19419 a_2151_4783.n1 a_2151_4783.n36 4.5005
R19420 a_2151_4783.n1 a_2151_4783.n15 4.5005
R19421 a_2151_4783.n28 a_2151_4783.n27 4.14168
R19422 a_2151_4783.n23 a_2151_4783.n22 4.14168
R19423 a_2151_4783.n15 a_2151_4783.n14 3.76521
R19424 a_2151_4783.n5 a_2151_4783.n52 3.42768
R19425 a_2151_4783.n12 a_2151_4783.n40 3.42683
R19426 a_2151_4783.n38 a_2151_4783.n37 3.38874
R19427 a_2151_4783.n32 a_2151_4783.t1 3.3065
R19428 a_2151_4783.n32 a_2151_4783.t0 3.3065
R19429 a_2151_4783.n16 a_2151_4783.t3 3.3065
R19430 a_2151_4783.n16 a_2151_4783.t2 3.3065
R19431 a_2151_4783.n36 a_2151_4783.n35 3.01226
R19432 a_2151_4783.n30 a_2151_4783.n29 2.25932
R19433 a_2151_4783.n19 a_2151_4783.n18 2.25932
R19434 a_2151_4783.n111 a_2151_4783.n1 1.50789
R19435 a_2151_4783.n17 a_2151_4783.n16 1.46878
R19436 a_2151_4783.n45 a_2151_4783.n44 0.994314
R19437 a_2151_4783.n101 a_2151_4783.n100 0.994314
R19438 a_2151_4783.n92 a_2151_4783.n91 0.994314
R19439 a_2151_4783.n79 a_2151_4783.n78 0.994314
R19440 a_2151_4783.n70 a_2151_4783.n69 0.994314
R19441 a_2151_4783.n57 a_2151_4783.n56 0.994314
R19442 a_2151_4783.n34 a_2151_4783.n25 0.920917
R19443 a_2151_4783.n46 a_2151_4783.n42 0.753441
R19444 a_2151_4783.n102 a_2151_4783.n98 0.753441
R19445 a_2151_4783.n93 a_2151_4783.n89 0.753441
R19446 a_2151_4783.n80 a_2151_4783.n76 0.753441
R19447 a_2151_4783.n71 a_2151_4783.n67 0.753441
R19448 a_2151_4783.n58 a_2151_4783.n54 0.753441
R19449 a_2151_4783.n13 a_2151_4783.n2 0.70141
R19450 a_2151_4783.n13 a_2151_4783.n34 0.700686
R19451 a_2151_4783.n2 a_2151_4783.n24 0.604067
R19452 a_2151_4783.n25 a_2151_4783.n33 0.594011
R19453 a_2151_4783.n4 a_2151_4783.n32 2.11687
R19454 a_2151_4783.n3 a_2151_4783.n17 0.555028
R19455 a_2151_4783.n9 a_2151_4783.n84 0.458354
R19456 a_2151_4783.n6 a_2151_4783.n62 0.458354
R19457 a_2151_4783.n1 a_2151_4783.n0 0.452411
R19458 a_2151_4783.n112 a_2151_4783.n111 0.400755
R19459 a_2151_4783.n28 a_2151_4783.n26 0.376971
R19460 a_2151_4783.n31 a_2151_4783.n30 0.376971
R19461 a_2151_4783.n23 a_2151_4783.n21 0.376971
R19462 a_2151_4783.n20 a_2151_4783.n19 0.376971
R19463 a_2151_4783.n2 a_2151_4783.n3 0.29091
R19464 a_2151_4783.n107 a_2151_4783.n50 0.229427
R19465 a_2151_4783.n107 a_2151_4783.n106 0.229427
R19466 a_2151_4783.n0 a_2151_4783.n107 0.215848
R19467 a_2151_4783.n25 a_2151_4783.n4 0.206871
R19468 a_2151_4783.n50 a_2151_4783.n12 0.205546
R19469 a_2151_4783.n106 a_2151_4783.n11 0.205546
R19470 a_2151_4783.n10 a_2151_4783.n9 0.205546
R19471 a_2151_4783.n84 a_2151_4783.n8 0.205546
R19472 a_2151_4783.n7 a_2151_4783.n6 0.205546
R19473 a_2151_4783.n62 a_2151_4783.n5 0.205546
R19474 a_2151_4783.n11 a_2151_4783.n96 0.190717
R19475 a_2151_4783.n96 a_2151_4783.n10 0.190717
R19476 a_2151_4783.n8 a_2151_4783.n74 0.190717
R19477 a_2151_4783.n74 a_2151_4783.n7 0.190717
R19478 a_2551_4880.n76 a_2551_4880.t2 60.2505
R19479 a_2551_4880.n53 a_2551_4880.t7 60.2505
R19480 a_2551_4880.n30 a_2551_4880.t6 60.2505
R19481 a_2551_4880.n90 a_2551_4880.t0 60.2505
R19482 a_2551_4880.n140 a_2551_4880.n10 10.3264
R19483 a_2551_4880.n140 a_2551_4880.n11 9.57347
R19484 a_2551_4880.n7 a_2551_4880.n98 9.3005
R19485 a_2551_4880.n100 a_2551_4880.n99 9.3005
R19486 a_2551_4880.n7 a_2551_4880.n97 9.3005
R19487 a_2551_4880.n97 a_2551_4880.n96 9.3005
R19488 a_2551_4880.n64 a_2551_4880.n63 9.3005
R19489 a_2551_4880.n1 a_2551_4880.n45 9.3005
R19490 a_2551_4880.n40 a_2551_4880.n39 9.3005
R19491 a_2551_4880.n0 a_2551_4880.n38 9.3005
R19492 a_2551_4880.n0 a_2551_4880.n37 9.3005
R19493 a_2551_4880.n37 a_2551_4880.n36 9.3005
R19494 a_2551_4880.n2 a_2551_4880.n46 9.3005
R19495 a_2551_4880.n2 a_2551_4880.n52 9.3005
R19496 a_2551_4880.n52 a_2551_4880.n51 9.3005
R19497 a_2551_4880.n3 a_2551_4880.n62 9.3005
R19498 a_2551_4880.n3 a_2551_4880.n61 9.3005
R19499 a_2551_4880.n61 a_2551_4880.n60 9.3005
R19500 a_2551_4880.n4 a_2551_4880.n68 9.3005
R19501 a_2551_4880.n5 a_2551_4880.n75 9.3005
R19502 a_2551_4880.n75 a_2551_4880.n74 9.3005
R19503 a_2551_4880.n5 a_2551_4880.n69 9.3005
R19504 a_2551_4880.n6 a_2551_4880.n84 9.3005
R19505 a_2551_4880.n84 a_2551_4880.n83 9.3005
R19506 a_2551_4880.n87 a_2551_4880.n86 9.3005
R19507 a_2551_4880.n6 a_2551_4880.n85 9.3005
R19508 a_2551_4880.n112 a_2551_4880.n113 9.3005
R19509 a_2551_4880.n110 a_2551_4880.n111 9.3005
R19510 a_2551_4880.n108 a_2551_4880.n109 9.3005
R19511 a_2551_4880.n106 a_2551_4880.n107 9.3005
R19512 a_2551_4880.n105 a_2551_4880.n104 9.3005
R19513 a_2551_4880.n54 a_2551_4880.n53 8.76429
R19514 a_2551_4880.n77 a_2551_4880.n76 8.76429
R19515 a_2551_4880.n35 a_2551_4880.n34 8.21641
R19516 a_2551_4880.n50 a_2551_4880.n49 8.21641
R19517 a_2551_4880.n59 a_2551_4880.n58 8.21641
R19518 a_2551_4880.n95 a_2551_4880.n94 8.21641
R19519 a_2551_4880.n73 a_2551_4880.n72 8.21641
R19520 a_2551_4880.n82 a_2551_4880.n81 8.21641
R19521 a_2551_4880.n140 a_2551_4880.n27 8.139
R19522 a_2551_4880.n140 a_2551_4880.n24 8.11104
R19523 a_2551_4880.n140 a_2551_4880.n21 8.08351
R19524 a_2551_4880.n140 a_2551_4880.n18 8.05639
R19525 a_2551_4880.n133 a_2551_4880.n132 8.0439
R19526 a_2551_4880.n140 a_2551_4880.n15 8.02969
R19527 a_2551_4880.n140 a_2551_4880.n12 8.00339
R19528 a_2551_4880.n31 a_2551_4880.n30 6.92242
R19529 a_2551_4880.n91 a_2551_4880.n90 6.92012
R19530 a_2551_4880.n33 a_2551_4880.n32 5.64756
R19531 a_2551_4880.n48 a_2551_4880.n47 5.64756
R19532 a_2551_4880.n57 a_2551_4880.n56 5.64756
R19533 a_2551_4880.n93 a_2551_4880.n92 5.64756
R19534 a_2551_4880.n71 a_2551_4880.n70 5.64756
R19535 a_2551_4880.n80 a_2551_4880.n79 5.64756
R19536 a_2551_4880.n122 a_2551_4880.n120 5.62996
R19537 a_2551_4880.n127 a_2551_4880.t4 5.5395
R19538 a_2551_4880.n127 a_2551_4880.t5 5.5395
R19539 a_2551_4880.n42 a_2551_4880.n41 4.76425
R19540 a_2551_4880.n44 a_2551_4880.n43 4.76425
R19541 a_2551_4880.n66 a_2551_4880.n65 4.76425
R19542 a_2551_4880.n101 a_2551_4880.n89 4.76425
R19543 a_2551_4880.n67 a_2551_4880.n29 4.76425
R19544 a_2551_4880.n88 a_2551_4880.n28 4.76425
R19545 a_2551_4880.n55 a_2551_4880.n54 4.6505
R19546 a_2551_4880.n78 a_2551_4880.n77 4.6505
R19547 a_2551_4880.n9 a_2551_4880.n130 4.5005
R19548 a_2551_4880.n8 a_2551_4880.n126 4.5005
R19549 a_2551_4880.n135 a_2551_4880.n137 4.5005
R19550 a_2551_4880.n134 a_2551_4880.n133 4.5005
R19551 a_2551_4880.n117 a_2551_4880.n118 4.5005
R19552 a_2551_4880.n114 a_2551_4880.n116 4.5005
R19553 a_2551_4880.n14 a_2551_4880.n13 4.14168
R19554 a_2551_4880.n130 a_2551_4880.n129 3.76521
R19555 a_2551_4880.n7 a_2551_4880.n91 3.47756
R19556 a_2551_4880.n0 a_2551_4880.n31 3.4767
R19557 a_2551_4880.n126 a_2551_4880.n123 3.38874
R19558 a_2551_4880.n17 a_2551_4880.n16 3.38874
R19559 a_2551_4880.t3 a_2551_4880.n140 3.3065
R19560 a_2551_4880.n140 a_2551_4880.t1 3.3065
R19561 a_2551_4880.n126 a_2551_4880.n125 3.01226
R19562 a_2551_4880.n130 a_2551_4880.n128 2.63579
R19563 a_2551_4880.n20 a_2551_4880.n19 2.63579
R19564 a_2551_4880.n137 a_2551_4880.n136 2.63579
R19565 a_2551_4880.n116 a_2551_4880.n115 2.25932
R19566 a_2551_4880.n9 a_2551_4880.n127 1.90814
R19567 a_2551_4880.n23 a_2551_4880.n22 1.88285
R19568 a_2551_4880.n140 a_2551_4880.n139 1.52638
R19569 a_2551_4880.n26 a_2551_4880.n25 1.12991
R19570 a_2551_4880.n36 a_2551_4880.n35 1.09595
R19571 a_2551_4880.n51 a_2551_4880.n50 1.09595
R19572 a_2551_4880.n60 a_2551_4880.n59 1.09595
R19573 a_2551_4880.n96 a_2551_4880.n95 1.09595
R19574 a_2551_4880.n74 a_2551_4880.n73 1.09595
R19575 a_2551_4880.n83 a_2551_4880.n82 1.09595
R19576 a_2551_4880.n139 a_2551_4880.n138 0.93881
R19577 a_2551_4880.n37 a_2551_4880.n33 0.753441
R19578 a_2551_4880.n52 a_2551_4880.n48 0.753441
R19579 a_2551_4880.n61 a_2551_4880.n57 0.753441
R19580 a_2551_4880.n97 a_2551_4880.n93 0.753441
R19581 a_2551_4880.n75 a_2551_4880.n71 0.753441
R19582 a_2551_4880.n84 a_2551_4880.n80 0.753441
R19583 a_2551_4880.n15 a_2551_4880.n14 0.461175
R19584 a_2551_4880.n44 a_2551_4880.n42 0.458354
R19585 a_2551_4880.n67 a_2551_4880.n66 0.458354
R19586 a_2551_4880.n18 a_2551_4880.n17 0.430121
R19587 a_2551_4880.n21 a_2551_4880.n20 0.398603
R19588 a_2551_4880.n24 a_2551_4880.n23 0.366615
R19589 a_2551_4880.n27 a_2551_4880.n26 0.334147
R19590 a_2551_4880.n119 a_2551_4880.n122 0.27883
R19591 a_2551_4880.n102 a_2551_4880.n88 0.229427
R19592 a_2551_4880.n102 a_2551_4880.n101 0.229427
R19593 a_2551_4880.n103 a_2551_4880.n102 0.191391
R19594 a_2551_4880.n106 a_2551_4880.n105 0.190717
R19595 a_2551_4880.n108 a_2551_4880.n106 0.190717
R19596 a_2551_4880.n110 a_2551_4880.n108 0.190717
R19597 a_2551_4880.n112 a_2551_4880.n110 0.190717
R19598 a_2551_4880.n55 a_2551_4880.n2 0.190717
R19599 a_2551_4880.n3 a_2551_4880.n55 0.190717
R19600 a_2551_4880.n78 a_2551_4880.n5 0.190717
R19601 a_2551_4880.n6 a_2551_4880.n78 0.190717
R19602 a_2551_4880.n114 a_2551_4880.n112 0.169023
R19603 a_2551_4880.n105 a_2551_4880.n103 0.164777
R19604 a_2551_4880.n120 a_2551_4880.n121 0.161367
R19605 a_2551_4880.n42 a_2551_4880.n40 0.15935
R19606 a_2551_4880.n1 a_2551_4880.n44 0.15935
R19607 a_2551_4880.n66 a_2551_4880.n64 0.15935
R19608 a_2551_4880.n4 a_2551_4880.n67 0.15935
R19609 a_2551_4880.n88 a_2551_4880.n87 0.15935
R19610 a_2551_4880.n101 a_2551_4880.n100 0.15935
R19611 a_2551_4880.n123 a_2551_4880.n124 0.150167
R19612 a_2551_4880.n9 a_2551_4880.n8 0.143833
R19613 a_2551_4880.n8 a_2551_4880.n119 0.1366
R19614 a_2551_4880.n100 a_2551_4880.n7 0.0466957
R19615 a_2551_4880.n87 a_2551_4880.n6 0.0466957
R19616 a_2551_4880.n5 a_2551_4880.n4 0.0466957
R19617 a_2551_4880.n64 a_2551_4880.n3 0.0466957
R19618 a_2551_4880.n2 a_2551_4880.n1 0.0466957
R19619 a_2551_4880.n40 a_2551_4880.n0 0.0466957
R19620 a_2551_4880.n134 a_2551_4880.n131 0.0456361
R19621 a_2551_4880.n117 a_2551_4880.n114 0.0454219
R19622 a_2551_4880.n135 a_2551_4880.n134 0.0454219
R19623 a_2551_4880.n131 a_2551_4880.n117 0.045375
R19624 a_2551_4880.n138 a_2551_4880.n135 0.0439417
R19625 a_2551_4880.n131 a_2551_4880.n9 7.51529
R19626 a_8881_1782.n109 a_8881_1782.t2 120.501
R19627 a_8881_1782.n21 a_8881_1782.t0 69.2068
R19628 a_8881_1782.n59 a_8881_1782.t3 60.2505
R19629 a_8881_1782.n46 a_8881_1782.n45 31.4488
R19630 a_8881_1782.n24 a_8881_1782.n23 27.5177
R19631 a_8881_1782.n7 a_8881_1782.n3 26.107
R19632 a_8881_1782.n35 a_8881_1782.n34 23.5867
R19633 a_8881_1782.n13 a_8881_1782.n12 19.6557
R19634 a_8881_1782.n3 a_8881_1782.n2 15.7246
R19635 a_8881_1782.n14 a_8881_1782.n13 13.7591
R19636 a_8881_1782.n36 a_8881_1782.n35 9.82809
R19637 a_8881_1782.n86 a_8881_1782.n85 9.3005
R19638 a_8881_1782.n69 a_8881_1782.n68 9.3005
R19639 a_8881_1782.n123 a_8881_1782.n122 9.3005
R19640 a_8881_1782.n104 a_8881_1782.n103 9.3005
R19641 a_8881_1782.n50 a_8881_1782.n52 9.3005
R19642 a_8881_1782.n15 a_8881_1782.n14 9.3005
R19643 a_8881_1782.n37 a_8881_1782.n36 9.3005
R19644 a_8881_1782.n28 a_8881_1782.n38 9.3005
R19645 a_8881_1782.n26 a_8881_1782.n25 9.3005
R19646 a_8881_1782.n39 a_8881_1782.n41 9.3005
R19647 a_8881_1782.n48 a_8881_1782.n47 9.3005
R19648 a_8881_1782.n1 a_8881_1782.n139 9.3005
R19649 a_8881_1782.n131 a_8881_1782.n146 9.3005
R19650 a_8881_1782.n1 a_8881_1782.n138 9.3005
R19651 a_8881_1782.n0 a_8881_1782.n134 9.3005
R19652 a_8881_1782.n131 a_8881_1782.n145 9.3005
R19653 a_8881_1782.n60 a_8881_1782.n59 8.76429
R19654 a_8881_1782.n110 a_8881_1782.n109 8.76429
R19655 a_8881_1782.n67 a_8881_1782.n66 8.21641
R19656 a_8881_1782.n84 a_8881_1782.n83 8.21641
R19657 a_8881_1782.n102 a_8881_1782.n101 7.45411
R19658 a_8881_1782.n121 a_8881_1782.n120 7.45411
R19659 a_8881_1782.n25 a_8881_1782.n24 5.89705
R19660 a_8881_1782.n150 a_8881_1782.n149 5.38095
R19661 a_8881_1782.n8 a_8881_1782.n7 5.20544
R19662 a_8881_1782.n56 a_8881_1782.n54 4.87224
R19663 a_8881_1782.n89 a_8881_1782.n74 4.86623
R19664 a_8881_1782.n92 a_8881_1782.n90 4.84151
R19665 a_8881_1782.n126 a_8881_1782.n108 4.83995
R19666 a_8881_1782.n111 a_8881_1782.n110 4.6505
R19667 a_8881_1782.n0 a_8881_1782.n133 4.5298
R19668 a_8881_1782.n30 a_8881_1782.n31 4.51815
R19669 a_8881_1782.n33 a_8881_1782.n32 4.51815
R19670 a_8881_1782.n55 a_8881_1782.n70 4.5005
R19671 a_8881_1782.n57 a_8881_1782.n63 4.5005
R19672 a_8881_1782.n77 a_8881_1782.n81 4.5005
R19673 a_8881_1782.n82 a_8881_1782.n88 4.5005
R19674 a_8881_1782.n91 a_8881_1782.n105 4.5005
R19675 a_8881_1782.n93 a_8881_1782.n98 4.5005
R19676 a_8881_1782.n114 a_8881_1782.n118 4.5005
R19677 a_8881_1782.n119 a_8881_1782.n125 4.5005
R19678 a_8881_1782.n8 a_8881_1782.n16 4.5005
R19679 a_8881_1782.n42 a_8881_1782.n49 4.5005
R19680 a_8881_1782.n29 a_8881_1782.n27 4.5005
R19681 a_8881_1782.n94 a_8881_1782.n95 4.5005
R19682 a_8881_1782.n113 a_8881_1782.n112 4.5005
R19683 a_8881_1782.n1 a_8881_1782.n137 4.5005
R19684 a_8881_1782.n130 a_8881_1782.n144 4.5005
R19685 a_8881_1782.n58 a_8881_1782.n60 4.14168
R19686 a_8881_1782.n76 a_8881_1782.n75 4.14168
R19687 a_8881_1782.n49 a_8881_1782.n43 4.14168
R19688 a_8881_1782.n88 a_8881_1782.n86 3.76521
R19689 a_8881_1782.n125 a_8881_1782.n123 3.76521
R19690 a_8881_1782.n16 a_8881_1782.n9 3.76521
R19691 a_8881_1782.n11 a_8881_1782.n10 3.76521
R19692 a_8881_1782.n70 a_8881_1782.n69 3.38874
R19693 a_8881_1782.n105 a_8881_1782.n104 3.38874
R19694 a_8881_1782.n6 a_8881_1782.n5 3.38874
R19695 a_8881_1782.n130 a_8881_1782.n141 3.17178
R19696 a_8881_1782.n70 a_8881_1782.n64 3.01226
R19697 a_8881_1782.n81 a_8881_1782.n80 3.01226
R19698 a_8881_1782.n105 a_8881_1782.n99 3.01226
R19699 a_8881_1782.n98 a_8881_1782.n96 3.01226
R19700 a_8881_1782.n5 a_8881_1782.n4 3.01226
R19701 a_8881_1782.t1 a_8881_1782.n151 2.77
R19702 a_8881_1782.n63 a_8881_1782.n61 2.63579
R19703 a_8881_1782.n88 a_8881_1782.n87 2.63579
R19704 a_8881_1782.n118 a_8881_1782.n117 2.63579
R19705 a_8881_1782.n125 a_8881_1782.n124 2.63579
R19706 a_8881_1782.n16 a_8881_1782.n15 2.63579
R19707 a_8881_1782.n15 a_8881_1782.n11 2.63579
R19708 a_8881_1782.n53 a_8881_1782.n21 2.41452
R19709 a_8881_1782.n107 a_8881_1782.n127 2.28493
R19710 a_8881_1782.n49 a_8881_1782.n48 2.25932
R19711 a_8881_1782.n52 a_8881_1782.n51 2.25932
R19712 a_8881_1782.n47 a_8881_1782.n46 1.96602
R19713 a_8881_1782.n30 a_8881_1782.n37 1.88285
R19714 a_8881_1782.n37 a_8881_1782.n33 1.88285
R19715 a_8881_1782.n151 a_8881_1782.n150 1.84417
R19716 a_8881_1782.n81 a_8881_1782.n78 1.50638
R19717 a_8881_1782.n118 a_8881_1782.n115 1.50638
R19718 a_8881_1782.n117 a_8881_1782.n116 1.50638
R19719 a_8881_1782.n27 a_8881_1782.n26 1.50638
R19720 a_8881_1782.n41 a_8881_1782.n40 1.50638
R19721 a_8881_1782.n151 a_8881_1782.n140 1.32032
R19722 a_8881_1782.n151 a_8881_1782.n148 1.29978
R19723 a_8881_1782.n18 a_8881_1782.n129 1.24675
R19724 a_8881_1782.n107 a_8881_1782.n92 1.21366
R19725 a_8881_1782.n71 a_8881_1782.n89 1.15702
R19726 a_8881_1782.n73 a_8881_1782.n56 1.21147
R19727 a_8881_1782.n106 a_8881_1782.n126 1.15482
R19728 a_8881_1782.n63 a_8881_1782.n62 1.12991
R19729 a_8881_1782.n80 a_8881_1782.n79 1.12991
R19730 a_8881_1782.n98 a_8881_1782.n97 1.12991
R19731 a_8881_1782.n26 a_8881_1782.n22 1.12991
R19732 a_8881_1782.n68 a_8881_1782.n67 1.09595
R19733 a_8881_1782.n85 a_8881_1782.n84 1.09595
R19734 a_8881_1782.n1 a_8881_1782.n132 1.04835
R19735 a_8881_1782.n147 a_8881_1782.n127 0.996877
R19736 a_8881_1782.n103 a_8881_1782.n102 0.994314
R19737 a_8881_1782.n122 a_8881_1782.n121 0.994314
R19738 a_8881_1782.n17 a_8881_1782.n53 0.994096
R19739 a_8881_1782.n72 a_8881_1782.n128 0.963
R19740 a_8881_1782.n69 a_8881_1782.n65 0.753441
R19741 a_8881_1782.n104 a_8881_1782.n100 0.753441
R19742 a_8881_1782.n137 a_8881_1782.n135 0.753441
R19743 a_8881_1782.n140 a_8881_1782.n1 0.418831
R19744 a_8881_1782.n148 a_8881_1782.n147 0.386668
R19745 a_8881_1782.n48 a_8881_1782.n44 0.376971
R19746 a_8881_1782.n144 a_8881_1782.n142 0.376971
R19747 a_8881_1782.n7 a_8881_1782.n6 0.319725
R19748 a_8881_1782.n135 a_8881_1782.n136 0.121922
R19749 a_8881_1782.n142 a_8881_1782.n143 0.110027
R19750 a_8881_1782.n147 a_8881_1782.n131 0.0843535
R19751 a_8881_1782.n53 a_8881_1782.n50 0.0827519
R19752 a_8881_1782.n107 a_8881_1782.n106 0.0590938
R19753 a_8881_1782.n42 a_8881_1782.n39 0.100109
R19754 a_8881_1782.n126 a_8881_1782.n119 0.0371012
R19755 a_8881_1782.n131 a_8881_1782.n130 0.0337031
R19756 a_8881_1782.n20 a_8881_1782.n18 0.0287031
R19757 a_8881_1782.n20 a_8881_1782.n19 0.028
R19758 a_8881_1782.n128 a_8881_1782.n107 0.028
R19759 a_8881_1782.n129 a_8881_1782.n73 0.028
R19760 a_8881_1782.n73 a_8881_1782.n72 0.0276737
R19761 a_8881_1782.n113 a_8881_1782.n111 0.0239375
R19762 a_8881_1782.n77 a_8881_1782.n76 4.5892
R19763 a_8881_1782.n114 a_8881_1782.n113 0.0892218
R19764 a_8881_1782.n93 a_8881_1782.n94 0.0883906
R19765 a_8881_1782.n57 a_8881_1782.n58 4.58839
R19766 a_8881_1782.n20 a_8881_1782.n17 0.119641
R19767 a_8881_1782.n28 a_8881_1782.n30 4.61452
R19768 a_8881_1782.n73 a_8881_1782.n71 0.0590938
R19769 a_8881_1782.n82 a_8881_1782.n77 0.0454219
R19770 a_8881_1782.n119 a_8881_1782.n114 0.0454219
R19771 a_8881_1782.n91 a_8881_1782.n93 0.0454219
R19772 a_8881_1782.n55 a_8881_1782.n57 0.0454219
R19773 a_8881_1782.n92 a_8881_1782.n91 0.0388205
R19774 a_8881_1782.n89 a_8881_1782.n82 0.0385721
R19775 a_8881_1782.n56 a_8881_1782.n55 0.0373496
R19776 a_8881_1782.n50 a_8881_1782.n42 0.0337031
R19777 a_8881_1782.n39 a_8881_1782.n29 0.0337031
R19778 a_8881_1782.n29 a_8881_1782.n28 0.0268395
R19779 a_8881_1782.n20 a_8881_1782.n8 1.5962
R19780 a_8881_1782.n1 a_8881_1782.n0 0.225375
R19781 DVSS.n749 DVSS.n616 234025
R19782 DVSS.n712 DVSS.n616 200023
R19783 DVSS.n3009 DVSS.n3008 109580
R19784 DVSS.n1271 DVSS.n713 69276.6
R19785 DVSS.n2609 DVSS.n748 39364.3
R19786 DVSS.n2611 DVSS.n748 33314.3
R19787 DVSS.n1753 DVSS.n1750 26823.1
R19788 DVSS.n2767 DVSS.n712 20457
R19789 DVSS.n661 DVSS.n621 18393.1
R19790 DVSS.n2691 DVSS.n2662 18000.5
R19791 DVSS.n1753 DVSS.n1752 17938.5
R19792 DVSS.n3009 DVSS.n616 17383.3
R19793 DVSS.n2821 DVSS.n2820 16981.8
R19794 DVSS.n2870 DVSS.n2869 14490.1
R19795 DVSS.n2516 DVSS.n1750 14342.3
R19796 DVSS.n3010 DVSS.n3009 12571
R19797 DVSS.n756 DVSS.n616 11429.2
R19798 DVSS.n712 DVSS.n621 9964.45
R19799 DVSS.n2856 DVSS.n2855 9138.82
R19800 DVSS.n2873 DVSS.n2872 8030
R19801 DVSS.n2794 DVSS.t94 8003.11
R19802 DVSS.n1916 DVSS.t43 8003.11
R19803 DVSS.t189 DVSS.n2568 8003.11
R19804 DVSS.t148 DVSS.n3038 8003.11
R19805 DVSS.t100 DVSS.t98 7626.67
R19806 DVSS.t96 DVSS.t94 7626.67
R19807 DVSS.t47 DVSS.t45 7626.67
R19808 DVSS.t43 DVSS.t51 7626.67
R19809 DVSS.t183 DVSS.t185 7626.67
R19810 DVSS.t189 DVSS.t181 7626.67
R19811 DVSS.t150 DVSS.t152 7626.67
R19812 DVSS.t146 DVSS.t148 7626.67
R19813 DVSS.n2856 DVSS.n631 7326.61
R19814 DVSS.n3053 DVSS.n22 7144.95
R19815 DVSS.n2440 DVSS.n1779 7104.59
R19816 DVSS.n2519 DVSS.n2518 6853.25
R19817 DVSS.n2427 DVSS.n1779 6723.32
R19818 DVSS.n3054 DVSS.n3053 6716.07
R19819 DVSS.n3010 DVSS.n615 6566.79
R19820 DVSS.n2834 DVSS.t126 6153.5
R19821 DVSS.t132 DVSS.n55 6153.5
R19822 DVSS.n2820 DVSS.n2819 5998.54
R19823 DVSS.n2855 DVSS.n2854 5096.51
R19824 DVSS.n3008 DVSS.n617 5078.3
R19825 DVSS.n3007 DVSS.n2870 4670.31
R19826 DVSS.n2869 DVSS.n2868 4655.91
R19827 DVSS.n3011 DVSS.n3010 4524.16
R19828 DVSS.n2873 DVSS.t33 4455
R19829 DVSS.n2440 DVSS.n2439 3438.1
R19830 DVSS.n2679 DVSS.n22 3438.1
R19831 DVSS.n1753 DVSS.n701 3433.78
R19832 DVSS.n1754 DVSS.n1753 3433.78
R19833 DVSS.n2662 DVSS.n2661 3276.86
R19834 DVSS.n2869 DVSS.n622 3274.06
R19835 DVSS.n2766 DVSS.n2765 3274.06
R19836 DVSS.n1836 DVSS.n631 3140.39
R19837 DVSS.n2717 DVSS.n748 2954.65
R19838 DVSS.n2597 DVSS.n748 2954.65
R19839 DVSS.n2427 DVSS.n9 2882.84
R19840 DVSS.n3055 DVSS.n3054 2865.59
R19841 DVSS.n1946 DVSS.n661 2607.41
R19842 DVSS.t30 DVSS.n618 2554.84
R19843 DVSS.t35 DVSS.t33 2310
R19844 DVSS.n2822 DVSS.n2821 2223.27
R19845 DVSS.n2692 DVSS.n2691 2223.27
R19846 DVSS.t14 DVSS.t16 2165.3
R19847 DVSS.n2821 DVSS.n660 1865.51
R19848 DVSS.n2691 DVSS.n2690 1865.51
R19849 DVSS.t118 DVSS.t120 1778.24
R19850 DVSS.t130 DVSS.t134 1778.24
R19851 DVSS.t120 DVSS.n1916 1652.85
R19852 DVSS.n3038 DVSS.t130 1652.85
R19853 DVSS.n2518 DVSS.n2517 1501.28
R19854 DVSS.n3007 DVSS.n3006 1366.89
R19855 DVSS.n2820 DVSS.n661 1280.42
R19856 DVSS.n2872 DVSS.t35 1265
R19857 DVSS.n2610 DVSS.n2609 1158.66
R19858 DVSS.n2609 DVSS.n1228 1114.67
R19859 DVSS.n1271 DVSS.t14 1068.77
R19860 DVSS.n384 DVSS.n247 1013.97
R19861 DVSS.n382 DVSS.n248 1013.97
R19862 DVSS.n374 DVSS.n373 1013.97
R19863 DVSS.n376 DVSS.n368 1013.97
R19864 DVSS.n2257 DVSS.n2120 1013.97
R19865 DVSS.n2255 DVSS.n2121 1013.97
R19866 DVSS.n2247 DVSS.n2246 1013.97
R19867 DVSS.n2249 DVSS.n2241 1013.97
R19868 DVSS.n1065 DVSS.n928 1013.97
R19869 DVSS.n1063 DVSS.n929 1013.97
R19870 DVSS.n1055 DVSS.n1054 1013.97
R19871 DVSS.n1057 DVSS.n1049 1013.97
R19872 DVSS.n1587 DVSS.n1450 1013.97
R19873 DVSS.n1585 DVSS.n1451 1013.97
R19874 DVSS.n1577 DVSS.n1576 1013.97
R19875 DVSS.n1579 DVSS.n1571 1013.97
R19876 DVSS.n3083 DVSS.n3082 947.086
R19877 DVSS.n3081 DVSS.n9 947.086
R19878 DVSS.n3069 DVSS.n3068 938.668
R19879 DVSS.n3067 DVSS.n3055 938.668
R19880 DVSS.n2854 DVSS.t90 878.028
R19881 DVSS.n1228 DVSS.t0 870.222
R19882 DVSS.t30 DVSS.n620 868.74
R19883 DVSS.n2822 DVSS.n653 823.393
R19884 DVSS.n2692 DVSS.n2610 823.393
R19885 DVSS.n2832 DVSS.n653 790.293
R19886 DVSS.n1837 DVSS.n1836 783.674
R19887 DVSS.n1849 DVSS.n1848 783.674
R19888 DVSS.n1862 DVSS.n1809 783.674
R19889 DVSS.n2853 DVSS.n633 783.674
R19890 DVSS.n2845 DVSS.n633 783.674
R19891 DVSS.n2843 DVSS.n642 783.674
R19892 DVSS.n2835 DVSS.n642 783.674
R19893 DVSS.n2833 DVSS.n2832 783.674
R19894 DVSS.n2532 DVSS.n1261 771.409
R19895 DVSS.n3008 DVSS.n3007 756.131
R19896 DVSS.n2654 DVSS.n2619 744.975
R19897 DVSS.n2653 DVSS.n2652 744.975
R19898 DVSS.n2652 DVSS.n2620 744.975
R19899 DVSS.n2644 DVSS.n2620 744.975
R19900 DVSS.n2644 DVSS.n2643 744.975
R19901 DVSS.n2643 DVSS.n2642 744.975
R19902 DVSS.n2642 DVSS.n2627 744.975
R19903 DVSS.n1889 DVSS.n1877 744.975
R19904 DVSS.n1891 DVSS.n1890 744.975
R19905 DVSS.n1891 DVSS.n1871 744.975
R19906 DVSS.n1899 DVSS.n1871 744.975
R19907 DVSS.n1900 DVSS.n1899 744.975
R19908 DVSS.n1901 DVSS.n1900 744.975
R19909 DVSS.n1901 DVSS.n1863 744.975
R19910 DVSS.n2764 DVSS.n715 744.975
R19911 DVSS.n2754 DVSS.n726 744.975
R19912 DVSS.n2754 DVSS.n2753 744.975
R19913 DVSS.n2753 DVSS.n2752 744.975
R19914 DVSS.n2752 DVSS.n727 744.975
R19915 DVSS.n2744 DVSS.n727 744.975
R19916 DVSS.n2816 DVSS.n2815 744.975
R19917 DVSS.n2814 DVSS.n665 744.975
R19918 DVSS.n679 DVSS.n665 744.975
R19919 DVSS.n2805 DVSS.n679 744.975
R19920 DVSS.n2805 DVSS.n2804 744.975
R19921 DVSS.n2804 DVSS.n2803 744.975
R19922 DVSS.n1915 DVSS.n1863 744.975
R19923 DVSS.n1808 DVSS.n1806 744.975
R19924 DVSS.n1917 DVSS.n1793 744.975
R19925 DVSS.n1944 DVSS.n1793 744.975
R19926 DVSS.n1945 DVSS.n1944 744.975
R19927 DVSS.n1946 DVSS.n1945 744.975
R19928 DVSS.n2634 DVSS.n2627 744.975
R19929 DVSS.n3037 DVSS.n42 744.975
R19930 DVSS.n3022 DVSS.n56 744.975
R19931 DVSS.n66 DVSS.n56 744.975
R19932 DVSS.n3012 DVSS.n66 744.975
R19933 DVSS.n3012 DVSS.n3011 744.975
R19934 DVSS.n263 DVSS.n255 728.663
R19935 DVSS.n404 DVSS.n229 728.663
R19936 DVSS.n2136 DVSS.n2128 728.663
R19937 DVSS.n2277 DVSS.n2102 728.663
R19938 DVSS.n944 DVSS.n936 728.663
R19939 DVSS.n1085 DVSS.n910 728.663
R19940 DVSS.n1466 DVSS.n1458 728.663
R19941 DVSS.n1607 DVSS.n1432 728.663
R19942 DVSS.n359 DVSS.n254 668.5
R19943 DVSS.n357 DVSS.n257 668.5
R19944 DVSS.n406 DVSS.n226 668.5
R19945 DVSS.n366 DVSS.n230 668.5
R19946 DVSS.n334 DVSS.n313 668.5
R19947 DVSS.n338 DVSS.n315 668.5
R19948 DVSS.n349 DVSS.n311 668.5
R19949 DVSS.n352 DVSS.n351 668.5
R19950 DVSS.n179 DVSS.n151 668.5
R19951 DVSS.n164 DVSS.n149 668.5
R19952 DVSS.n521 DVSS.n520 668.5
R19953 DVSS.n536 DVSS.n535 668.5
R19954 DVSS.n2232 DVSS.n2127 668.5
R19955 DVSS.n2230 DVSS.n2130 668.5
R19956 DVSS.n2279 DVSS.n2099 668.5
R19957 DVSS.n2239 DVSS.n2103 668.5
R19958 DVSS.n2207 DVSS.n2186 668.5
R19959 DVSS.n2211 DVSS.n2188 668.5
R19960 DVSS.n2222 DVSS.n2184 668.5
R19961 DVSS.n2225 DVSS.n2224 668.5
R19962 DVSS.n2052 DVSS.n2024 668.5
R19963 DVSS.n2037 DVSS.n2022 668.5
R19964 DVSS.n2394 DVSS.n2393 668.5
R19965 DVSS.n2409 DVSS.n2408 668.5
R19966 DVSS.n1040 DVSS.n935 668.5
R19967 DVSS.n1038 DVSS.n938 668.5
R19968 DVSS.n1087 DVSS.n907 668.5
R19969 DVSS.n1047 DVSS.n911 668.5
R19970 DVSS.n1015 DVSS.n994 668.5
R19971 DVSS.n1019 DVSS.n996 668.5
R19972 DVSS.n1030 DVSS.n992 668.5
R19973 DVSS.n1033 DVSS.n1032 668.5
R19974 DVSS.n860 DVSS.n832 668.5
R19975 DVSS.n845 DVSS.n830 668.5
R19976 DVSS.n1202 DVSS.n1201 668.5
R19977 DVSS.n1217 DVSS.n1216 668.5
R19978 DVSS.n1562 DVSS.n1457 668.5
R19979 DVSS.n1560 DVSS.n1460 668.5
R19980 DVSS.n1609 DVSS.n1429 668.5
R19981 DVSS.n1569 DVSS.n1433 668.5
R19982 DVSS.n1537 DVSS.n1516 668.5
R19983 DVSS.n1541 DVSS.n1518 668.5
R19984 DVSS.n1552 DVSS.n1514 668.5
R19985 DVSS.n1555 DVSS.n1554 668.5
R19986 DVSS.n1382 DVSS.n1354 668.5
R19987 DVSS.n1367 DVSS.n1352 668.5
R19988 DVSS.n1724 DVSS.n1723 668.5
R19989 DVSS.n1739 DVSS.n1738 668.5
R19990 DVSS.t120 DVSS.n1807 667.372
R19991 DVSS.t130 DVSS.n41 667.372
R19992 DVSS.n2661 DVSS.t92 659.612
R19993 DVSS.t176 DVSS.n622 659.612
R19994 DVSS.n2765 DVSS.t88 659.612
R19995 DVSS.n2819 DVSS.t140 659.612
R19996 DVSS.n2855 DVSS.n2853 653.062
R19997 DVSS.n2870 DVSS.n621 648.317
R19998 DVSS.n2872 DVSS.t4 643.51
R19999 DVSS.n1850 DVSS.t49 636.567
R20000 DVSS.n1838 DVSS.t51 622.577
R20001 DVSS.n2835 DVSS.n2834 587.755
R20002 DVSS.n448 DVSS.n113 562.173
R20003 DVSS.n496 DVSS.n97 562.173
R20004 DVSS.n2321 DVSS.n1986 562.173
R20005 DVSS.n2369 DVSS.n1970 562.173
R20006 DVSS.n1129 DVSS.n794 562.173
R20007 DVSS.n1177 DVSS.n778 562.173
R20008 DVSS.n1651 DVSS.n1316 562.173
R20009 DVSS.n1699 DVSS.n1300 562.173
R20010 DVSS.n2518 DVSS.n2516 550
R20011 DVSS.t122 DVSS.n1807 543.211
R20012 DVSS.n41 DVSS.t138 543.211
R20013 DVSS.n2988 DVSS.n2987 539.294
R20014 DVSS.n2984 DVSS.n2983 539.294
R20015 DVSS.n2975 DVSS.n2974 539.294
R20016 DVSS.n2971 DVSS.n2970 539.294
R20017 DVSS.n2689 DVSS.n2663 539.294
R20018 DVSS.n2682 DVSS.n2663 539.294
R20019 DVSS.n2682 DVSS.n2681 539.294
R20020 DVSS.n2681 DVSS.n2678 539.294
R20021 DVSS.n3051 DVSS.n24 539.294
R20022 DVSS.n3051 DVSS.n25 539.294
R20023 DVSS.n34 DVSS.n25 539.294
R20024 DVSS.n3042 DVSS.n34 539.294
R20025 DVSS.n3042 DVSS.n35 539.294
R20026 DVSS.n37 DVSS.n35 539.294
R20027 DVSS.n567 DVSS.n37 539.294
R20028 DVSS.n568 DVSS.n567 539.294
R20029 DVSS.n568 DVSS.n556 539.294
R20030 DVSS.n576 DVSS.n556 539.294
R20031 DVSS.n576 DVSS.n555 539.294
R20032 DVSS.n581 DVSS.n555 539.294
R20033 DVSS.n581 DVSS.n549 539.294
R20034 DVSS.n595 DVSS.n549 539.294
R20035 DVSS.n595 DVSS.n547 539.294
R20036 DVSS.n599 DVSS.n547 539.294
R20037 DVSS.n600 DVSS.n599 539.294
R20038 DVSS.n603 DVSS.n600 539.294
R20039 DVSS.n603 DVSS.n68 539.294
R20040 DVSS.n614 DVSS.n68 539.294
R20041 DVSS.n2660 DVSS.n2612 539.294
R20042 DVSS.n2655 DVSS.n2612 539.294
R20043 DVSS.n2655 DVSS.n2618 539.294
R20044 DVSS.n2651 DVSS.n2618 539.294
R20045 DVSS.n2651 DVSS.n2621 539.294
R20046 DVSS.n2645 DVSS.n2621 539.294
R20047 DVSS.n2645 DVSS.n2626 539.294
R20048 DVSS.n2641 DVSS.n2626 539.294
R20049 DVSS.n2641 DVSS.n2628 539.294
R20050 DVSS.n2635 DVSS.n2628 539.294
R20051 DVSS.n2635 DVSS.n43 539.294
R20052 DVSS.n3036 DVSS.n43 539.294
R20053 DVSS.n3036 DVSS.n44 539.294
R20054 DVSS.n53 DVSS.n44 539.294
R20055 DVSS.n3026 DVSS.n53 539.294
R20056 DVSS.n3026 DVSS.n54 539.294
R20057 DVSS.n3021 DVSS.n54 539.294
R20058 DVSS.n3021 DVSS.n57 539.294
R20059 DVSS.n64 DVSS.n57 539.294
R20060 DVSS.n3013 DVSS.n64 539.294
R20061 DVSS.n3013 DVSS.n65 539.294
R20062 DVSS.n3070 DVSS.n16 539.294
R20063 DVSS.n3070 DVSS.n19 539.294
R20064 DVSS.n3066 DVSS.n19 539.294
R20065 DVSS.n3066 DVSS.n3056 539.294
R20066 DVSS.n2425 DVSS.n2424 539.294
R20067 DVSS.n2429 DVSS.n2425 539.294
R20068 DVSS.n2429 DVSS.n1783 539.294
R20069 DVSS.n2438 DVSS.n1783 539.294
R20070 DVSS.n2866 DVSS.n623 539.294
R20071 DVSS.n2866 DVSS.n625 539.294
R20072 DVSS.n2859 DVSS.n625 539.294
R20073 DVSS.n2859 DVSS.n630 539.294
R20074 DVSS.n1880 DVSS.n1878 539.294
R20075 DVSS.n1888 DVSS.n1878 539.294
R20076 DVSS.n1888 DVSS.n1876 539.294
R20077 DVSS.n1892 DVSS.n1876 539.294
R20078 DVSS.n1892 DVSS.n1872 539.294
R20079 DVSS.n1898 DVSS.n1872 539.294
R20080 DVSS.n1898 DVSS.n1870 539.294
R20081 DVSS.n1902 DVSS.n1870 539.294
R20082 DVSS.n1902 DVSS.n1864 539.294
R20083 DVSS.n1914 DVSS.n1864 539.294
R20084 DVSS.n1914 DVSS.n1865 539.294
R20085 DVSS.n1906 DVSS.n1865 539.294
R20086 DVSS.n1906 DVSS.n1804 539.294
R20087 DVSS.n1927 DVSS.n1804 539.294
R20088 DVSS.n1927 DVSS.n1805 539.294
R20089 DVSS.n1923 DVSS.n1805 539.294
R20090 DVSS.n1923 DVSS.n1918 539.294
R20091 DVSS.n1918 DVSS.n1794 539.294
R20092 DVSS.n1943 DVSS.n1794 539.294
R20093 DVSS.n1943 DVSS.n1792 539.294
R20094 DVSS.n1947 DVSS.n1792 539.294
R20095 DVSS.n1835 DVSS.n1823 539.294
R20096 DVSS.n1835 DVSS.n1821 539.294
R20097 DVSS.n1851 DVSS.n1821 539.294
R20098 DVSS.n1851 DVSS.n1822 539.294
R20099 DVSS.n1847 DVSS.n1822 539.294
R20100 DVSS.n1847 DVSS.n1839 539.294
R20101 DVSS.n1839 DVSS.n1810 539.294
R20102 DVSS.n1861 DVSS.n1810 539.294
R20103 DVSS.n1861 DVSS.n634 539.294
R20104 DVSS.n2852 DVSS.n634 539.294
R20105 DVSS.n2852 DVSS.n635 539.294
R20106 DVSS.n2846 DVSS.n635 539.294
R20107 DVSS.n2846 DVSS.n641 539.294
R20108 DVSS.n2842 DVSS.n641 539.294
R20109 DVSS.n2842 DVSS.n643 539.294
R20110 DVSS.n2836 DVSS.n643 539.294
R20111 DVSS.n2836 DVSS.n652 539.294
R20112 DVSS.n2831 DVSS.n652 539.294
R20113 DVSS.n2831 DVSS.n654 539.294
R20114 DVSS.n2823 DVSS.n654 539.294
R20115 DVSS.n2763 DVSS.n714 539.294
R20116 DVSS.n2763 DVSS.n716 539.294
R20117 DVSS.n724 DVSS.n716 539.294
R20118 DVSS.n2755 DVSS.n724 539.294
R20119 DVSS.n2755 DVSS.n725 539.294
R20120 DVSS.n2751 DVSS.n725 539.294
R20121 DVSS.n2751 DVSS.n728 539.294
R20122 DVSS.n2745 DVSS.n728 539.294
R20123 DVSS.n2745 DVSS.n732 539.294
R20124 DVSS.n2741 DVSS.n732 539.294
R20125 DVSS.n2741 DVSS.n733 539.294
R20126 DVSS.n2733 DVSS.n733 539.294
R20127 DVSS.n2733 DVSS.n740 539.294
R20128 DVSS.n2729 DVSS.n740 539.294
R20129 DVSS.n2729 DVSS.n742 539.294
R20130 DVSS.n2720 DVSS.n742 539.294
R20131 DVSS.n2720 DVSS.n747 539.294
R20132 DVSS.n2715 DVSS.n747 539.294
R20133 DVSS.n2715 DVSS.n750 539.294
R20134 DVSS.n2708 DVSS.n750 539.294
R20135 DVSS.n2544 DVSS.n1262 539.294
R20136 DVSS.n2544 DVSS.n1260 539.294
R20137 DVSS.n2548 DVSS.n1260 539.294
R20138 DVSS.n2548 DVSS.n1253 539.294
R20139 DVSS.n2564 DVSS.n1253 539.294
R20140 DVSS.n2564 DVSS.n1254 539.294
R20141 DVSS.n1254 DVSS.n1250 539.294
R20142 DVSS.n1250 DVSS.n1248 539.294
R20143 DVSS.n2570 DVSS.n1248 539.294
R20144 DVSS.n2570 DVSS.n1242 539.294
R20145 DVSS.n2578 DVSS.n1242 539.294
R20146 DVSS.n2578 DVSS.n1240 539.294
R20147 DVSS.n2583 DVSS.n1240 539.294
R20148 DVSS.n2583 DVSS.n1235 539.294
R20149 DVSS.n2594 DVSS.n1235 539.294
R20150 DVSS.n2594 DVSS.n1234 539.294
R20151 DVSS.n2599 DVSS.n1234 539.294
R20152 DVSS.n2599 DVSS.n1230 539.294
R20153 DVSS.n2607 DVSS.n1230 539.294
R20154 DVSS.n2607 DVSS.n1227 539.294
R20155 DVSS.n2693 DVSS.n1227 539.294
R20156 DVSS.n2529 DVSS.n1272 539.294
R20157 DVSS.n2529 DVSS.n1269 539.294
R20158 DVSS.n2534 DVSS.n1269 539.294
R20159 DVSS.n2534 DVSS.n1270 539.294
R20160 DVSS.n2447 DVSS.n1780 539.294
R20161 DVSS.n2447 DVSS.n1777 539.294
R20162 DVSS.n2469 DVSS.n1777 539.294
R20163 DVSS.n2469 DVSS.n1778 539.294
R20164 DVSS.n2465 DVSS.n1778 539.294
R20165 DVSS.n2465 DVSS.n2450 539.294
R20166 DVSS.n2457 DVSS.n2450 539.294
R20167 DVSS.n2457 DVSS.n1767 539.294
R20168 DVSS.n2479 DVSS.n1767 539.294
R20169 DVSS.n2479 DVSS.n1766 539.294
R20170 DVSS.n2484 DVSS.n1766 539.294
R20171 DVSS.n2484 DVSS.n1762 539.294
R20172 DVSS.n2496 DVSS.n1762 539.294
R20173 DVSS.n2496 DVSS.n1761 539.294
R20174 DVSS.n2501 DVSS.n1761 539.294
R20175 DVSS.n2501 DVSS.n1755 539.294
R20176 DVSS.n2514 DVSS.n1755 539.294
R20177 DVSS.n2514 DVSS.n1756 539.294
R20178 DVSS.n1756 DVSS.n1749 539.294
R20179 DVSS.n2818 DVSS.n2817 539.294
R20180 DVSS.n2817 DVSS.n663 539.294
R20181 DVSS.n2813 DVSS.n663 539.294
R20182 DVSS.n2813 DVSS.n666 539.294
R20183 DVSS.n677 DVSS.n666 539.294
R20184 DVSS.n2806 DVSS.n677 539.294
R20185 DVSS.n2806 DVSS.n678 539.294
R20186 DVSS.n2802 DVSS.n678 539.294
R20187 DVSS.n2802 DVSS.n681 539.294
R20188 DVSS.n2796 DVSS.n681 539.294
R20189 DVSS.n2796 DVSS.n685 539.294
R20190 DVSS.n2791 DVSS.n685 539.294
R20191 DVSS.n2791 DVSS.n687 539.294
R20192 DVSS.n698 DVSS.n687 539.294
R20193 DVSS.n2781 DVSS.n698 539.294
R20194 DVSS.n2781 DVSS.n699 539.294
R20195 DVSS.n2777 DVSS.n699 539.294
R20196 DVSS.n2777 DVSS.n702 539.294
R20197 DVSS.n709 DVSS.n702 539.294
R20198 DVSS.n2769 DVSS.n2768 539.294
R20199 DVSS.n3084 DVSS.n7 539.294
R20200 DVSS.n3084 DVSS.n8 539.294
R20201 DVSS.n3080 DVSS.n8 539.294
R20202 DVSS.n3080 DVSS.n10 539.294
R20203 DVSS.n2914 DVSS.n2912 539.294
R20204 DVSS.n2918 DVSS.n2912 539.294
R20205 DVSS.n2922 DVSS.n2920 539.294
R20206 DVSS.n2931 DVSS.n2908 539.294
R20207 DVSS.n2935 DVSS.n2933 539.294
R20208 DVSS.n2944 DVSS.n2904 539.294
R20209 DVSS.n2948 DVSS.n2946 539.294
R20210 DVSS.n2958 DVSS.n2900 539.294
R20211 DVSS.n3006 DVSS.t166 538.777
R20212 DVSS.n375 DVSS.n371 535.801
R20213 DVSS.n2248 DVSS.n2244 535.801
R20214 DVSS.n1056 DVSS.n1052 535.801
R20215 DVSS.n1578 DVSS.n1574 535.801
R20216 DVSS.n2744 DVSS.n2743 534.384
R20217 DVSS.n2803 DVSS.n680 534.384
R20218 DVSS.n619 DVSS.n617 534.009
R20219 DVSS.n3082 DVSS.t9 522.87
R20220 DVSS.n2439 DVSS.n1782 522.126
R20221 DVSS.n2680 DVSS.n2679 522.126
R20222 DVSS.n336 DVSS.n314 518.471
R20223 DVSS.n350 DVSS.n263 518.471
R20224 DVSS.n358 DVSS.n255 518.471
R20225 DVSS.n404 DVSS.n228 518.471
R20226 DVSS.n2209 DVSS.n2187 518.471
R20227 DVSS.n2223 DVSS.n2136 518.471
R20228 DVSS.n2231 DVSS.n2128 518.471
R20229 DVSS.n2277 DVSS.n2101 518.471
R20230 DVSS.n1017 DVSS.n995 518.471
R20231 DVSS.n1031 DVSS.n944 518.471
R20232 DVSS.n1039 DVSS.n936 518.471
R20233 DVSS.n1085 DVSS.n909 518.471
R20234 DVSS.n1539 DVSS.n1517 518.471
R20235 DVSS.n1553 DVSS.n1466 518.471
R20236 DVSS.n1561 DVSS.n1458 518.471
R20237 DVSS.n1607 DVSS.n1431 518.471
R20238 DVSS.n3068 DVSS.t2 518.222
R20239 DVSS.n178 DVSS.n150 491.349
R20240 DVSS.n434 DVSS.n113 491.349
R20241 DVSS.n97 DVSS.n88 491.349
R20242 DVSS.n518 DVSS.n82 491.349
R20243 DVSS.n2051 DVSS.n2023 491.349
R20244 DVSS.n2307 DVSS.n1986 491.349
R20245 DVSS.n1970 DVSS.n1961 491.349
R20246 DVSS.n2391 DVSS.n1955 491.349
R20247 DVSS.n859 DVSS.n831 491.349
R20248 DVSS.n1115 DVSS.n794 491.349
R20249 DVSS.n778 DVSS.n769 491.349
R20250 DVSS.n1199 DVSS.n763 491.349
R20251 DVSS.n1381 DVSS.n1353 491.349
R20252 DVSS.n1637 DVSS.n1316 491.349
R20253 DVSS.n1300 DVSS.n1291 491.349
R20254 DVSS.n1721 DVSS.n1285 491.349
R20255 DVSS.n3007 DVSS.n619 489.507
R20256 DVSS.t160 DVSS.n660 484.055
R20257 DVSS.n2690 DVSS.t68 484.055
R20258 DVSS.n2845 DVSS.t124 481.634
R20259 DVSS.n1838 DVSS.t45 468.682
R20260 DVSS.n1850 DVSS.t47 454.69
R20261 DVSS.n2654 DVSS.t76 450.089
R20262 DVSS.t86 DVSS.n1889 450.089
R20263 DVSS.t37 DVSS.n715 450.089
R20264 DVSS.n2815 DVSS.t56 450.089
R20265 DVSS.n370 DVSS.n229 448.409
R20266 DVSS.n2243 DVSS.n2102 448.409
R20267 DVSS.n1051 DVSS.n910 448.409
R20268 DVSS.n1573 DVSS.n1432 448.409
R20269 DVSS.n1926 DVSS.n1925 443.233
R20270 DVSS.n3025 DVSS.n3024 443.233
R20271 DVSS.n2795 DVSS.n680 443.233
R20272 DVSS.n2792 DVSS.n686 443.233
R20273 DVSS.n2780 DVSS.n700 443.233
R20274 DVSS.n2743 DVSS.n2742 443.233
R20275 DVSS.n2732 DVSS.n2731 443.233
R20276 DVSS.n2730 DVSS.n741 443.233
R20277 DVSS.n2716 DVSS.n749 443.233
R20278 DVSS.t43 DVSS.n1862 432.654
R20279 DVSS.t9 DVSS.n3081 424.216
R20280 DVSS.t2 DVSS.n3067 420.445
R20281 DVSS.n2844 DVSS.t78 400
R20282 DVSS.n2793 DVSS.t24 397.062
R20283 DVSS.n2567 DVSS.t112 397.062
R20284 DVSS.t58 DVSS.t164 394.712
R20285 DVSS.n368 DVSS.n248 394
R20286 DVSS.n2241 DVSS.n2121 394
R20287 DVSS.n1049 DVSS.n929 394
R20288 DVSS.n1571 DVSS.n1451 394
R20289 DVSS.n2611 DVSS.n756 391.668
R20290 DVSS.t30 DVSS.t169 390.324
R20291 DVSS.t118 DVSS.n1806 388.007
R20292 DVSS.n42 DVSS.t134 388.007
R20293 DVSS.t78 DVSS.n2843 383.673
R20294 DVSS.t116 DVSS.n1924 378.594
R20295 DVSS.t128 DVSS.n3023 378.594
R20296 DVSS.t22 DVSS.n2779 378.594
R20297 DVSS.n2719 DVSS.t110 378.594
R20298 DVSS.n472 DVSS.n95 366.841
R20299 DVSS.n487 DVSS.n99 366.841
R20300 DVSS.n126 DVSS.n112 366.841
R20301 DVSS.n142 DVSS.n115 366.841
R20302 DVSS.n2345 DVSS.n1968 366.841
R20303 DVSS.n2360 DVSS.n1972 366.841
R20304 DVSS.n1999 DVSS.n1985 366.841
R20305 DVSS.n2015 DVSS.n1988 366.841
R20306 DVSS.n1153 DVSS.n776 366.841
R20307 DVSS.n1168 DVSS.n780 366.841
R20308 DVSS.n807 DVSS.n793 366.841
R20309 DVSS.n823 DVSS.n796 366.841
R20310 DVSS.n1675 DVSS.n1298 366.841
R20311 DVSS.n1690 DVSS.n1302 366.841
R20312 DVSS.n1329 DVSS.n1315 366.841
R20313 DVSS.n1345 DVSS.n1318 366.841
R20314 DVSS.n2857 DVSS.n2856 357.685
R20315 DVSS.t43 DVSS.n632 351.021
R20316 DVSS.n1751 DVSS.n701 350.892
R20317 DVSS.t164 DVSS.n2873 349.909
R20318 DVSS.n2767 DVSS.n2766 343.353
R20319 DVSS.n1924 DVSS.t126 341.659
R20320 DVSS.n3023 DVSS.t132 341.659
R20321 DVSS.n2779 DVSS.t20 341.659
R20322 DVSS.n2719 DVSS.t106 341.659
R20323 DVSS.n1752 DVSS.n1751 332.425
R20324 DVSS.n344 DVSS.n314 317.623
R20325 DVSS.n350 DVSS.n262 317.623
R20326 DVSS.n358 DVSS.n256 317.623
R20327 DVSS.n364 DVSS.n228 317.623
R20328 DVSS.n2217 DVSS.n2187 317.623
R20329 DVSS.n2223 DVSS.n2135 317.623
R20330 DVSS.n2231 DVSS.n2129 317.623
R20331 DVSS.n2237 DVSS.n2101 317.623
R20332 DVSS.n1025 DVSS.n995 317.623
R20333 DVSS.n1031 DVSS.n943 317.623
R20334 DVSS.n1039 DVSS.n937 317.623
R20335 DVSS.n1045 DVSS.n909 317.623
R20336 DVSS.n1547 DVSS.n1517 317.623
R20337 DVSS.n1553 DVSS.n1465 317.623
R20338 DVSS.n1561 DVSS.n1459 317.623
R20339 DVSS.n1567 DVSS.n1431 317.623
R20340 DVSS.n447 DVSS.n115 306.26
R20341 DVSS.n495 DVSS.n99 306.26
R20342 DVSS.n449 DVSS.n112 306.26
R20343 DVSS.n497 DVSS.n95 306.26
R20344 DVSS.n2320 DVSS.n1988 306.26
R20345 DVSS.n2368 DVSS.n1972 306.26
R20346 DVSS.n2322 DVSS.n1985 306.26
R20347 DVSS.n2370 DVSS.n1968 306.26
R20348 DVSS.n1128 DVSS.n796 306.26
R20349 DVSS.n1176 DVSS.n780 306.26
R20350 DVSS.n1130 DVSS.n793 306.26
R20351 DVSS.n1178 DVSS.n776 306.26
R20352 DVSS.n1650 DVSS.n1318 306.26
R20353 DVSS.n1698 DVSS.n1302 306.26
R20354 DVSS.n1652 DVSS.n1315 306.26
R20355 DVSS.n1700 DVSS.n1298 306.26
R20356 DVSS.t124 DVSS.n2844 302.041
R20357 DVSS.n428 DVSS.n150 301.007
R20358 DVSS.n434 DVSS.n146 301.007
R20359 DVSS.n448 DVSS.n114 301.007
R20360 DVSS.n455 DVSS.n108 301.007
R20361 DVSS.n496 DVSS.n96 301.007
R20362 DVSS.n526 DVSS.n88 301.007
R20363 DVSS.n90 DVSS.n82 301.007
R20364 DVSS.n2301 DVSS.n2023 301.007
R20365 DVSS.n2307 DVSS.n2019 301.007
R20366 DVSS.n2321 DVSS.n1987 301.007
R20367 DVSS.n2328 DVSS.n1981 301.007
R20368 DVSS.n2369 DVSS.n1969 301.007
R20369 DVSS.n2399 DVSS.n1961 301.007
R20370 DVSS.n1963 DVSS.n1955 301.007
R20371 DVSS.n1109 DVSS.n831 301.007
R20372 DVSS.n1115 DVSS.n827 301.007
R20373 DVSS.n1129 DVSS.n795 301.007
R20374 DVSS.n1136 DVSS.n789 301.007
R20375 DVSS.n1177 DVSS.n777 301.007
R20376 DVSS.n1207 DVSS.n769 301.007
R20377 DVSS.n771 DVSS.n763 301.007
R20378 DVSS.n1631 DVSS.n1353 301.007
R20379 DVSS.n1637 DVSS.n1349 301.007
R20380 DVSS.n1651 DVSS.n1317 301.007
R20381 DVSS.n1658 DVSS.n1311 301.007
R20382 DVSS.n1699 DVSS.n1299 301.007
R20383 DVSS.n1729 DVSS.n1291 301.007
R20384 DVSS.n1293 DVSS.n1285 301.007
R20385 DVSS.t76 DVSS.n2653 294.885
R20386 DVSS.n1890 DVSS.t86 294.885
R20387 DVSS.n726 DVSS.t37 294.885
R20388 DVSS.t56 DVSS.n2814 294.885
R20389 DVSS.n351 DVSS.n258 292.5
R20390 DVSS.n351 DVSS.n350 292.5
R20391 DVSS.n367 DVSS.n366 292.5
R20392 DVSS.n366 DVSS.n228 292.5
R20393 DVSS.n334 DVSS.n333 292.5
R20394 DVSS.n332 DVSS.n321 292.5
R20395 DVSS.n331 DVSS.n330 292.5
R20396 DVSS.n329 DVSS.n328 292.5
R20397 DVSS.n327 DVSS.n326 292.5
R20398 DVSS.n325 DVSS.n324 292.5
R20399 DVSS.n323 DVSS.n322 292.5
R20400 DVSS.n317 DVSS.n316 292.5
R20401 DVSS.n365 DVSS.n250 292.5
R20402 DVSS.n365 DVSS.n364 292.5
R20403 DVSS.n355 DVSS.n251 292.5
R20404 DVSS.n256 DVSS.n251 292.5
R20405 DVSS.n343 DVSS.n342 292.5
R20406 DVSS.n344 DVSS.n343 292.5
R20407 DVSS.n341 DVSS.n261 292.5
R20408 DVSS.n262 DVSS.n261 292.5
R20409 DVSS.n357 DVSS.n356 292.5
R20410 DVSS.n358 DVSS.n357 292.5
R20411 DVSS.n339 DVSS.n338 292.5
R20412 DVSS.n340 DVSS.n315 292.5
R20413 DVSS.n315 DVSS.n314 292.5
R20414 DVSS.n378 DVSS.n368 292.5
R20415 DVSS.n371 DVSS.n368 292.5
R20416 DVSS.n379 DVSS.n248 292.5
R20417 DVSS.n370 DVSS.n248 292.5
R20418 DVSS.n377 DVSS.n376 292.5
R20419 DVSS.n374 DVSS.n369 292.5
R20420 DVSS.n385 DVSS.n384 292.5
R20421 DVSS.n387 DVSS.n386 292.5
R20422 DVSS.n249 DVSS.n230 292.5
R20423 DVSS.n404 DVSS.n230 292.5
R20424 DVSS.n382 DVSS.n381 292.5
R20425 DVSS.n373 DVSS.n371 292.5
R20426 DVSS.n370 DVSS.n247 292.5
R20427 DVSS.n245 DVSS.n244 292.5
R20428 DVSS.n393 DVSS.n392 292.5
R20429 DVSS.n396 DVSS.n395 292.5
R20430 DVSS.n239 DVSS.n238 292.5
R20431 DVSS.n402 DVSS.n401 292.5
R20432 DVSS.n236 DVSS.n227 292.5
R20433 DVSS.n407 DVSS.n406 292.5
R20434 DVSS.n226 DVSS.n224 292.5
R20435 DVSS.n228 DVSS.n226 292.5
R20436 DVSS.n363 DVSS.n362 292.5
R20437 DVSS.n364 DVSS.n363 292.5
R20438 DVSS.n361 DVSS.n252 292.5
R20439 DVSS.n256 DVSS.n252 292.5
R20440 DVSS.n360 DVSS.n359 292.5
R20441 DVSS.n359 DVSS.n358 292.5
R20442 DVSS.n313 DVSS.n312 292.5
R20443 DVSS.n314 DVSS.n313 292.5
R20444 DVSS.n346 DVSS.n345 292.5
R20445 DVSS.n345 DVSS.n344 292.5
R20446 DVSS.n347 DVSS.n264 292.5
R20447 DVSS.n264 DVSS.n262 292.5
R20448 DVSS.n349 DVSS.n348 292.5
R20449 DVSS.n350 DVSS.n349 292.5
R20450 DVSS.n353 DVSS.n257 292.5
R20451 DVSS.n311 DVSS.n310 292.5
R20452 DVSS.n310 DVSS.n254 292.5
R20453 DVSS.n269 DVSS.n267 292.5
R20454 DVSS.n274 DVSS.n267 292.5
R20455 DVSS.n305 DVSS.n271 292.5
R20456 DVSS.n305 DVSS.n304 292.5
R20457 DVSS.n279 DVSS.n276 292.5
R20458 DVSS.n303 DVSS.n276 292.5
R20459 DVSS.n300 DVSS.n281 292.5
R20460 DVSS.n301 DVSS.n300 292.5
R20461 DVSS.n286 DVSS.n282 292.5
R20462 DVSS.n282 DVSS.n277 292.5
R20463 DVSS.n295 DVSS.n288 292.5
R20464 DVSS.n295 DVSS.n294 292.5
R20465 DVSS.n293 DVSS.n291 292.5
R20466 DVSS.n291 DVSS.n290 292.5
R20467 DVSS.n353 DVSS.n352 292.5
R20468 DVSS.n165 DVSS.n164 292.5
R20469 DVSS.n156 DVSS.n155 292.5
R20470 DVSS.n168 DVSS.n167 292.5
R20471 DVSS.n170 DVSS.n169 292.5
R20472 DVSS.n172 DVSS.n171 292.5
R20473 DVSS.n174 DVSS.n173 292.5
R20474 DVSS.n176 DVSS.n175 292.5
R20475 DVSS.n166 DVSS.n163 292.5
R20476 DVSS.n180 DVSS.n179 292.5
R20477 DVSS.n179 DVSS.n178 292.5
R20478 DVSS.n472 DVSS.n92 292.5
R20479 DVSS.n472 DVSS.n97 292.5
R20480 DVSS.n485 DVSS.n468 292.5
R20481 DVSS.n484 DVSS.n483 292.5
R20482 DVSS.n482 DVSS.n481 292.5
R20483 DVSS.n480 DVSS.n470 292.5
R20484 DVSS.n478 DVSS.n477 292.5
R20485 DVSS.n476 DVSS.n471 292.5
R20486 DVSS.n475 DVSS.n474 292.5
R20487 DVSS.n488 DVSS.n487 292.5
R20488 DVSS.n128 DVSS.n124 292.5
R20489 DVSS.n141 DVSS.n120 292.5
R20490 DVSS.n139 DVSS.n138 292.5
R20491 DVSS.n137 DVSS.n136 292.5
R20492 DVSS.n134 DVSS.n122 292.5
R20493 DVSS.n132 DVSS.n131 292.5
R20494 DVSS.n130 DVSS.n129 292.5
R20495 DVSS.n143 DVSS.n142 292.5
R20496 DVSS.n142 DVSS.n113 292.5
R20497 DVSS.n126 DVSS.n125 292.5
R20498 DVSS.n522 DVSS.n521 292.5
R20499 DVSS.n521 DVSS.n82 292.5
R20500 DVSS.n523 DVSS.n91 292.5
R20501 DVSS.n91 DVSS.n90 292.5
R20502 DVSS.n525 DVSS.n524 292.5
R20503 DVSS.n526 DVSS.n525 292.5
R20504 DVSS.n500 DVSS.n89 292.5
R20505 DVSS.n89 DVSS.n88 292.5
R20506 DVSS.n498 DVSS.n497 292.5
R20507 DVSS.n497 DVSS.n496 292.5
R20508 DVSS.n94 DVSS.n93 292.5
R20509 DVSS.n96 DVSS.n94 292.5
R20510 DVSS.n452 DVSS.n110 292.5
R20511 DVSS.n110 DVSS.n108 292.5
R20512 DVSS.n454 DVSS.n453 292.5
R20513 DVSS.n455 DVSS.n454 292.5
R20514 DVSS.n451 DVSS.n109 292.5
R20515 DVSS.n114 DVSS.n109 292.5
R20516 DVSS.n450 DVSS.n449 292.5
R20517 DVSS.n449 DVSS.n448 292.5
R20518 DVSS.n433 DVSS.n432 292.5
R20519 DVSS.n434 DVSS.n433 292.5
R20520 DVSS.n431 DVSS.n147 292.5
R20521 DVSS.n147 DVSS.n146 292.5
R20522 DVSS.n430 DVSS.n429 292.5
R20523 DVSS.n429 DVSS.n428 292.5
R20524 DVSS.n149 DVSS.n148 292.5
R20525 DVSS.n150 DVSS.n149 292.5
R20526 DVSS.n520 DVSS.n501 292.5
R20527 DVSS.n506 DVSS.n502 292.5
R20528 DVSS.n516 DVSS.n515 292.5
R20529 DVSS.n514 DVSS.n505 292.5
R20530 DVSS.n513 DVSS.n512 292.5
R20531 DVSS.n511 DVSS.n510 292.5
R20532 DVSS.n509 DVSS.n508 292.5
R20533 DVSS.n507 DVSS.n79 292.5
R20534 DVSS.n537 DVSS.n536 292.5
R20535 DVSS.n2224 DVSS.n2131 292.5
R20536 DVSS.n2224 DVSS.n2223 292.5
R20537 DVSS.n2240 DVSS.n2239 292.5
R20538 DVSS.n2239 DVSS.n2101 292.5
R20539 DVSS.n2207 DVSS.n2206 292.5
R20540 DVSS.n2205 DVSS.n2194 292.5
R20541 DVSS.n2204 DVSS.n2203 292.5
R20542 DVSS.n2202 DVSS.n2201 292.5
R20543 DVSS.n2200 DVSS.n2199 292.5
R20544 DVSS.n2198 DVSS.n2197 292.5
R20545 DVSS.n2196 DVSS.n2195 292.5
R20546 DVSS.n2190 DVSS.n2189 292.5
R20547 DVSS.n2238 DVSS.n2123 292.5
R20548 DVSS.n2238 DVSS.n2237 292.5
R20549 DVSS.n2228 DVSS.n2124 292.5
R20550 DVSS.n2129 DVSS.n2124 292.5
R20551 DVSS.n2216 DVSS.n2215 292.5
R20552 DVSS.n2217 DVSS.n2216 292.5
R20553 DVSS.n2214 DVSS.n2134 292.5
R20554 DVSS.n2135 DVSS.n2134 292.5
R20555 DVSS.n2230 DVSS.n2229 292.5
R20556 DVSS.n2231 DVSS.n2230 292.5
R20557 DVSS.n2212 DVSS.n2211 292.5
R20558 DVSS.n2213 DVSS.n2188 292.5
R20559 DVSS.n2188 DVSS.n2187 292.5
R20560 DVSS.n2251 DVSS.n2241 292.5
R20561 DVSS.n2244 DVSS.n2241 292.5
R20562 DVSS.n2252 DVSS.n2121 292.5
R20563 DVSS.n2243 DVSS.n2121 292.5
R20564 DVSS.n2250 DVSS.n2249 292.5
R20565 DVSS.n2247 DVSS.n2242 292.5
R20566 DVSS.n2258 DVSS.n2257 292.5
R20567 DVSS.n2260 DVSS.n2259 292.5
R20568 DVSS.n2122 DVSS.n2103 292.5
R20569 DVSS.n2277 DVSS.n2103 292.5
R20570 DVSS.n2255 DVSS.n2254 292.5
R20571 DVSS.n2246 DVSS.n2244 292.5
R20572 DVSS.n2243 DVSS.n2120 292.5
R20573 DVSS.n2118 DVSS.n2117 292.5
R20574 DVSS.n2266 DVSS.n2265 292.5
R20575 DVSS.n2269 DVSS.n2268 292.5
R20576 DVSS.n2112 DVSS.n2111 292.5
R20577 DVSS.n2275 DVSS.n2274 292.5
R20578 DVSS.n2109 DVSS.n2100 292.5
R20579 DVSS.n2280 DVSS.n2279 292.5
R20580 DVSS.n2099 DVSS.n2097 292.5
R20581 DVSS.n2101 DVSS.n2099 292.5
R20582 DVSS.n2236 DVSS.n2235 292.5
R20583 DVSS.n2237 DVSS.n2236 292.5
R20584 DVSS.n2234 DVSS.n2125 292.5
R20585 DVSS.n2129 DVSS.n2125 292.5
R20586 DVSS.n2233 DVSS.n2232 292.5
R20587 DVSS.n2232 DVSS.n2231 292.5
R20588 DVSS.n2186 DVSS.n2185 292.5
R20589 DVSS.n2187 DVSS.n2186 292.5
R20590 DVSS.n2219 DVSS.n2218 292.5
R20591 DVSS.n2218 DVSS.n2217 292.5
R20592 DVSS.n2220 DVSS.n2137 292.5
R20593 DVSS.n2137 DVSS.n2135 292.5
R20594 DVSS.n2222 DVSS.n2221 292.5
R20595 DVSS.n2223 DVSS.n2222 292.5
R20596 DVSS.n2226 DVSS.n2130 292.5
R20597 DVSS.n2184 DVSS.n2183 292.5
R20598 DVSS.n2183 DVSS.n2127 292.5
R20599 DVSS.n2142 DVSS.n2140 292.5
R20600 DVSS.n2147 DVSS.n2140 292.5
R20601 DVSS.n2178 DVSS.n2144 292.5
R20602 DVSS.n2178 DVSS.n2177 292.5
R20603 DVSS.n2152 DVSS.n2149 292.5
R20604 DVSS.n2176 DVSS.n2149 292.5
R20605 DVSS.n2173 DVSS.n2154 292.5
R20606 DVSS.n2174 DVSS.n2173 292.5
R20607 DVSS.n2159 DVSS.n2155 292.5
R20608 DVSS.n2155 DVSS.n2150 292.5
R20609 DVSS.n2168 DVSS.n2161 292.5
R20610 DVSS.n2168 DVSS.n2167 292.5
R20611 DVSS.n2166 DVSS.n2164 292.5
R20612 DVSS.n2164 DVSS.n2163 292.5
R20613 DVSS.n2226 DVSS.n2225 292.5
R20614 DVSS.n2038 DVSS.n2037 292.5
R20615 DVSS.n2029 DVSS.n2028 292.5
R20616 DVSS.n2041 DVSS.n2040 292.5
R20617 DVSS.n2043 DVSS.n2042 292.5
R20618 DVSS.n2045 DVSS.n2044 292.5
R20619 DVSS.n2047 DVSS.n2046 292.5
R20620 DVSS.n2049 DVSS.n2048 292.5
R20621 DVSS.n2039 DVSS.n2036 292.5
R20622 DVSS.n2053 DVSS.n2052 292.5
R20623 DVSS.n2052 DVSS.n2051 292.5
R20624 DVSS.n2345 DVSS.n1965 292.5
R20625 DVSS.n2345 DVSS.n1970 292.5
R20626 DVSS.n2358 DVSS.n2341 292.5
R20627 DVSS.n2357 DVSS.n2356 292.5
R20628 DVSS.n2355 DVSS.n2354 292.5
R20629 DVSS.n2353 DVSS.n2343 292.5
R20630 DVSS.n2351 DVSS.n2350 292.5
R20631 DVSS.n2349 DVSS.n2344 292.5
R20632 DVSS.n2348 DVSS.n2347 292.5
R20633 DVSS.n2361 DVSS.n2360 292.5
R20634 DVSS.n2001 DVSS.n1997 292.5
R20635 DVSS.n2014 DVSS.n1993 292.5
R20636 DVSS.n2012 DVSS.n2011 292.5
R20637 DVSS.n2010 DVSS.n2009 292.5
R20638 DVSS.n2007 DVSS.n1995 292.5
R20639 DVSS.n2005 DVSS.n2004 292.5
R20640 DVSS.n2003 DVSS.n2002 292.5
R20641 DVSS.n2016 DVSS.n2015 292.5
R20642 DVSS.n2015 DVSS.n1986 292.5
R20643 DVSS.n1999 DVSS.n1998 292.5
R20644 DVSS.n2395 DVSS.n2394 292.5
R20645 DVSS.n2394 DVSS.n1955 292.5
R20646 DVSS.n2396 DVSS.n1964 292.5
R20647 DVSS.n1964 DVSS.n1963 292.5
R20648 DVSS.n2398 DVSS.n2397 292.5
R20649 DVSS.n2399 DVSS.n2398 292.5
R20650 DVSS.n2373 DVSS.n1962 292.5
R20651 DVSS.n1962 DVSS.n1961 292.5
R20652 DVSS.n2371 DVSS.n2370 292.5
R20653 DVSS.n2370 DVSS.n2369 292.5
R20654 DVSS.n1967 DVSS.n1966 292.5
R20655 DVSS.n1969 DVSS.n1967 292.5
R20656 DVSS.n2325 DVSS.n1983 292.5
R20657 DVSS.n1983 DVSS.n1981 292.5
R20658 DVSS.n2327 DVSS.n2326 292.5
R20659 DVSS.n2328 DVSS.n2327 292.5
R20660 DVSS.n2324 DVSS.n1982 292.5
R20661 DVSS.n1987 DVSS.n1982 292.5
R20662 DVSS.n2323 DVSS.n2322 292.5
R20663 DVSS.n2322 DVSS.n2321 292.5
R20664 DVSS.n2306 DVSS.n2305 292.5
R20665 DVSS.n2307 DVSS.n2306 292.5
R20666 DVSS.n2304 DVSS.n2020 292.5
R20667 DVSS.n2020 DVSS.n2019 292.5
R20668 DVSS.n2303 DVSS.n2302 292.5
R20669 DVSS.n2302 DVSS.n2301 292.5
R20670 DVSS.n2022 DVSS.n2021 292.5
R20671 DVSS.n2023 DVSS.n2022 292.5
R20672 DVSS.n2393 DVSS.n2374 292.5
R20673 DVSS.n2379 DVSS.n2375 292.5
R20674 DVSS.n2389 DVSS.n2388 292.5
R20675 DVSS.n2387 DVSS.n2378 292.5
R20676 DVSS.n2386 DVSS.n2385 292.5
R20677 DVSS.n2384 DVSS.n2383 292.5
R20678 DVSS.n2382 DVSS.n2381 292.5
R20679 DVSS.n2380 DVSS.n1952 292.5
R20680 DVSS.n2410 DVSS.n2409 292.5
R20681 DVSS.n1032 DVSS.n939 292.5
R20682 DVSS.n1032 DVSS.n1031 292.5
R20683 DVSS.n1048 DVSS.n1047 292.5
R20684 DVSS.n1047 DVSS.n909 292.5
R20685 DVSS.n1015 DVSS.n1014 292.5
R20686 DVSS.n1013 DVSS.n1002 292.5
R20687 DVSS.n1012 DVSS.n1011 292.5
R20688 DVSS.n1010 DVSS.n1009 292.5
R20689 DVSS.n1008 DVSS.n1007 292.5
R20690 DVSS.n1006 DVSS.n1005 292.5
R20691 DVSS.n1004 DVSS.n1003 292.5
R20692 DVSS.n998 DVSS.n997 292.5
R20693 DVSS.n1046 DVSS.n931 292.5
R20694 DVSS.n1046 DVSS.n1045 292.5
R20695 DVSS.n1036 DVSS.n932 292.5
R20696 DVSS.n937 DVSS.n932 292.5
R20697 DVSS.n1024 DVSS.n1023 292.5
R20698 DVSS.n1025 DVSS.n1024 292.5
R20699 DVSS.n1022 DVSS.n942 292.5
R20700 DVSS.n943 DVSS.n942 292.5
R20701 DVSS.n1038 DVSS.n1037 292.5
R20702 DVSS.n1039 DVSS.n1038 292.5
R20703 DVSS.n1020 DVSS.n1019 292.5
R20704 DVSS.n1021 DVSS.n996 292.5
R20705 DVSS.n996 DVSS.n995 292.5
R20706 DVSS.n1059 DVSS.n1049 292.5
R20707 DVSS.n1052 DVSS.n1049 292.5
R20708 DVSS.n1060 DVSS.n929 292.5
R20709 DVSS.n1051 DVSS.n929 292.5
R20710 DVSS.n1058 DVSS.n1057 292.5
R20711 DVSS.n1055 DVSS.n1050 292.5
R20712 DVSS.n1066 DVSS.n1065 292.5
R20713 DVSS.n1068 DVSS.n1067 292.5
R20714 DVSS.n930 DVSS.n911 292.5
R20715 DVSS.n1085 DVSS.n911 292.5
R20716 DVSS.n1063 DVSS.n1062 292.5
R20717 DVSS.n1054 DVSS.n1052 292.5
R20718 DVSS.n1051 DVSS.n928 292.5
R20719 DVSS.n926 DVSS.n925 292.5
R20720 DVSS.n1074 DVSS.n1073 292.5
R20721 DVSS.n1077 DVSS.n1076 292.5
R20722 DVSS.n920 DVSS.n919 292.5
R20723 DVSS.n1083 DVSS.n1082 292.5
R20724 DVSS.n917 DVSS.n908 292.5
R20725 DVSS.n1088 DVSS.n1087 292.5
R20726 DVSS.n907 DVSS.n905 292.5
R20727 DVSS.n909 DVSS.n907 292.5
R20728 DVSS.n1044 DVSS.n1043 292.5
R20729 DVSS.n1045 DVSS.n1044 292.5
R20730 DVSS.n1042 DVSS.n933 292.5
R20731 DVSS.n937 DVSS.n933 292.5
R20732 DVSS.n1041 DVSS.n1040 292.5
R20733 DVSS.n1040 DVSS.n1039 292.5
R20734 DVSS.n994 DVSS.n993 292.5
R20735 DVSS.n995 DVSS.n994 292.5
R20736 DVSS.n1027 DVSS.n1026 292.5
R20737 DVSS.n1026 DVSS.n1025 292.5
R20738 DVSS.n1028 DVSS.n945 292.5
R20739 DVSS.n945 DVSS.n943 292.5
R20740 DVSS.n1030 DVSS.n1029 292.5
R20741 DVSS.n1031 DVSS.n1030 292.5
R20742 DVSS.n1034 DVSS.n938 292.5
R20743 DVSS.n992 DVSS.n991 292.5
R20744 DVSS.n991 DVSS.n935 292.5
R20745 DVSS.n950 DVSS.n948 292.5
R20746 DVSS.n955 DVSS.n948 292.5
R20747 DVSS.n986 DVSS.n952 292.5
R20748 DVSS.n986 DVSS.n985 292.5
R20749 DVSS.n960 DVSS.n957 292.5
R20750 DVSS.n984 DVSS.n957 292.5
R20751 DVSS.n981 DVSS.n962 292.5
R20752 DVSS.n982 DVSS.n981 292.5
R20753 DVSS.n967 DVSS.n963 292.5
R20754 DVSS.n963 DVSS.n958 292.5
R20755 DVSS.n976 DVSS.n969 292.5
R20756 DVSS.n976 DVSS.n975 292.5
R20757 DVSS.n974 DVSS.n972 292.5
R20758 DVSS.n972 DVSS.n971 292.5
R20759 DVSS.n1034 DVSS.n1033 292.5
R20760 DVSS.n846 DVSS.n845 292.5
R20761 DVSS.n837 DVSS.n836 292.5
R20762 DVSS.n849 DVSS.n848 292.5
R20763 DVSS.n851 DVSS.n850 292.5
R20764 DVSS.n853 DVSS.n852 292.5
R20765 DVSS.n855 DVSS.n854 292.5
R20766 DVSS.n857 DVSS.n856 292.5
R20767 DVSS.n847 DVSS.n844 292.5
R20768 DVSS.n861 DVSS.n860 292.5
R20769 DVSS.n860 DVSS.n859 292.5
R20770 DVSS.n1153 DVSS.n773 292.5
R20771 DVSS.n1153 DVSS.n778 292.5
R20772 DVSS.n1166 DVSS.n1149 292.5
R20773 DVSS.n1165 DVSS.n1164 292.5
R20774 DVSS.n1163 DVSS.n1162 292.5
R20775 DVSS.n1161 DVSS.n1151 292.5
R20776 DVSS.n1159 DVSS.n1158 292.5
R20777 DVSS.n1157 DVSS.n1152 292.5
R20778 DVSS.n1156 DVSS.n1155 292.5
R20779 DVSS.n1169 DVSS.n1168 292.5
R20780 DVSS.n809 DVSS.n805 292.5
R20781 DVSS.n822 DVSS.n801 292.5
R20782 DVSS.n820 DVSS.n819 292.5
R20783 DVSS.n818 DVSS.n817 292.5
R20784 DVSS.n815 DVSS.n803 292.5
R20785 DVSS.n813 DVSS.n812 292.5
R20786 DVSS.n811 DVSS.n810 292.5
R20787 DVSS.n824 DVSS.n823 292.5
R20788 DVSS.n823 DVSS.n794 292.5
R20789 DVSS.n807 DVSS.n806 292.5
R20790 DVSS.n1203 DVSS.n1202 292.5
R20791 DVSS.n1202 DVSS.n763 292.5
R20792 DVSS.n1204 DVSS.n772 292.5
R20793 DVSS.n772 DVSS.n771 292.5
R20794 DVSS.n1206 DVSS.n1205 292.5
R20795 DVSS.n1207 DVSS.n1206 292.5
R20796 DVSS.n1181 DVSS.n770 292.5
R20797 DVSS.n770 DVSS.n769 292.5
R20798 DVSS.n1179 DVSS.n1178 292.5
R20799 DVSS.n1178 DVSS.n1177 292.5
R20800 DVSS.n775 DVSS.n774 292.5
R20801 DVSS.n777 DVSS.n775 292.5
R20802 DVSS.n1133 DVSS.n791 292.5
R20803 DVSS.n791 DVSS.n789 292.5
R20804 DVSS.n1135 DVSS.n1134 292.5
R20805 DVSS.n1136 DVSS.n1135 292.5
R20806 DVSS.n1132 DVSS.n790 292.5
R20807 DVSS.n795 DVSS.n790 292.5
R20808 DVSS.n1131 DVSS.n1130 292.5
R20809 DVSS.n1130 DVSS.n1129 292.5
R20810 DVSS.n1114 DVSS.n1113 292.5
R20811 DVSS.n1115 DVSS.n1114 292.5
R20812 DVSS.n1112 DVSS.n828 292.5
R20813 DVSS.n828 DVSS.n827 292.5
R20814 DVSS.n1111 DVSS.n1110 292.5
R20815 DVSS.n1110 DVSS.n1109 292.5
R20816 DVSS.n830 DVSS.n829 292.5
R20817 DVSS.n831 DVSS.n830 292.5
R20818 DVSS.n1201 DVSS.n1182 292.5
R20819 DVSS.n1187 DVSS.n1183 292.5
R20820 DVSS.n1197 DVSS.n1196 292.5
R20821 DVSS.n1195 DVSS.n1186 292.5
R20822 DVSS.n1194 DVSS.n1193 292.5
R20823 DVSS.n1192 DVSS.n1191 292.5
R20824 DVSS.n1190 DVSS.n1189 292.5
R20825 DVSS.n1188 DVSS.n760 292.5
R20826 DVSS.n1218 DVSS.n1217 292.5
R20827 DVSS.n1554 DVSS.n1461 292.5
R20828 DVSS.n1554 DVSS.n1553 292.5
R20829 DVSS.n1570 DVSS.n1569 292.5
R20830 DVSS.n1569 DVSS.n1431 292.5
R20831 DVSS.n1537 DVSS.n1536 292.5
R20832 DVSS.n1535 DVSS.n1524 292.5
R20833 DVSS.n1534 DVSS.n1533 292.5
R20834 DVSS.n1532 DVSS.n1531 292.5
R20835 DVSS.n1530 DVSS.n1529 292.5
R20836 DVSS.n1528 DVSS.n1527 292.5
R20837 DVSS.n1526 DVSS.n1525 292.5
R20838 DVSS.n1520 DVSS.n1519 292.5
R20839 DVSS.n1568 DVSS.n1453 292.5
R20840 DVSS.n1568 DVSS.n1567 292.5
R20841 DVSS.n1558 DVSS.n1454 292.5
R20842 DVSS.n1459 DVSS.n1454 292.5
R20843 DVSS.n1546 DVSS.n1545 292.5
R20844 DVSS.n1547 DVSS.n1546 292.5
R20845 DVSS.n1544 DVSS.n1464 292.5
R20846 DVSS.n1465 DVSS.n1464 292.5
R20847 DVSS.n1560 DVSS.n1559 292.5
R20848 DVSS.n1561 DVSS.n1560 292.5
R20849 DVSS.n1542 DVSS.n1541 292.5
R20850 DVSS.n1543 DVSS.n1518 292.5
R20851 DVSS.n1518 DVSS.n1517 292.5
R20852 DVSS.n1581 DVSS.n1571 292.5
R20853 DVSS.n1574 DVSS.n1571 292.5
R20854 DVSS.n1582 DVSS.n1451 292.5
R20855 DVSS.n1573 DVSS.n1451 292.5
R20856 DVSS.n1580 DVSS.n1579 292.5
R20857 DVSS.n1577 DVSS.n1572 292.5
R20858 DVSS.n1588 DVSS.n1587 292.5
R20859 DVSS.n1590 DVSS.n1589 292.5
R20860 DVSS.n1452 DVSS.n1433 292.5
R20861 DVSS.n1607 DVSS.n1433 292.5
R20862 DVSS.n1585 DVSS.n1584 292.5
R20863 DVSS.n1576 DVSS.n1574 292.5
R20864 DVSS.n1573 DVSS.n1450 292.5
R20865 DVSS.n1448 DVSS.n1447 292.5
R20866 DVSS.n1596 DVSS.n1595 292.5
R20867 DVSS.n1599 DVSS.n1598 292.5
R20868 DVSS.n1442 DVSS.n1441 292.5
R20869 DVSS.n1605 DVSS.n1604 292.5
R20870 DVSS.n1439 DVSS.n1430 292.5
R20871 DVSS.n1610 DVSS.n1609 292.5
R20872 DVSS.n1429 DVSS.n1427 292.5
R20873 DVSS.n1431 DVSS.n1429 292.5
R20874 DVSS.n1566 DVSS.n1565 292.5
R20875 DVSS.n1567 DVSS.n1566 292.5
R20876 DVSS.n1564 DVSS.n1455 292.5
R20877 DVSS.n1459 DVSS.n1455 292.5
R20878 DVSS.n1563 DVSS.n1562 292.5
R20879 DVSS.n1562 DVSS.n1561 292.5
R20880 DVSS.n1516 DVSS.n1515 292.5
R20881 DVSS.n1517 DVSS.n1516 292.5
R20882 DVSS.n1549 DVSS.n1548 292.5
R20883 DVSS.n1548 DVSS.n1547 292.5
R20884 DVSS.n1550 DVSS.n1467 292.5
R20885 DVSS.n1467 DVSS.n1465 292.5
R20886 DVSS.n1552 DVSS.n1551 292.5
R20887 DVSS.n1553 DVSS.n1552 292.5
R20888 DVSS.n1556 DVSS.n1460 292.5
R20889 DVSS.n1514 DVSS.n1513 292.5
R20890 DVSS.n1513 DVSS.n1457 292.5
R20891 DVSS.n1472 DVSS.n1470 292.5
R20892 DVSS.n1477 DVSS.n1470 292.5
R20893 DVSS.n1508 DVSS.n1474 292.5
R20894 DVSS.n1508 DVSS.n1507 292.5
R20895 DVSS.n1482 DVSS.n1479 292.5
R20896 DVSS.n1506 DVSS.n1479 292.5
R20897 DVSS.n1503 DVSS.n1484 292.5
R20898 DVSS.n1504 DVSS.n1503 292.5
R20899 DVSS.n1489 DVSS.n1485 292.5
R20900 DVSS.n1485 DVSS.n1480 292.5
R20901 DVSS.n1498 DVSS.n1491 292.5
R20902 DVSS.n1498 DVSS.n1497 292.5
R20903 DVSS.n1496 DVSS.n1494 292.5
R20904 DVSS.n1494 DVSS.n1493 292.5
R20905 DVSS.n1556 DVSS.n1555 292.5
R20906 DVSS.n1368 DVSS.n1367 292.5
R20907 DVSS.n1359 DVSS.n1358 292.5
R20908 DVSS.n1371 DVSS.n1370 292.5
R20909 DVSS.n1373 DVSS.n1372 292.5
R20910 DVSS.n1375 DVSS.n1374 292.5
R20911 DVSS.n1377 DVSS.n1376 292.5
R20912 DVSS.n1379 DVSS.n1378 292.5
R20913 DVSS.n1369 DVSS.n1366 292.5
R20914 DVSS.n1383 DVSS.n1382 292.5
R20915 DVSS.n1382 DVSS.n1381 292.5
R20916 DVSS.n1675 DVSS.n1295 292.5
R20917 DVSS.n1675 DVSS.n1300 292.5
R20918 DVSS.n1688 DVSS.n1671 292.5
R20919 DVSS.n1687 DVSS.n1686 292.5
R20920 DVSS.n1685 DVSS.n1684 292.5
R20921 DVSS.n1683 DVSS.n1673 292.5
R20922 DVSS.n1681 DVSS.n1680 292.5
R20923 DVSS.n1679 DVSS.n1674 292.5
R20924 DVSS.n1678 DVSS.n1677 292.5
R20925 DVSS.n1691 DVSS.n1690 292.5
R20926 DVSS.n1331 DVSS.n1327 292.5
R20927 DVSS.n1344 DVSS.n1323 292.5
R20928 DVSS.n1342 DVSS.n1341 292.5
R20929 DVSS.n1340 DVSS.n1339 292.5
R20930 DVSS.n1337 DVSS.n1325 292.5
R20931 DVSS.n1335 DVSS.n1334 292.5
R20932 DVSS.n1333 DVSS.n1332 292.5
R20933 DVSS.n1346 DVSS.n1345 292.5
R20934 DVSS.n1345 DVSS.n1316 292.5
R20935 DVSS.n1329 DVSS.n1328 292.5
R20936 DVSS.n1725 DVSS.n1724 292.5
R20937 DVSS.n1724 DVSS.n1285 292.5
R20938 DVSS.n1726 DVSS.n1294 292.5
R20939 DVSS.n1294 DVSS.n1293 292.5
R20940 DVSS.n1728 DVSS.n1727 292.5
R20941 DVSS.n1729 DVSS.n1728 292.5
R20942 DVSS.n1703 DVSS.n1292 292.5
R20943 DVSS.n1292 DVSS.n1291 292.5
R20944 DVSS.n1701 DVSS.n1700 292.5
R20945 DVSS.n1700 DVSS.n1699 292.5
R20946 DVSS.n1297 DVSS.n1296 292.5
R20947 DVSS.n1299 DVSS.n1297 292.5
R20948 DVSS.n1655 DVSS.n1313 292.5
R20949 DVSS.n1313 DVSS.n1311 292.5
R20950 DVSS.n1657 DVSS.n1656 292.5
R20951 DVSS.n1658 DVSS.n1657 292.5
R20952 DVSS.n1654 DVSS.n1312 292.5
R20953 DVSS.n1317 DVSS.n1312 292.5
R20954 DVSS.n1653 DVSS.n1652 292.5
R20955 DVSS.n1652 DVSS.n1651 292.5
R20956 DVSS.n1636 DVSS.n1635 292.5
R20957 DVSS.n1637 DVSS.n1636 292.5
R20958 DVSS.n1634 DVSS.n1350 292.5
R20959 DVSS.n1350 DVSS.n1349 292.5
R20960 DVSS.n1633 DVSS.n1632 292.5
R20961 DVSS.n1632 DVSS.n1631 292.5
R20962 DVSS.n1352 DVSS.n1351 292.5
R20963 DVSS.n1353 DVSS.n1352 292.5
R20964 DVSS.n1723 DVSS.n1704 292.5
R20965 DVSS.n1709 DVSS.n1705 292.5
R20966 DVSS.n1719 DVSS.n1718 292.5
R20967 DVSS.n1717 DVSS.n1708 292.5
R20968 DVSS.n1716 DVSS.n1715 292.5
R20969 DVSS.n1714 DVSS.n1713 292.5
R20970 DVSS.n1712 DVSS.n1711 292.5
R20971 DVSS.n1710 DVSS.n1282 292.5
R20972 DVSS.n1740 DVSS.n1739 292.5
R20973 DVSS.n615 DVSS.n67 288.92
R20974 DVSS.n2428 DVSS.t162 288.257
R20975 DVSS.t66 DVSS.n21 288.257
R20976 DVSS.n2531 DVSS.n2530 284.829
R20977 DVSS.n2533 DVSS.n2531 284.829
R20978 DVSS.n2533 DVSS.n2532 284.829
R20979 DVSS.n2545 DVSS.n1261 284.829
R20980 DVSS.n602 DVSS.n67 284.712
R20981 DVSS.n2449 DVSS.n2448 284.637
R20982 DVSS.n2467 DVSS.n2466 284.637
R20983 DVSS.n2456 DVSS.n2455 284.637
R20984 DVSS.n2481 DVSS.n2480 284.637
R20985 DVSS.n2483 DVSS.n2481 284.637
R20986 DVSS.n2483 DVSS.n2482 284.637
R20987 DVSS.n2500 DVSS.n2498 284.637
R20988 DVSS.n2500 DVSS.n2499 284.637
R20989 DVSS.n3052 DVSS.n23 283.872
R20990 DVSS.n3041 DVSS.n3040 283.872
R20991 DVSS.n39 DVSS.n38 283.872
R20992 DVSS.n577 DVSS.n40 283.872
R20993 DVSS.n578 DVSS.n577 283.872
R20994 DVSS.n580 DVSS.n578 283.872
R20995 DVSS.n597 DVSS.n596 283.872
R20996 DVSS.n598 DVSS.n597 283.872
R20997 DVSS.n602 DVSS.n601 283.872
R20998 DVSS.n2546 DVSS.n2545 280.329
R20999 DVSS.n2547 DVSS.n2546 279.921
R21000 DVSS.n2565 DVSS.n1251 279.921
R21001 DVSS.n2569 DVSS.n1249 279.921
R21002 DVSS.n2579 DVSS.n1241 279.921
R21003 DVSS.n2580 DVSS.n2579 279.921
R21004 DVSS.n2582 DVSS.n2580 279.921
R21005 DVSS.n2596 DVSS.n2595 279.921
R21006 DVSS.n2598 DVSS.n2596 279.921
R21007 DVSS.n2608 DVSS.n1229 279.921
R21008 DVSS.n3005 DVSS.n2884 278.344
R21009 DVSS.n2960 DVSS.n2959 278.344
R21010 DVSS.n2794 DVSS.n2793 272.404
R21011 DVSS.n2568 DVSS.n2567 272.404
R21012 DVSS.n435 DVSS.n115 270.034
R21013 DVSS.n95 DVSS.n89 270.034
R21014 DVSS.n99 DVSS.n87 270.034
R21015 DVSS.n433 DVSS.n112 270.034
R21016 DVSS.n2308 DVSS.n1988 270.034
R21017 DVSS.n1968 DVSS.n1962 270.034
R21018 DVSS.n1972 DVSS.n1960 270.034
R21019 DVSS.n2306 DVSS.n1985 270.034
R21020 DVSS.n1116 DVSS.n796 270.034
R21021 DVSS.n776 DVSS.n770 270.034
R21022 DVSS.n780 DVSS.n768 270.034
R21023 DVSS.n1114 DVSS.n793 270.034
R21024 DVSS.n1638 DVSS.n1318 270.034
R21025 DVSS.n1298 DVSS.n1292 270.034
R21026 DVSS.n1302 DVSS.n1290 270.034
R21027 DVSS.n1636 DVSS.n1315 270.034
R21028 DVSS.n2427 DVSS.n2426 261.063
R21029 DVSS.n2428 DVSS.n2427 261.063
R21030 DVSS.n3054 DVSS.n20 261.063
R21031 DVSS.n3054 DVSS.n21 261.063
R21032 DVSS.n2448 DVSS.n1779 260.916
R21033 DVSS.n3053 DVSS.n3052 260.216
R21034 DVSS.n2468 DVSS.t102 254.385
R21035 DVSS.n36 DVSS.t154 253.739
R21036 DVSS.t47 DVSS.n1849 253.061
R21037 DVSS.t187 DVSS.n1252 250.407
R21038 DVSS.n2530 DVSS.n1271 249.226
R21039 DVSS.t96 DVSS.n2454 248.793
R21040 DVSS.n121 DVSS.n113 248.683
R21041 DVSS.n135 DVSS.n113 248.683
R21042 DVSS.n133 DVSS.n113 248.683
R21043 DVSS.n1994 DVSS.n1986 248.683
R21044 DVSS.n2008 DVSS.n1986 248.683
R21045 DVSS.n2006 DVSS.n1986 248.683
R21046 DVSS.n802 DVSS.n794 248.683
R21047 DVSS.n816 DVSS.n794 248.683
R21048 DVSS.n814 DVSS.n794 248.683
R21049 DVSS.n1324 DVSS.n1316 248.683
R21050 DVSS.n1338 DVSS.n1316 248.683
R21051 DVSS.n1336 DVSS.n1316 248.683
R21052 DVSS.n3039 DVSS.t146 248.163
R21053 DVSS.n404 DVSS.n232 245.512
R21054 DVSS.n404 DVSS.n233 245.512
R21055 DVSS.n404 DVSS.n234 245.512
R21056 DVSS.n404 DVSS.n235 245.512
R21057 DVSS.n404 DVSS.n403 245.512
R21058 DVSS.n178 DVSS.n159 245.512
R21059 DVSS.n178 DVSS.n160 245.512
R21060 DVSS.n178 DVSS.n161 245.512
R21061 DVSS.n178 DVSS.n162 245.512
R21062 DVSS.n178 DVSS.n177 245.512
R21063 DVSS.n2277 DVSS.n2105 245.512
R21064 DVSS.n2277 DVSS.n2106 245.512
R21065 DVSS.n2277 DVSS.n2107 245.512
R21066 DVSS.n2277 DVSS.n2108 245.512
R21067 DVSS.n2277 DVSS.n2276 245.512
R21068 DVSS.n2051 DVSS.n2032 245.512
R21069 DVSS.n2051 DVSS.n2033 245.512
R21070 DVSS.n2051 DVSS.n2034 245.512
R21071 DVSS.n2051 DVSS.n2035 245.512
R21072 DVSS.n2051 DVSS.n2050 245.512
R21073 DVSS.n1085 DVSS.n913 245.512
R21074 DVSS.n1085 DVSS.n914 245.512
R21075 DVSS.n1085 DVSS.n915 245.512
R21076 DVSS.n1085 DVSS.n916 245.512
R21077 DVSS.n1085 DVSS.n1084 245.512
R21078 DVSS.n859 DVSS.n840 245.512
R21079 DVSS.n859 DVSS.n841 245.512
R21080 DVSS.n859 DVSS.n842 245.512
R21081 DVSS.n859 DVSS.n843 245.512
R21082 DVSS.n859 DVSS.n858 245.512
R21083 DVSS.n1607 DVSS.n1435 245.512
R21084 DVSS.n1607 DVSS.n1436 245.512
R21085 DVSS.n1607 DVSS.n1437 245.512
R21086 DVSS.n1607 DVSS.n1438 245.512
R21087 DVSS.n1607 DVSS.n1606 245.512
R21088 DVSS.n1381 DVSS.n1362 245.512
R21089 DVSS.n1381 DVSS.n1363 245.512
R21090 DVSS.n1381 DVSS.n1364 245.512
R21091 DVSS.n1381 DVSS.n1365 245.512
R21092 DVSS.n1381 DVSS.n1380 245.512
R21093 DVSS.t181 DVSS.n2566 244.905
R21094 DVSS.n2717 DVSS.n2716 240.084
R21095 DVSS.n1848 DVSS.t45 236.736
R21096 DVSS.n2867 DVSS.n624 235.19
R21097 DVSS.n2858 DVSS.n2857 235.19
R21098 DVSS.t162 DVSS.n1782 233.869
R21099 DVSS.n2680 DVSS.t66 233.869
R21100 DVSS.t18 DVSS.n686 230.851
R21101 DVSS.n2731 DVSS.t108 230.851
R21102 DVSS.n2515 DVSS.n1754 225.338
R21103 DVSS.n3007 DVSS.n618 224.732
R21104 DVSS.n304 DVSS.n303 223.931
R21105 DVSS.n301 DVSS.n277 223.931
R21106 DVSS.n294 DVSS.n293 223.931
R21107 DVSS.n359 DVSS.n252 223.931
R21108 DVSS.n363 DVSS.n252 223.931
R21109 DVSS.n363 DVSS.n226 223.931
R21110 DVSS.n386 DVSS.n230 223.931
R21111 DVSS.n357 DVSS.n251 223.931
R21112 DVSS.n365 DVSS.n251 223.931
R21113 DVSS.n366 DVSS.n365 223.931
R21114 DVSS.n330 DVSS.n329 223.931
R21115 DVSS.n326 DVSS.n325 223.931
R21116 DVSS.n322 DVSS.n317 223.931
R21117 DVSS.n345 DVSS.n313 223.931
R21118 DVSS.n345 DVSS.n264 223.931
R21119 DVSS.n349 DVSS.n264 223.931
R21120 DVSS.n279 DVSS.n271 223.931
R21121 DVSS.n286 DVSS.n281 223.931
R21122 DVSS.n290 DVSS.n288 223.931
R21123 DVSS.n343 DVSS.n315 223.931
R21124 DVSS.n343 DVSS.n261 223.931
R21125 DVSS.n351 DVSS.n261 223.931
R21126 DVSS.n427 DVSS.n151 223.931
R21127 DVSS.n427 DVSS.n145 223.931
R21128 DVSS.n435 DVSS.n145 223.931
R21129 DVSS.n179 DVSS.n156 223.931
R21130 DVSS.n525 DVSS.n89 223.931
R21131 DVSS.n525 DVSS.n91 223.931
R21132 DVSS.n521 DVSS.n91 223.931
R21133 DVSS.n516 DVSS.n505 223.931
R21134 DVSS.n512 DVSS.n511 223.931
R21135 DVSS.n508 DVSS.n507 223.931
R21136 DVSS.n527 DVSS.n87 223.931
R21137 DVSS.n527 DVSS.n81 223.931
R21138 DVSS.n535 DVSS.n81 223.931
R21139 DVSS.n447 DVSS.n106 223.931
R21140 DVSS.n456 DVSS.n106 223.931
R21141 DVSS.n456 DVSS.n107 223.931
R21142 DVSS.n107 DVSS.n98 223.931
R21143 DVSS.n495 DVSS.n98 223.931
R21144 DVSS.n449 DVSS.n109 223.931
R21145 DVSS.n454 DVSS.n109 223.931
R21146 DVSS.n454 DVSS.n110 223.931
R21147 DVSS.n110 DVSS.n94 223.931
R21148 DVSS.n497 DVSS.n94 223.931
R21149 DVSS.n429 DVSS.n149 223.931
R21150 DVSS.n429 DVSS.n147 223.931
R21151 DVSS.n433 DVSS.n147 223.931
R21152 DVSS.n2177 DVSS.n2176 223.931
R21153 DVSS.n2174 DVSS.n2150 223.931
R21154 DVSS.n2167 DVSS.n2166 223.931
R21155 DVSS.n2232 DVSS.n2125 223.931
R21156 DVSS.n2236 DVSS.n2125 223.931
R21157 DVSS.n2236 DVSS.n2099 223.931
R21158 DVSS.n2259 DVSS.n2103 223.931
R21159 DVSS.n2230 DVSS.n2124 223.931
R21160 DVSS.n2238 DVSS.n2124 223.931
R21161 DVSS.n2239 DVSS.n2238 223.931
R21162 DVSS.n2203 DVSS.n2202 223.931
R21163 DVSS.n2199 DVSS.n2198 223.931
R21164 DVSS.n2195 DVSS.n2190 223.931
R21165 DVSS.n2218 DVSS.n2186 223.931
R21166 DVSS.n2218 DVSS.n2137 223.931
R21167 DVSS.n2222 DVSS.n2137 223.931
R21168 DVSS.n2152 DVSS.n2144 223.931
R21169 DVSS.n2159 DVSS.n2154 223.931
R21170 DVSS.n2163 DVSS.n2161 223.931
R21171 DVSS.n2216 DVSS.n2188 223.931
R21172 DVSS.n2216 DVSS.n2134 223.931
R21173 DVSS.n2224 DVSS.n2134 223.931
R21174 DVSS.n2300 DVSS.n2024 223.931
R21175 DVSS.n2300 DVSS.n2018 223.931
R21176 DVSS.n2308 DVSS.n2018 223.931
R21177 DVSS.n2052 DVSS.n2029 223.931
R21178 DVSS.n2398 DVSS.n1962 223.931
R21179 DVSS.n2398 DVSS.n1964 223.931
R21180 DVSS.n2394 DVSS.n1964 223.931
R21181 DVSS.n2389 DVSS.n2378 223.931
R21182 DVSS.n2385 DVSS.n2384 223.931
R21183 DVSS.n2381 DVSS.n2380 223.931
R21184 DVSS.n2400 DVSS.n1960 223.931
R21185 DVSS.n2400 DVSS.n1954 223.931
R21186 DVSS.n2408 DVSS.n1954 223.931
R21187 DVSS.n2320 DVSS.n1979 223.931
R21188 DVSS.n2329 DVSS.n1979 223.931
R21189 DVSS.n2329 DVSS.n1980 223.931
R21190 DVSS.n1980 DVSS.n1971 223.931
R21191 DVSS.n2368 DVSS.n1971 223.931
R21192 DVSS.n2322 DVSS.n1982 223.931
R21193 DVSS.n2327 DVSS.n1982 223.931
R21194 DVSS.n2327 DVSS.n1983 223.931
R21195 DVSS.n1983 DVSS.n1967 223.931
R21196 DVSS.n2370 DVSS.n1967 223.931
R21197 DVSS.n2302 DVSS.n2022 223.931
R21198 DVSS.n2302 DVSS.n2020 223.931
R21199 DVSS.n2306 DVSS.n2020 223.931
R21200 DVSS.n985 DVSS.n984 223.931
R21201 DVSS.n982 DVSS.n958 223.931
R21202 DVSS.n975 DVSS.n974 223.931
R21203 DVSS.n1040 DVSS.n933 223.931
R21204 DVSS.n1044 DVSS.n933 223.931
R21205 DVSS.n1044 DVSS.n907 223.931
R21206 DVSS.n1067 DVSS.n911 223.931
R21207 DVSS.n1038 DVSS.n932 223.931
R21208 DVSS.n1046 DVSS.n932 223.931
R21209 DVSS.n1047 DVSS.n1046 223.931
R21210 DVSS.n1011 DVSS.n1010 223.931
R21211 DVSS.n1007 DVSS.n1006 223.931
R21212 DVSS.n1003 DVSS.n998 223.931
R21213 DVSS.n1026 DVSS.n994 223.931
R21214 DVSS.n1026 DVSS.n945 223.931
R21215 DVSS.n1030 DVSS.n945 223.931
R21216 DVSS.n960 DVSS.n952 223.931
R21217 DVSS.n967 DVSS.n962 223.931
R21218 DVSS.n971 DVSS.n969 223.931
R21219 DVSS.n1024 DVSS.n996 223.931
R21220 DVSS.n1024 DVSS.n942 223.931
R21221 DVSS.n1032 DVSS.n942 223.931
R21222 DVSS.n1108 DVSS.n832 223.931
R21223 DVSS.n1108 DVSS.n826 223.931
R21224 DVSS.n1116 DVSS.n826 223.931
R21225 DVSS.n860 DVSS.n837 223.931
R21226 DVSS.n1206 DVSS.n770 223.931
R21227 DVSS.n1206 DVSS.n772 223.931
R21228 DVSS.n1202 DVSS.n772 223.931
R21229 DVSS.n1197 DVSS.n1186 223.931
R21230 DVSS.n1193 DVSS.n1192 223.931
R21231 DVSS.n1189 DVSS.n1188 223.931
R21232 DVSS.n1208 DVSS.n768 223.931
R21233 DVSS.n1208 DVSS.n762 223.931
R21234 DVSS.n1216 DVSS.n762 223.931
R21235 DVSS.n1128 DVSS.n787 223.931
R21236 DVSS.n1137 DVSS.n787 223.931
R21237 DVSS.n1137 DVSS.n788 223.931
R21238 DVSS.n788 DVSS.n779 223.931
R21239 DVSS.n1176 DVSS.n779 223.931
R21240 DVSS.n1130 DVSS.n790 223.931
R21241 DVSS.n1135 DVSS.n790 223.931
R21242 DVSS.n1135 DVSS.n791 223.931
R21243 DVSS.n791 DVSS.n775 223.931
R21244 DVSS.n1178 DVSS.n775 223.931
R21245 DVSS.n1110 DVSS.n830 223.931
R21246 DVSS.n1110 DVSS.n828 223.931
R21247 DVSS.n1114 DVSS.n828 223.931
R21248 DVSS.n1507 DVSS.n1506 223.931
R21249 DVSS.n1504 DVSS.n1480 223.931
R21250 DVSS.n1497 DVSS.n1496 223.931
R21251 DVSS.n1562 DVSS.n1455 223.931
R21252 DVSS.n1566 DVSS.n1455 223.931
R21253 DVSS.n1566 DVSS.n1429 223.931
R21254 DVSS.n1589 DVSS.n1433 223.931
R21255 DVSS.n1560 DVSS.n1454 223.931
R21256 DVSS.n1568 DVSS.n1454 223.931
R21257 DVSS.n1569 DVSS.n1568 223.931
R21258 DVSS.n1533 DVSS.n1532 223.931
R21259 DVSS.n1529 DVSS.n1528 223.931
R21260 DVSS.n1525 DVSS.n1520 223.931
R21261 DVSS.n1548 DVSS.n1516 223.931
R21262 DVSS.n1548 DVSS.n1467 223.931
R21263 DVSS.n1552 DVSS.n1467 223.931
R21264 DVSS.n1482 DVSS.n1474 223.931
R21265 DVSS.n1489 DVSS.n1484 223.931
R21266 DVSS.n1493 DVSS.n1491 223.931
R21267 DVSS.n1546 DVSS.n1518 223.931
R21268 DVSS.n1546 DVSS.n1464 223.931
R21269 DVSS.n1554 DVSS.n1464 223.931
R21270 DVSS.n1630 DVSS.n1354 223.931
R21271 DVSS.n1630 DVSS.n1348 223.931
R21272 DVSS.n1638 DVSS.n1348 223.931
R21273 DVSS.n1382 DVSS.n1359 223.931
R21274 DVSS.n1728 DVSS.n1292 223.931
R21275 DVSS.n1728 DVSS.n1294 223.931
R21276 DVSS.n1724 DVSS.n1294 223.931
R21277 DVSS.n1719 DVSS.n1708 223.931
R21278 DVSS.n1715 DVSS.n1714 223.931
R21279 DVSS.n1711 DVSS.n1710 223.931
R21280 DVSS.n1730 DVSS.n1290 223.931
R21281 DVSS.n1730 DVSS.n1284 223.931
R21282 DVSS.n1738 DVSS.n1284 223.931
R21283 DVSS.n1650 DVSS.n1309 223.931
R21284 DVSS.n1659 DVSS.n1309 223.931
R21285 DVSS.n1659 DVSS.n1310 223.931
R21286 DVSS.n1310 DVSS.n1301 223.931
R21287 DVSS.n1698 DVSS.n1301 223.931
R21288 DVSS.n1652 DVSS.n1312 223.931
R21289 DVSS.n1657 DVSS.n1312 223.931
R21290 DVSS.n1657 DVSS.n1313 223.931
R21291 DVSS.n1313 DVSS.n1297 223.931
R21292 DVSS.n1700 DVSS.n1297 223.931
R21293 DVSS.n1632 DVSS.n1352 223.931
R21294 DVSS.n1632 DVSS.n1350 223.931
R21295 DVSS.n1636 DVSS.n1350 223.931
R21296 DVSS.n2868 DVSS.t70 218.041
R21297 DVSS.n2516 DVSS.n2515 213.477
R21298 DVSS.n598 DVSS.n55 212.904
R21299 DVSS.n1926 DVSS.t118 212.382
R21300 DVSS.n3024 DVSS.t134 212.382
R21301 DVSS.n700 DVSS.t18 212.382
R21302 DVSS.t108 DVSS.n2730 212.382
R21303 DVSS.n474 DVSS.n472 206.16
R21304 DVSS.n478 DVSS.n471 206.16
R21305 DVSS.n481 DVSS.n480 206.16
R21306 DVSS.n485 DVSS.n484 206.16
R21307 DVSS.n129 DVSS.n128 206.16
R21308 DVSS.n142 DVSS.n141 206.16
R21309 DVSS.n2347 DVSS.n2345 206.16
R21310 DVSS.n2351 DVSS.n2344 206.16
R21311 DVSS.n2354 DVSS.n2353 206.16
R21312 DVSS.n2358 DVSS.n2357 206.16
R21313 DVSS.n2002 DVSS.n2001 206.16
R21314 DVSS.n2015 DVSS.n2014 206.16
R21315 DVSS.n1155 DVSS.n1153 206.16
R21316 DVSS.n1159 DVSS.n1152 206.16
R21317 DVSS.n1162 DVSS.n1161 206.16
R21318 DVSS.n1166 DVSS.n1165 206.16
R21319 DVSS.n810 DVSS.n809 206.16
R21320 DVSS.n823 DVSS.n822 206.16
R21321 DVSS.n1677 DVSS.n1675 206.16
R21322 DVSS.n1681 DVSS.n1674 206.16
R21323 DVSS.n1684 DVSS.n1683 206.16
R21324 DVSS.n1688 DVSS.n1687 206.16
R21325 DVSS.n1332 DVSS.n1331 206.16
R21326 DVSS.n1345 DVSS.n1344 206.16
R21327 DVSS.n2718 DVSS.n2717 203.149
R21328 DVSS.t122 DVSS.n1915 201.764
R21329 DVSS.n2634 DVSS.t138 201.764
R21330 DVSS.n3006 DVSS.n2878 200.215
R21331 DVSS.n3006 DVSS.n2880 200.215
R21332 DVSS.n3006 DVSS.n2882 200.215
R21333 DVSS.n455 DVSS.t39 199.196
R21334 DVSS.n108 DVSS.t40 199.196
R21335 DVSS.n2328 DVSS.t63 199.196
R21336 DVSS.n1981 DVSS.t62 199.196
R21337 DVSS.n1136 DVSS.t172 199.196
R21338 DVSS.n789 DVSS.t173 199.196
R21339 DVSS.n1658 DVSS.t145 199.196
R21340 DVSS.n1311 DVSS.t144 199.196
R21341 DVSS.n2834 DVSS.n2833 195.918
R21342 DVSS.n2454 DVSS.t98 187.294
R21343 DVSS.t150 DVSS.n3039 186.82
R21344 DVSS.n218 DVSS.n205 185
R21345 DVSS.n220 DVSS.n219 185
R21346 DVSS.n197 DVSS.n184 185
R21347 DVSS.n199 DVSS.n198 185
R21348 DVSS.n2091 DVSS.n2078 185
R21349 DVSS.n2093 DVSS.n2092 185
R21350 DVSS.n2070 DVSS.n2057 185
R21351 DVSS.n2072 DVSS.n2071 185
R21352 DVSS.n899 DVSS.n886 185
R21353 DVSS.n901 DVSS.n900 185
R21354 DVSS.n878 DVSS.n865 185
R21355 DVSS.n880 DVSS.n879 185
R21356 DVSS.n1421 DVSS.n1408 185
R21357 DVSS.n1423 DVSS.n1422 185
R21358 DVSS.n1400 DVSS.n1387 185
R21359 DVSS.n1402 DVSS.n1401 185
R21360 DVSS.n2999 DVSS.n2882 184.572
R21361 DVSS.n2887 DVSS.n2880 184.572
R21362 DVSS.n2990 DVSS.n2878 184.572
R21363 DVSS.n2992 DVSS.n2878 184.572
R21364 DVSS.n2997 DVSS.n2880 184.572
R21365 DVSS.n3001 DVSS.n2882 184.572
R21366 DVSS.n2566 DVSS.t183 184.367
R21367 DVSS.n2468 DVSS.t100 181.703
R21368 DVSS.t152 DVSS.n36 181.244
R21369 DVSS.t185 DVSS.n1252 178.863
R21370 DVSS.n2482 DVSS.t28 174.934
R21371 DVSS.n580 DVSS.t136 174.463
R21372 DVSS.n2582 DVSS.t104 172.035
R21373 DVSS.n1917 DVSS.t126 170.724
R21374 DVSS.t132 DVSS.n3022 170.724
R21375 DVSS.n344 DVSS.t178 158.811
R21376 DVSS.t178 DVSS.n262 158.811
R21377 DVSS.n256 DVSS.t41 158.811
R21378 DVSS.n364 DVSS.t41 158.811
R21379 DVSS.t180 DVSS.n370 158.811
R21380 DVSS.n371 DVSS.t180 158.811
R21381 DVSS.n2217 DVSS.t11 158.811
R21382 DVSS.t11 DVSS.n2135 158.811
R21383 DVSS.n2129 DVSS.t64 158.811
R21384 DVSS.n2237 DVSS.t64 158.811
R21385 DVSS.t13 DVSS.n2243 158.811
R21386 DVSS.n2244 DVSS.t13 158.811
R21387 DVSS.n1025 DVSS.t53 158.811
R21388 DVSS.t53 DVSS.n943 158.811
R21389 DVSS.n937 DVSS.t174 158.811
R21390 DVSS.n1045 DVSS.t174 158.811
R21391 DVSS.t55 DVSS.n1051 158.811
R21392 DVSS.n1052 DVSS.t55 158.811
R21393 DVSS.n1547 DVSS.t6 158.811
R21394 DVSS.t6 DVSS.n1465 158.811
R21395 DVSS.n1459 DVSS.t142 158.811
R21396 DVSS.n1567 DVSS.t142 158.811
R21397 DVSS.t8 DVSS.n1573 158.811
R21398 DVSS.n1574 DVSS.t8 158.811
R21399 DVSS.n123 DVSS.n113 157.904
R21400 DVSS.n1996 DVSS.n1986 157.904
R21401 DVSS.n804 DVSS.n794 157.904
R21402 DVSS.n1326 DVSS.n1316 157.904
R21403 DVSS.n140 DVSS.n113 157.904
R21404 DVSS.n2013 DVSS.n1986 157.904
R21405 DVSS.n821 DVSS.n794 157.904
R21406 DVSS.n1343 DVSS.n1316 157.904
R21407 DVSS.n2455 DVSS.t94 157.143
R21408 DVSS.t148 DVSS.n39 156.72
R21409 DVSS.n405 DVSS.n404 155.356
R21410 DVSS.n2278 DVSS.n2277 155.356
R21411 DVSS.n1086 DVSS.n1085 155.356
R21412 DVSS.n1608 DVSS.n1607 155.356
R21413 DVSS.n336 DVSS.n335 155.356
R21414 DVSS.n336 DVSS.n320 155.356
R21415 DVSS.n404 DVSS.n231 155.356
R21416 DVSS.n265 DVSS.n263 155.356
R21417 DVSS.n273 DVSS.n255 155.356
R21418 DVSS.n270 DVSS.n263 155.356
R21419 DVSS.n275 DVSS.n255 155.356
R21420 DVSS.n178 DVSS.n157 155.356
R21421 DVSS.n178 DVSS.n158 155.356
R21422 DVSS.n519 DVSS.n518 155.356
R21423 DVSS.n518 DVSS.n517 155.356
R21424 DVSS.n2209 DVSS.n2208 155.356
R21425 DVSS.n2209 DVSS.n2193 155.356
R21426 DVSS.n2277 DVSS.n2104 155.356
R21427 DVSS.n2138 DVSS.n2136 155.356
R21428 DVSS.n2146 DVSS.n2128 155.356
R21429 DVSS.n2143 DVSS.n2136 155.356
R21430 DVSS.n2148 DVSS.n2128 155.356
R21431 DVSS.n2051 DVSS.n2030 155.356
R21432 DVSS.n2051 DVSS.n2031 155.356
R21433 DVSS.n2392 DVSS.n2391 155.356
R21434 DVSS.n2391 DVSS.n2390 155.356
R21435 DVSS.n1017 DVSS.n1016 155.356
R21436 DVSS.n1017 DVSS.n1001 155.356
R21437 DVSS.n1085 DVSS.n912 155.356
R21438 DVSS.n946 DVSS.n944 155.356
R21439 DVSS.n954 DVSS.n936 155.356
R21440 DVSS.n951 DVSS.n944 155.356
R21441 DVSS.n956 DVSS.n936 155.356
R21442 DVSS.n859 DVSS.n838 155.356
R21443 DVSS.n859 DVSS.n839 155.356
R21444 DVSS.n1200 DVSS.n1199 155.356
R21445 DVSS.n1199 DVSS.n1198 155.356
R21446 DVSS.n1539 DVSS.n1538 155.356
R21447 DVSS.n1539 DVSS.n1523 155.356
R21448 DVSS.n1607 DVSS.n1434 155.356
R21449 DVSS.n1468 DVSS.n1466 155.356
R21450 DVSS.n1476 DVSS.n1458 155.356
R21451 DVSS.n1473 DVSS.n1466 155.356
R21452 DVSS.n1478 DVSS.n1458 155.356
R21453 DVSS.n1381 DVSS.n1360 155.356
R21454 DVSS.n1381 DVSS.n1361 155.356
R21455 DVSS.n1722 DVSS.n1721 155.356
R21456 DVSS.n1721 DVSS.n1720 155.356
R21457 DVSS.n2569 DVSS.t189 154.54
R21458 DVSS.n2597 DVSS.n1229 151.625
R21459 DVSS.n428 DVSS.t75 150.504
R21460 DVSS.t75 DVSS.n146 150.504
R21461 DVSS.n526 DVSS.t74 150.504
R21462 DVSS.n90 DVSS.t74 150.504
R21463 DVSS.n2301 DVSS.t156 150.504
R21464 DVSS.t156 DVSS.n2019 150.504
R21465 DVSS.n2399 DVSS.t157 150.504
R21466 DVSS.n1963 DVSS.t157 150.504
R21467 DVSS.n1109 DVSS.t81 150.504
R21468 DVSS.t81 DVSS.n827 150.504
R21469 DVSS.n1207 DVSS.t80 150.504
R21470 DVSS.n771 DVSS.t80 150.504
R21471 DVSS.n1631 DVSS.t84 150.504
R21472 DVSS.t84 DVSS.n1349 150.504
R21473 DVSS.n1729 DVSS.t85 150.504
R21474 DVSS.n1293 DVSS.t85 150.504
R21475 DVSS.t158 DVSS.n2497 145.284
R21476 DVSS.n579 DVSS.t60 144.893
R21477 DVSS.n2581 DVSS.t82 142.876
R21478 DVSS.n2498 DVSS.t158 139.353
R21479 DVSS.n596 DVSS.t60 138.98
R21480 DVSS.n2595 DVSS.t82 137.044
R21481 DVSS.n1924 DVSS.n1923 131.416
R21482 DVSS.n3023 DVSS.n54 131.416
R21483 DVSS.n2855 DVSS.n632 130.613
R21484 DVSS.t72 DVSS.n624 129.845
R21485 DVSS.n2598 DVSS.n2597 128.298
R21486 DVSS.n2480 DVSS.t94 127.493
R21487 DVSS.t148 DVSS.n40 127.151
R21488 DVSS.n1916 DVSS.t122 125.389
R21489 DVSS.n3038 DVSS.t138 125.389
R21490 DVSS.t189 DVSS.n1241 125.382
R21491 DVSS.n2795 DVSS.t26 120.043
R21492 DVSS.n2742 DVSS.t114 120.043
R21493 DVSS.n213 DVSS.t42 119.998
R21494 DVSS.n192 DVSS.t179 119.998
R21495 DVSS.n2086 DVSS.t65 119.998
R21496 DVSS.n2065 DVSS.t12 119.998
R21497 DVSS.n894 DVSS.t175 119.998
R21498 DVSS.n873 DVSS.t54 119.998
R21499 DVSS.n1416 DVSS.t143 119.998
R21500 DVSS.n1395 DVSS.t7 119.998
R21501 DVSS.n405 DVSS.n227 118.938
R21502 DVSS.n2278 DVSS.n2100 118.938
R21503 DVSS.n1086 DVSS.n908 118.938
R21504 DVSS.n1608 DVSS.n1430 118.938
R21505 DVSS.n335 DVSS.n321 118.936
R21506 DVSS.n321 DVSS.n320 118.936
R21507 DVSS.n244 DVSS.n231 118.936
R21508 DVSS.n269 DVSS.n265 118.936
R21509 DVSS.n274 DVSS.n273 118.936
R21510 DVSS.n270 DVSS.n269 118.936
R21511 DVSS.n275 DVSS.n274 118.936
R21512 DVSS.n163 DVSS.n157 118.936
R21513 DVSS.n167 DVSS.n158 118.936
R21514 DVSS.n519 DVSS.n502 118.936
R21515 DVSS.n517 DVSS.n502 118.936
R21516 DVSS.n2208 DVSS.n2194 118.936
R21517 DVSS.n2194 DVSS.n2193 118.936
R21518 DVSS.n2117 DVSS.n2104 118.936
R21519 DVSS.n2142 DVSS.n2138 118.936
R21520 DVSS.n2147 DVSS.n2146 118.936
R21521 DVSS.n2143 DVSS.n2142 118.936
R21522 DVSS.n2148 DVSS.n2147 118.936
R21523 DVSS.n2036 DVSS.n2030 118.936
R21524 DVSS.n2040 DVSS.n2031 118.936
R21525 DVSS.n2392 DVSS.n2375 118.936
R21526 DVSS.n2390 DVSS.n2375 118.936
R21527 DVSS.n1016 DVSS.n1002 118.936
R21528 DVSS.n1002 DVSS.n1001 118.936
R21529 DVSS.n925 DVSS.n912 118.936
R21530 DVSS.n950 DVSS.n946 118.936
R21531 DVSS.n955 DVSS.n954 118.936
R21532 DVSS.n951 DVSS.n950 118.936
R21533 DVSS.n956 DVSS.n955 118.936
R21534 DVSS.n844 DVSS.n838 118.936
R21535 DVSS.n848 DVSS.n839 118.936
R21536 DVSS.n1200 DVSS.n1183 118.936
R21537 DVSS.n1198 DVSS.n1183 118.936
R21538 DVSS.n1538 DVSS.n1524 118.936
R21539 DVSS.n1524 DVSS.n1523 118.936
R21540 DVSS.n1447 DVSS.n1434 118.936
R21541 DVSS.n1472 DVSS.n1468 118.936
R21542 DVSS.n1477 DVSS.n1476 118.936
R21543 DVSS.n1473 DVSS.n1472 118.936
R21544 DVSS.n1478 DVSS.n1477 118.936
R21545 DVSS.n1366 DVSS.n1360 118.936
R21546 DVSS.n1370 DVSS.n1361 118.936
R21547 DVSS.n1722 DVSS.n1705 118.936
R21548 DVSS.n1720 DVSS.n1705 118.936
R21549 DVSS.n376 DVSS.n375 117.719
R21550 DVSS.n384 DVSS.n383 117.719
R21551 DVSS.n373 DVSS.n372 117.719
R21552 DVSS.n2249 DVSS.n2248 117.719
R21553 DVSS.n2257 DVSS.n2256 117.719
R21554 DVSS.n2246 DVSS.n2245 117.719
R21555 DVSS.n1057 DVSS.n1056 117.719
R21556 DVSS.n1065 DVSS.n1064 117.719
R21557 DVSS.n1054 DVSS.n1053 117.719
R21558 DVSS.n1579 DVSS.n1578 117.719
R21559 DVSS.n1587 DVSS.n1586 117.719
R21560 DVSS.n1576 DVSS.n1575 117.719
R21561 DVSS.n383 DVSS.n382 117.719
R21562 DVSS.n372 DVSS.n247 117.719
R21563 DVSS.n2256 DVSS.n2255 117.719
R21564 DVSS.n2245 DVSS.n2120 117.719
R21565 DVSS.n1064 DVSS.n1063 117.719
R21566 DVSS.n1053 DVSS.n928 117.719
R21567 DVSS.n1586 DVSS.n1585 117.719
R21568 DVSS.n1575 DVSS.n1450 117.719
R21569 DVSS.n375 DVSS.n374 117.719
R21570 DVSS.n2248 DVSS.n2247 117.719
R21571 DVSS.n1056 DVSS.n1055 117.719
R21572 DVSS.n1578 DVSS.n1577 117.719
R21573 DVSS.n2980 DVSS.t165 115.689
R21574 DVSS.n2686 DVSS.t69 114.245
R21575 DVSS.n2525 DVSS.t15 114.245
R21576 DVSS.n15 DVSS.t1 114.245
R21577 DVSS.n2421 DVSS.t161 114.245
R21578 DVSS.n2 DVSS.t71 114.245
R21579 DVSS.n3087 DVSS.t91 114.245
R21580 DVSS.n2939 DVSS.t34 113.74
R21581 DVSS.n221 DVSS.n220 112.831
R21582 DVSS.n200 DVSS.n199 112.831
R21583 DVSS.n2094 DVSS.n2093 112.831
R21584 DVSS.n2073 DVSS.n2072 112.831
R21585 DVSS.n902 DVSS.n901 112.831
R21586 DVSS.n881 DVSS.n880 112.831
R21587 DVSS.n1424 DVSS.n1423 112.831
R21588 DVSS.n1403 DVSS.n1402 112.831
R21589 DVSS.n132 DVSS.n123 111.293
R21590 DVSS.n2005 DVSS.n1996 111.293
R21591 DVSS.n813 DVSS.n804 111.293
R21592 DVSS.n1335 DVSS.n1326 111.293
R21593 DVSS.n140 DVSS.n139 111.293
R21594 DVSS.n2013 DVSS.n2012 111.293
R21595 DVSS.n821 DVSS.n820 111.293
R21596 DVSS.n1343 DVSS.n1342 111.293
R21597 DVSS.n2611 DVSS.n749 110.808
R21598 DVSS.n2497 DVSS.t28 109.704
R21599 DVSS.t136 DVSS.n579 109.409
R21600 DVSS.n127 DVSS.n113 108.141
R21601 DVSS.n2000 DVSS.n1986 108.141
R21602 DVSS.n808 DVSS.n794 108.141
R21603 DVSS.n1330 DVSS.n1316 108.141
R21604 DVSS.n473 DVSS.n97 108.141
R21605 DVSS.n479 DVSS.n97 108.141
R21606 DVSS.n469 DVSS.n97 108.141
R21607 DVSS.n486 DVSS.n97 108.141
R21608 DVSS.n2346 DVSS.n1970 108.141
R21609 DVSS.n2352 DVSS.n1970 108.141
R21610 DVSS.n2342 DVSS.n1970 108.141
R21611 DVSS.n2359 DVSS.n1970 108.141
R21612 DVSS.n1154 DVSS.n778 108.141
R21613 DVSS.n1160 DVSS.n778 108.141
R21614 DVSS.n1150 DVSS.n778 108.141
R21615 DVSS.n1167 DVSS.n778 108.141
R21616 DVSS.n1676 DVSS.n1300 108.141
R21617 DVSS.n1682 DVSS.n1300 108.141
R21618 DVSS.n1672 DVSS.n1300 108.141
R21619 DVSS.n1689 DVSS.n1300 108.141
R21620 DVSS.n2926 DVSS.t5 108.037
R21621 DVSS.t104 DVSS.n2581 107.886
R21622 DVSS.n292 DVSS.n255 105.766
R21623 DVSS.n2165 DVSS.n2128 105.766
R21624 DVSS.n973 DVSS.n936 105.766
R21625 DVSS.n1495 DVSS.n1458 105.766
R21626 DVSS.n336 DVSS.n319 105.766
R21627 DVSS.n336 DVSS.n318 105.766
R21628 DVSS.n337 DVSS.n336 105.766
R21629 DVSS.n280 DVSS.n263 105.766
R21630 DVSS.n302 DVSS.n255 105.766
R21631 DVSS.n287 DVSS.n263 105.766
R21632 DVSS.n289 DVSS.n255 105.766
R21633 DVSS.n263 DVSS.n260 105.766
R21634 DVSS.n518 DVSS.n504 105.766
R21635 DVSS.n518 DVSS.n503 105.766
R21636 DVSS.n518 DVSS.n80 105.766
R21637 DVSS.n2209 DVSS.n2192 105.766
R21638 DVSS.n2209 DVSS.n2191 105.766
R21639 DVSS.n2210 DVSS.n2209 105.766
R21640 DVSS.n2153 DVSS.n2136 105.766
R21641 DVSS.n2175 DVSS.n2128 105.766
R21642 DVSS.n2160 DVSS.n2136 105.766
R21643 DVSS.n2162 DVSS.n2128 105.766
R21644 DVSS.n2136 DVSS.n2133 105.766
R21645 DVSS.n2391 DVSS.n2377 105.766
R21646 DVSS.n2391 DVSS.n2376 105.766
R21647 DVSS.n2391 DVSS.n1953 105.766
R21648 DVSS.n1017 DVSS.n1000 105.766
R21649 DVSS.n1017 DVSS.n999 105.766
R21650 DVSS.n1018 DVSS.n1017 105.766
R21651 DVSS.n961 DVSS.n944 105.766
R21652 DVSS.n983 DVSS.n936 105.766
R21653 DVSS.n968 DVSS.n944 105.766
R21654 DVSS.n970 DVSS.n936 105.766
R21655 DVSS.n944 DVSS.n941 105.766
R21656 DVSS.n1199 DVSS.n1185 105.766
R21657 DVSS.n1199 DVSS.n1184 105.766
R21658 DVSS.n1199 DVSS.n761 105.766
R21659 DVSS.n1539 DVSS.n1522 105.766
R21660 DVSS.n1539 DVSS.n1521 105.766
R21661 DVSS.n1540 DVSS.n1539 105.766
R21662 DVSS.n1483 DVSS.n1466 105.766
R21663 DVSS.n1505 DVSS.n1458 105.766
R21664 DVSS.n1490 DVSS.n1466 105.766
R21665 DVSS.n1492 DVSS.n1458 105.766
R21666 DVSS.n1466 DVSS.n1463 105.766
R21667 DVSS.n1721 DVSS.n1707 105.766
R21668 DVSS.n1721 DVSS.n1706 105.766
R21669 DVSS.n1721 DVSS.n1283 105.766
R21670 DVSS.n2858 DVSS.t72 105.346
R21671 DVSS.n216 DVSS.n215 104.172
R21672 DVSS.n195 DVSS.n194 104.172
R21673 DVSS.n2089 DVSS.n2088 104.172
R21674 DVSS.n2068 DVSS.n2067 104.172
R21675 DVSS.n897 DVSS.n896 104.172
R21676 DVSS.n876 DVSS.n875 104.172
R21677 DVSS.n1419 DVSS.n1418 104.172
R21678 DVSS.n1398 DVSS.n1397 104.172
R21679 DVSS.n114 DVSS.t39 101.811
R21680 DVSS.t40 DVSS.n96 101.811
R21681 DVSS.n1987 DVSS.t63 101.811
R21682 DVSS.t62 DVSS.n1969 101.811
R21683 DVSS.n795 DVSS.t172 101.811
R21684 DVSS.t173 DVSS.n777 101.811
R21685 DVSS.n1317 DVSS.t145 101.811
R21686 DVSS.t144 DVSS.n1299 101.811
R21687 DVSS.t20 DVSS.n2778 101.575
R21688 DVSS.t106 DVSS.n2718 101.575
R21689 DVSS.n2669 DVSS.t67 101.038
R21690 DVSS.n2538 DVSS.t17 101.038
R21691 DVSS.n3060 DVSS.t3 101.038
R21692 DVSS.n2434 DVSS.t163 101.038
R21693 DVSS.n628 DVSS.t73 101.038
R21694 DVSS.n13 DVSS.t10 101.038
R21695 DVSS.n403 DVSS.n402 93.9796
R21696 DVSS.n238 DVSS.n235 93.9796
R21697 DVSS.n395 DVSS.n234 93.9796
R21698 DVSS.n392 DVSS.n233 93.9796
R21699 DVSS.n244 DVSS.n232 93.9796
R21700 DVSS.n392 DVSS.n232 93.9796
R21701 DVSS.n395 DVSS.n233 93.9796
R21702 DVSS.n238 DVSS.n234 93.9796
R21703 DVSS.n402 DVSS.n235 93.9796
R21704 DVSS.n403 DVSS.n227 93.9796
R21705 DVSS.n177 DVSS.n176 93.9796
R21706 DVSS.n173 DVSS.n162 93.9796
R21707 DVSS.n171 DVSS.n161 93.9796
R21708 DVSS.n169 DVSS.n160 93.9796
R21709 DVSS.n167 DVSS.n159 93.9796
R21710 DVSS.n176 DVSS.n162 93.9796
R21711 DVSS.n173 DVSS.n161 93.9796
R21712 DVSS.n171 DVSS.n160 93.9796
R21713 DVSS.n169 DVSS.n159 93.9796
R21714 DVSS.n177 DVSS.n163 93.9796
R21715 DVSS.n2276 DVSS.n2275 93.9796
R21716 DVSS.n2111 DVSS.n2108 93.9796
R21717 DVSS.n2268 DVSS.n2107 93.9796
R21718 DVSS.n2265 DVSS.n2106 93.9796
R21719 DVSS.n2117 DVSS.n2105 93.9796
R21720 DVSS.n2265 DVSS.n2105 93.9796
R21721 DVSS.n2268 DVSS.n2106 93.9796
R21722 DVSS.n2111 DVSS.n2107 93.9796
R21723 DVSS.n2275 DVSS.n2108 93.9796
R21724 DVSS.n2276 DVSS.n2100 93.9796
R21725 DVSS.n2050 DVSS.n2049 93.9796
R21726 DVSS.n2046 DVSS.n2035 93.9796
R21727 DVSS.n2044 DVSS.n2034 93.9796
R21728 DVSS.n2042 DVSS.n2033 93.9796
R21729 DVSS.n2040 DVSS.n2032 93.9796
R21730 DVSS.n2049 DVSS.n2035 93.9796
R21731 DVSS.n2046 DVSS.n2034 93.9796
R21732 DVSS.n2044 DVSS.n2033 93.9796
R21733 DVSS.n2042 DVSS.n2032 93.9796
R21734 DVSS.n2050 DVSS.n2036 93.9796
R21735 DVSS.n1084 DVSS.n1083 93.9796
R21736 DVSS.n919 DVSS.n916 93.9796
R21737 DVSS.n1076 DVSS.n915 93.9796
R21738 DVSS.n1073 DVSS.n914 93.9796
R21739 DVSS.n925 DVSS.n913 93.9796
R21740 DVSS.n1073 DVSS.n913 93.9796
R21741 DVSS.n1076 DVSS.n914 93.9796
R21742 DVSS.n919 DVSS.n915 93.9796
R21743 DVSS.n1083 DVSS.n916 93.9796
R21744 DVSS.n1084 DVSS.n908 93.9796
R21745 DVSS.n858 DVSS.n857 93.9796
R21746 DVSS.n854 DVSS.n843 93.9796
R21747 DVSS.n852 DVSS.n842 93.9796
R21748 DVSS.n850 DVSS.n841 93.9796
R21749 DVSS.n848 DVSS.n840 93.9796
R21750 DVSS.n857 DVSS.n843 93.9796
R21751 DVSS.n854 DVSS.n842 93.9796
R21752 DVSS.n852 DVSS.n841 93.9796
R21753 DVSS.n850 DVSS.n840 93.9796
R21754 DVSS.n858 DVSS.n844 93.9796
R21755 DVSS.n1606 DVSS.n1605 93.9796
R21756 DVSS.n1441 DVSS.n1438 93.9796
R21757 DVSS.n1598 DVSS.n1437 93.9796
R21758 DVSS.n1595 DVSS.n1436 93.9796
R21759 DVSS.n1447 DVSS.n1435 93.9796
R21760 DVSS.n1595 DVSS.n1435 93.9796
R21761 DVSS.n1598 DVSS.n1436 93.9796
R21762 DVSS.n1441 DVSS.n1437 93.9796
R21763 DVSS.n1605 DVSS.n1438 93.9796
R21764 DVSS.n1606 DVSS.n1430 93.9796
R21765 DVSS.n1380 DVSS.n1379 93.9796
R21766 DVSS.n1376 DVSS.n1365 93.9796
R21767 DVSS.n1374 DVSS.n1364 93.9796
R21768 DVSS.n1372 DVSS.n1363 93.9796
R21769 DVSS.n1370 DVSS.n1362 93.9796
R21770 DVSS.n1379 DVSS.n1365 93.9796
R21771 DVSS.n1376 DVSS.n1364 93.9796
R21772 DVSS.n1374 DVSS.n1363 93.9796
R21773 DVSS.n1372 DVSS.n1362 93.9796
R21774 DVSS.n1380 DVSS.n1366 93.9796
R21775 DVSS.n215 DVSS.n214 92.5005
R21776 DVSS.n194 DVSS.n193 92.5005
R21777 DVSS.n2088 DVSS.n2087 92.5005
R21778 DVSS.n2067 DVSS.n2066 92.5005
R21779 DVSS.n896 DVSS.n895 92.5005
R21780 DVSS.n875 DVSS.n874 92.5005
R21781 DVSS.n1418 DVSS.n1417 92.5005
R21782 DVSS.n1397 DVSS.n1396 92.5005
R21783 DVSS.n2778 DVSS.n701 92.3405
R21784 DVSS.t100 DVSS.n2467 91.9142
R21785 DVSS.n3041 DVSS.t152 91.6672
R21786 DVSS.n2940 DVSS.t31 91.1965
R21787 DVSS.n2939 DVSS.t36 91.1965
R21788 DVSS.n2574 DVSS.t190 90.704
R21789 DVSS.n572 DVSS.t149 90.704
R21790 DVSS.n2475 DVSS.t95 90.704
R21791 DVSS.n1857 DVSS.t44 90.704
R21792 DVSS.n60 DVSS.t133 90.703
R21793 DVSS.n1933 DVSS.t127 90.703
R21794 DVSS.n752 DVSS.t107 90.703
R21795 DVSS.n705 DVSS.t21 90.703
R21796 DVSS.t185 DVSS.n2565 90.3915
R21797 DVSS.n134 DVSS.n133 87.6383
R21798 DVSS.n136 DVSS.n135 87.6383
R21799 DVSS.n139 DVSS.n121 87.6383
R21800 DVSS.n133 DVSS.n132 87.6383
R21801 DVSS.n135 DVSS.n134 87.6383
R21802 DVSS.n136 DVSS.n121 87.6383
R21803 DVSS.n2007 DVSS.n2006 87.6383
R21804 DVSS.n2009 DVSS.n2008 87.6383
R21805 DVSS.n2012 DVSS.n1994 87.6383
R21806 DVSS.n2006 DVSS.n2005 87.6383
R21807 DVSS.n2008 DVSS.n2007 87.6383
R21808 DVSS.n2009 DVSS.n1994 87.6383
R21809 DVSS.n815 DVSS.n814 87.6383
R21810 DVSS.n817 DVSS.n816 87.6383
R21811 DVSS.n820 DVSS.n802 87.6383
R21812 DVSS.n814 DVSS.n813 87.6383
R21813 DVSS.n816 DVSS.n815 87.6383
R21814 DVSS.n817 DVSS.n802 87.6383
R21815 DVSS.n1337 DVSS.n1336 87.6383
R21816 DVSS.n1339 DVSS.n1338 87.6383
R21817 DVSS.n1342 DVSS.n1324 87.6383
R21818 DVSS.n1336 DVSS.n1335 87.6383
R21819 DVSS.n1338 DVSS.n1337 87.6383
R21820 DVSS.n1339 DVSS.n1324 87.6383
R21821 DVSS.n383 DVSS.n229 87.3927
R21822 DVSS.n372 DVSS.n242 87.3927
R21823 DVSS.n2256 DVSS.n2102 87.3927
R21824 DVSS.n2245 DVSS.n2115 87.3927
R21825 DVSS.n1064 DVSS.n910 87.3927
R21826 DVSS.n1053 DVSS.n923 87.3927
R21827 DVSS.n1586 DVSS.n1432 87.3927
R21828 DVSS.n1575 DVSS.n1445 87.3927
R21829 DVSS.n2466 DVSS.t98 85.9843
R21830 DVSS.n3040 DVSS.t150 85.7532
R21831 DVSS.n2619 DVSS.t92 85.3621
R21832 DVSS.n1877 DVSS.t176 85.3621
R21833 DVSS.t88 DVSS.n2764 85.3621
R21834 DVSS.n2816 DVSS.t140 85.3621
R21835 DVSS.t183 DVSS.n1251 84.5598
R21836 DVSS.t166 DVSS.t58 82.3134
R21837 DVSS.n292 DVSS.n257 80.9725
R21838 DVSS.n2165 DVSS.n2130 80.9725
R21839 DVSS.n973 DVSS.n938 80.9725
R21840 DVSS.n1495 DVSS.n1460 80.9725
R21841 DVSS.n293 DVSS.n292 80.9721
R21842 DVSS.n2166 DVSS.n2165 80.9721
R21843 DVSS.n974 DVSS.n973 80.9721
R21844 DVSS.n1496 DVSS.n1495 80.9721
R21845 DVSS.n302 DVSS.n301 80.9719
R21846 DVSS.n294 DVSS.n289 80.9719
R21847 DVSS.n326 DVSS.n319 80.9719
R21848 DVSS.n322 DVSS.n318 80.9719
R21849 DVSS.n338 DVSS.n337 80.9719
R21850 DVSS.n281 DVSS.n280 80.9719
R21851 DVSS.n288 DVSS.n287 80.9719
R21852 DVSS.n352 DVSS.n260 80.9719
R21853 DVSS.n329 DVSS.n319 80.9719
R21854 DVSS.n325 DVSS.n318 80.9719
R21855 DVSS.n337 DVSS.n317 80.9719
R21856 DVSS.n280 DVSS.n279 80.9719
R21857 DVSS.n303 DVSS.n302 80.9719
R21858 DVSS.n287 DVSS.n286 80.9719
R21859 DVSS.n289 DVSS.n277 80.9719
R21860 DVSS.n290 DVSS.n260 80.9719
R21861 DVSS.n512 DVSS.n504 80.9719
R21862 DVSS.n508 DVSS.n503 80.9719
R21863 DVSS.n536 DVSS.n80 80.9719
R21864 DVSS.n505 DVSS.n504 80.9719
R21865 DVSS.n511 DVSS.n503 80.9719
R21866 DVSS.n507 DVSS.n80 80.9719
R21867 DVSS.n2175 DVSS.n2174 80.9719
R21868 DVSS.n2167 DVSS.n2162 80.9719
R21869 DVSS.n2199 DVSS.n2192 80.9719
R21870 DVSS.n2195 DVSS.n2191 80.9719
R21871 DVSS.n2211 DVSS.n2210 80.9719
R21872 DVSS.n2154 DVSS.n2153 80.9719
R21873 DVSS.n2161 DVSS.n2160 80.9719
R21874 DVSS.n2225 DVSS.n2133 80.9719
R21875 DVSS.n2202 DVSS.n2192 80.9719
R21876 DVSS.n2198 DVSS.n2191 80.9719
R21877 DVSS.n2210 DVSS.n2190 80.9719
R21878 DVSS.n2153 DVSS.n2152 80.9719
R21879 DVSS.n2176 DVSS.n2175 80.9719
R21880 DVSS.n2160 DVSS.n2159 80.9719
R21881 DVSS.n2162 DVSS.n2150 80.9719
R21882 DVSS.n2163 DVSS.n2133 80.9719
R21883 DVSS.n2385 DVSS.n2377 80.9719
R21884 DVSS.n2381 DVSS.n2376 80.9719
R21885 DVSS.n2409 DVSS.n1953 80.9719
R21886 DVSS.n2378 DVSS.n2377 80.9719
R21887 DVSS.n2384 DVSS.n2376 80.9719
R21888 DVSS.n2380 DVSS.n1953 80.9719
R21889 DVSS.n983 DVSS.n982 80.9719
R21890 DVSS.n975 DVSS.n970 80.9719
R21891 DVSS.n1007 DVSS.n1000 80.9719
R21892 DVSS.n1003 DVSS.n999 80.9719
R21893 DVSS.n1019 DVSS.n1018 80.9719
R21894 DVSS.n962 DVSS.n961 80.9719
R21895 DVSS.n969 DVSS.n968 80.9719
R21896 DVSS.n1033 DVSS.n941 80.9719
R21897 DVSS.n1010 DVSS.n1000 80.9719
R21898 DVSS.n1006 DVSS.n999 80.9719
R21899 DVSS.n1018 DVSS.n998 80.9719
R21900 DVSS.n961 DVSS.n960 80.9719
R21901 DVSS.n984 DVSS.n983 80.9719
R21902 DVSS.n968 DVSS.n967 80.9719
R21903 DVSS.n970 DVSS.n958 80.9719
R21904 DVSS.n971 DVSS.n941 80.9719
R21905 DVSS.n1193 DVSS.n1185 80.9719
R21906 DVSS.n1189 DVSS.n1184 80.9719
R21907 DVSS.n1217 DVSS.n761 80.9719
R21908 DVSS.n1186 DVSS.n1185 80.9719
R21909 DVSS.n1192 DVSS.n1184 80.9719
R21910 DVSS.n1188 DVSS.n761 80.9719
R21911 DVSS.n1505 DVSS.n1504 80.9719
R21912 DVSS.n1497 DVSS.n1492 80.9719
R21913 DVSS.n1529 DVSS.n1522 80.9719
R21914 DVSS.n1525 DVSS.n1521 80.9719
R21915 DVSS.n1541 DVSS.n1540 80.9719
R21916 DVSS.n1484 DVSS.n1483 80.9719
R21917 DVSS.n1491 DVSS.n1490 80.9719
R21918 DVSS.n1555 DVSS.n1463 80.9719
R21919 DVSS.n1532 DVSS.n1522 80.9719
R21920 DVSS.n1528 DVSS.n1521 80.9719
R21921 DVSS.n1540 DVSS.n1520 80.9719
R21922 DVSS.n1483 DVSS.n1482 80.9719
R21923 DVSS.n1506 DVSS.n1505 80.9719
R21924 DVSS.n1490 DVSS.n1489 80.9719
R21925 DVSS.n1492 DVSS.n1480 80.9719
R21926 DVSS.n1493 DVSS.n1463 80.9719
R21927 DVSS.n1715 DVSS.n1707 80.9719
R21928 DVSS.n1711 DVSS.n1706 80.9719
R21929 DVSS.n1739 DVSS.n1283 80.9719
R21930 DVSS.n1708 DVSS.n1707 80.9719
R21931 DVSS.n1714 DVSS.n1706 80.9719
R21932 DVSS.n1710 DVSS.n1283 80.9719
R21933 DVSS.t120 DVSS.n1808 77.6019
R21934 DVSS.t130 DVSS.n3037 77.6019
R21935 DVSS.n2574 DVSS.n1245 76.7239
R21936 DVSS.n2552 DVSS.n1245 76.7239
R21937 DVSS.n3046 DVSS.n31 76.7239
R21938 DVSS.n572 DVSS.n31 76.7239
R21939 DVSS.n2632 DVSS.n49 76.7239
R21940 DVSS.n60 DVSS.n49 76.7239
R21941 DVSS.n2475 DVSS.n2474 76.7239
R21942 DVSS.n2474 DVSS.n2473 76.7239
R21943 DVSS.n1857 DVSS.n1856 76.7239
R21944 DVSS.n1856 DVSS.n1855 76.7239
R21945 DVSS.n1932 DVSS.n1798 76.7239
R21946 DVSS.n1933 DVSS.n1932 76.7239
R21947 DVSS.n2737 DVSS.n736 76.7239
R21948 DVSS.n752 DVSS.n736 76.7239
R21949 DVSS.n694 DVSS.n693 76.7239
R21950 DVSS.n705 DVSS.n694 76.7239
R21951 DVSS.n3007 DVSS.n620 76.4173
R21952 DVSS.n128 DVSS.n127 76.2208
R21953 DVSS.n2001 DVSS.n2000 76.2208
R21954 DVSS.n809 DVSS.n808 76.2208
R21955 DVSS.n1331 DVSS.n1330 76.2208
R21956 DVSS.n127 DVSS.n126 76.2204
R21957 DVSS.n2000 DVSS.n1999 76.2204
R21958 DVSS.n808 DVSS.n807 76.2204
R21959 DVSS.n1330 DVSS.n1329 76.2204
R21960 DVSS.n473 DVSS.n471 76.2201
R21961 DVSS.n480 DVSS.n479 76.2201
R21962 DVSS.n484 DVSS.n469 76.2201
R21963 DVSS.n487 DVSS.n486 76.2201
R21964 DVSS.n474 DVSS.n473 76.2201
R21965 DVSS.n479 DVSS.n478 76.2201
R21966 DVSS.n481 DVSS.n469 76.2201
R21967 DVSS.n486 DVSS.n485 76.2201
R21968 DVSS.n2346 DVSS.n2344 76.2201
R21969 DVSS.n2353 DVSS.n2352 76.2201
R21970 DVSS.n2357 DVSS.n2342 76.2201
R21971 DVSS.n2360 DVSS.n2359 76.2201
R21972 DVSS.n2347 DVSS.n2346 76.2201
R21973 DVSS.n2352 DVSS.n2351 76.2201
R21974 DVSS.n2354 DVSS.n2342 76.2201
R21975 DVSS.n2359 DVSS.n2358 76.2201
R21976 DVSS.n1154 DVSS.n1152 76.2201
R21977 DVSS.n1161 DVSS.n1160 76.2201
R21978 DVSS.n1165 DVSS.n1150 76.2201
R21979 DVSS.n1168 DVSS.n1167 76.2201
R21980 DVSS.n1155 DVSS.n1154 76.2201
R21981 DVSS.n1160 DVSS.n1159 76.2201
R21982 DVSS.n1162 DVSS.n1150 76.2201
R21983 DVSS.n1167 DVSS.n1166 76.2201
R21984 DVSS.n1676 DVSS.n1674 76.2201
R21985 DVSS.n1683 DVSS.n1682 76.2201
R21986 DVSS.n1687 DVSS.n1672 76.2201
R21987 DVSS.n1690 DVSS.n1689 76.2201
R21988 DVSS.n1677 DVSS.n1676 76.2201
R21989 DVSS.n1682 DVSS.n1681 76.2201
R21990 DVSS.n1684 DVSS.n1672 76.2201
R21991 DVSS.n1689 DVSS.n1688 76.2201
R21992 DVSS.n601 DVSS.n55 70.9682
R21993 DVSS.n2609 DVSS.n2608 69.9806
R21994 DVSS.n2589 DVSS.n2588 69.3226
R21995 DVSS.n587 DVSS.n586 69.3226
R21996 DVSS.n2490 DVSS.n2489 69.3226
R21997 DVSS.n648 DVSS.n647 69.3226
R21998 DVSS.n3083 DVSS.t90 69.0588
R21999 DVSS.n3069 DVSS.t0 68.4449
R22000 DVSS.n215 DVSS.t42 66.8281
R22001 DVSS.n194 DVSS.t179 66.8281
R22002 DVSS.n2088 DVSS.t65 66.8281
R22003 DVSS.n2067 DVSS.t12 66.8281
R22004 DVSS.n896 DVSS.t175 66.8281
R22005 DVSS.n875 DVSS.t54 66.8281
R22006 DVSS.n1418 DVSS.t143 66.8281
R22007 DVSS.n1397 DVSS.t7 66.8281
R22008 DVSS.n1925 DVSS.t116 64.639
R22009 DVSS.n3025 DVSS.t128 64.639
R22010 DVSS.n2780 DVSS.t22 64.6385
R22011 DVSS.t110 DVSS.n741 64.6385
R22012 DVSS.n406 DVSS.n405 59.4692
R22013 DVSS.n2279 DVSS.n2278 59.4692
R22014 DVSS.n1087 DVSS.n1086 59.4692
R22015 DVSS.n1609 DVSS.n1608 59.4692
R22016 DVSS.n273 DVSS.n254 59.4689
R22017 DVSS.n304 DVSS.n275 59.4689
R22018 DVSS.n386 DVSS.n231 59.4689
R22019 DVSS.n335 DVSS.n334 59.4689
R22020 DVSS.n330 DVSS.n320 59.4689
R22021 DVSS.n311 DVSS.n265 59.4689
R22022 DVSS.n271 DVSS.n270 59.4689
R22023 DVSS.n164 DVSS.n157 59.4689
R22024 DVSS.n158 DVSS.n156 59.4689
R22025 DVSS.n520 DVSS.n519 59.4689
R22026 DVSS.n517 DVSS.n516 59.4689
R22027 DVSS.n2146 DVSS.n2127 59.4689
R22028 DVSS.n2177 DVSS.n2148 59.4689
R22029 DVSS.n2259 DVSS.n2104 59.4689
R22030 DVSS.n2208 DVSS.n2207 59.4689
R22031 DVSS.n2203 DVSS.n2193 59.4689
R22032 DVSS.n2184 DVSS.n2138 59.4689
R22033 DVSS.n2144 DVSS.n2143 59.4689
R22034 DVSS.n2037 DVSS.n2030 59.4689
R22035 DVSS.n2031 DVSS.n2029 59.4689
R22036 DVSS.n2393 DVSS.n2392 59.4689
R22037 DVSS.n2390 DVSS.n2389 59.4689
R22038 DVSS.n954 DVSS.n935 59.4689
R22039 DVSS.n985 DVSS.n956 59.4689
R22040 DVSS.n1067 DVSS.n912 59.4689
R22041 DVSS.n1016 DVSS.n1015 59.4689
R22042 DVSS.n1011 DVSS.n1001 59.4689
R22043 DVSS.n992 DVSS.n946 59.4689
R22044 DVSS.n952 DVSS.n951 59.4689
R22045 DVSS.n845 DVSS.n838 59.4689
R22046 DVSS.n839 DVSS.n837 59.4689
R22047 DVSS.n1201 DVSS.n1200 59.4689
R22048 DVSS.n1198 DVSS.n1197 59.4689
R22049 DVSS.n1476 DVSS.n1457 59.4689
R22050 DVSS.n1507 DVSS.n1478 59.4689
R22051 DVSS.n1589 DVSS.n1434 59.4689
R22052 DVSS.n1538 DVSS.n1537 59.4689
R22053 DVSS.n1533 DVSS.n1523 59.4689
R22054 DVSS.n1514 DVSS.n1468 59.4689
R22055 DVSS.n1474 DVSS.n1473 59.4689
R22056 DVSS.n1367 DVSS.n1360 59.4689
R22057 DVSS.n1361 DVSS.n1359 59.4689
R22058 DVSS.n1723 DVSS.n1722 59.4689
R22059 DVSS.n1720 DVSS.n1719 59.4689
R22060 DVSS.n2954 DVSS.n2953 59.3519
R22061 DVSS.n2897 DVSS.n2896 59.3519
R22062 DVSS.n2499 DVSS.n1754 59.2997
R22063 DVSS.n1809 DVSS.t51 57.1434
R22064 DVSS.n129 DVSS.n123 55.6474
R22065 DVSS.n2002 DVSS.n1996 55.6474
R22066 DVSS.n810 DVSS.n804 55.6474
R22067 DVSS.n1332 DVSS.n1326 55.6474
R22068 DVSS.n141 DVSS.n140 55.6471
R22069 DVSS.n2014 DVSS.n2013 55.6471
R22070 DVSS.n822 DVSS.n821 55.6471
R22071 DVSS.n1344 DVSS.n1343 55.6471
R22072 DVSS.n2766 DVSS.n713 54.6435
R22073 DVSS.n1851 DVSS.n1850 53.4435
R22074 DVSS.n2615 DVSS.n2614 52.3069
R22075 DVSS.n1884 DVSS.n1883 52.3069
R22076 DVSS.n721 DVSS.n720 52.3069
R22077 DVSS.n671 DVSS.n670 52.3069
R22078 DVSS.t26 DVSS.n2794 50.7875
R22079 DVSS.n2568 DVSS.t114 50.7875
R22080 DVSS.n1925 DVSS.n1805 47.1783
R22081 DVSS.n3026 DVSS.n3025 47.1783
R22082 DVSS.t24 DVSS.n2792 46.1705
R22083 DVSS.n2732 DVSS.t112 46.1705
R22084 DVSS.n333 DVSS.n312 45.5782
R22085 DVSS.n340 DVSS.n339 45.5782
R22086 DVSS.n2206 DVSS.n2185 45.5782
R22087 DVSS.n2213 DVSS.n2212 45.5782
R22088 DVSS.n1014 DVSS.n993 45.5782
R22089 DVSS.n1021 DVSS.n1020 45.5782
R22090 DVSS.n1536 DVSS.n1515 45.5782
R22091 DVSS.n1543 DVSS.n1542 45.5782
R22092 DVSS.n2980 DVSS.n2979 43.8838
R22093 DVSS.n378 DVSS.n377 42.4097
R22094 DVSS.n2251 DVSS.n2250 42.4097
R22095 DVSS.n1059 DVSS.n1058 42.4097
R22096 DVSS.n1581 DVSS.n1580 42.4097
R22097 DVSS.t49 DVSS.n1837 40.8168
R22098 DVSS.n3089 DVSS.n1 39.8886
R22099 DVSS.n2662 DVSS.n2611 38.7626
R22100 DVSS.n2426 DVSS.t160 38.0722
R22101 DVSS.t68 DVSS.n20 38.0722
R22102 DVSS.n408 DVSS.n224 36.7611
R22103 DVSS.n2281 DVSS.n2097 36.7611
R22104 DVSS.n1089 DVSS.n905 36.7611
R22105 DVSS.n1611 DVSS.n1427 36.7611
R22106 DVSS.t4 DVSS.t30 36.1979
R22107 DVSS.n3002 DVSS.n2885 36.1417
R22108 DVSS.n3002 DVSS.n3000 36.1417
R22109 DVSS.n3000 DVSS.n2998 36.1417
R22110 DVSS.n2998 DVSS.n2888 36.1417
R22111 DVSS.n2993 DVSS.n2888 36.1417
R22112 DVSS.n2993 DVSS.n2991 36.1417
R22113 DVSS.n2991 DVSS.n2989 36.1417
R22114 DVSS.n2989 DVSS.n2986 36.1417
R22115 DVSS.n2986 DVSS.n2985 36.1417
R22116 DVSS.n2985 DVSS.n2892 36.1417
R22117 DVSS.n2976 DVSS.n2892 36.1417
R22118 DVSS.n2976 DVSS.n2973 36.1417
R22119 DVSS.n2973 DVSS.n2972 36.1417
R22120 DVSS.n2972 DVSS.n2894 36.1417
R22121 DVSS.n2965 DVSS.n2894 36.1417
R22122 DVSS.n2688 DVSS.n2664 36.1417
R22123 DVSS.n2683 DVSS.n2664 36.1417
R22124 DVSS.n2683 DVSS.n2666 36.1417
R22125 DVSS.n2677 DVSS.n2666 36.1417
R22126 DVSS.n2673 DVSS.n26 36.1417
R22127 DVSS.n3050 DVSS.n26 36.1417
R22128 DVSS.n3050 DVSS.n3049 36.1417
R22129 DVSS.n3049 DVSS.n28 36.1417
R22130 DVSS.n3043 DVSS.n28 36.1417
R22131 DVSS.n3043 DVSS.n33 36.1417
R22132 DVSS.n565 DVSS.n33 36.1417
R22133 DVSS.n566 DVSS.n565 36.1417
R22134 DVSS.n569 DVSS.n566 36.1417
R22135 DVSS.n569 DVSS.n557 36.1417
R22136 DVSS.n575 DVSS.n557 36.1417
R22137 DVSS.n575 DVSS.n554 36.1417
R22138 DVSS.n582 DVSS.n554 36.1417
R22139 DVSS.n582 DVSS.n550 36.1417
R22140 DVSS.n594 DVSS.n550 36.1417
R22141 DVSS.n594 DVSS.n551 36.1417
R22142 DVSS.n551 DVSS.n548 36.1417
R22143 DVSS.n548 DVSS.n545 36.1417
R22144 DVSS.n604 DVSS.n545 36.1417
R22145 DVSS.n2656 DVSS.n2613 36.1417
R22146 DVSS.n2656 DVSS.n2617 36.1417
R22147 DVSS.n2650 DVSS.n2617 36.1417
R22148 DVSS.n2650 DVSS.n2622 36.1417
R22149 DVSS.n2646 DVSS.n2622 36.1417
R22150 DVSS.n2646 DVSS.n2625 36.1417
R22151 DVSS.n2640 DVSS.n2625 36.1417
R22152 DVSS.n2640 DVSS.n2629 36.1417
R22153 DVSS.n2636 DVSS.n2629 36.1417
R22154 DVSS.n2636 DVSS.n45 36.1417
R22155 DVSS.n3035 DVSS.n45 36.1417
R22156 DVSS.n3035 DVSS.n46 36.1417
R22157 DVSS.n51 DVSS.n46 36.1417
R22158 DVSS.n3027 DVSS.n51 36.1417
R22159 DVSS.n3027 DVSS.n52 36.1417
R22160 DVSS.n3020 DVSS.n52 36.1417
R22161 DVSS.n3020 DVSS.n3019 36.1417
R22162 DVSS.n3019 DVSS.n59 36.1417
R22163 DVSS.n3072 DVSS.n3071 36.1417
R22164 DVSS.n3071 DVSS.n17 36.1417
R22165 DVSS.n3065 DVSS.n17 36.1417
R22166 DVSS.n3065 DVSS.n3057 36.1417
R22167 DVSS.n2423 DVSS.n1787 36.1417
R22168 DVSS.n2430 DVSS.n1787 36.1417
R22169 DVSS.n2430 DVSS.n1784 36.1417
R22170 DVSS.n2437 DVSS.n1784 36.1417
R22171 DVSS.n2865 DVSS.n626 36.1417
R22172 DVSS.n2865 DVSS.n627 36.1417
R22173 DVSS.n2860 DVSS.n627 36.1417
R22174 DVSS.n2860 DVSS.n629 36.1417
R22175 DVSS.n1887 DVSS.n1879 36.1417
R22176 DVSS.n1887 DVSS.n1875 36.1417
R22177 DVSS.n1893 DVSS.n1875 36.1417
R22178 DVSS.n1893 DVSS.n1873 36.1417
R22179 DVSS.n1897 DVSS.n1873 36.1417
R22180 DVSS.n1897 DVSS.n1869 36.1417
R22181 DVSS.n1903 DVSS.n1869 36.1417
R22182 DVSS.n1903 DVSS.n1866 36.1417
R22183 DVSS.n1913 DVSS.n1866 36.1417
R22184 DVSS.n1913 DVSS.n1867 36.1417
R22185 DVSS.n1907 DVSS.n1867 36.1417
R22186 DVSS.n1907 DVSS.n1802 36.1417
R22187 DVSS.n1928 DVSS.n1802 36.1417
R22188 DVSS.n1928 DVSS.n1803 36.1417
R22189 DVSS.n1922 DVSS.n1803 36.1417
R22190 DVSS.n1922 DVSS.n1919 36.1417
R22191 DVSS.n1919 DVSS.n1795 36.1417
R22192 DVSS.n1942 DVSS.n1795 36.1417
R22193 DVSS.n1829 DVSS.n1824 36.1417
R22194 DVSS.n1834 DVSS.n1824 36.1417
R22195 DVSS.n1834 DVSS.n1819 36.1417
R22196 DVSS.n1852 DVSS.n1819 36.1417
R22197 DVSS.n1852 DVSS.n1820 36.1417
R22198 DVSS.n1846 DVSS.n1820 36.1417
R22199 DVSS.n1846 DVSS.n1840 36.1417
R22200 DVSS.n1840 DVSS.n1811 36.1417
R22201 DVSS.n1860 DVSS.n1811 36.1417
R22202 DVSS.n1860 DVSS.n636 36.1417
R22203 DVSS.n2851 DVSS.n636 36.1417
R22204 DVSS.n2851 DVSS.n637 36.1417
R22205 DVSS.n2847 DVSS.n637 36.1417
R22206 DVSS.n2847 DVSS.n640 36.1417
R22207 DVSS.n2841 DVSS.n640 36.1417
R22208 DVSS.n2841 DVSS.n644 36.1417
R22209 DVSS.n2837 DVSS.n644 36.1417
R22210 DVSS.n2837 DVSS.n651 36.1417
R22211 DVSS.n2830 DVSS.n651 36.1417
R22212 DVSS.n2762 DVSS.n2761 36.1417
R22213 DVSS.n2761 DVSS.n718 36.1417
R22214 DVSS.n2756 DVSS.n718 36.1417
R22215 DVSS.n2756 DVSS.n723 36.1417
R22216 DVSS.n2750 DVSS.n723 36.1417
R22217 DVSS.n2750 DVSS.n729 36.1417
R22218 DVSS.n2746 DVSS.n729 36.1417
R22219 DVSS.n2746 DVSS.n731 36.1417
R22220 DVSS.n2740 DVSS.n731 36.1417
R22221 DVSS.n2740 DVSS.n734 36.1417
R22222 DVSS.n2734 DVSS.n734 36.1417
R22223 DVSS.n2734 DVSS.n739 36.1417
R22224 DVSS.n2728 DVSS.n739 36.1417
R22225 DVSS.n2728 DVSS.n743 36.1417
R22226 DVSS.n2721 DVSS.n743 36.1417
R22227 DVSS.n2721 DVSS.n746 36.1417
R22228 DVSS.n2714 DVSS.n746 36.1417
R22229 DVSS.n2714 DVSS.n751 36.1417
R22230 DVSS.n2543 DVSS.n1263 36.1417
R22231 DVSS.n2543 DVSS.n1259 36.1417
R22232 DVSS.n2549 DVSS.n1259 36.1417
R22233 DVSS.n2549 DVSS.n1255 36.1417
R22234 DVSS.n2563 DVSS.n1255 36.1417
R22235 DVSS.n2563 DVSS.n2562 36.1417
R22236 DVSS.n2562 DVSS.n2555 36.1417
R22237 DVSS.n2555 DVSS.n1247 36.1417
R22238 DVSS.n2571 DVSS.n1247 36.1417
R22239 DVSS.n2571 DVSS.n1243 36.1417
R22240 DVSS.n2577 DVSS.n1243 36.1417
R22241 DVSS.n2577 DVSS.n1239 36.1417
R22242 DVSS.n2584 DVSS.n1239 36.1417
R22243 DVSS.n2584 DVSS.n1236 36.1417
R22244 DVSS.n2593 DVSS.n1236 36.1417
R22245 DVSS.n2593 DVSS.n1233 36.1417
R22246 DVSS.n2600 DVSS.n1233 36.1417
R22247 DVSS.n2600 DVSS.n1231 36.1417
R22248 DVSS.n2606 DVSS.n1231 36.1417
R22249 DVSS.n2528 DVSS.n1273 36.1417
R22250 DVSS.n2528 DVSS.n1267 36.1417
R22251 DVSS.n2535 DVSS.n1267 36.1417
R22252 DVSS.n2535 DVSS.n1268 36.1417
R22253 DVSS.n2442 DVSS.n1781 36.1417
R22254 DVSS.n2446 DVSS.n1781 36.1417
R22255 DVSS.n2446 DVSS.n1775 36.1417
R22256 DVSS.n2470 DVSS.n1775 36.1417
R22257 DVSS.n2470 DVSS.n1776 36.1417
R22258 DVSS.n2464 DVSS.n1776 36.1417
R22259 DVSS.n2464 DVSS.n2451 36.1417
R22260 DVSS.n2458 DVSS.n2451 36.1417
R22261 DVSS.n2458 DVSS.n1768 36.1417
R22262 DVSS.n2478 DVSS.n1768 36.1417
R22263 DVSS.n2478 DVSS.n1765 36.1417
R22264 DVSS.n2485 DVSS.n1765 36.1417
R22265 DVSS.n2485 DVSS.n1763 36.1417
R22266 DVSS.n2495 DVSS.n1763 36.1417
R22267 DVSS.n2495 DVSS.n1760 36.1417
R22268 DVSS.n2502 DVSS.n1760 36.1417
R22269 DVSS.n2502 DVSS.n1757 36.1417
R22270 DVSS.n2513 DVSS.n1757 36.1417
R22271 DVSS.n2513 DVSS.n1758 36.1417
R22272 DVSS.n667 DVSS.n664 36.1417
R22273 DVSS.n2812 DVSS.n667 36.1417
R22274 DVSS.n2812 DVSS.n2811 36.1417
R22275 DVSS.n2811 DVSS.n674 36.1417
R22276 DVSS.n2807 DVSS.n674 36.1417
R22277 DVSS.n2807 DVSS.n676 36.1417
R22278 DVSS.n2801 DVSS.n676 36.1417
R22279 DVSS.n2801 DVSS.n682 36.1417
R22280 DVSS.n2797 DVSS.n682 36.1417
R22281 DVSS.n2797 DVSS.n684 36.1417
R22282 DVSS.n2790 DVSS.n684 36.1417
R22283 DVSS.n2790 DVSS.n688 36.1417
R22284 DVSS.n696 DVSS.n688 36.1417
R22285 DVSS.n2782 DVSS.n696 36.1417
R22286 DVSS.n2782 DVSS.n697 36.1417
R22287 DVSS.n2776 DVSS.n697 36.1417
R22288 DVSS.n2776 DVSS.n2775 36.1417
R22289 DVSS.n2775 DVSS.n704 36.1417
R22290 DVSS.n3085 DVSS.n4 36.1417
R22291 DVSS.n3085 DVSS.n6 36.1417
R22292 DVSS.n3079 DVSS.n6 36.1417
R22293 DVSS.n3079 DVSS.n11 36.1417
R22294 DVSS.n2917 DVSS.n2913 36.1417
R22295 DVSS.n2917 DVSS.n2911 36.1417
R22296 DVSS.n2923 DVSS.n2911 36.1417
R22297 DVSS.n2923 DVSS.n2909 36.1417
R22298 DVSS.n2930 DVSS.n2909 36.1417
R22299 DVSS.n2930 DVSS.n2907 36.1417
R22300 DVSS.n2936 DVSS.n2907 36.1417
R22301 DVSS.n2936 DVSS.n2905 36.1417
R22302 DVSS.n2943 DVSS.n2905 36.1417
R22303 DVSS.n2943 DVSS.n2903 36.1417
R22304 DVSS.n2949 DVSS.n2903 36.1417
R22305 DVSS.n2949 DVSS.n2901 36.1417
R22306 DVSS.n2957 DVSS.n2901 36.1417
R22307 DVSS.n2957 DVSS.n2899 36.1417
R22308 DVSS.n2962 DVSS.n2899 36.1417
R22309 DVSS.n2517 DVSS.n1271 35.604
R22310 DVSS.n605 DVSS.n604 35.3887
R22311 DVSS.n356 DVSS.n354 35.3887
R22312 DVSS.n380 DVSS.n367 35.3887
R22313 DVSS.n354 DVSS.n258 35.3887
R22314 DVSS.n360 DVSS.n253 35.3887
R22315 DVSS.n348 DVSS.n253 35.3887
R22316 DVSS.n2229 DVSS.n2227 35.3887
R22317 DVSS.n2253 DVSS.n2240 35.3887
R22318 DVSS.n2227 DVSS.n2131 35.3887
R22319 DVSS.n2233 DVSS.n2126 35.3887
R22320 DVSS.n2221 DVSS.n2126 35.3887
R22321 DVSS.n2830 DVSS.n655 35.3887
R22322 DVSS.n1037 DVSS.n1035 35.3887
R22323 DVSS.n1061 DVSS.n1048 35.3887
R22324 DVSS.n1035 DVSS.n939 35.3887
R22325 DVSS.n1041 DVSS.n934 35.3887
R22326 DVSS.n1029 DVSS.n934 35.3887
R22327 DVSS.n2606 DVSS.n2605 35.3887
R22328 DVSS.n2509 DVSS.n1758 35.3887
R22329 DVSS.n1559 DVSS.n1557 35.3887
R22330 DVSS.n1583 DVSS.n1570 35.3887
R22331 DVSS.n1557 DVSS.n1461 35.3887
R22332 DVSS.n1563 DVSS.n1456 35.3887
R22333 DVSS.n1551 DVSS.n1456 35.3887
R22334 DVSS.n2953 DVSS.t170 35.0689
R22335 DVSS.n2896 DVSS.t59 35.0689
R22336 DVSS.n3015 DVSS.n59 35.0123
R22337 DVSS.n1942 DVSS.n1941 35.0123
R22338 DVSS.n2710 DVSS.n751 35.0123
R22339 DVSS.n2771 DVSS.n704 35.0123
R22340 DVSS.n499 DVSS.n92 34.1338
R22341 DVSS.n125 DVSS.n111 34.1338
R22342 DVSS.n2372 DVSS.n1965 34.1338
R22343 DVSS.n1998 DVSS.n1984 34.1338
R22344 DVSS.n1180 DVSS.n773 34.1338
R22345 DVSS.n806 DVSS.n792 34.1338
R22346 DVSS.n1702 DVSS.n1295 34.1338
R22347 DVSS.n1328 DVSS.n1314 34.1338
R22348 DVSS.n2559 DVSS.n2557 33.5205
R22349 DVSS.n2552 DVSS.n1257 33.5205
R22350 DVSS.n3046 DVSS.n30 33.5205
R22351 DVSS.n562 DVSS.n561 33.5205
R22352 DVSS.n2632 DVSS.n2631 33.5205
R22353 DVSS.n3031 DVSS.n3030 33.5205
R22354 DVSS.n1771 DVSS.n1770 33.5205
R22355 DVSS.n2473 DVSS.n1772 33.5205
R22356 DVSS.n1815 DVSS.n1814 33.5205
R22357 DVSS.n1855 DVSS.n1816 33.5205
R22358 DVSS.n1798 DVSS.n1797 33.5205
R22359 DVSS.n1931 DVSS.n1800 33.5205
R22360 DVSS.n2737 DVSS.n737 33.5205
R22361 DVSS.n2725 DVSS.n2724 33.5205
R22362 DVSS.n693 DVSS.n692 33.5205
R22363 DVSS.n2786 DVSS.n2785 33.5205
R22364 DVSS.n2523 DVSS.n14 32.3755
R22365 DVSS.n75 DVSS.n63 30.8711
R22366 DVSS.n1948 DVSS.n1791 30.8711
R22367 DVSS.n2706 DVSS.n755 30.8711
R22368 DVSS.n711 DVSS.n708 30.8711
R22369 DVSS.n2940 DVSS.n2939 30.5709
R22370 DVSS.n613 DVSS.n69 30.4946
R22371 DVSS.n2825 DVSS.n2824 30.4946
R22372 DVSS.n2695 DVSS.n2694 30.4946
R22373 DVSS.n2520 DVSS.n1748 30.4946
R22374 DVSS.n380 DVSS.n379 29.7417
R22375 DVSS.n2253 DVSS.n2252 29.7417
R22376 DVSS.n1061 DVSS.n1060 29.7417
R22377 DVSS.n1583 DVSS.n1582 29.7417
R22378 DVSS.n216 DVSS.n205 29.4833
R22379 DVSS.n195 DVSS.n184 29.4833
R22380 DVSS.n2089 DVSS.n2078 29.4833
R22381 DVSS.n2068 DVSS.n2057 29.4833
R22382 DVSS.n897 DVSS.n886 29.4833
R22383 DVSS.n876 DVSS.n865 29.4833
R22384 DVSS.n1419 DVSS.n1408 29.4833
R22385 DVSS.n1398 DVSS.n1387 29.4833
R22386 DVSS.n165 DVSS.n148 29.1989
R22387 DVSS.n522 DVSS.n501 29.1989
R22388 DVSS.n2038 DVSS.n2021 29.1989
R22389 DVSS.n2395 DVSS.n2374 29.1989
R22390 DVSS.n846 DVSS.n829 29.1989
R22391 DVSS.n1203 DVSS.n1182 29.1989
R22392 DVSS.n1368 DVSS.n1351 29.1989
R22393 DVSS.n1725 DVSS.n1704 29.1989
R22394 DVSS.n1839 DVSS.n1838 29.0014
R22395 DVSS.n1927 DVSS.n1926 28.2515
R22396 DVSS.n3024 DVSS.n53 28.2515
R22397 DVSS.n2614 DVSS.t77 28.1205
R22398 DVSS.n1883 DVSS.t87 28.1205
R22399 DVSS.n720 DVSS.t38 28.1205
R22400 DVSS.n670 DVSS.t57 28.1205
R22401 DVSS DVSS.n3089 26.5398
R22402 DVSS.n356 DVSS.n355 25.6005
R22403 DVSS.n355 DVSS.n250 25.6005
R22404 DVSS.n367 DVSS.n250 25.6005
R22405 DVSS.n342 DVSS.n340 25.6005
R22406 DVSS.n342 DVSS.n341 25.6005
R22407 DVSS.n341 DVSS.n258 25.6005
R22408 DVSS.n379 DVSS.n378 25.6005
R22409 DVSS.n361 DVSS.n360 25.6005
R22410 DVSS.n362 DVSS.n361 25.6005
R22411 DVSS.n362 DVSS.n224 25.6005
R22412 DVSS.n346 DVSS.n312 25.6005
R22413 DVSS.n347 DVSS.n346 25.6005
R22414 DVSS.n348 DVSS.n347 25.6005
R22415 DVSS.n2229 DVSS.n2228 25.6005
R22416 DVSS.n2228 DVSS.n2123 25.6005
R22417 DVSS.n2240 DVSS.n2123 25.6005
R22418 DVSS.n2215 DVSS.n2213 25.6005
R22419 DVSS.n2215 DVSS.n2214 25.6005
R22420 DVSS.n2214 DVSS.n2131 25.6005
R22421 DVSS.n2252 DVSS.n2251 25.6005
R22422 DVSS.n2234 DVSS.n2233 25.6005
R22423 DVSS.n2235 DVSS.n2234 25.6005
R22424 DVSS.n2235 DVSS.n2097 25.6005
R22425 DVSS.n2219 DVSS.n2185 25.6005
R22426 DVSS.n2220 DVSS.n2219 25.6005
R22427 DVSS.n2221 DVSS.n2220 25.6005
R22428 DVSS.n1037 DVSS.n1036 25.6005
R22429 DVSS.n1036 DVSS.n931 25.6005
R22430 DVSS.n1048 DVSS.n931 25.6005
R22431 DVSS.n1023 DVSS.n1021 25.6005
R22432 DVSS.n1023 DVSS.n1022 25.6005
R22433 DVSS.n1022 DVSS.n939 25.6005
R22434 DVSS.n1060 DVSS.n1059 25.6005
R22435 DVSS.n1042 DVSS.n1041 25.6005
R22436 DVSS.n1043 DVSS.n1042 25.6005
R22437 DVSS.n1043 DVSS.n905 25.6005
R22438 DVSS.n1027 DVSS.n993 25.6005
R22439 DVSS.n1028 DVSS.n1027 25.6005
R22440 DVSS.n1029 DVSS.n1028 25.6005
R22441 DVSS.n1559 DVSS.n1558 25.6005
R22442 DVSS.n1558 DVSS.n1453 25.6005
R22443 DVSS.n1570 DVSS.n1453 25.6005
R22444 DVSS.n1545 DVSS.n1543 25.6005
R22445 DVSS.n1545 DVSS.n1544 25.6005
R22446 DVSS.n1544 DVSS.n1461 25.6005
R22447 DVSS.n1582 DVSS.n1581 25.6005
R22448 DVSS.n1564 DVSS.n1563 25.6005
R22449 DVSS.n1565 DVSS.n1564 25.6005
R22450 DVSS.n1565 DVSS.n1427 25.6005
R22451 DVSS.n1549 DVSS.n1515 25.6005
R22452 DVSS.n1550 DVSS.n1549 25.6005
R22453 DVSS.n1551 DVSS.n1550 25.6005
R22454 DVSS.n475 DVSS.n92 22.3184
R22455 DVSS.n476 DVSS.n475 22.3184
R22456 DVSS.n477 DVSS.n476 22.3184
R22457 DVSS.n477 DVSS.n470 22.3184
R22458 DVSS.n482 DVSS.n470 22.3184
R22459 DVSS.n483 DVSS.n482 22.3184
R22460 DVSS.n483 DVSS.n468 22.3184
R22461 DVSS.n488 DVSS.n468 22.3184
R22462 DVSS.n125 DVSS.n124 22.3184
R22463 DVSS.n130 DVSS.n124 22.3184
R22464 DVSS.n131 DVSS.n130 22.3184
R22465 DVSS.n131 DVSS.n122 22.3184
R22466 DVSS.n137 DVSS.n122 22.3184
R22467 DVSS.n138 DVSS.n137 22.3184
R22468 DVSS.n138 DVSS.n120 22.3184
R22469 DVSS.n143 DVSS.n120 22.3184
R22470 DVSS.n2348 DVSS.n1965 22.3184
R22471 DVSS.n2349 DVSS.n2348 22.3184
R22472 DVSS.n2350 DVSS.n2349 22.3184
R22473 DVSS.n2350 DVSS.n2343 22.3184
R22474 DVSS.n2355 DVSS.n2343 22.3184
R22475 DVSS.n2356 DVSS.n2355 22.3184
R22476 DVSS.n2356 DVSS.n2341 22.3184
R22477 DVSS.n2361 DVSS.n2341 22.3184
R22478 DVSS.n1998 DVSS.n1997 22.3184
R22479 DVSS.n2003 DVSS.n1997 22.3184
R22480 DVSS.n2004 DVSS.n2003 22.3184
R22481 DVSS.n2004 DVSS.n1995 22.3184
R22482 DVSS.n2010 DVSS.n1995 22.3184
R22483 DVSS.n2011 DVSS.n2010 22.3184
R22484 DVSS.n2011 DVSS.n1993 22.3184
R22485 DVSS.n2016 DVSS.n1993 22.3184
R22486 DVSS.n1156 DVSS.n773 22.3184
R22487 DVSS.n1157 DVSS.n1156 22.3184
R22488 DVSS.n1158 DVSS.n1157 22.3184
R22489 DVSS.n1158 DVSS.n1151 22.3184
R22490 DVSS.n1163 DVSS.n1151 22.3184
R22491 DVSS.n1164 DVSS.n1163 22.3184
R22492 DVSS.n1164 DVSS.n1149 22.3184
R22493 DVSS.n1169 DVSS.n1149 22.3184
R22494 DVSS.n806 DVSS.n805 22.3184
R22495 DVSS.n811 DVSS.n805 22.3184
R22496 DVSS.n812 DVSS.n811 22.3184
R22497 DVSS.n812 DVSS.n803 22.3184
R22498 DVSS.n818 DVSS.n803 22.3184
R22499 DVSS.n819 DVSS.n818 22.3184
R22500 DVSS.n819 DVSS.n801 22.3184
R22501 DVSS.n824 DVSS.n801 22.3184
R22502 DVSS.n1678 DVSS.n1295 22.3184
R22503 DVSS.n1679 DVSS.n1678 22.3184
R22504 DVSS.n1680 DVSS.n1679 22.3184
R22505 DVSS.n1680 DVSS.n1673 22.3184
R22506 DVSS.n1685 DVSS.n1673 22.3184
R22507 DVSS.n1686 DVSS.n1685 22.3184
R22508 DVSS.n1686 DVSS.n1671 22.3184
R22509 DVSS.n1691 DVSS.n1671 22.3184
R22510 DVSS.n1328 DVSS.n1327 22.3184
R22511 DVSS.n1333 DVSS.n1327 22.3184
R22512 DVSS.n1334 DVSS.n1333 22.3184
R22513 DVSS.n1334 DVSS.n1325 22.3184
R22514 DVSS.n1340 DVSS.n1325 22.3184
R22515 DVSS.n1341 DVSS.n1340 22.3184
R22516 DVSS.n1341 DVSS.n1323 22.3184
R22517 DVSS.n1346 DVSS.n1323 22.3184
R22518 DVSS.n2953 DVSS.t32 22.2377
R22519 DVSS.n2896 DVSS.t171 22.2377
R22520 DVSS.n2979 DVSS.t167 21.2805
R22521 DVSS.n2979 DVSS.t168 21.2805
R22522 DVSS.n2614 DVSS.t93 21.2805
R22523 DVSS.n1883 DVSS.t177 21.2805
R22524 DVSS.n720 DVSS.t89 21.2805
R22525 DVSS.n670 DVSS.t141 21.2805
R22526 DVSS.n2456 DVSS.t96 20.7552
R22527 DVSS.t146 DVSS.n38 20.6994
R22528 DVSS.t181 DVSS.n1249 20.4114
R22529 DVSS.n489 DVSS.n488 20.3492
R22530 DVSS.n144 DVSS.n143 20.3492
R22531 DVSS.n2362 DVSS.n2361 20.3492
R22532 DVSS.n2017 DVSS.n2016 20.3492
R22533 DVSS.n1170 DVSS.n1169 20.3492
R22534 DVSS.n825 DVSS.n824 20.3492
R22535 DVSS.n1692 DVSS.n1691 20.3492
R22536 DVSS.n1347 DVSS.n1346 20.3492
R22537 DVSS.n2588 DVSS.t105 20.0005
R22538 DVSS.n2588 DVSS.t83 20.0005
R22539 DVSS.n586 DVSS.t137 20.0005
R22540 DVSS.n586 DVSS.t61 20.0005
R22541 DVSS.n2489 DVSS.t29 20.0005
R22542 DVSS.n2489 DVSS.t159 20.0005
R22543 DVSS.n647 DVSS.t125 20.0005
R22544 DVSS.n647 DVSS.t79 20.0005
R22545 DVSS.n2442 DVSS.n2441 18.0103
R22546 DVSS.n2707 DVSS.n2706 18.0103
R22547 DVSS.n2673 DVSS.n2672 18.0103
R22548 DVSS.n2965 DVSS.n2874 18.0093
R22549 DVSS.n1829 DVSS.n1828 18.0093
R22550 DVSS.n2520 DVSS.n2519 18.0093
R22551 DVSS.n2962 DVSS.n2961 18.007
R22552 DVSS.n3005 DVSS.n3004 17.2422
R22553 DVSS.n2591 DVSS.n2590 17.1722
R22554 DVSS.n2590 DVSS.n2587 17.1722
R22555 DVSS.n589 DVSS.n588 17.1722
R22556 DVSS.n588 DVSS.n585 17.1722
R22557 DVSS.n2492 DVSS.n2491 17.1722
R22558 DVSS.n2491 DVSS.n2488 17.1722
R22559 DVSS.n650 DVSS.n649 17.1722
R22560 DVSS.n649 DVSS.n639 17.1722
R22561 DVSS.t70 DVSS.n2867 17.1497
R22562 DVSS.n499 DVSS.n498 17.0218
R22563 DVSS.n2372 DVSS.n2371 17.0218
R22564 DVSS.n1180 DVSS.n1179 17.0218
R22565 DVSS.n1702 DVSS.n1701 17.0218
R22566 DVSS.n450 DVSS.n111 16.8856
R22567 DVSS.n2323 DVSS.n1984 16.8856
R22568 DVSS.n1131 DVSS.n792 16.8856
R22569 DVSS.n1653 DVSS.n1314 16.8856
R22570 DVSS.n2469 DVSS.n2468 15.5836
R22571 DVSS.n36 DVSS.n34 15.5501
R22572 DVSS.n432 DVSS.n111 15.5239
R22573 DVSS.n2305 DVSS.n1984 15.5239
R22574 DVSS.n1113 DVSS.n792 15.5239
R22575 DVSS.n1635 DVSS.n1314 15.5239
R22576 DVSS.n214 DVSS.n213 15.463
R22577 DVSS.n193 DVSS.n192 15.463
R22578 DVSS.n2087 DVSS.n2086 15.463
R22579 DVSS.n2066 DVSS.n2065 15.463
R22580 DVSS.n895 DVSS.n894 15.463
R22581 DVSS.n874 DVSS.n873 15.463
R22582 DVSS.n1417 DVSS.n1416 15.463
R22583 DVSS.n1396 DVSS.n1395 15.463
R22584 DVSS.n500 DVSS.n499 15.3877
R22585 DVSS.n2373 DVSS.n2372 15.3877
R22586 DVSS.n1181 DVSS.n1180 15.3877
R22587 DVSS.n1703 DVSS.n1702 15.3877
R22588 DVSS.n1253 DVSS.n1252 15.3783
R22589 DVSS.n3058 DVSS 15.0005
R22590 DVSS.t102 DVSS.n2449 14.8253
R22591 DVSS.t154 DVSS.n23 14.7854
R22592 DVSS.n2547 DVSS.t187 14.5797
R22593 DVSS.n2941 DVSS.n2940 14.4554
R22594 DVSS.n2981 DVSS.n2980 14.4288
R22595 DVSS.n219 DVSS.n206 13.5534
R22596 DVSS.n214 DVSS.n210 13.5534
R22597 DVSS.n198 DVSS.n185 13.5534
R22598 DVSS.n193 DVSS.n189 13.5534
R22599 DVSS.n2092 DVSS.n2079 13.5534
R22600 DVSS.n2087 DVSS.n2083 13.5534
R22601 DVSS.n2071 DVSS.n2058 13.5534
R22602 DVSS.n2066 DVSS.n2062 13.5534
R22603 DVSS.n900 DVSS.n887 13.5534
R22604 DVSS.n895 DVSS.n891 13.5534
R22605 DVSS.n879 DVSS.n866 13.5534
R22606 DVSS.n874 DVSS.n870 13.5534
R22607 DVSS.n1422 DVSS.n1409 13.5534
R22608 DVSS.n1417 DVSS.n1413 13.5534
R22609 DVSS.n1401 DVSS.n1388 13.5534
R22610 DVSS.n1396 DVSS.n1392 13.5534
R22611 DVSS.n2660 DVSS.n2659 12.8977
R22612 DVSS.n1881 DVSS.n1880 12.8977
R22613 DVSS.n717 DVSS.n714 12.8977
R22614 DVSS.n2818 DVSS.n662 12.8977
R22615 DVSS.n2915 DVSS.n2914 12.8862
R22616 DVSS.n2454 DVSS.n2450 12.036
R22617 DVSS.n3039 DVSS.n37 12.021
R22618 DVSS.n2566 DVSS.n1250 11.944
R22619 DVSS.n1257 DVSS.t188 10.6405
R22620 DVSS.n1257 DVSS.t186 10.6405
R22621 DVSS.n2557 DVSS.t184 10.6405
R22622 DVSS.n2557 DVSS.t182 10.6405
R22623 DVSS.n30 DVSS.t155 10.6405
R22624 DVSS.n30 DVSS.t153 10.6405
R22625 DVSS.n561 DVSS.t151 10.6405
R22626 DVSS.n561 DVSS.t147 10.6405
R22627 DVSS.n2631 DVSS.t139 10.6405
R22628 DVSS.n2631 DVSS.t131 10.6405
R22629 DVSS.n3030 DVSS.t135 10.6405
R22630 DVSS.n3030 DVSS.t129 10.6405
R22631 DVSS.n1772 DVSS.t103 10.6405
R22632 DVSS.n1772 DVSS.t101 10.6405
R22633 DVSS.n1770 DVSS.t99 10.6405
R22634 DVSS.n1770 DVSS.t97 10.6405
R22635 DVSS.n1816 DVSS.t50 10.6405
R22636 DVSS.n1816 DVSS.t48 10.6405
R22637 DVSS.n1814 DVSS.t46 10.6405
R22638 DVSS.n1814 DVSS.t52 10.6405
R22639 DVSS.n1797 DVSS.t123 10.6405
R22640 DVSS.n1797 DVSS.t121 10.6405
R22641 DVSS.n1800 DVSS.t119 10.6405
R22642 DVSS.n1800 DVSS.t117 10.6405
R22643 DVSS.n737 DVSS.t115 10.6405
R22644 DVSS.n737 DVSS.t113 10.6405
R22645 DVSS.n2724 DVSS.t109 10.6405
R22646 DVSS.n2724 DVSS.t111 10.6405
R22647 DVSS.n692 DVSS.t27 10.6405
R22648 DVSS.n692 DVSS.t25 10.6405
R22649 DVSS.n2785 DVSS.t19 10.6405
R22650 DVSS.n2785 DVSS.t23 10.6405
R22651 DVSS.n369 DVSS.n246 10.4252
R22652 DVSS.n2242 DVSS.n2119 10.4252
R22653 DVSS.n1050 DVSS.n927 10.4252
R22654 DVSS.n1572 DVSS.n1449 10.4252
R22655 DVSS.n539 DVSS.n538 9.31763
R22656 DVSS.n2412 DVSS.n2411 9.31763
R22657 DVSS.n1220 DVSS.n1219 9.31763
R22658 DVSS.n1742 DVSS.n1741 9.31763
R22659 DVSS.n3016 DVSS.n3015 9.3005
R22660 DVSS.n204 DVSS.n203 9.3005
R22661 DVSS.n211 DVSS.n207 9.3005
R22662 DVSS.n212 DVSS.n210 9.3005
R22663 DVSS.n217 DVSS.n209 9.3005
R22664 DVSS.n217 DVSS.n216 9.3005
R22665 DVSS.n208 DVSS.n206 9.3005
R22666 DVSS.n222 DVSS.n221 9.3005
R22667 DVSS.n183 DVSS.n182 9.3005
R22668 DVSS.n190 DVSS.n186 9.3005
R22669 DVSS.n191 DVSS.n189 9.3005
R22670 DVSS.n196 DVSS.n188 9.3005
R22671 DVSS.n196 DVSS.n195 9.3005
R22672 DVSS.n187 DVSS.n185 9.3005
R22673 DVSS.n201 DVSS.n200 9.3005
R22674 DVSS.n417 DVSS.n416 9.3005
R22675 DVSS.n420 DVSS.n419 9.3005
R22676 DVSS.n421 DVSS.n152 9.3005
R22677 DVSS.n426 DVSS.n425 9.3005
R22678 DVSS.n424 DVSS.n153 9.3005
R22679 DVSS.n423 DVSS.n422 9.3005
R22680 DVSS.n119 DVSS.n118 9.3005
R22681 DVSS.n437 DVSS.n436 9.3005
R22682 DVSS.n438 DVSS.n116 9.3005
R22683 DVSS.n446 DVSS.n445 9.3005
R22684 DVSS.n444 DVSS.n117 9.3005
R22685 DVSS.n441 DVSS.n440 9.3005
R22686 DVSS.n439 DVSS.n105 9.3005
R22687 DVSS.n457 DVSS.n104 9.3005
R22688 DVSS.n459 DVSS.n458 9.3005
R22689 DVSS.n460 DVSS.n103 9.3005
R22690 DVSS.n463 DVSS.n102 9.3005
R22691 DVSS.n465 DVSS.n464 9.3005
R22692 DVSS.n466 DVSS.n100 9.3005
R22693 DVSS.n494 DVSS.n493 9.3005
R22694 DVSS.n492 DVSS.n101 9.3005
R22695 DVSS.n491 DVSS.n490 9.3005
R22696 DVSS.n467 DVSS.n85 9.3005
R22697 DVSS.n528 DVSS.n86 9.3005
R22698 DVSS.n529 DVSS.n84 9.3005
R22699 DVSS.n531 DVSS.n530 9.3005
R22700 DVSS.n532 DVSS.n83 9.3005
R22701 DVSS.n534 DVSS.n533 9.3005
R22702 DVSS.n605 DVSS.n544 9.3005
R22703 DVSS.n607 DVSS.n606 9.3005
R22704 DVSS.n2077 DVSS.n2076 9.3005
R22705 DVSS.n2084 DVSS.n2080 9.3005
R22706 DVSS.n2085 DVSS.n2083 9.3005
R22707 DVSS.n2090 DVSS.n2082 9.3005
R22708 DVSS.n2090 DVSS.n2089 9.3005
R22709 DVSS.n2081 DVSS.n2079 9.3005
R22710 DVSS.n2095 DVSS.n2094 9.3005
R22711 DVSS.n2056 DVSS.n2055 9.3005
R22712 DVSS.n2063 DVSS.n2059 9.3005
R22713 DVSS.n2064 DVSS.n2062 9.3005
R22714 DVSS.n2069 DVSS.n2061 9.3005
R22715 DVSS.n2069 DVSS.n2068 9.3005
R22716 DVSS.n2060 DVSS.n2058 9.3005
R22717 DVSS.n2074 DVSS.n2073 9.3005
R22718 DVSS.n2290 DVSS.n2289 9.3005
R22719 DVSS.n2293 DVSS.n2292 9.3005
R22720 DVSS.n2294 DVSS.n2025 9.3005
R22721 DVSS.n2299 DVSS.n2298 9.3005
R22722 DVSS.n2297 DVSS.n2026 9.3005
R22723 DVSS.n2296 DVSS.n2295 9.3005
R22724 DVSS.n1992 DVSS.n1991 9.3005
R22725 DVSS.n2310 DVSS.n2309 9.3005
R22726 DVSS.n2311 DVSS.n1989 9.3005
R22727 DVSS.n2319 DVSS.n2318 9.3005
R22728 DVSS.n2317 DVSS.n1990 9.3005
R22729 DVSS.n2314 DVSS.n2313 9.3005
R22730 DVSS.n2312 DVSS.n1978 9.3005
R22731 DVSS.n2330 DVSS.n1977 9.3005
R22732 DVSS.n2332 DVSS.n2331 9.3005
R22733 DVSS.n2333 DVSS.n1976 9.3005
R22734 DVSS.n2336 DVSS.n1975 9.3005
R22735 DVSS.n2338 DVSS.n2337 9.3005
R22736 DVSS.n2339 DVSS.n1973 9.3005
R22737 DVSS.n2367 DVSS.n2366 9.3005
R22738 DVSS.n2365 DVSS.n1974 9.3005
R22739 DVSS.n2364 DVSS.n2363 9.3005
R22740 DVSS.n2340 DVSS.n1958 9.3005
R22741 DVSS.n2401 DVSS.n1959 9.3005
R22742 DVSS.n2402 DVSS.n1957 9.3005
R22743 DVSS.n2404 DVSS.n2403 9.3005
R22744 DVSS.n2405 DVSS.n1956 9.3005
R22745 DVSS.n2407 DVSS.n2406 9.3005
R22746 DVSS.n1941 DVSS.n1940 9.3005
R22747 DVSS.n885 DVSS.n884 9.3005
R22748 DVSS.n892 DVSS.n888 9.3005
R22749 DVSS.n893 DVSS.n891 9.3005
R22750 DVSS.n898 DVSS.n890 9.3005
R22751 DVSS.n898 DVSS.n897 9.3005
R22752 DVSS.n889 DVSS.n887 9.3005
R22753 DVSS.n903 DVSS.n902 9.3005
R22754 DVSS.n864 DVSS.n863 9.3005
R22755 DVSS.n871 DVSS.n867 9.3005
R22756 DVSS.n872 DVSS.n870 9.3005
R22757 DVSS.n877 DVSS.n869 9.3005
R22758 DVSS.n877 DVSS.n876 9.3005
R22759 DVSS.n868 DVSS.n866 9.3005
R22760 DVSS.n882 DVSS.n881 9.3005
R22761 DVSS.n1098 DVSS.n1097 9.3005
R22762 DVSS.n1101 DVSS.n1100 9.3005
R22763 DVSS.n1102 DVSS.n833 9.3005
R22764 DVSS.n1107 DVSS.n1106 9.3005
R22765 DVSS.n1105 DVSS.n834 9.3005
R22766 DVSS.n1104 DVSS.n1103 9.3005
R22767 DVSS.n800 DVSS.n799 9.3005
R22768 DVSS.n1118 DVSS.n1117 9.3005
R22769 DVSS.n1119 DVSS.n797 9.3005
R22770 DVSS.n1127 DVSS.n1126 9.3005
R22771 DVSS.n1125 DVSS.n798 9.3005
R22772 DVSS.n1122 DVSS.n1121 9.3005
R22773 DVSS.n1120 DVSS.n786 9.3005
R22774 DVSS.n1138 DVSS.n785 9.3005
R22775 DVSS.n1140 DVSS.n1139 9.3005
R22776 DVSS.n1141 DVSS.n784 9.3005
R22777 DVSS.n1144 DVSS.n783 9.3005
R22778 DVSS.n1146 DVSS.n1145 9.3005
R22779 DVSS.n1147 DVSS.n781 9.3005
R22780 DVSS.n1175 DVSS.n1174 9.3005
R22781 DVSS.n1173 DVSS.n782 9.3005
R22782 DVSS.n1172 DVSS.n1171 9.3005
R22783 DVSS.n1148 DVSS.n766 9.3005
R22784 DVSS.n1209 DVSS.n767 9.3005
R22785 DVSS.n1210 DVSS.n765 9.3005
R22786 DVSS.n1212 DVSS.n1211 9.3005
R22787 DVSS.n1213 DVSS.n764 9.3005
R22788 DVSS.n1215 DVSS.n1214 9.3005
R22789 DVSS.n2711 DVSS.n2710 9.3005
R22790 DVSS.n1407 DVSS.n1406 9.3005
R22791 DVSS.n1414 DVSS.n1410 9.3005
R22792 DVSS.n1415 DVSS.n1413 9.3005
R22793 DVSS.n1420 DVSS.n1412 9.3005
R22794 DVSS.n1420 DVSS.n1419 9.3005
R22795 DVSS.n1411 DVSS.n1409 9.3005
R22796 DVSS.n1425 DVSS.n1424 9.3005
R22797 DVSS.n1386 DVSS.n1385 9.3005
R22798 DVSS.n1393 DVSS.n1389 9.3005
R22799 DVSS.n1394 DVSS.n1392 9.3005
R22800 DVSS.n1399 DVSS.n1391 9.3005
R22801 DVSS.n1399 DVSS.n1398 9.3005
R22802 DVSS.n1390 DVSS.n1388 9.3005
R22803 DVSS.n1404 DVSS.n1403 9.3005
R22804 DVSS.n1620 DVSS.n1619 9.3005
R22805 DVSS.n1623 DVSS.n1622 9.3005
R22806 DVSS.n1624 DVSS.n1355 9.3005
R22807 DVSS.n1629 DVSS.n1628 9.3005
R22808 DVSS.n1627 DVSS.n1356 9.3005
R22809 DVSS.n1626 DVSS.n1625 9.3005
R22810 DVSS.n1322 DVSS.n1321 9.3005
R22811 DVSS.n1640 DVSS.n1639 9.3005
R22812 DVSS.n1641 DVSS.n1319 9.3005
R22813 DVSS.n1649 DVSS.n1648 9.3005
R22814 DVSS.n1647 DVSS.n1320 9.3005
R22815 DVSS.n1644 DVSS.n1643 9.3005
R22816 DVSS.n1642 DVSS.n1308 9.3005
R22817 DVSS.n1660 DVSS.n1307 9.3005
R22818 DVSS.n1662 DVSS.n1661 9.3005
R22819 DVSS.n1663 DVSS.n1306 9.3005
R22820 DVSS.n1666 DVSS.n1305 9.3005
R22821 DVSS.n1668 DVSS.n1667 9.3005
R22822 DVSS.n1669 DVSS.n1303 9.3005
R22823 DVSS.n1697 DVSS.n1696 9.3005
R22824 DVSS.n1695 DVSS.n1304 9.3005
R22825 DVSS.n1694 DVSS.n1693 9.3005
R22826 DVSS.n1670 DVSS.n1288 9.3005
R22827 DVSS.n1731 DVSS.n1289 9.3005
R22828 DVSS.n1732 DVSS.n1287 9.3005
R22829 DVSS.n1734 DVSS.n1733 9.3005
R22830 DVSS.n1735 DVSS.n1286 9.3005
R22831 DVSS.n1737 DVSS.n1736 9.3005
R22832 DVSS.n2770 DVSS.n707 9.3005
R22833 DVSS.n2772 DVSS.n2771 9.3005
R22834 DVSS.n1939 DVSS.n1937 9.3005
R22835 DVSS.n2828 DVSS.n655 9.3005
R22836 DVSS.n2827 DVSS.n2826 9.3005
R22837 DVSS.n2510 DVSS.n2509 9.3005
R22838 DVSS.n2508 DVSS.n2507 9.3005
R22839 DVSS.n2605 DVSS.n2604 9.3005
R22840 DVSS.n1225 DVSS.n1224 9.3005
R22841 DVSS.n2709 DVSS.n754 9.3005
R22842 DVSS.n3014 DVSS.n62 9.3005
R22843 DVSS.n430 DVSS.n148 9.26007
R22844 DVSS.n431 DVSS.n430 9.26007
R22845 DVSS.n432 DVSS.n431 9.26007
R22846 DVSS.n451 DVSS.n450 9.26007
R22847 DVSS.n453 DVSS.n451 9.26007
R22848 DVSS.n453 DVSS.n452 9.26007
R22849 DVSS.n452 DVSS.n93 9.26007
R22850 DVSS.n498 DVSS.n93 9.26007
R22851 DVSS.n524 DVSS.n500 9.26007
R22852 DVSS.n524 DVSS.n523 9.26007
R22853 DVSS.n523 DVSS.n522 9.26007
R22854 DVSS.n2303 DVSS.n2021 9.26007
R22855 DVSS.n2304 DVSS.n2303 9.26007
R22856 DVSS.n2305 DVSS.n2304 9.26007
R22857 DVSS.n2324 DVSS.n2323 9.26007
R22858 DVSS.n2326 DVSS.n2324 9.26007
R22859 DVSS.n2326 DVSS.n2325 9.26007
R22860 DVSS.n2325 DVSS.n1966 9.26007
R22861 DVSS.n2371 DVSS.n1966 9.26007
R22862 DVSS.n2397 DVSS.n2373 9.26007
R22863 DVSS.n2397 DVSS.n2396 9.26007
R22864 DVSS.n2396 DVSS.n2395 9.26007
R22865 DVSS.n1111 DVSS.n829 9.26007
R22866 DVSS.n1112 DVSS.n1111 9.26007
R22867 DVSS.n1113 DVSS.n1112 9.26007
R22868 DVSS.n1132 DVSS.n1131 9.26007
R22869 DVSS.n1134 DVSS.n1132 9.26007
R22870 DVSS.n1134 DVSS.n1133 9.26007
R22871 DVSS.n1133 DVSS.n774 9.26007
R22872 DVSS.n1179 DVSS.n774 9.26007
R22873 DVSS.n1205 DVSS.n1181 9.26007
R22874 DVSS.n1205 DVSS.n1204 9.26007
R22875 DVSS.n1204 DVSS.n1203 9.26007
R22876 DVSS.n1633 DVSS.n1351 9.26007
R22877 DVSS.n1634 DVSS.n1633 9.26007
R22878 DVSS.n1635 DVSS.n1634 9.26007
R22879 DVSS.n1654 DVSS.n1653 9.26007
R22880 DVSS.n1656 DVSS.n1654 9.26007
R22881 DVSS.n1656 DVSS.n1655 9.26007
R22882 DVSS.n1655 DVSS.n1296 9.26007
R22883 DVSS.n1701 DVSS.n1296 9.26007
R22884 DVSS.n1727 DVSS.n1703 9.26007
R22885 DVSS.n1727 DVSS.n1726 9.26007
R22886 DVSS.n1726 DVSS.n1725 9.26007
R22887 DVSS.n606 DVSS.n68 9.15497
R22888 DVSS.n68 DVSS.n67 9.15497
R22889 DVSS.n2661 DVSS.n2660 9.15497
R22890 DVSS.n2613 DVSS.n2612 9.15497
R22891 DVSS.n2619 DVSS.n2612 9.15497
R22892 DVSS.n2656 DVSS.n2655 9.15497
R22893 DVSS.n2655 DVSS.n2654 9.15497
R22894 DVSS.n2618 DVSS.n2617 9.15497
R22895 DVSS.n2653 DVSS.n2618 9.15497
R22896 DVSS.n2651 DVSS.n2650 9.15497
R22897 DVSS.n2652 DVSS.n2651 9.15497
R22898 DVSS.n2622 DVSS.n2621 9.15497
R22899 DVSS.n2621 DVSS.n2620 9.15497
R22900 DVSS.n2646 DVSS.n2645 9.15497
R22901 DVSS.n2645 DVSS.n2644 9.15497
R22902 DVSS.n2626 DVSS.n2625 9.15497
R22903 DVSS.n2643 DVSS.n2626 9.15497
R22904 DVSS.n2641 DVSS.n2640 9.15497
R22905 DVSS.n2642 DVSS.n2641 9.15497
R22906 DVSS.n614 DVSS.n613 9.15497
R22907 DVSS.n615 DVSS.n614 9.15497
R22908 DVSS.n3057 DVSS.n3056 9.15497
R22909 DVSS.n3056 DVSS.n3055 9.15497
R22910 DVSS.n1880 DVSS.n622 9.15497
R22911 DVSS.n1879 DVSS.n1878 9.15497
R22912 DVSS.n1878 DVSS.n1877 9.15497
R22913 DVSS.n1888 DVSS.n1887 9.15497
R22914 DVSS.n1889 DVSS.n1888 9.15497
R22915 DVSS.n1876 DVSS.n1875 9.15497
R22916 DVSS.n1890 DVSS.n1876 9.15497
R22917 DVSS.n1893 DVSS.n1892 9.15497
R22918 DVSS.n1892 DVSS.n1891 9.15497
R22919 DVSS.n1873 DVSS.n1872 9.15497
R22920 DVSS.n1872 DVSS.n1871 9.15497
R22921 DVSS.n1898 DVSS.n1897 9.15497
R22922 DVSS.n1899 DVSS.n1898 9.15497
R22923 DVSS.n1870 DVSS.n1869 9.15497
R22924 DVSS.n1900 DVSS.n1870 9.15497
R22925 DVSS.n1903 DVSS.n1902 9.15497
R22926 DVSS.n1902 DVSS.n1901 9.15497
R22927 DVSS.n626 DVSS.n623 9.15497
R22928 DVSS.n2868 DVSS.n623 9.15497
R22929 DVSS.n1824 DVSS.n1823 9.15497
R22930 DVSS.n2824 DVSS.n2823 9.15497
R22931 DVSS.n2765 DVSS.n714 9.15497
R22932 DVSS.n2763 DVSS.n2762 9.15497
R22933 DVSS.n2764 DVSS.n2763 9.15497
R22934 DVSS.n2761 DVSS.n716 9.15497
R22935 DVSS.n716 DVSS.n715 9.15497
R22936 DVSS.n724 DVSS.n718 9.15497
R22937 DVSS.n726 DVSS.n724 9.15497
R22938 DVSS.n2756 DVSS.n2755 9.15497
R22939 DVSS.n2755 DVSS.n2754 9.15497
R22940 DVSS.n725 DVSS.n723 9.15497
R22941 DVSS.n2753 DVSS.n725 9.15497
R22942 DVSS.n2751 DVSS.n2750 9.15497
R22943 DVSS.n2752 DVSS.n2751 9.15497
R22944 DVSS.n729 DVSS.n728 9.15497
R22945 DVSS.n728 DVSS.n727 9.15497
R22946 DVSS.n2746 DVSS.n2745 9.15497
R22947 DVSS.n2745 DVSS.n2744 9.15497
R22948 DVSS.n2508 DVSS.n1749 9.15497
R22949 DVSS.n1273 DVSS.n1272 9.15497
R22950 DVSS.n2517 DVSS.n1272 9.15497
R22951 DVSS.n2544 DVSS.n2543 9.15497
R22952 DVSS.n2545 DVSS.n2544 9.15497
R22953 DVSS.n2768 DVSS.n711 9.15497
R22954 DVSS.n2768 DVSS.n2767 9.15497
R22955 DVSS.n709 DVSS.n704 9.15497
R22956 DVSS.n2770 DVSS.n2769 9.15497
R22957 DVSS.n2819 DVSS.n2818 9.15497
R22958 DVSS.n2817 DVSS.n664 9.15497
R22959 DVSS.n2817 DVSS.n2816 9.15497
R22960 DVSS.n667 DVSS.n663 9.15497
R22961 DVSS.n2815 DVSS.n663 9.15497
R22962 DVSS.n2813 DVSS.n2812 9.15497
R22963 DVSS.n2814 DVSS.n2813 9.15497
R22964 DVSS.n2811 DVSS.n666 9.15497
R22965 DVSS.n666 DVSS.n665 9.15497
R22966 DVSS.n677 DVSS.n674 9.15497
R22967 DVSS.n679 DVSS.n677 9.15497
R22968 DVSS.n2807 DVSS.n2806 9.15497
R22969 DVSS.n2806 DVSS.n2805 9.15497
R22970 DVSS.n678 DVSS.n676 9.15497
R22971 DVSS.n2804 DVSS.n678 9.15497
R22972 DVSS.n2802 DVSS.n2801 9.15497
R22973 DVSS.n2803 DVSS.n2802 9.15497
R22974 DVSS.n682 DVSS.n681 9.15497
R22975 DVSS.n681 DVSS.n680 9.15497
R22976 DVSS.n2797 DVSS.n2796 9.15497
R22977 DVSS.n2796 DVSS.n2795 9.15497
R22978 DVSS.n685 DVSS.n684 9.15497
R22979 DVSS.n2793 DVSS.n685 9.15497
R22980 DVSS.n2791 DVSS.n2790 9.15497
R22981 DVSS.n2792 DVSS.n2791 9.15497
R22982 DVSS.n688 DVSS.n687 9.15497
R22983 DVSS.n687 DVSS.n686 9.15497
R22984 DVSS.n698 DVSS.n696 9.15497
R22985 DVSS.n700 DVSS.n698 9.15497
R22986 DVSS.n2782 DVSS.n2781 9.15497
R22987 DVSS.n2781 DVSS.n2780 9.15497
R22988 DVSS.n699 DVSS.n697 9.15497
R22989 DVSS.n2779 DVSS.n699 9.15497
R22990 DVSS.n2777 DVSS.n2776 9.15497
R22991 DVSS.n2778 DVSS.n2777 9.15497
R22992 DVSS.n2775 DVSS.n702 9.15497
R22993 DVSS.n1751 DVSS.n702 9.15497
R22994 DVSS.n2424 DVSS.n2423 9.15497
R22995 DVSS.n2424 DVSS.n660 9.15497
R22996 DVSS.n1948 DVSS.n1947 9.15497
R22997 DVSS.n1947 DVSS.n1946 9.15497
R22998 DVSS.n1866 DVSS.n1864 9.15497
R22999 DVSS.n1864 DVSS.n1863 9.15497
R23000 DVSS.n1914 DVSS.n1913 9.15497
R23001 DVSS.n1915 DVSS.n1914 9.15497
R23002 DVSS.n1867 DVSS.n1865 9.15497
R23003 DVSS.n1865 DVSS.n1807 9.15497
R23004 DVSS.n1907 DVSS.n1906 9.15497
R23005 DVSS.n1906 DVSS.n1808 9.15497
R23006 DVSS.n1804 DVSS.n1802 9.15497
R23007 DVSS.n1806 DVSS.n1804 9.15497
R23008 DVSS.n1928 DVSS.n1927 9.15497
R23009 DVSS.n1805 DVSS.n1803 9.15497
R23010 DVSS.n1923 DVSS.n1922 9.15497
R23011 DVSS.n1919 DVSS.n1918 9.15497
R23012 DVSS.n1918 DVSS.n1917 9.15497
R23013 DVSS.n1795 DVSS.n1794 9.15497
R23014 DVSS.n1794 DVSS.n1793 9.15497
R23015 DVSS.n1943 DVSS.n1942 9.15497
R23016 DVSS.n1944 DVSS.n1943 9.15497
R23017 DVSS.n1937 DVSS.n1792 9.15497
R23018 DVSS.n1945 DVSS.n1792 9.15497
R23019 DVSS.n7 DVSS.n4 9.15497
R23020 DVSS.n2854 DVSS.n7 9.15497
R23021 DVSS.n3085 DVSS.n3084 9.15497
R23022 DVSS.n3084 DVSS.n3083 9.15497
R23023 DVSS.n8 DVSS.n6 9.15497
R23024 DVSS.n3082 DVSS.n8 9.15497
R23025 DVSS.n3080 DVSS.n3079 9.15497
R23026 DVSS.n3081 DVSS.n3080 9.15497
R23027 DVSS.n11 DVSS.n10 9.15497
R23028 DVSS.n10 DVSS.n9 9.15497
R23029 DVSS.n2866 DVSS.n2865 9.15497
R23030 DVSS.n2867 DVSS.n2866 9.15497
R23031 DVSS.n627 DVSS.n625 9.15497
R23032 DVSS.n625 DVSS.n624 9.15497
R23033 DVSS.n2860 DVSS.n2859 9.15497
R23034 DVSS.n2859 DVSS.n2858 9.15497
R23035 DVSS.n630 DVSS.n629 9.15497
R23036 DVSS.n2857 DVSS.n630 9.15497
R23037 DVSS.n652 DVSS.n651 9.15497
R23038 DVSS.n2833 DVSS.n652 9.15497
R23039 DVSS.n2837 DVSS.n2836 9.15497
R23040 DVSS.n2836 DVSS.n2835 9.15497
R23041 DVSS.n644 DVSS.n643 9.15497
R23042 DVSS.n643 DVSS.n642 9.15497
R23043 DVSS.n2842 DVSS.n2841 9.15497
R23044 DVSS.n2843 DVSS.n2842 9.15497
R23045 DVSS.n641 DVSS.n640 9.15497
R23046 DVSS.n2844 DVSS.n641 9.15497
R23047 DVSS.n2847 DVSS.n2846 9.15497
R23048 DVSS.n2846 DVSS.n2845 9.15497
R23049 DVSS.n637 DVSS.n635 9.15497
R23050 DVSS.n635 DVSS.n633 9.15497
R23051 DVSS.n2852 DVSS.n2851 9.15497
R23052 DVSS.n2853 DVSS.n2852 9.15497
R23053 DVSS.n636 DVSS.n634 9.15497
R23054 DVSS.n634 DVSS.n632 9.15497
R23055 DVSS.n1861 DVSS.n1860 9.15497
R23056 DVSS.n1862 DVSS.n1861 9.15497
R23057 DVSS.n1811 DVSS.n1810 9.15497
R23058 DVSS.n1810 DVSS.n1809 9.15497
R23059 DVSS.n1840 DVSS.n1839 9.15497
R23060 DVSS.n1847 DVSS.n1846 9.15497
R23061 DVSS.n1848 DVSS.n1847 9.15497
R23062 DVSS.n1822 DVSS.n1820 9.15497
R23063 DVSS.n1849 DVSS.n1822 9.15497
R23064 DVSS.n1852 DVSS.n1851 9.15497
R23065 DVSS.n1821 DVSS.n1819 9.15497
R23066 DVSS.n1837 DVSS.n1821 9.15497
R23067 DVSS.n1835 DVSS.n1834 9.15497
R23068 DVSS.n1836 DVSS.n1835 9.15497
R23069 DVSS.n2823 DVSS.n2822 9.15497
R23070 DVSS.n2826 DVSS.n654 9.15497
R23071 DVSS.n654 DVSS.n653 9.15497
R23072 DVSS.n2831 DVSS.n2830 9.15497
R23073 DVSS.n2832 DVSS.n2831 9.15497
R23074 DVSS.n2425 DVSS.n1787 9.15497
R23075 DVSS.n2426 DVSS.n2425 9.15497
R23076 DVSS.n2430 DVSS.n2429 9.15497
R23077 DVSS.n2429 DVSS.n2428 9.15497
R23078 DVSS.n1784 DVSS.n1783 9.15497
R23079 DVSS.n1783 DVSS.n1782 9.15497
R23080 DVSS.n2438 DVSS.n2437 9.15497
R23081 DVSS.n2439 DVSS.n2438 9.15497
R23082 DVSS.n1781 DVSS.n1780 9.15497
R23083 DVSS.n2447 DVSS.n2446 9.15497
R23084 DVSS.n2448 DVSS.n2447 9.15497
R23085 DVSS.n1777 DVSS.n1775 9.15497
R23086 DVSS.n2449 DVSS.n1777 9.15497
R23087 DVSS.n2470 DVSS.n2469 9.15497
R23088 DVSS.n1778 DVSS.n1776 9.15497
R23089 DVSS.n2467 DVSS.n1778 9.15497
R23090 DVSS.n2465 DVSS.n2464 9.15497
R23091 DVSS.n2466 DVSS.n2465 9.15497
R23092 DVSS.n2451 DVSS.n2450 9.15497
R23093 DVSS.n2458 DVSS.n2457 9.15497
R23094 DVSS.n2457 DVSS.n2456 9.15497
R23095 DVSS.n1768 DVSS.n1767 9.15497
R23096 DVSS.n2455 DVSS.n1767 9.15497
R23097 DVSS.n2479 DVSS.n2478 9.15497
R23098 DVSS.n2480 DVSS.n2479 9.15497
R23099 DVSS.n1766 DVSS.n1765 9.15497
R23100 DVSS.n2481 DVSS.n1766 9.15497
R23101 DVSS.n2485 DVSS.n2484 9.15497
R23102 DVSS.n2484 DVSS.n2483 9.15497
R23103 DVSS.n1763 DVSS.n1762 9.15497
R23104 DVSS.n2482 DVSS.n1762 9.15497
R23105 DVSS.n2496 DVSS.n2495 9.15497
R23106 DVSS.n2497 DVSS.n2496 9.15497
R23107 DVSS.n1761 DVSS.n1760 9.15497
R23108 DVSS.n2498 DVSS.n1761 9.15497
R23109 DVSS.n2502 DVSS.n2501 9.15497
R23110 DVSS.n2501 DVSS.n2500 9.15497
R23111 DVSS.n1757 DVSS.n1755 9.15497
R23112 DVSS.n2499 DVSS.n1755 9.15497
R23113 DVSS.n2514 DVSS.n2513 9.15497
R23114 DVSS.n2515 DVSS.n2514 9.15497
R23115 DVSS.n1758 DVSS.n1756 9.15497
R23116 DVSS.n1756 DVSS.n1750 9.15497
R23117 DVSS.n3066 DVSS.n3065 9.15497
R23118 DVSS.n3067 DVSS.n3066 9.15497
R23119 DVSS.n19 DVSS.n17 9.15497
R23120 DVSS.n3068 DVSS.n19 9.15497
R23121 DVSS.n3071 DVSS.n3070 9.15497
R23122 DVSS.n3070 DVSS.n3069 9.15497
R23123 DVSS.n3072 DVSS.n16 9.15497
R23124 DVSS.n1228 DVSS.n16 9.15497
R23125 DVSS.n2529 DVSS.n2528 9.15497
R23126 DVSS.n2530 DVSS.n2529 9.15497
R23127 DVSS.n1269 DVSS.n1267 9.15497
R23128 DVSS.n2531 DVSS.n1269 9.15497
R23129 DVSS.n2535 DVSS.n2534 9.15497
R23130 DVSS.n2534 DVSS.n2533 9.15497
R23131 DVSS.n1270 DVSS.n1268 9.15497
R23132 DVSS.n2532 DVSS.n1270 9.15497
R23133 DVSS.n1263 DVSS.n1262 9.15497
R23134 DVSS.n1262 DVSS.n1261 9.15497
R23135 DVSS.n2694 DVSS.n2693 9.15497
R23136 DVSS.n2693 DVSS.n2692 9.15497
R23137 DVSS.n1227 DVSS.n1225 9.15497
R23138 DVSS.n2610 DVSS.n1227 9.15497
R23139 DVSS.n2607 DVSS.n2606 9.15497
R23140 DVSS.n2608 DVSS.n2607 9.15497
R23141 DVSS.n1231 DVSS.n1230 9.15497
R23142 DVSS.n1230 DVSS.n1229 9.15497
R23143 DVSS.n2600 DVSS.n2599 9.15497
R23144 DVSS.n2599 DVSS.n2598 9.15497
R23145 DVSS.n1234 DVSS.n1233 9.15497
R23146 DVSS.n2596 DVSS.n1234 9.15497
R23147 DVSS.n2594 DVSS.n2593 9.15497
R23148 DVSS.n2595 DVSS.n2594 9.15497
R23149 DVSS.n1236 DVSS.n1235 9.15497
R23150 DVSS.n2581 DVSS.n1235 9.15497
R23151 DVSS.n2584 DVSS.n2583 9.15497
R23152 DVSS.n2583 DVSS.n2582 9.15497
R23153 DVSS.n1240 DVSS.n1239 9.15497
R23154 DVSS.n2580 DVSS.n1240 9.15497
R23155 DVSS.n2578 DVSS.n2577 9.15497
R23156 DVSS.n2579 DVSS.n2578 9.15497
R23157 DVSS.n1243 DVSS.n1242 9.15497
R23158 DVSS.n1242 DVSS.n1241 9.15497
R23159 DVSS.n2571 DVSS.n2570 9.15497
R23160 DVSS.n2570 DVSS.n2569 9.15497
R23161 DVSS.n1248 DVSS.n1247 9.15497
R23162 DVSS.n1249 DVSS.n1248 9.15497
R23163 DVSS.n2555 DVSS.n1250 9.15497
R23164 DVSS.n2562 DVSS.n1254 9.15497
R23165 DVSS.n1254 DVSS.n1251 9.15497
R23166 DVSS.n2564 DVSS.n2563 9.15497
R23167 DVSS.n2565 DVSS.n2564 9.15497
R23168 DVSS.n1255 DVSS.n1253 9.15497
R23169 DVSS.n2549 DVSS.n2548 9.15497
R23170 DVSS.n2548 DVSS.n2547 9.15497
R23171 DVSS.n1260 DVSS.n1259 9.15497
R23172 DVSS.n2546 DVSS.n1260 9.15497
R23173 DVSS.n732 DVSS.n731 9.15497
R23174 DVSS.n2743 DVSS.n732 9.15497
R23175 DVSS.n2741 DVSS.n2740 9.15497
R23176 DVSS.n2742 DVSS.n2741 9.15497
R23177 DVSS.n734 DVSS.n733 9.15497
R23178 DVSS.n2567 DVSS.n733 9.15497
R23179 DVSS.n2734 DVSS.n2733 9.15497
R23180 DVSS.n2733 DVSS.n2732 9.15497
R23181 DVSS.n740 DVSS.n739 9.15497
R23182 DVSS.n2731 DVSS.n740 9.15497
R23183 DVSS.n2729 DVSS.n2728 9.15497
R23184 DVSS.n2730 DVSS.n2729 9.15497
R23185 DVSS.n743 DVSS.n742 9.15497
R23186 DVSS.n742 DVSS.n741 9.15497
R23187 DVSS.n2721 DVSS.n2720 9.15497
R23188 DVSS.n2720 DVSS.n2719 9.15497
R23189 DVSS.n747 DVSS.n746 9.15497
R23190 DVSS.n2718 DVSS.n747 9.15497
R23191 DVSS.n2715 DVSS.n2714 9.15497
R23192 DVSS.n2716 DVSS.n2715 9.15497
R23193 DVSS.n750 DVSS.n749 9.15497
R23194 DVSS.n751 DVSS.n750 9.15497
R23195 DVSS.n2709 DVSS.n2708 9.15497
R23196 DVSS.n2689 DVSS.n2688 9.15497
R23197 DVSS.n2690 DVSS.n2689 9.15497
R23198 DVSS.n2664 DVSS.n2663 9.15497
R23199 DVSS.n2663 DVSS.n20 9.15497
R23200 DVSS.n2683 DVSS.n2682 9.15497
R23201 DVSS.n2682 DVSS.n21 9.15497
R23202 DVSS.n2681 DVSS.n2666 9.15497
R23203 DVSS.n2681 DVSS.n2680 9.15497
R23204 DVSS.n2678 DVSS.n2677 9.15497
R23205 DVSS.n2679 DVSS.n2678 9.15497
R23206 DVSS.n26 DVSS.n24 9.15497
R23207 DVSS.n3051 DVSS.n3050 9.15497
R23208 DVSS.n3052 DVSS.n3051 9.15497
R23209 DVSS.n3049 DVSS.n25 9.15497
R23210 DVSS.n25 DVSS.n23 9.15497
R23211 DVSS.n34 DVSS.n28 9.15497
R23212 DVSS.n3043 DVSS.n3042 9.15497
R23213 DVSS.n3042 DVSS.n3041 9.15497
R23214 DVSS.n35 DVSS.n33 9.15497
R23215 DVSS.n3040 DVSS.n35 9.15497
R23216 DVSS.n565 DVSS.n37 9.15497
R23217 DVSS.n567 DVSS.n566 9.15497
R23218 DVSS.n567 DVSS.n38 9.15497
R23219 DVSS.n569 DVSS.n568 9.15497
R23220 DVSS.n568 DVSS.n39 9.15497
R23221 DVSS.n557 DVSS.n556 9.15497
R23222 DVSS.n556 DVSS.n40 9.15497
R23223 DVSS.n576 DVSS.n575 9.15497
R23224 DVSS.n577 DVSS.n576 9.15497
R23225 DVSS.n555 DVSS.n554 9.15497
R23226 DVSS.n578 DVSS.n555 9.15497
R23227 DVSS.n582 DVSS.n581 9.15497
R23228 DVSS.n581 DVSS.n580 9.15497
R23229 DVSS.n550 DVSS.n549 9.15497
R23230 DVSS.n579 DVSS.n549 9.15497
R23231 DVSS.n595 DVSS.n594 9.15497
R23232 DVSS.n596 DVSS.n595 9.15497
R23233 DVSS.n551 DVSS.n547 9.15497
R23234 DVSS.n597 DVSS.n547 9.15497
R23235 DVSS.n599 DVSS.n548 9.15497
R23236 DVSS.n599 DVSS.n598 9.15497
R23237 DVSS.n600 DVSS.n545 9.15497
R23238 DVSS.n601 DVSS.n600 9.15497
R23239 DVSS.n604 DVSS.n603 9.15497
R23240 DVSS.n603 DVSS.n602 9.15497
R23241 DVSS.n75 DVSS.n65 9.15497
R23242 DVSS.n3011 DVSS.n65 9.15497
R23243 DVSS.n2629 DVSS.n2628 9.15497
R23244 DVSS.n2628 DVSS.n2627 9.15497
R23245 DVSS.n2636 DVSS.n2635 9.15497
R23246 DVSS.n2635 DVSS.n2634 9.15497
R23247 DVSS.n45 DVSS.n43 9.15497
R23248 DVSS.n43 DVSS.n41 9.15497
R23249 DVSS.n3036 DVSS.n3035 9.15497
R23250 DVSS.n3037 DVSS.n3036 9.15497
R23251 DVSS.n46 DVSS.n44 9.15497
R23252 DVSS.n44 DVSS.n42 9.15497
R23253 DVSS.n53 DVSS.n51 9.15497
R23254 DVSS.n3027 DVSS.n3026 9.15497
R23255 DVSS.n54 DVSS.n52 9.15497
R23256 DVSS.n3021 DVSS.n3020 9.15497
R23257 DVSS.n3022 DVSS.n3021 9.15497
R23258 DVSS.n3019 DVSS.n57 9.15497
R23259 DVSS.n57 DVSS.n56 9.15497
R23260 DVSS.n64 DVSS.n59 9.15497
R23261 DVSS.n66 DVSS.n64 9.15497
R23262 DVSS.n3014 DVSS.n3013 9.15497
R23263 DVSS.n3013 DVSS.n3012 9.15497
R23264 DVSS.n2989 DVSS.n2988 9.15497
R23265 DVSS.n2991 DVSS.n2990 9.15497
R23266 DVSS.n2993 DVSS.n2992 9.15497
R23267 DVSS.n2888 DVSS.n2887 9.15497
R23268 DVSS.n2998 DVSS.n2997 9.15497
R23269 DVSS.n3000 DVSS.n2999 9.15497
R23270 DVSS.n3002 DVSS.n3001 9.15497
R23271 DVSS.n2885 DVSS.n2884 9.15497
R23272 DVSS.n2987 DVSS.n2986 9.15497
R23273 DVSS.n2970 DVSS.n2894 9.15497
R23274 DVSS.n2972 DVSS.n2971 9.15497
R23275 DVSS.n2974 DVSS.n2973 9.15497
R23276 DVSS.n2976 DVSS.n2975 9.15497
R23277 DVSS.n2983 DVSS.n2892 9.15497
R23278 DVSS.n2985 DVSS.n2984 9.15497
R23279 DVSS.n2913 DVSS.n2912 9.15497
R23280 DVSS.n2912 DVSS.n619 9.15497
R23281 DVSS.n2918 DVSS.n2917 9.15497
R23282 DVSS.n2920 DVSS.n2911 9.15497
R23283 DVSS.n2923 DVSS.n2922 9.15497
R23284 DVSS.n2909 DVSS.n2908 9.15497
R23285 DVSS.n2931 DVSS.n2930 9.15497
R23286 DVSS.n2933 DVSS.n2907 9.15497
R23287 DVSS.n2936 DVSS.n2935 9.15497
R23288 DVSS.n2905 DVSS.n2904 9.15497
R23289 DVSS.n2944 DVSS.n2943 9.15497
R23290 DVSS.n2946 DVSS.n2903 9.15497
R23291 DVSS.n2949 DVSS.n2948 9.15497
R23292 DVSS.n2901 DVSS.n2900 9.15497
R23293 DVSS.n2958 DVSS.n2957 9.15497
R23294 DVSS.n2960 DVSS.n2899 9.15497
R23295 DVSS.n2914 DVSS.n617 9.15497
R23296 DVSS.n535 DVSS.n82 9.01392
R23297 DVSS.n90 DVSS.n81 9.01392
R23298 DVSS.n527 DVSS.n526 9.01392
R23299 DVSS.n88 DVSS.n87 9.01392
R23300 DVSS.n496 DVSS.n495 9.01392
R23301 DVSS.n98 DVSS.n96 9.01392
R23302 DVSS.n108 DVSS.n107 9.01392
R23303 DVSS.n456 DVSS.n455 9.01392
R23304 DVSS.n114 DVSS.n106 9.01392
R23305 DVSS.n448 DVSS.n447 9.01392
R23306 DVSS.n435 DVSS.n434 9.01392
R23307 DVSS.n146 DVSS.n145 9.01392
R23308 DVSS.n428 DVSS.n427 9.01392
R23309 DVSS.n151 DVSS.n150 9.01392
R23310 DVSS.n2408 DVSS.n1955 9.01392
R23311 DVSS.n1963 DVSS.n1954 9.01392
R23312 DVSS.n2400 DVSS.n2399 9.01392
R23313 DVSS.n1961 DVSS.n1960 9.01392
R23314 DVSS.n2369 DVSS.n2368 9.01392
R23315 DVSS.n1971 DVSS.n1969 9.01392
R23316 DVSS.n1981 DVSS.n1980 9.01392
R23317 DVSS.n2329 DVSS.n2328 9.01392
R23318 DVSS.n1987 DVSS.n1979 9.01392
R23319 DVSS.n2321 DVSS.n2320 9.01392
R23320 DVSS.n2308 DVSS.n2307 9.01392
R23321 DVSS.n2019 DVSS.n2018 9.01392
R23322 DVSS.n2301 DVSS.n2300 9.01392
R23323 DVSS.n2024 DVSS.n2023 9.01392
R23324 DVSS.n1216 DVSS.n763 9.01392
R23325 DVSS.n771 DVSS.n762 9.01392
R23326 DVSS.n1208 DVSS.n1207 9.01392
R23327 DVSS.n769 DVSS.n768 9.01392
R23328 DVSS.n1177 DVSS.n1176 9.01392
R23329 DVSS.n779 DVSS.n777 9.01392
R23330 DVSS.n789 DVSS.n788 9.01392
R23331 DVSS.n1137 DVSS.n1136 9.01392
R23332 DVSS.n795 DVSS.n787 9.01392
R23333 DVSS.n1129 DVSS.n1128 9.01392
R23334 DVSS.n1116 DVSS.n1115 9.01392
R23335 DVSS.n827 DVSS.n826 9.01392
R23336 DVSS.n1109 DVSS.n1108 9.01392
R23337 DVSS.n832 DVSS.n831 9.01392
R23338 DVSS.n1738 DVSS.n1285 9.01392
R23339 DVSS.n1293 DVSS.n1284 9.01392
R23340 DVSS.n1730 DVSS.n1729 9.01392
R23341 DVSS.n1291 DVSS.n1290 9.01392
R23342 DVSS.n1699 DVSS.n1698 9.01392
R23343 DVSS.n1301 DVSS.n1299 9.01392
R23344 DVSS.n1311 DVSS.n1310 9.01392
R23345 DVSS.n1659 DVSS.n1658 9.01392
R23346 DVSS.n1317 DVSS.n1309 9.01392
R23347 DVSS.n1651 DVSS.n1650 9.01392
R23348 DVSS.n1638 DVSS.n1637 9.01392
R23349 DVSS.n1349 DVSS.n1348 9.01392
R23350 DVSS.n1631 DVSS.n1630 9.01392
R23351 DVSS.n1354 DVSS.n1353 9.01392
R23352 DVSS.n419 DVSS.n151 9.01392
R23353 DVSS.n427 DVSS.n426 9.01392
R23354 DVSS.n422 DVSS.n145 9.01392
R23355 DVSS.n436 DVSS.n435 9.01392
R23356 DVSS.n447 DVSS.n446 9.01392
R23357 DVSS.n441 DVSS.n106 9.01392
R23358 DVSS.n457 DVSS.n456 9.01392
R23359 DVSS.n107 DVSS.n103 9.01392
R23360 DVSS.n464 DVSS.n98 9.01392
R23361 DVSS.n495 DVSS.n494 9.01392
R23362 DVSS.n490 DVSS.n87 9.01392
R23363 DVSS.n528 DVSS.n527 9.01392
R23364 DVSS.n530 DVSS.n81 9.01392
R23365 DVSS.n535 DVSS.n534 9.01392
R23366 DVSS.n2292 DVSS.n2024 9.01392
R23367 DVSS.n2300 DVSS.n2299 9.01392
R23368 DVSS.n2295 DVSS.n2018 9.01392
R23369 DVSS.n2309 DVSS.n2308 9.01392
R23370 DVSS.n2320 DVSS.n2319 9.01392
R23371 DVSS.n2314 DVSS.n1979 9.01392
R23372 DVSS.n2330 DVSS.n2329 9.01392
R23373 DVSS.n1980 DVSS.n1976 9.01392
R23374 DVSS.n2337 DVSS.n1971 9.01392
R23375 DVSS.n2368 DVSS.n2367 9.01392
R23376 DVSS.n2363 DVSS.n1960 9.01392
R23377 DVSS.n2401 DVSS.n2400 9.01392
R23378 DVSS.n2403 DVSS.n1954 9.01392
R23379 DVSS.n2408 DVSS.n2407 9.01392
R23380 DVSS.n1100 DVSS.n832 9.01392
R23381 DVSS.n1108 DVSS.n1107 9.01392
R23382 DVSS.n1103 DVSS.n826 9.01392
R23383 DVSS.n1117 DVSS.n1116 9.01392
R23384 DVSS.n1128 DVSS.n1127 9.01392
R23385 DVSS.n1122 DVSS.n787 9.01392
R23386 DVSS.n1138 DVSS.n1137 9.01392
R23387 DVSS.n788 DVSS.n784 9.01392
R23388 DVSS.n1145 DVSS.n779 9.01392
R23389 DVSS.n1176 DVSS.n1175 9.01392
R23390 DVSS.n1171 DVSS.n768 9.01392
R23391 DVSS.n1209 DVSS.n1208 9.01392
R23392 DVSS.n1211 DVSS.n762 9.01392
R23393 DVSS.n1216 DVSS.n1215 9.01392
R23394 DVSS.n1622 DVSS.n1354 9.01392
R23395 DVSS.n1630 DVSS.n1629 9.01392
R23396 DVSS.n1625 DVSS.n1348 9.01392
R23397 DVSS.n1639 DVSS.n1638 9.01392
R23398 DVSS.n1650 DVSS.n1649 9.01392
R23399 DVSS.n1644 DVSS.n1309 9.01392
R23400 DVSS.n1660 DVSS.n1659 9.01392
R23401 DVSS.n1310 DVSS.n1306 9.01392
R23402 DVSS.n1667 DVSS.n1301 9.01392
R23403 DVSS.n1698 DVSS.n1697 9.01392
R23404 DVSS.n1693 DVSS.n1290 9.01392
R23405 DVSS.n1731 DVSS.n1730 9.01392
R23406 DVSS.n1733 DVSS.n1284 9.01392
R23407 DVSS.n1738 DVSS.n1737 9.01392
R23408 DVSS.n2990 DVSS.n2871 8.99329
R23409 DVSS.n2961 DVSS.n2960 8.99329
R23410 DVSS.n3001 DVSS.n2883 8.99094
R23411 DVSS.n2997 DVSS.n2881 8.99094
R23412 DVSS.n2992 DVSS.n2879 8.99094
R23413 DVSS.n2887 DVSS.n2879 8.99094
R23414 DVSS.n2999 DVSS.n2881 8.99094
R23415 DVSS.n2884 DVSS.n2883 8.99094
R23416 DVSS.n377 DVSS.n369 8.9737
R23417 DVSS.n2250 DVSS.n2242 8.9737
R23418 DVSS.n1058 DVSS.n1050 8.9737
R23419 DVSS.n1580 DVSS.n1572 8.9737
R23420 DVSS.n417 DVSS.n180 8.8706
R23421 DVSS.n2290 DVSS.n2053 8.8706
R23422 DVSS.n1098 DVSS.n861 8.8706
R23423 DVSS.n1620 DVSS.n1383 8.8706
R23424 DVSS.n2519 DVSS.n1749 8.85585
R23425 DVSS.n2919 DVSS.n2918 8.85585
R23426 DVSS.n2984 DVSS.n2877 8.85488
R23427 DVSS.n2975 DVSS.n2876 8.85488
R23428 DVSS.n2971 DVSS.n2875 8.85488
R23429 DVSS.n1828 DVSS.n1823 8.85488
R23430 DVSS.n2769 DVSS.n710 8.85488
R23431 DVSS.n710 DVSS.n709 8.85488
R23432 DVSS.n2987 DVSS.n2877 8.85488
R23433 DVSS.n2970 DVSS.n2874 8.85488
R23434 DVSS.n2974 DVSS.n2875 8.85488
R23435 DVSS.n2983 DVSS.n2876 8.85488
R23436 DVSS.n2921 DVSS.n2908 8.85488
R23437 DVSS.n2933 DVSS.n2932 8.85488
R23438 DVSS.n2934 DVSS.n2904 8.85488
R23439 DVSS.n2946 DVSS.n2945 8.85488
R23440 DVSS.n2947 DVSS.n2900 8.85488
R23441 DVSS.n2922 DVSS.n2921 8.85488
R23442 DVSS.n2932 DVSS.n2931 8.85488
R23443 DVSS.n2935 DVSS.n2934 8.85488
R23444 DVSS.n2945 DVSS.n2944 8.85488
R23445 DVSS.n2948 DVSS.n2947 8.85488
R23446 DVSS.n2441 DVSS.n1780 8.85487
R23447 DVSS.n2708 DVSS.n2707 8.85487
R23448 DVSS.n2672 DVSS.n24 8.85487
R23449 DVSS.n2920 DVSS.n2919 8.85487
R23450 DVSS.n2988 DVSS.n2871 8.85257
R23451 DVSS.n354 DVSS.n353 8.15208
R23452 DVSS.n2227 DVSS.n2226 8.15208
R23453 DVSS.n1035 DVSS.n1034 8.15208
R23454 DVSS.n1557 DVSS.n1556 8.15208
R23455 DVSS.n166 DVSS.n165 7.5692
R23456 DVSS.n175 DVSS.n166 7.5692
R23457 DVSS.n175 DVSS.n174 7.5692
R23458 DVSS.n174 DVSS.n172 7.5692
R23459 DVSS.n172 DVSS.n170 7.5692
R23460 DVSS.n170 DVSS.n168 7.5692
R23461 DVSS.n168 DVSS.n155 7.5692
R23462 DVSS.n180 DVSS.n155 7.5692
R23463 DVSS.n506 DVSS.n501 7.5692
R23464 DVSS.n515 DVSS.n506 7.5692
R23465 DVSS.n515 DVSS.n514 7.5692
R23466 DVSS.n514 DVSS.n513 7.5692
R23467 DVSS.n513 DVSS.n510 7.5692
R23468 DVSS.n510 DVSS.n509 7.5692
R23469 DVSS.n509 DVSS.n79 7.5692
R23470 DVSS.n537 DVSS.n79 7.5692
R23471 DVSS.n2039 DVSS.n2038 7.5692
R23472 DVSS.n2048 DVSS.n2039 7.5692
R23473 DVSS.n2048 DVSS.n2047 7.5692
R23474 DVSS.n2047 DVSS.n2045 7.5692
R23475 DVSS.n2045 DVSS.n2043 7.5692
R23476 DVSS.n2043 DVSS.n2041 7.5692
R23477 DVSS.n2041 DVSS.n2028 7.5692
R23478 DVSS.n2053 DVSS.n2028 7.5692
R23479 DVSS.n2379 DVSS.n2374 7.5692
R23480 DVSS.n2388 DVSS.n2379 7.5692
R23481 DVSS.n2388 DVSS.n2387 7.5692
R23482 DVSS.n2387 DVSS.n2386 7.5692
R23483 DVSS.n2386 DVSS.n2383 7.5692
R23484 DVSS.n2383 DVSS.n2382 7.5692
R23485 DVSS.n2382 DVSS.n1952 7.5692
R23486 DVSS.n2410 DVSS.n1952 7.5692
R23487 DVSS.n847 DVSS.n846 7.5692
R23488 DVSS.n856 DVSS.n847 7.5692
R23489 DVSS.n856 DVSS.n855 7.5692
R23490 DVSS.n855 DVSS.n853 7.5692
R23491 DVSS.n853 DVSS.n851 7.5692
R23492 DVSS.n851 DVSS.n849 7.5692
R23493 DVSS.n849 DVSS.n836 7.5692
R23494 DVSS.n861 DVSS.n836 7.5692
R23495 DVSS.n1187 DVSS.n1182 7.5692
R23496 DVSS.n1196 DVSS.n1187 7.5692
R23497 DVSS.n1196 DVSS.n1195 7.5692
R23498 DVSS.n1195 DVSS.n1194 7.5692
R23499 DVSS.n1194 DVSS.n1191 7.5692
R23500 DVSS.n1191 DVSS.n1190 7.5692
R23501 DVSS.n1190 DVSS.n760 7.5692
R23502 DVSS.n1218 DVSS.n760 7.5692
R23503 DVSS.n1369 DVSS.n1368 7.5692
R23504 DVSS.n1378 DVSS.n1369 7.5692
R23505 DVSS.n1378 DVSS.n1377 7.5692
R23506 DVSS.n1377 DVSS.n1375 7.5692
R23507 DVSS.n1375 DVSS.n1373 7.5692
R23508 DVSS.n1373 DVSS.n1371 7.5692
R23509 DVSS.n1371 DVSS.n1358 7.5692
R23510 DVSS.n1383 DVSS.n1358 7.5692
R23511 DVSS.n1709 DVSS.n1704 7.5692
R23512 DVSS.n1718 DVSS.n1709 7.5692
R23513 DVSS.n1718 DVSS.n1717 7.5692
R23514 DVSS.n1717 DVSS.n1716 7.5692
R23515 DVSS.n1716 DVSS.n1713 7.5692
R23516 DVSS.n1713 DVSS.n1712 7.5692
R23517 DVSS.n1712 DVSS.n1282 7.5692
R23518 DVSS.n1740 DVSS.n1282 7.5692
R23519 DVSS.n538 DVSS.n537 7.1358
R23520 DVSS.n2411 DVSS.n2410 7.1358
R23521 DVSS.n1219 DVSS.n1218 7.1358
R23522 DVSS.n1741 DVSS.n1740 7.1358
R23523 DVSS.n538 DVSS.n78 6.65838
R23524 DVSS.n2411 DVSS.n1951 6.65838
R23525 DVSS.n1219 DVSS.n759 6.65838
R23526 DVSS.n1741 DVSS.n1281 6.65838
R23527 DVSS.n381 DVSS.n380 6.46787
R23528 DVSS.n2254 DVSS.n2253 6.46787
R23529 DVSS.n1062 DVSS.n1061 6.46787
R23530 DVSS.n1584 DVSS.n1583 6.46787
R23531 DVSS.n333 DVSS.n332 5.72682
R23532 DVSS.n332 DVSS.n331 5.72682
R23533 DVSS.n331 DVSS.n328 5.72682
R23534 DVSS.n328 DVSS.n327 5.72682
R23535 DVSS.n327 DVSS.n324 5.72682
R23536 DVSS.n324 DVSS.n323 5.72682
R23537 DVSS.n323 DVSS.n316 5.72682
R23538 DVSS.n339 DVSS.n316 5.72682
R23539 DVSS.n2206 DVSS.n2205 5.72682
R23540 DVSS.n2205 DVSS.n2204 5.72682
R23541 DVSS.n2204 DVSS.n2201 5.72682
R23542 DVSS.n2201 DVSS.n2200 5.72682
R23543 DVSS.n2200 DVSS.n2197 5.72682
R23544 DVSS.n2197 DVSS.n2196 5.72682
R23545 DVSS.n2196 DVSS.n2189 5.72682
R23546 DVSS.n2212 DVSS.n2189 5.72682
R23547 DVSS.n1014 DVSS.n1013 5.72682
R23548 DVSS.n1013 DVSS.n1012 5.72682
R23549 DVSS.n1012 DVSS.n1009 5.72682
R23550 DVSS.n1009 DVSS.n1008 5.72682
R23551 DVSS.n1008 DVSS.n1005 5.72682
R23552 DVSS.n1005 DVSS.n1004 5.72682
R23553 DVSS.n1004 DVSS.n997 5.72682
R23554 DVSS.n1020 DVSS.n997 5.72682
R23555 DVSS.n1536 DVSS.n1535 5.72682
R23556 DVSS.n1535 DVSS.n1534 5.72682
R23557 DVSS.n1534 DVSS.n1531 5.72682
R23558 DVSS.n1531 DVSS.n1530 5.72682
R23559 DVSS.n1530 DVSS.n1527 5.72682
R23560 DVSS.n1527 DVSS.n1526 5.72682
R23561 DVSS.n1526 DVSS.n1519 5.72682
R23562 DVSS.n1542 DVSS.n1519 5.72682
R23563 DVSS.n606 DVSS.n69 5.64756
R23564 DVSS.n218 DVSS.n217 5.64756
R23565 DVSS.n217 DVSS.n207 5.64756
R23566 DVSS.n197 DVSS.n196 5.64756
R23567 DVSS.n196 DVSS.n186 5.64756
R23568 DVSS.n2091 DVSS.n2090 5.64756
R23569 DVSS.n2090 DVSS.n2080 5.64756
R23570 DVSS.n2070 DVSS.n2069 5.64756
R23571 DVSS.n2069 DVSS.n2059 5.64756
R23572 DVSS.n2826 DVSS.n2825 5.64756
R23573 DVSS.n899 DVSS.n898 5.64756
R23574 DVSS.n898 DVSS.n888 5.64756
R23575 DVSS.n878 DVSS.n877 5.64756
R23576 DVSS.n877 DVSS.n867 5.64756
R23577 DVSS.n2695 DVSS.n1225 5.64756
R23578 DVSS.n2508 DVSS.n1748 5.64756
R23579 DVSS.n1421 DVSS.n1420 5.64756
R23580 DVSS.n1420 DVSS.n1410 5.64756
R23581 DVSS.n1400 DVSS.n1399 5.64756
R23582 DVSS.n1399 DVSS.n1389 5.64756
R23583 DVSS.n446 DVSS.n116 5.57999
R23584 DVSS.n494 DVSS.n101 5.57999
R23585 DVSS.n2319 DVSS.n1989 5.57999
R23586 DVSS.n2367 DVSS.n1974 5.57999
R23587 DVSS.n1127 DVSS.n797 5.57999
R23588 DVSS.n1175 DVSS.n782 5.57999
R23589 DVSS.n1649 DVSS.n1319 5.57999
R23590 DVSS.n1697 DVSS.n1304 5.57999
R23591 DVSS.n436 DVSS.n144 5.34556
R23592 DVSS.n2309 DVSS.n2017 5.34556
R23593 DVSS.n1117 DVSS.n825 5.34556
R23594 DVSS.n1639 DVSS.n1347 5.34556
R23595 DVSS.n490 DVSS.n489 5.29867
R23596 DVSS.n2363 DVSS.n2362 5.29867
R23597 DVSS.n1171 DVSS.n1170 5.29867
R23598 DVSS.n1693 DVSS.n1692 5.29867
R23599 DVSS.n3014 DVSS.n63 5.27109
R23600 DVSS.n1937 DVSS.n1791 5.27109
R23601 DVSS.n2709 DVSS.n755 5.27109
R23602 DVSS.n2770 DVSS.n708 5.27109
R23603 DVSS.n221 DVSS.n204 4.89462
R23604 DVSS.n200 DVSS.n183 4.89462
R23605 DVSS.n2094 DVSS.n2077 4.89462
R23606 DVSS.n2073 DVSS.n2056 4.89462
R23607 DVSS.n902 DVSS.n885 4.89462
R23608 DVSS.n881 DVSS.n864 4.89462
R23609 DVSS.n1424 DVSS.n1407 4.89462
R23610 DVSS.n1403 DVSS.n1386 4.89462
R23611 DVSS.n389 DVSS.n243 4.74328
R23612 DVSS.n284 DVSS.n259 4.74328
R23613 DVSS.n2262 DVSS.n2116 4.74328
R23614 DVSS.n2157 DVSS.n2132 4.74328
R23615 DVSS.n1070 DVSS.n924 4.74328
R23616 DVSS.n965 DVSS.n940 4.74328
R23617 DVSS.n1592 DVSS.n1446 4.74328
R23618 DVSS.n1487 DVSS.n1462 4.74328
R23619 DVSS.n2959 DVSS.n618 4.72584
R23620 DVSS.n3006 DVSS.n3005 4.72584
R23621 DVSS.n2968 DVSS.n2897 4.6505
R23622 DVSS.n2897 DVSS.n2895 4.6505
R23623 DVSS.n2966 DVSS.n2965 4.6505
R23624 DVSS.n2989 DVSS.n2890 4.6505
R23625 DVSS.n3031 DVSS.n3029 4.6505
R23626 DVSS.n3032 DVSS.n3031 4.6505
R23627 DVSS.n2632 DVSS.n47 4.6505
R23628 DVSS.n2633 DVSS.n2632 4.6505
R23629 DVSS.n2616 DVSS.n2615 4.6505
R23630 DVSS.n2658 DVSS.n2615 4.6505
R23631 DVSS.n2657 DVSS.n2656 4.6505
R23632 DVSS.n2623 DVSS.n2617 4.6505
R23633 DVSS.n2650 DVSS.n2649 4.6505
R23634 DVSS.n2648 DVSS.n2622 4.6505
R23635 DVSS.n2647 DVSS.n2646 4.6505
R23636 DVSS.n2625 DVSS.n2624 4.6505
R23637 DVSS.n2640 DVSS.n2639 4.6505
R23638 DVSS.n389 DVSS.n388 4.6505
R23639 DVSS.n409 DVSS.n408 4.6505
R23640 DVSS.n391 DVSS.n390 4.6505
R23641 DVSS.n394 DVSS.n241 4.6505
R23642 DVSS.n398 DVSS.n397 4.6505
R23643 DVSS.n400 DVSS.n399 4.6505
R23644 DVSS.n240 DVSS.n237 4.6505
R23645 DVSS.n225 DVSS.n223 4.6505
R23646 DVSS.n266 DVSS.n202 4.6505
R23647 DVSS.n297 DVSS.n296 4.6505
R23648 DVSS.n299 DVSS.n298 4.6505
R23649 DVSS.n283 DVSS.n278 4.6505
R23650 DVSS.n272 DVSS.n268 4.6505
R23651 DVSS.n307 DVSS.n306 4.6505
R23652 DVSS.n309 DVSS.n308 4.6505
R23653 DVSS.n285 DVSS.n284 4.6505
R23654 DVSS.n587 DVSS.n552 4.6505
R23655 DVSS.n573 DVSS.n572 4.6505
R23656 DVSS.n572 DVSS.n571 4.6505
R23657 DVSS.n3046 DVSS.n3045 4.6505
R23658 DVSS.n562 DVSS.n560 4.6505
R23659 DVSS.n563 DVSS.n562 4.6505
R23660 DVSS.n3047 DVSS.n3046 4.6505
R23661 DVSS.n2670 DVSS.n26 4.6505
R23662 DVSS.n2688 DVSS.n2687 4.6505
R23663 DVSS.n2669 DVSS.n2665 4.6505
R23664 DVSS.n2669 DVSS.n2668 4.6505
R23665 DVSS.n2675 DVSS.n2669 4.6505
R23666 DVSS.n1931 DVSS.n1799 4.6505
R23667 DVSS.n1931 DVSS.n1930 4.6505
R23668 DVSS.n1909 DVSS.n1798 4.6505
R23669 DVSS.n1911 DVSS.n1798 4.6505
R23670 DVSS.n1885 DVSS.n1884 4.6505
R23671 DVSS.n1884 DVSS.n1882 4.6505
R23672 DVSS.n2262 DVSS.n2261 4.6505
R23673 DVSS.n2282 DVSS.n2281 4.6505
R23674 DVSS.n2264 DVSS.n2263 4.6505
R23675 DVSS.n2267 DVSS.n2114 4.6505
R23676 DVSS.n2271 DVSS.n2270 4.6505
R23677 DVSS.n2273 DVSS.n2272 4.6505
R23678 DVSS.n2113 DVSS.n2110 4.6505
R23679 DVSS.n2098 DVSS.n2096 4.6505
R23680 DVSS.n2139 DVSS.n2075 4.6505
R23681 DVSS.n2170 DVSS.n2169 4.6505
R23682 DVSS.n2172 DVSS.n2171 4.6505
R23683 DVSS.n2156 DVSS.n2151 4.6505
R23684 DVSS.n2145 DVSS.n2141 4.6505
R23685 DVSS.n2180 DVSS.n2179 4.6505
R23686 DVSS.n2182 DVSS.n2181 4.6505
R23687 DVSS.n2158 DVSS.n2157 4.6505
R23688 DVSS.n1887 DVSS.n1886 4.6505
R23689 DVSS.n1875 DVSS.n1874 4.6505
R23690 DVSS.n1894 DVSS.n1893 4.6505
R23691 DVSS.n1895 DVSS.n1873 4.6505
R23692 DVSS.n1897 DVSS.n1896 4.6505
R23693 DVSS.n1869 DVSS.n1868 4.6505
R23694 DVSS.n1904 DVSS.n1903 4.6505
R23695 DVSS.n2726 DVSS.n2725 4.6505
R23696 DVSS.n2725 DVSS.n744 4.6505
R23697 DVSS.n2737 DVSS.n2736 4.6505
R23698 DVSS.n2738 DVSS.n2737 4.6505
R23699 DVSS.n2759 DVSS.n721 4.6505
R23700 DVSS.n721 DVSS.n719 4.6505
R23701 DVSS.n1070 DVSS.n1069 4.6505
R23702 DVSS.n1090 DVSS.n1089 4.6505
R23703 DVSS.n1072 DVSS.n1071 4.6505
R23704 DVSS.n1075 DVSS.n922 4.6505
R23705 DVSS.n1079 DVSS.n1078 4.6505
R23706 DVSS.n1081 DVSS.n1080 4.6505
R23707 DVSS.n921 DVSS.n918 4.6505
R23708 DVSS.n906 DVSS.n904 4.6505
R23709 DVSS.n947 DVSS.n883 4.6505
R23710 DVSS.n978 DVSS.n977 4.6505
R23711 DVSS.n980 DVSS.n979 4.6505
R23712 DVSS.n964 DVSS.n959 4.6505
R23713 DVSS.n953 DVSS.n949 4.6505
R23714 DVSS.n988 DVSS.n987 4.6505
R23715 DVSS.n990 DVSS.n989 4.6505
R23716 DVSS.n966 DVSS.n965 4.6505
R23717 DVSS.n2761 DVSS.n2760 4.6505
R23718 DVSS.n2758 DVSS.n718 4.6505
R23719 DVSS.n2757 DVSS.n2756 4.6505
R23720 DVSS.n723 DVSS.n722 4.6505
R23721 DVSS.n2750 DVSS.n2749 4.6505
R23722 DVSS.n2748 DVSS.n729 4.6505
R23723 DVSS.n2747 DVSS.n2746 4.6505
R23724 DVSS.n2786 DVSS.n2784 4.6505
R23725 DVSS.n2787 DVSS.n2786 4.6505
R23726 DVSS.n693 DVSS.n690 4.6505
R23727 DVSS.n693 DVSS.n683 4.6505
R23728 DVSS.n672 DVSS.n671 4.6505
R23729 DVSS.n671 DVSS.n669 4.6505
R23730 DVSS.n1592 DVSS.n1591 4.6505
R23731 DVSS.n1612 DVSS.n1611 4.6505
R23732 DVSS.n1594 DVSS.n1593 4.6505
R23733 DVSS.n1597 DVSS.n1444 4.6505
R23734 DVSS.n1601 DVSS.n1600 4.6505
R23735 DVSS.n1603 DVSS.n1602 4.6505
R23736 DVSS.n1443 DVSS.n1440 4.6505
R23737 DVSS.n1428 DVSS.n1426 4.6505
R23738 DVSS.n1469 DVSS.n1405 4.6505
R23739 DVSS.n1500 DVSS.n1499 4.6505
R23740 DVSS.n1502 DVSS.n1501 4.6505
R23741 DVSS.n1486 DVSS.n1481 4.6505
R23742 DVSS.n1475 DVSS.n1471 4.6505
R23743 DVSS.n1510 DVSS.n1509 4.6505
R23744 DVSS.n1512 DVSS.n1511 4.6505
R23745 DVSS.n1488 DVSS.n1487 4.6505
R23746 DVSS.n2773 DVSS.n704 4.6505
R23747 DVSS.n668 DVSS.n667 4.6505
R23748 DVSS.n2812 DVSS.n673 4.6505
R23749 DVSS.n2811 DVSS.n2810 4.6505
R23750 DVSS.n2809 DVSS.n674 4.6505
R23751 DVSS.n2808 DVSS.n2807 4.6505
R23752 DVSS.n676 DVSS.n675 4.6505
R23753 DVSS.n2801 DVSS.n2800 4.6505
R23754 DVSS.n2799 DVSS.n682 4.6505
R23755 DVSS.n2798 DVSS.n2797 4.6505
R23756 DVSS.n689 DVSS.n684 4.6505
R23757 DVSS.n2790 DVSS.n2789 4.6505
R23758 DVSS.n2788 DVSS.n688 4.6505
R23759 DVSS.n696 DVSS.n691 4.6505
R23760 DVSS.n2783 DVSS.n2782 4.6505
R23761 DVSS.n697 DVSS.n695 4.6505
R23762 DVSS.n2776 DVSS.n703 4.6505
R23763 DVSS.n2775 DVSS.n2774 4.6505
R23764 DVSS.n1905 DVSS.n1866 4.6505
R23765 DVSS.n1913 DVSS.n1912 4.6505
R23766 DVSS.n1910 DVSS.n1867 4.6505
R23767 DVSS.n1908 DVSS.n1907 4.6505
R23768 DVSS.n1802 DVSS.n1801 4.6505
R23769 DVSS.n1929 DVSS.n1928 4.6505
R23770 DVSS.n1920 DVSS.n1803 4.6505
R23771 DVSS.n1922 DVSS.n1921 4.6505
R23772 DVSS.n1919 DVSS.n1796 4.6505
R23773 DVSS.n1935 DVSS.n1795 4.6505
R23774 DVSS.n1942 DVSS.n1936 4.6505
R23775 DVSS.n3088 DVSS.n4 4.6505
R23776 DVSS.n3086 DVSS.n3085 4.6505
R23777 DVSS.n6 DVSS.n5 4.6505
R23778 DVSS.n3079 DVSS.n3078 4.6505
R23779 DVSS.n3076 DVSS.n11 4.6505
R23780 DVSS.n3077 DVSS.n13 4.6505
R23781 DVSS.n3075 DVSS.n13 4.6505
R23782 DVSS.n13 DVSS.n12 4.6505
R23783 DVSS.n626 DVSS.n1 4.6505
R23784 DVSS.n2865 DVSS.n2864 4.6505
R23785 DVSS.n2863 DVSS.n627 4.6505
R23786 DVSS.n2861 DVSS.n2860 4.6505
R23787 DVSS.n1826 DVSS.n629 4.6505
R23788 DVSS.n2862 DVSS.n628 4.6505
R23789 DVSS.n1825 DVSS.n628 4.6505
R23790 DVSS.n1827 DVSS.n628 4.6505
R23791 DVSS.n1830 DVSS.n1829 4.6505
R23792 DVSS.n1855 DVSS.n1854 4.6505
R23793 DVSS.n1855 DVSS.n1817 4.6505
R23794 DVSS.n1844 DVSS.n1815 4.6505
R23795 DVSS.n1842 DVSS.n1815 4.6505
R23796 DVSS.n1858 DVSS.n1857 4.6505
R23797 DVSS.n1857 DVSS.n638 4.6505
R23798 DVSS.n648 DVSS.n646 4.6505
R23799 DVSS.n656 DVSS.n651 4.6505
R23800 DVSS.n2838 DVSS.n2837 4.6505
R23801 DVSS.n2839 DVSS.n644 4.6505
R23802 DVSS.n2841 DVSS.n2840 4.6505
R23803 DVSS.n645 DVSS.n640 4.6505
R23804 DVSS.n2848 DVSS.n2847 4.6505
R23805 DVSS.n2849 DVSS.n637 4.6505
R23806 DVSS.n2851 DVSS.n2850 4.6505
R23807 DVSS.n1813 DVSS.n636 4.6505
R23808 DVSS.n1860 DVSS.n1859 4.6505
R23809 DVSS.n1812 DVSS.n1811 4.6505
R23810 DVSS.n1843 DVSS.n1840 4.6505
R23811 DVSS.n1846 DVSS.n1845 4.6505
R23812 DVSS.n1841 DVSS.n1820 4.6505
R23813 DVSS.n1853 DVSS.n1852 4.6505
R23814 DVSS.n1819 DVSS.n1818 4.6505
R23815 DVSS.n1834 DVSS.n1833 4.6505
R23816 DVSS.n1832 DVSS.n1824 4.6505
R23817 DVSS.n2830 DVSS.n2829 4.6505
R23818 DVSS.n2423 DVSS.n2422 4.6505
R23819 DVSS.n1787 DVSS.n1786 4.6505
R23820 DVSS.n2431 DVSS.n2430 4.6505
R23821 DVSS.n2432 DVSS.n1784 4.6505
R23822 DVSS.n2437 DVSS.n2436 4.6505
R23823 DVSS.n2434 DVSS.n2433 4.6505
R23824 DVSS.n2434 DVSS.n1785 4.6505
R23825 DVSS.n2435 DVSS.n2434 4.6505
R23826 DVSS.n2493 DVSS.n2490 4.6505
R23827 DVSS.n2473 DVSS.n2472 4.6505
R23828 DVSS.n2473 DVSS.n1773 4.6505
R23829 DVSS.n2462 DVSS.n1771 4.6505
R23830 DVSS.n2460 DVSS.n1771 4.6505
R23831 DVSS.n2475 DVSS.n1769 4.6505
R23832 DVSS.n2476 DVSS.n2475 4.6505
R23833 DVSS.n2443 DVSS.n2442 4.6505
R23834 DVSS.n2444 DVSS.n1781 4.6505
R23835 DVSS.n2446 DVSS.n2445 4.6505
R23836 DVSS.n1775 DVSS.n1774 4.6505
R23837 DVSS.n2471 DVSS.n2470 4.6505
R23838 DVSS.n2452 DVSS.n1776 4.6505
R23839 DVSS.n2464 DVSS.n2463 4.6505
R23840 DVSS.n2461 DVSS.n2451 4.6505
R23841 DVSS.n2459 DVSS.n2458 4.6505
R23842 DVSS.n2453 DVSS.n1768 4.6505
R23843 DVSS.n2478 DVSS.n2477 4.6505
R23844 DVSS.n1765 DVSS.n1764 4.6505
R23845 DVSS.n2486 DVSS.n2485 4.6505
R23846 DVSS.n2487 DVSS.n1763 4.6505
R23847 DVSS.n2495 DVSS.n2494 4.6505
R23848 DVSS.n1760 DVSS.n1759 4.6505
R23849 DVSS.n2503 DVSS.n2502 4.6505
R23850 DVSS.n2504 DVSS.n1757 4.6505
R23851 DVSS.n2513 DVSS.n2512 4.6505
R23852 DVSS.n2511 DVSS.n1758 4.6505
R23853 DVSS.n3062 DVSS.n3057 4.6505
R23854 DVSS.n3065 DVSS.n3064 4.6505
R23855 DVSS.n3058 DVSS.n17 4.6505
R23856 DVSS.n3071 DVSS.n18 4.6505
R23857 DVSS.n3073 DVSS.n3072 4.6505
R23858 DVSS.n3063 DVSS.n3060 4.6505
R23859 DVSS.n3061 DVSS.n3060 4.6505
R23860 DVSS.n3060 DVSS.n3059 4.6505
R23861 DVSS.n2524 DVSS.n1273 4.6505
R23862 DVSS.n2528 DVSS.n2527 4.6505
R23863 DVSS.n1267 DVSS.n1266 4.6505
R23864 DVSS.n2536 DVSS.n2535 4.6505
R23865 DVSS.n1268 DVSS.n1264 4.6505
R23866 DVSS.n2538 DVSS.n2537 4.6505
R23867 DVSS.n2538 DVSS.n1265 4.6505
R23868 DVSS.n2539 DVSS.n2538 4.6505
R23869 DVSS.n2540 DVSS.n1263 4.6505
R23870 DVSS.n2553 DVSS.n2552 4.6505
R23871 DVSS.n2589 DVSS.n1237 4.6505
R23872 DVSS.n2543 DVSS.n2542 4.6505
R23873 DVSS.n2560 DVSS.n2559 4.6505
R23874 DVSS.n2559 DVSS.n2558 4.6505
R23875 DVSS.n2574 DVSS.n2573 4.6505
R23876 DVSS.n2575 DVSS.n2574 4.6505
R23877 DVSS.n2552 DVSS.n2551 4.6505
R23878 DVSS.n2606 DVSS.n2603 4.6505
R23879 DVSS.n2602 DVSS.n1231 4.6505
R23880 DVSS.n2601 DVSS.n2600 4.6505
R23881 DVSS.n1233 DVSS.n1232 4.6505
R23882 DVSS.n2593 DVSS.n2592 4.6505
R23883 DVSS.n2586 DVSS.n1236 4.6505
R23884 DVSS.n2585 DVSS.n2584 4.6505
R23885 DVSS.n1239 DVSS.n1238 4.6505
R23886 DVSS.n2577 DVSS.n2576 4.6505
R23887 DVSS.n1244 DVSS.n1243 4.6505
R23888 DVSS.n2572 DVSS.n2571 4.6505
R23889 DVSS.n1247 DVSS.n1246 4.6505
R23890 DVSS.n2556 DVSS.n2555 4.6505
R23891 DVSS.n2562 DVSS.n2561 4.6505
R23892 DVSS.n2563 DVSS.n2554 4.6505
R23893 DVSS.n1256 DVSS.n1255 4.6505
R23894 DVSS.n2550 DVSS.n2549 4.6505
R23895 DVSS.n1259 DVSS.n1258 4.6505
R23896 DVSS.n731 DVSS.n730 4.6505
R23897 DVSS.n2740 DVSS.n2739 4.6505
R23898 DVSS.n735 DVSS.n734 4.6505
R23899 DVSS.n2735 DVSS.n2734 4.6505
R23900 DVSS.n739 DVSS.n738 4.6505
R23901 DVSS.n2728 DVSS.n2727 4.6505
R23902 DVSS.n2723 DVSS.n743 4.6505
R23903 DVSS.n2722 DVSS.n2721 4.6505
R23904 DVSS.n746 DVSS.n745 4.6505
R23905 DVSS.n2714 DVSS.n2713 4.6505
R23906 DVSS.n2712 DVSS.n751 4.6505
R23907 DVSS.n2685 DVSS.n2664 4.6505
R23908 DVSS.n2684 DVSS.n2683 4.6505
R23909 DVSS.n2667 DVSS.n2666 4.6505
R23910 DVSS.n2677 DVSS.n2676 4.6505
R23911 DVSS.n2674 DVSS.n2673 4.6505
R23912 DVSS.n3050 DVSS.n27 4.6505
R23913 DVSS.n3049 DVSS.n3048 4.6505
R23914 DVSS.n29 DVSS.n28 4.6505
R23915 DVSS.n3044 DVSS.n3043 4.6505
R23916 DVSS.n33 DVSS.n32 4.6505
R23917 DVSS.n565 DVSS.n564 4.6505
R23918 DVSS.n566 DVSS.n559 4.6505
R23919 DVSS.n570 DVSS.n569 4.6505
R23920 DVSS.n558 DVSS.n557 4.6505
R23921 DVSS.n575 DVSS.n574 4.6505
R23922 DVSS.n554 DVSS.n553 4.6505
R23923 DVSS.n583 DVSS.n582 4.6505
R23924 DVSS.n584 DVSS.n550 4.6505
R23925 DVSS.n594 DVSS.n593 4.6505
R23926 DVSS.n592 DVSS.n551 4.6505
R23927 DVSS.n591 DVSS.n548 4.6505
R23928 DVSS.n590 DVSS.n545 4.6505
R23929 DVSS.n604 DVSS.n546 4.6505
R23930 DVSS.n2638 DVSS.n2629 4.6505
R23931 DVSS.n2637 DVSS.n2636 4.6505
R23932 DVSS.n2630 DVSS.n45 4.6505
R23933 DVSS.n3035 DVSS.n3034 4.6505
R23934 DVSS.n3033 DVSS.n46 4.6505
R23935 DVSS.n51 DVSS.n48 4.6505
R23936 DVSS.n3028 DVSS.n3027 4.6505
R23937 DVSS.n52 DVSS.n50 4.6505
R23938 DVSS.n3020 DVSS.n58 4.6505
R23939 DVSS.n3019 DVSS.n3018 4.6505
R23940 DVSS.n3017 DVSS.n59 4.6505
R23941 DVSS.n2991 DVSS.n2889 4.6505
R23942 DVSS.n2994 DVSS.n2993 4.6505
R23943 DVSS.n2995 DVSS.n2888 4.6505
R23944 DVSS.n2998 DVSS.n2996 4.6505
R23945 DVSS.n3000 DVSS.n2886 4.6505
R23946 DVSS.n3003 DVSS.n3002 4.6505
R23947 DVSS.n2986 DVSS.n2891 4.6505
R23948 DVSS.n2967 DVSS.n2894 4.6505
R23949 DVSS.n2972 DVSS.n2969 4.6505
R23950 DVSS.n2973 DVSS.n2893 4.6505
R23951 DVSS.n2977 DVSS.n2976 4.6505
R23952 DVSS.n2978 DVSS.n2892 4.6505
R23953 DVSS.n2985 DVSS.n2982 4.6505
R23954 DVSS.n2928 DVSS.n2926 4.6505
R23955 DVSS.n2926 DVSS.n2906 4.6505
R23956 DVSS.n2954 DVSS.n2952 4.6505
R23957 DVSS.n2955 DVSS.n2954 4.6505
R23958 DVSS.n2917 DVSS.n2916 4.6505
R23959 DVSS.n2911 DVSS.n2910 4.6505
R23960 DVSS.n2924 DVSS.n2923 4.6505
R23961 DVSS.n2925 DVSS.n2909 4.6505
R23962 DVSS.n2930 DVSS.n2929 4.6505
R23963 DVSS.n2927 DVSS.n2907 4.6505
R23964 DVSS.n2937 DVSS.n2936 4.6505
R23965 DVSS.n2938 DVSS.n2905 4.6505
R23966 DVSS.n2943 DVSS.n2942 4.6505
R23967 DVSS.n2903 DVSS.n2902 4.6505
R23968 DVSS.n2950 DVSS.n2949 4.6505
R23969 DVSS.n2951 DVSS.n2901 4.6505
R23970 DVSS.n2957 DVSS.n2956 4.6505
R23971 DVSS.n2899 DVSS.n2898 4.6505
R23972 DVSS.n2963 DVSS.n2962 4.6505
R23973 DVSS.n413 DVSS.n181 4.5005
R23974 DVSS.n72 DVSS.n63 4.5005
R23975 DVSS.n541 DVSS.n540 4.5005
R23976 DVSS.n608 DVSS.n69 4.5005
R23977 DVSS.n2286 DVSS.n2054 4.5005
R23978 DVSS.n2414 DVSS.n2413 4.5005
R23979 DVSS.n1938 DVSS.n1791 4.5005
R23980 DVSS.n1094 DVSS.n862 4.5005
R23981 DVSS.n1221 DVSS.n757 4.5005
R23982 DVSS.n2701 DVSS.n755 4.5005
R23983 DVSS.n1616 DVSS.n1384 4.5005
R23984 DVSS.n1744 DVSS.n1743 4.5005
R23985 DVSS.n1276 DVSS.n708 4.5005
R23986 DVSS.n2825 DVSS.n658 4.5005
R23987 DVSS.n2506 DVSS.n1748 4.5005
R23988 DVSS.n2696 DVSS.n2695 4.5005
R23989 DVSS.n419 DVSS.n418 4.40783
R23990 DVSS.n2292 DVSS.n2291 4.40783
R23991 DVSS.n1100 DVSS.n1099 4.40783
R23992 DVSS.n1622 DVSS.n1621 4.40783
R23993 DVSS.n2959 DVSS.n2958 4.35669
R23994 DVSS.n310 DVSS.n266 4.31208
R23995 DVSS.n2183 DVSS.n2139 4.31208
R23996 DVSS.n991 DVSS.n947 4.31208
R23997 DVSS.n1513 DVSS.n1469 4.31208
R23998 DVSS.n309 DVSS.n267 4.04261
R23999 DVSS.n2182 DVSS.n2140 4.04261
R24000 DVSS.n990 DVSS.n948 4.04261
R24001 DVSS.n1512 DVSS.n1470 4.04261
R24002 DVSS.n220 DVSS.n205 3.93153
R24003 DVSS.n199 DVSS.n184 3.93153
R24004 DVSS.n2093 DVSS.n2078 3.93153
R24005 DVSS.n2072 DVSS.n2057 3.93153
R24006 DVSS.n901 DVSS.n886 3.93153
R24007 DVSS.n880 DVSS.n865 3.93153
R24008 DVSS.n1423 DVSS.n1408 3.93153
R24009 DVSS.n1402 DVSS.n1387 3.93153
R24010 DVSS.n266 DVSS.n253 3.8405
R24011 DVSS.n2139 DVSS.n2126 3.8405
R24012 DVSS.n947 DVSS.n934 3.8405
R24013 DVSS.n1469 DVSS.n1456 3.8405
R24014 DVSS.n306 DVSS.n305 3.77313
R24015 DVSS.n2179 DVSS.n2178 3.77313
R24016 DVSS.n987 DVSS.n986 3.77313
R24017 DVSS.n1509 DVSS.n1508 3.77313
R24018 DVSS.n3004 DVSS.n2885 3.69566
R24019 DVSS.n2915 DVSS.n2913 3.69563
R24020 DVSS.n2659 DVSS.n2613 3.69446
R24021 DVSS.n1881 DVSS.n1879 3.69446
R24022 DVSS.n2762 DVSS.n717 3.69446
R24023 DVSS.n664 DVSS.n662 3.69446
R24024 DVSS.n2559 DVSS.n1245 3.68864
R24025 DVSS.n562 DVSS.n31 3.68864
R24026 DVSS.n3031 DVSS.n49 3.68864
R24027 DVSS.n2474 DVSS.n1771 3.68864
R24028 DVSS.n1856 DVSS.n1815 3.68864
R24029 DVSS.n1932 DVSS.n1931 3.68864
R24030 DVSS.n2725 DVSS.n736 3.68864
R24031 DVSS.n2786 DVSS.n694 3.68864
R24032 DVSS.n276 DVSS.n272 3.50366
R24033 DVSS.n2149 DVSS.n2145 3.50366
R24034 DVSS.n957 DVSS.n953 3.50366
R24035 DVSS.n1479 DVSS.n1475 3.50366
R24036 DVSS.n300 DVSS.n278 3.23418
R24037 DVSS.n2173 DVSS.n2151 3.23418
R24038 DVSS.n981 DVSS.n959 3.23418
R24039 DVSS.n1503 DVSS.n1481 3.23418
R24040 DVSS.n414 DVSS.n412 3.20387
R24041 DVSS.n2287 DVSS.n2285 3.20387
R24042 DVSS.n1095 DVSS.n1093 3.20387
R24043 DVSS.n1617 DVSS.n1615 3.20387
R24044 DVSS.n613 DVSS.n612 3.03311
R24045 DVSS.n1279 DVSS.n711 3.03311
R24046 DVSS.n1949 DVSS.n1948 3.03311
R24047 DVSS.n2824 DVSS.n659 3.03311
R24048 DVSS.n2521 DVSS.n2520 3.03311
R24049 DVSS.n2694 DVSS.n1226 3.03311
R24050 DVSS.n2706 DVSS.n2705 3.03311
R24051 DVSS.n76 DVSS.n75 3.03311
R24052 DVSS.n299 DVSS.n282 2.96471
R24053 DVSS.n2172 DVSS.n2155 2.96471
R24054 DVSS.n980 DVSS.n963 2.96471
R24055 DVSS.n1502 DVSS.n1485 2.96471
R24056 DVSS.n2590 DVSS.n2589 2.84494
R24057 DVSS.n588 DVSS.n587 2.84494
R24058 DVSS.n2491 DVSS.n2490 2.84494
R24059 DVSS.n649 DVSS.n648 2.84494
R24060 DVSS DVSS.n3074 2.78465
R24061 DVSS.n296 DVSS.n295 2.69524
R24062 DVSS.n2169 DVSS.n2168 2.69524
R24063 DVSS.n977 DVSS.n976 2.69524
R24064 DVSS.n1499 DVSS.n1498 2.69524
R24065 DVSS.n388 DVSS.n387 2.5605
R24066 DVSS.n2261 DVSS.n2260 2.5605
R24067 DVSS.n1069 DVSS.n1068 2.5605
R24068 DVSS.n1591 DVSS.n1590 2.5605
R24069 DVSS.n291 DVSS.n285 2.42576
R24070 DVSS.n291 DVSS.n259 2.42576
R24071 DVSS.n2164 DVSS.n2158 2.42576
R24072 DVSS.n2164 DVSS.n2132 2.42576
R24073 DVSS.n972 DVSS.n966 2.42576
R24074 DVSS.n972 DVSS.n940 2.42576
R24075 DVSS.n1494 DVSS.n1488 2.42576
R24076 DVSS.n1494 DVSS.n1462 2.42576
R24077 DVSS.n2524 DVSS.n2523 2.38846
R24078 DVSS.n61 DVSS.n60 2.31469
R24079 DVSS.n1934 DVSS.n1933 2.31469
R24080 DVSS.n753 DVSS.n752 2.31469
R24081 DVSS.n706 DVSS.n705 2.31469
R24082 DVSS.n249 DVSS.n243 2.29103
R24083 DVSS.n2122 DVSS.n2116 2.29103
R24084 DVSS.n930 DVSS.n924 2.29103
R24085 DVSS.n1452 DVSS.n1446 2.29103
R24086 DVSS.n2420 DVSS.n2419 2.24741
R24087 DVSS.n2698 DVSS.n1223 2.24741
R24088 DVSS.n2522 DVSS.n1274 2.24725
R24089 DVSS.n74 DVSS.n71 2.24722
R24090 DVSS.n1790 DVSS.n1788 2.24722
R24091 DVSS.n2704 DVSS.n2703 2.24722
R24092 DVSS.n1278 DVSS.n1275 2.24722
R24093 DVSS.n611 DVSS.n610 2.24702
R24094 DVSS.n2419 DVSS.n2418 2.24626
R24095 DVSS.n73 DVSS.n71 2.24565
R24096 DVSS.n1789 DVSS.n1788 2.24565
R24097 DVSS.n2703 DVSS.n2702 2.24565
R24098 DVSS.n1277 DVSS.n1275 2.24565
R24099 DVSS.n295 DVSS.n285 2.15629
R24100 DVSS.n353 DVSS.n259 2.15629
R24101 DVSS.n2168 DVSS.n2158 2.15629
R24102 DVSS.n2226 DVSS.n2132 2.15629
R24103 DVSS.n976 DVSS.n966 2.15629
R24104 DVSS.n1034 DVSS.n940 2.15629
R24105 DVSS.n1498 DVSS.n1488 2.15629
R24106 DVSS.n1556 DVSS.n1462 2.15629
R24107 DVSS.n3089 DVSS.n3088 2.01072
R24108 DVSS.n3090 DVSS 1.96635
R24109 DVSS.n3074 DVSS.n3073 1.93608
R24110 DVSS.n296 DVSS.n282 1.88682
R24111 DVSS.n2169 DVSS.n2155 1.88682
R24112 DVSS.n977 DVSS.n963 1.88682
R24113 DVSS.n1499 DVSS.n1485 1.88682
R24114 DVSS.n387 DVSS.n385 1.68471
R24115 DVSS.n381 DVSS.n249 1.68471
R24116 DVSS.n2260 DVSS.n2258 1.68471
R24117 DVSS.n2254 DVSS.n2122 1.68471
R24118 DVSS.n1068 DVSS.n1066 1.68471
R24119 DVSS.n1062 DVSS.n930 1.68471
R24120 DVSS.n1590 DVSS.n1588 1.68471
R24121 DVSS.n1584 DVSS.n1452 1.68471
R24122 DVSS.n408 DVSS.n407 1.64728
R24123 DVSS.n2281 DVSS.n2280 1.64728
R24124 DVSS.n1089 DVSS.n1088 1.64728
R24125 DVSS.n1611 DVSS.n1610 1.64728
R24126 DVSS.n300 DVSS.n299 1.61734
R24127 DVSS.n2173 DVSS.n2172 1.61734
R24128 DVSS.n981 DVSS.n980 1.61734
R24129 DVSS.n1503 DVSS.n1502 1.61734
R24130 DVSS.n419 DVSS.n152 1.59464
R24131 DVSS.n426 DVSS.n152 1.59464
R24132 DVSS.n426 DVSS.n153 1.59464
R24133 DVSS.n422 DVSS.n153 1.59464
R24134 DVSS.n422 DVSS.n119 1.59464
R24135 DVSS.n436 DVSS.n119 1.59464
R24136 DVSS.n446 DVSS.n117 1.59464
R24137 DVSS.n441 DVSS.n105 1.59464
R24138 DVSS.n457 DVSS.n105 1.59464
R24139 DVSS.n458 DVSS.n457 1.59464
R24140 DVSS.n458 DVSS.n103 1.59464
R24141 DVSS.n464 DVSS.n463 1.59464
R24142 DVSS.n464 DVSS.n100 1.59464
R24143 DVSS.n494 DVSS.n100 1.59464
R24144 DVSS.n490 DVSS.n85 1.59464
R24145 DVSS.n528 DVSS.n85 1.59464
R24146 DVSS.n529 DVSS.n528 1.59464
R24147 DVSS.n530 DVSS.n529 1.59464
R24148 DVSS.n530 DVSS.n83 1.59464
R24149 DVSS.n534 DVSS.n83 1.59464
R24150 DVSS.n2292 DVSS.n2025 1.59464
R24151 DVSS.n2299 DVSS.n2025 1.59464
R24152 DVSS.n2299 DVSS.n2026 1.59464
R24153 DVSS.n2295 DVSS.n2026 1.59464
R24154 DVSS.n2295 DVSS.n1992 1.59464
R24155 DVSS.n2309 DVSS.n1992 1.59464
R24156 DVSS.n2319 DVSS.n1990 1.59464
R24157 DVSS.n2314 DVSS.n1978 1.59464
R24158 DVSS.n2330 DVSS.n1978 1.59464
R24159 DVSS.n2331 DVSS.n2330 1.59464
R24160 DVSS.n2331 DVSS.n1976 1.59464
R24161 DVSS.n2337 DVSS.n2336 1.59464
R24162 DVSS.n2337 DVSS.n1973 1.59464
R24163 DVSS.n2367 DVSS.n1973 1.59464
R24164 DVSS.n2363 DVSS.n1958 1.59464
R24165 DVSS.n2401 DVSS.n1958 1.59464
R24166 DVSS.n2402 DVSS.n2401 1.59464
R24167 DVSS.n2403 DVSS.n2402 1.59464
R24168 DVSS.n2403 DVSS.n1956 1.59464
R24169 DVSS.n2407 DVSS.n1956 1.59464
R24170 DVSS.n1100 DVSS.n833 1.59464
R24171 DVSS.n1107 DVSS.n833 1.59464
R24172 DVSS.n1107 DVSS.n834 1.59464
R24173 DVSS.n1103 DVSS.n834 1.59464
R24174 DVSS.n1103 DVSS.n800 1.59464
R24175 DVSS.n1117 DVSS.n800 1.59464
R24176 DVSS.n1127 DVSS.n798 1.59464
R24177 DVSS.n1122 DVSS.n786 1.59464
R24178 DVSS.n1138 DVSS.n786 1.59464
R24179 DVSS.n1139 DVSS.n1138 1.59464
R24180 DVSS.n1139 DVSS.n784 1.59464
R24181 DVSS.n1145 DVSS.n1144 1.59464
R24182 DVSS.n1145 DVSS.n781 1.59464
R24183 DVSS.n1175 DVSS.n781 1.59464
R24184 DVSS.n1171 DVSS.n766 1.59464
R24185 DVSS.n1209 DVSS.n766 1.59464
R24186 DVSS.n1210 DVSS.n1209 1.59464
R24187 DVSS.n1211 DVSS.n1210 1.59464
R24188 DVSS.n1211 DVSS.n764 1.59464
R24189 DVSS.n1215 DVSS.n764 1.59464
R24190 DVSS.n1622 DVSS.n1355 1.59464
R24191 DVSS.n1629 DVSS.n1355 1.59464
R24192 DVSS.n1629 DVSS.n1356 1.59464
R24193 DVSS.n1625 DVSS.n1356 1.59464
R24194 DVSS.n1625 DVSS.n1322 1.59464
R24195 DVSS.n1639 DVSS.n1322 1.59464
R24196 DVSS.n1649 DVSS.n1320 1.59464
R24197 DVSS.n1644 DVSS.n1308 1.59464
R24198 DVSS.n1660 DVSS.n1308 1.59464
R24199 DVSS.n1661 DVSS.n1660 1.59464
R24200 DVSS.n1661 DVSS.n1306 1.59464
R24201 DVSS.n1667 DVSS.n1666 1.59464
R24202 DVSS.n1667 DVSS.n1303 1.59464
R24203 DVSS.n1697 DVSS.n1303 1.59464
R24204 DVSS.n1693 DVSS.n1288 1.59464
R24205 DVSS.n1731 DVSS.n1288 1.59464
R24206 DVSS.n1732 DVSS.n1731 1.59464
R24207 DVSS.n1733 DVSS.n1732 1.59464
R24208 DVSS.n1733 DVSS.n1286 1.59464
R24209 DVSS.n1737 DVSS.n1286 1.59464
R24210 DVSS.n236 DVSS.n225 1.54748
R24211 DVSS.n2109 DVSS.n2098 1.54748
R24212 DVSS.n917 DVSS.n906 1.54748
R24213 DVSS.n1439 DVSS.n1428 1.54748
R24214 DVSS.n206 DVSS.n204 1.50638
R24215 DVSS.n185 DVSS.n183 1.50638
R24216 DVSS.n2079 DVSS.n2077 1.50638
R24217 DVSS.n2058 DVSS.n2056 1.50638
R24218 DVSS.n887 DVSS.n885 1.50638
R24219 DVSS.n866 DVSS.n864 1.50638
R24220 DVSS.n1409 DVSS.n1407 1.50638
R24221 DVSS.n1388 DVSS.n1386 1.50638
R24222 DVSS.n2698 DVSS.n2697 1.49558
R24223 DVSS.n2505 DVSS.n1274 1.49528
R24224 DVSS.n610 DVSS.n609 1.49482
R24225 DVSS.n463 DVSS.n462 1.45398
R24226 DVSS.n2336 DVSS.n2335 1.45398
R24227 DVSS.n1144 DVSS.n1143 1.45398
R24228 DVSS.n1666 DVSS.n1665 1.45398
R24229 DVSS.n213 DVSS.n212 1.45108
R24230 DVSS.n192 DVSS.n191 1.45108
R24231 DVSS.n2086 DVSS.n2085 1.45108
R24232 DVSS.n2065 DVSS.n2064 1.45108
R24233 DVSS.n894 DVSS.n893 1.45108
R24234 DVSS.n873 DVSS.n872 1.45108
R24235 DVSS.n1416 DVSS.n1415 1.45108
R24236 DVSS.n1395 DVSS.n1394 1.45108
R24237 DVSS.n401 DVSS.n237 1.44767
R24238 DVSS.n2274 DVSS.n2110 1.44767
R24239 DVSS.n1082 DVSS.n918 1.44767
R24240 DVSS.n1604 DVSS.n1440 1.44767
R24241 DVSS.n2964 DVSS 1.39202
R24242 DVSS DVSS.n2964 1.39044
R24243 DVSS.n400 DVSS.n239 1.34787
R24244 DVSS.n278 DVSS.n276 1.34787
R24245 DVSS.n2273 DVSS.n2112 1.34787
R24246 DVSS.n2151 DVSS.n2149 1.34787
R24247 DVSS.n1081 DVSS.n920 1.34787
R24248 DVSS.n959 DVSS.n957 1.34787
R24249 DVSS.n1603 DVSS.n1442 1.34787
R24250 DVSS.n1481 DVSS.n1479 1.34787
R24251 DVSS.n442 DVSS.n441 1.26643
R24252 DVSS.n2315 DVSS.n2314 1.26643
R24253 DVSS.n1123 DVSS.n1122 1.26643
R24254 DVSS.n1645 DVSS.n1644 1.26643
R24255 DVSS.n2671 DVSS 1.2505
R24256 DVSS.n397 DVSS.n396 1.24806
R24257 DVSS.n2270 DVSS.n2269 1.24806
R24258 DVSS.n1078 DVSS.n1077 1.24806
R24259 DVSS.n1600 DVSS.n1599 1.24806
R24260 DVSS.n1831 DVSS 1.15435
R24261 DVSS.n394 DVSS.n393 1.14826
R24262 DVSS.n2267 DVSS.n2266 1.14826
R24263 DVSS.n1075 DVSS.n1074 1.14826
R24264 DVSS.n1597 DVSS.n1596 1.14826
R24265 DVSS.n2541 DVSS 1.13383
R24266 DVSS.n3015 DVSS.n3014 1.12991
R24267 DVSS.n1941 DVSS.n1937 1.12991
R24268 DVSS.n2710 DVSS.n2709 1.12991
R24269 DVSS.n2771 DVSS.n2770 1.12991
R24270 DVSS.n2416 DVSS.n2415 1.10812
R24271 DVSS.n543 DVSS.n542 1.10762
R24272 DVSS.n2700 DVSS.n2699 1.10762
R24273 DVSS.n1746 DVSS.n1745 1.10762
R24274 DVSS.n388 DVSS.n246 1.07839
R24275 DVSS.n305 DVSS.n272 1.07839
R24276 DVSS.n2261 DVSS.n2119 1.07839
R24277 DVSS.n2178 DVSS.n2145 1.07839
R24278 DVSS.n1069 DVSS.n927 1.07839
R24279 DVSS.n986 DVSS.n953 1.07839
R24280 DVSS.n1591 DVSS.n1449 1.07839
R24281 DVSS.n1508 DVSS.n1475 1.07839
R24282 DVSS.n391 DVSS.n242 0.973599
R24283 DVSS.n2264 DVSS.n2115 0.973599
R24284 DVSS.n1072 DVSS.n923 0.973599
R24285 DVSS.n1594 DVSS.n1445 0.973599
R24286 DVSS.n306 DVSS.n267 0.808921
R24287 DVSS.n2179 DVSS.n2140 0.808921
R24288 DVSS.n987 DVSS.n948 0.808921
R24289 DVSS.n1509 DVSS.n1470 0.808921
R24290 DVSS.n606 DVSS.n605 0.753441
R24291 DVSS.n219 DVSS.n218 0.753441
R24292 DVSS.n210 DVSS.n207 0.753441
R24293 DVSS.n198 DVSS.n197 0.753441
R24294 DVSS.n189 DVSS.n186 0.753441
R24295 DVSS.n2092 DVSS.n2091 0.753441
R24296 DVSS.n2083 DVSS.n2080 0.753441
R24297 DVSS.n2071 DVSS.n2070 0.753441
R24298 DVSS.n2062 DVSS.n2059 0.753441
R24299 DVSS.n2826 DVSS.n655 0.753441
R24300 DVSS.n900 DVSS.n899 0.753441
R24301 DVSS.n891 DVSS.n888 0.753441
R24302 DVSS.n879 DVSS.n878 0.753441
R24303 DVSS.n870 DVSS.n867 0.753441
R24304 DVSS.n2605 DVSS.n1225 0.753441
R24305 DVSS.n2509 DVSS.n2508 0.753441
R24306 DVSS.n1422 DVSS.n1421 0.753441
R24307 DVSS.n1413 DVSS.n1410 0.753441
R24308 DVSS.n1401 DVSS.n1400 0.753441
R24309 DVSS.n1392 DVSS.n1389 0.753441
R24310 DVSS.n393 DVSS.n391 0.649233
R24311 DVSS.n2266 DVSS.n2264 0.649233
R24312 DVSS.n1074 DVSS.n1072 0.649233
R24313 DVSS.n1596 DVSS.n1594 0.649233
R24314 DVSS.n385 DVSS.n243 0.606816
R24315 DVSS.n2258 DVSS.n2116 0.606816
R24316 DVSS.n1066 DVSS.n924 0.606816
R24317 DVSS.n1588 DVSS.n1446 0.606816
R24318 DVSS.n418 DVSS.n417 0.563137
R24319 DVSS.n2291 DVSS.n2290 0.563137
R24320 DVSS.n1099 DVSS.n1098 0.563137
R24321 DVSS.n1621 DVSS.n1620 0.563137
R24322 DVSS.n396 DVSS.n394 0.549428
R24323 DVSS.n2269 DVSS.n2267 0.549428
R24324 DVSS.n1077 DVSS.n1075 0.549428
R24325 DVSS.n1599 DVSS.n1597 0.549428
R24326 DVSS.n310 DVSS.n309 0.539447
R24327 DVSS.n2183 DVSS.n2182 0.539447
R24328 DVSS.n991 DVSS.n990 0.539447
R24329 DVSS.n1513 DVSS.n1512 0.539447
R24330 DVSS.n2916 DVSS.n2915 0.526461
R24331 DVSS.n3004 DVSS.n3003 0.526088
R24332 DVSS.n2659 DVSS.n2658 0.502212
R24333 DVSS.n1882 DVSS.n1881 0.502212
R24334 DVSS.n719 DVSS.n717 0.502212
R24335 DVSS.n669 DVSS.n662 0.502212
R24336 DVSS.n397 DVSS.n239 0.449623
R24337 DVSS.n2270 DVSS.n2112 0.449623
R24338 DVSS.n1078 DVSS.n920 0.449623
R24339 DVSS.n1600 DVSS.n1442 0.449623
R24340 DVSS.n1752 DVSS.n713 0.441318
R24341 DVSS.n401 DVSS.n400 0.349818
R24342 DVSS.n246 DVSS.n245 0.349818
R24343 DVSS.n2274 DVSS.n2273 0.349818
R24344 DVSS.n2119 DVSS.n2118 0.349818
R24345 DVSS.n1082 DVSS.n1081 0.349818
R24346 DVSS.n927 DVSS.n926 0.349818
R24347 DVSS.n1604 DVSS.n1603 0.349818
R24348 DVSS.n1449 DVSS.n1448 0.349818
R24349 DVSS.n410 DVSS.n222 0.337926
R24350 DVSS.n412 DVSS.n201 0.337926
R24351 DVSS.n2283 DVSS.n2095 0.337926
R24352 DVSS.n2285 DVSS.n2074 0.337926
R24353 DVSS.n1091 DVSS.n903 0.337926
R24354 DVSS.n1093 DVSS.n882 0.337926
R24355 DVSS.n1613 DVSS.n1425 0.337926
R24356 DVSS.n1615 DVSS.n1404 0.337926
R24357 DVSS.n442 DVSS.n117 0.328705
R24358 DVSS.n2315 DVSS.n1990 0.328705
R24359 DVSS.n1123 DVSS.n798 0.328705
R24360 DVSS.n1645 DVSS.n1320 0.328705
R24361 DVSS.n2523 DVSS 0.316512
R24362 DVSS DVSS.n3090 0.300422
R24363 DVSS.n489 DVSS.n101 0.281819
R24364 DVSS.n2362 DVSS.n1974 0.281819
R24365 DVSS.n1170 DVSS.n782 0.281819
R24366 DVSS.n1692 DVSS.n1304 0.281819
R24367 DVSS.n3089 DVSS.n3 0.256648
R24368 DVSS.n237 DVSS.n236 0.250013
R24369 DVSS.n2110 DVSS.n2109 0.250013
R24370 DVSS.n918 DVSS.n917 0.250013
R24371 DVSS.n1440 DVSS.n1439 0.250013
R24372 DVSS DVSS.n539 0.249718
R24373 DVSS DVSS.n2412 0.249718
R24374 DVSS DVSS.n1220 0.249718
R24375 DVSS DVSS.n1742 0.249718
R24376 DVSS.n144 DVSS.n116 0.234932
R24377 DVSS.n2017 DVSS.n1989 0.234932
R24378 DVSS.n825 DVSS.n797 0.234932
R24379 DVSS.n1347 DVSS.n1319 0.234932
R24380 DVSS.n2526 DVSS.n14 0.213615
R24381 DVSS.n3074 DVSS.n14 0.211531
R24382 DVSS.n410 DVSS.n409 0.198603
R24383 DVSS.n2283 DVSS.n2282 0.198603
R24384 DVSS.n1091 DVSS.n1090 0.198603
R24385 DVSS.n1613 DVSS.n1612 0.198603
R24386 DVSS.n412 DVSS.n411 0.196998
R24387 DVSS.n2285 DVSS.n2284 0.196998
R24388 DVSS.n1093 DVSS.n1092 0.196998
R24389 DVSS.n1615 DVSS.n1614 0.196998
R24390 DVSS.n657 DVSS 0.18712
R24391 DVSS.n0 DVSS 0.17755
R24392 DVSS.n3006 DVSS.n2879 0.156029
R24393 DVSS.n3006 DVSS.n2881 0.156029
R24394 DVSS.n3006 DVSS.n2883 0.156029
R24395 DVSS.n3006 DVSS.n2871 0.153643
R24396 DVSS.n2961 DVSS.n618 0.153643
R24397 DVSS.n2441 DVSS.n2440 0.151309
R24398 DVSS.n2707 DVSS.n756 0.151309
R24399 DVSS.n2672 DVSS.n22 0.151309
R24400 DVSS.n2919 DVSS.n620 0.151309
R24401 DVSS.n1828 DVSS.n631 0.151294
R24402 DVSS.n2767 DVSS.n710 0.151294
R24403 DVSS.n3006 DVSS.n2874 0.151294
R24404 DVSS.n3006 DVSS.n2875 0.151294
R24405 DVSS.n3006 DVSS.n2876 0.151294
R24406 DVSS.n3006 DVSS.n2877 0.151294
R24407 DVSS.n2921 DVSS.n620 0.151294
R24408 DVSS.n2932 DVSS.n620 0.151294
R24409 DVSS.n2934 DVSS.n620 0.151294
R24410 DVSS.n2945 DVSS.n620 0.151294
R24411 DVSS.n2947 DVSS.n620 0.151294
R24412 DVSS.n407 DVSS.n225 0.150208
R24413 DVSS.n2280 DVSS.n2098 0.150208
R24414 DVSS.n1088 DVSS.n906 0.150208
R24415 DVSS.n1610 DVSS.n1428 0.150208
R24416 DVSS.n540 DVSS 0.147302
R24417 DVSS.n2413 DVSS 0.147302
R24418 DVSS.n1221 DVSS 0.147302
R24419 DVSS.n1743 DVSS 0.147302
R24420 DVSS.n2687 DVSS 0.146353
R24421 DVSS.n2422 DVSS 0.143808
R24422 DVSS.n462 DVSS.n103 0.141159
R24423 DVSS.n2335 DVSS.n1976 0.141159
R24424 DVSS.n1143 DVSS.n784 0.141159
R24425 DVSS.n1665 DVSS.n1306 0.141159
R24426 DVSS.n3090 DVSS.n0 0.126683
R24427 DVSS.n534 DVSS.n78 0.0942729
R24428 DVSS.n2407 DVSS.n1951 0.0942729
R24429 DVSS.n1215 DVSS.n759 0.0942729
R24430 DVSS.n1737 DVSS.n1281 0.0942729
R24431 DVSS.n409 DVSS.n223 0.0932835
R24432 DVSS.n240 DVSS.n223 0.0932835
R24433 DVSS.n399 DVSS.n240 0.0932835
R24434 DVSS.n399 DVSS.n398 0.0932835
R24435 DVSS.n398 DVSS.n241 0.0932835
R24436 DVSS.n390 DVSS.n241 0.0932835
R24437 DVSS.n390 DVSS.n389 0.0932835
R24438 DVSS.n308 DVSS.n202 0.0932835
R24439 DVSS.n308 DVSS.n307 0.0932835
R24440 DVSS.n307 DVSS.n268 0.0932835
R24441 DVSS.n283 DVSS.n268 0.0932835
R24442 DVSS.n298 DVSS.n283 0.0932835
R24443 DVSS.n298 DVSS.n297 0.0932835
R24444 DVSS.n297 DVSS.n284 0.0932835
R24445 DVSS.n2282 DVSS.n2096 0.0932835
R24446 DVSS.n2113 DVSS.n2096 0.0932835
R24447 DVSS.n2272 DVSS.n2113 0.0932835
R24448 DVSS.n2272 DVSS.n2271 0.0932835
R24449 DVSS.n2271 DVSS.n2114 0.0932835
R24450 DVSS.n2263 DVSS.n2114 0.0932835
R24451 DVSS.n2263 DVSS.n2262 0.0932835
R24452 DVSS.n2181 DVSS.n2075 0.0932835
R24453 DVSS.n2181 DVSS.n2180 0.0932835
R24454 DVSS.n2180 DVSS.n2141 0.0932835
R24455 DVSS.n2156 DVSS.n2141 0.0932835
R24456 DVSS.n2171 DVSS.n2156 0.0932835
R24457 DVSS.n2171 DVSS.n2170 0.0932835
R24458 DVSS.n2170 DVSS.n2157 0.0932835
R24459 DVSS.n1090 DVSS.n904 0.0932835
R24460 DVSS.n921 DVSS.n904 0.0932835
R24461 DVSS.n1080 DVSS.n921 0.0932835
R24462 DVSS.n1080 DVSS.n1079 0.0932835
R24463 DVSS.n1079 DVSS.n922 0.0932835
R24464 DVSS.n1071 DVSS.n922 0.0932835
R24465 DVSS.n1071 DVSS.n1070 0.0932835
R24466 DVSS.n989 DVSS.n883 0.0932835
R24467 DVSS.n989 DVSS.n988 0.0932835
R24468 DVSS.n988 DVSS.n949 0.0932835
R24469 DVSS.n964 DVSS.n949 0.0932835
R24470 DVSS.n979 DVSS.n964 0.0932835
R24471 DVSS.n979 DVSS.n978 0.0932835
R24472 DVSS.n978 DVSS.n965 0.0932835
R24473 DVSS.n1612 DVSS.n1426 0.0932835
R24474 DVSS.n1443 DVSS.n1426 0.0932835
R24475 DVSS.n1602 DVSS.n1443 0.0932835
R24476 DVSS.n1602 DVSS.n1601 0.0932835
R24477 DVSS.n1601 DVSS.n1444 0.0932835
R24478 DVSS.n1593 DVSS.n1444 0.0932835
R24479 DVSS.n1593 DVSS.n1592 0.0932835
R24480 DVSS.n1511 DVSS.n1405 0.0932835
R24481 DVSS.n1511 DVSS.n1510 0.0932835
R24482 DVSS.n1510 DVSS.n1471 0.0932835
R24483 DVSS.n1486 DVSS.n1471 0.0932835
R24484 DVSS.n1501 DVSS.n1486 0.0932835
R24485 DVSS.n1501 DVSS.n1500 0.0932835
R24486 DVSS.n1500 DVSS.n1487 0.0932835
R24487 DVSS.n411 DVSS.n410 0.0870759
R24488 DVSS.n2284 DVSS.n2283 0.0870759
R24489 DVSS.n1092 DVSS.n1091 0.0870759
R24490 DVSS.n1614 DVSS.n1613 0.0870759
R24491 DVSS DVSS.n2674 0.0854216
R24492 DVSS.n2443 DVSS 0.0843846
R24493 DVSS.n1830 DVSS 0.0802544
R24494 DVSS.n209 DVSS.n208 0.0793691
R24495 DVSS.n188 DVSS.n187 0.0793691
R24496 DVSS.n2082 DVSS.n2081 0.0793691
R24497 DVSS.n2061 DVSS.n2060 0.0793691
R24498 DVSS.n890 DVSS.n889 0.0793691
R24499 DVSS.n869 DVSS.n868 0.0793691
R24500 DVSS.n1412 DVSS.n1411 0.0793691
R24501 DVSS.n1391 DVSS.n1390 0.0793691
R24502 DVSS.n2540 DVSS 0.0791394
R24503 DVSS.n245 DVSS.n242 0.0753538
R24504 DVSS.n2118 DVSS.n2115 0.0753538
R24505 DVSS.n926 DVSS.n923 0.0753538
R24506 DVSS.n1448 DVSS.n1445 0.0753538
R24507 DVSS.n3058 DVSS.n18 0.0736707
R24508 DVSS.n3086 DVSS.n5 0.0719286
R24509 DVSS.n438 DVSS.n437 0.0637979
R24510 DVSS.n445 DVSS.n438 0.0637979
R24511 DVSS.n493 DVSS.n492 0.0637979
R24512 DVSS.n492 DVSS.n491 0.0637979
R24513 DVSS.n2311 DVSS.n2310 0.0637979
R24514 DVSS.n2318 DVSS.n2311 0.0637979
R24515 DVSS.n2366 DVSS.n2365 0.0637979
R24516 DVSS.n2365 DVSS.n2364 0.0637979
R24517 DVSS.n1119 DVSS.n1118 0.0637979
R24518 DVSS.n1126 DVSS.n1119 0.0637979
R24519 DVSS.n1174 DVSS.n1173 0.0637979
R24520 DVSS.n1173 DVSS.n1172 0.0637979
R24521 DVSS.n1641 DVSS.n1640 0.0637979
R24522 DVSS.n1648 DVSS.n1641 0.0637979
R24523 DVSS.n1696 DVSS.n1695 0.0637979
R24524 DVSS.n1695 DVSS.n1694 0.0637979
R24525 DVSS.n18 DVSS.n15 0.0637622
R24526 DVSS.n3087 DVSS.n3086 0.062256
R24527 DVSS.n2670 DVSS.n27 0.0617245
R24528 DVSS.n3048 DVSS.n27 0.0617245
R24529 DVSS.n3044 DVSS.n32 0.0617245
R24530 DVSS.n570 DVSS.n559 0.0617245
R24531 DVSS.n574 DVSS.n553 0.0617245
R24532 DVSS.n583 DVSS.n553 0.0617245
R24533 DVSS.n593 DVSS.n592 0.0617245
R24534 DVSS.n592 DVSS.n591 0.0617245
R24535 DVSS.n590 DVSS.n546 0.0617245
R24536 DVSS.n2649 DVSS.n2623 0.0611061
R24537 DVSS.n2649 DVSS.n2648 0.0611061
R24538 DVSS.n2648 DVSS.n2647 0.0611061
R24539 DVSS.n2647 DVSS.n2624 0.0611061
R24540 DVSS.n2639 DVSS.n2624 0.0611061
R24541 DVSS.n2639 DVSS.n2638 0.0611061
R24542 DVSS.n2638 DVSS.n2637 0.0611061
R24543 DVSS.n3034 DVSS.n3033 0.0611061
R24544 DVSS.n3028 DVSS.n50 0.0611061
R24545 DVSS.n58 DVSS.n50 0.0611061
R24546 DVSS.n3018 DVSS.n3017 0.0611061
R24547 DVSS.n1894 DVSS.n1874 0.0611061
R24548 DVSS.n1895 DVSS.n1894 0.0611061
R24549 DVSS.n1896 DVSS.n1895 0.0611061
R24550 DVSS.n1896 DVSS.n1868 0.0611061
R24551 DVSS.n1904 DVSS.n1868 0.0611061
R24552 DVSS.n1905 DVSS.n1904 0.0611061
R24553 DVSS.n1912 DVSS.n1905 0.0611061
R24554 DVSS.n1908 DVSS.n1801 0.0611061
R24555 DVSS.n1921 DVSS.n1920 0.0611061
R24556 DVSS.n1921 DVSS.n1796 0.0611061
R24557 DVSS.n1936 DVSS.n1935 0.0611061
R24558 DVSS.n2758 DVSS.n2757 0.0611061
R24559 DVSS.n2757 DVSS.n722 0.0611061
R24560 DVSS.n2749 DVSS.n722 0.0611061
R24561 DVSS.n2749 DVSS.n2748 0.0611061
R24562 DVSS.n2748 DVSS.n2747 0.0611061
R24563 DVSS.n2747 DVSS.n730 0.0611061
R24564 DVSS.n2739 DVSS.n730 0.0611061
R24565 DVSS.n2735 DVSS.n738 0.0611061
R24566 DVSS.n2723 DVSS.n2722 0.0611061
R24567 DVSS.n2722 DVSS.n745 0.0611061
R24568 DVSS.n2713 DVSS.n2712 0.0611061
R24569 DVSS.n2810 DVSS.n673 0.0611061
R24570 DVSS.n2810 DVSS.n2809 0.0611061
R24571 DVSS.n2809 DVSS.n2808 0.0611061
R24572 DVSS.n2808 DVSS.n675 0.0611061
R24573 DVSS.n2800 DVSS.n675 0.0611061
R24574 DVSS.n2800 DVSS.n2799 0.0611061
R24575 DVSS.n2799 DVSS.n2798 0.0611061
R24576 DVSS.n2789 DVSS.n2788 0.0611061
R24577 DVSS.n2783 DVSS.n695 0.0611061
R24578 DVSS.n703 DVSS.n695 0.0611061
R24579 DVSS.n2774 DVSS.n2773 0.0611061
R24580 DVSS.n571 DVSS.n570 0.0610867
R24581 DVSS.n546 DVSS.n544 0.060449
R24582 DVSS.n3017 DVSS.n3016 0.0592121
R24583 DVSS.n1940 DVSS.n1936 0.0592121
R24584 DVSS.n2712 DVSS.n2711 0.0592121
R24585 DVSS.n2773 DVSS.n2772 0.0592121
R24586 DVSS.n3033 DVSS.n3032 0.0585808
R24587 DVSS.n1930 DVSS.n1801 0.0585808
R24588 DVSS.n744 DVSS.n738 0.0585808
R24589 DVSS.n2788 DVSS.n2787 0.0585808
R24590 DVSS.n2444 DVSS.n2443 0.0581923
R24591 DVSS.n2445 DVSS.n2444 0.0581923
R24592 DVSS.n2445 DVSS.n1774 0.0581923
R24593 DVSS.n2463 DVSS.n2452 0.0581923
R24594 DVSS.n2459 DVSS.n2453 0.0581923
R24595 DVSS.n2486 DVSS.n1764 0.0581923
R24596 DVSS.n2487 DVSS.n2486 0.0581923
R24597 DVSS.n2503 DVSS.n1759 0.0581923
R24598 DVSS.n2504 DVSS.n2503 0.0581923
R24599 DVSS.n2512 DVSS.n2511 0.0581923
R24600 DVSS.n2453 DVSS.n1769 0.0575913
R24601 DVSS.n2511 DVSS.n2510 0.0569904
R24602 DVSS.n1833 DVSS.n1832 0.056838
R24603 DVSS.n1833 DVSS.n1818 0.056838
R24604 DVSS.n1845 DVSS.n1841 0.056838
R24605 DVSS.n1859 DVSS.n1812 0.056838
R24606 DVSS.n2850 DVSS.n2849 0.056838
R24607 DVSS.n2849 DVSS.n2848 0.056838
R24608 DVSS.n2840 DVSS.n2839 0.056838
R24609 DVSS.n2839 DVSS.n2838 0.056838
R24610 DVSS.n2623 DVSS.n2616 0.0566869
R24611 DVSS.n1885 DVSS.n1874 0.0566869
R24612 DVSS.n2759 DVSS.n2758 0.0566869
R24613 DVSS.n673 DVSS.n672 0.0566869
R24614 DVSS.n1859 DVSS.n1858 0.0562512
R24615 DVSS.n2542 DVSS.n1258 0.0557995
R24616 DVSS.n2550 DVSS.n1258 0.0557995
R24617 DVSS.n2561 DVSS.n2554 0.0557995
R24618 DVSS.n2572 DVSS.n1246 0.0557995
R24619 DVSS.n2576 DVSS.n1238 0.0557995
R24620 DVSS.n2585 DVSS.n1238 0.0557995
R24621 DVSS.n2592 DVSS.n1232 0.0557995
R24622 DVSS.n2601 DVSS.n1232 0.0557995
R24623 DVSS.n2603 DVSS.n2602 0.0557995
R24624 DVSS.n2573 DVSS.n2572 0.0552235
R24625 DVSS.n415 DVSS.n181 0.0547553
R24626 DVSS.n2288 DVSS.n2054 0.0547553
R24627 DVSS.n1096 DVSS.n862 0.0547553
R24628 DVSS.n1618 DVSS.n1384 0.0547553
R24629 DVSS.n2829 DVSS.n2828 0.0546475
R24630 DVSS.n2604 DVSS.n2603 0.0546475
R24631 DVSS.n420 DVSS.n154 0.0505
R24632 DVSS.n2293 DVSS.n2027 0.0505
R24633 DVSS.n1101 DVSS.n835 0.0505
R24634 DVSS.n1623 DVSS.n1357 0.0505
R24635 DVSS.n591 DVSS 0.0476939
R24636 DVSS.n3045 DVSS.n3044 0.0470561
R24637 DVSS.n2671 DVSS.n2670 0.0464184
R24638 DVSS.n589 DVSS.n552 0.0464184
R24639 DVSS.n2916 DVSS.n2910 0.0459545
R24640 DVSS.n2924 DVSS.n2910 0.0459545
R24641 DVSS.n2925 DVSS.n2924 0.0459545
R24642 DVSS.n2929 DVSS.n2925 0.0459545
R24643 DVSS.n2938 DVSS.n2937 0.0459545
R24644 DVSS.n2942 DVSS.n2938 0.0459545
R24645 DVSS.n2950 DVSS.n2902 0.0459545
R24646 DVSS.n2951 DVSS.n2950 0.0459545
R24647 DVSS.n2963 DVSS.n2898 0.0459545
R24648 DVSS.n560 DVSS.n32 0.0457806
R24649 DVSS.n573 DVSS.n558 0.0457806
R24650 DVSS.n3003 DVSS.n2886 0.0456128
R24651 DVSS.n2996 DVSS.n2886 0.0456128
R24652 DVSS.n2996 DVSS.n2995 0.0456128
R24653 DVSS.n2995 DVSS.n2994 0.0456128
R24654 DVSS.n2994 DVSS.n2889 0.0456128
R24655 DVSS.n2890 DVSS.n2889 0.0456128
R24656 DVSS.n2891 DVSS.n2890 0.0456128
R24657 DVSS.n2982 DVSS.n2891 0.0456128
R24658 DVSS.n2978 DVSS.n2977 0.0456128
R24659 DVSS.n2977 DVSS.n2893 0.0456128
R24660 DVSS.n2967 DVSS.n2966 0.0456128
R24661 DVSS.n2829 DVSS.n657 0.0454309
R24662 DVSS DVSS.n2504 0.0449712
R24663 DVSS.n2452 DVSS.n1773 0.0443702
R24664 DVSS.n3059 DVSS.n3058 0.0439451
R24665 DVSS.n2838 DVSS 0.0439272
R24666 DVSS.n2493 DVSS.n2492 0.0437692
R24667 DVSS.n2637 DVSS.n2633 0.0434293
R24668 DVSS.n3029 DVSS.n48 0.0434293
R24669 DVSS.n1912 DVSS.n1911 0.0434293
R24670 DVSS.n1929 DVSS.n1799 0.0434293
R24671 DVSS.n2739 DVSS.n2738 0.0434293
R24672 DVSS.n2727 DVSS.n2726 0.0434293
R24673 DVSS.n2798 DVSS.n683 0.0434293
R24674 DVSS.n2784 DVSS.n691 0.0434293
R24675 DVSS.n1841 DVSS.n1817 0.0433404
R24676 DVSS.n2463 DVSS.n2462 0.0431683
R24677 DVSS.n2477 DVSS.n2476 0.0431683
R24678 DVSS DVSS.n2601 0.0431267
R24679 DVSS.n12 DVSS.n5 0.0429107
R24680 DVSS.n1832 DVSS.n1831 0.0427535
R24681 DVSS.n650 DVSS.n646 0.0427535
R24682 DVSS.n585 DVSS.n584 0.0425918
R24683 DVSS.n2554 DVSS.n2553 0.0425507
R24684 DVSS.n3063 DVSS 0.0424207
R24685 DVSS.n1845 DVSS.n1844 0.0421667
R24686 DVSS.n1813 DVSS.n638 0.0421667
R24687 DVSS.n2542 DVSS.n2541 0.0419747
R24688 DVSS.n2591 DVSS.n1237 0.0419747
R24689 DVSS.n2929 DVSS.n2928 0.0416932
R24690 DVSS.n2658 DVSS.n2657 0.0415354
R24691 DVSS.n1886 DVSS.n1882 0.0415354
R24692 DVSS.n2760 DVSS.n719 0.0415354
R24693 DVSS.n669 DVSS.n668 0.0415354
R24694 DVSS.n3077 DVSS 0.0414226
R24695 DVSS.n2561 DVSS.n2560 0.0413986
R24696 DVSS.n2575 DVSS.n1244 0.0413986
R24697 DVSS.n539 DVSS.n77 0.0401852
R24698 DVSS.n2412 DVSS.n1950 0.0401852
R24699 DVSS.n1220 DVSS.n758 0.0401852
R24700 DVSS.n1742 DVSS.n1280 0.0401852
R24701 DVSS.n2494 DVSS.n2488 0.0401635
R24702 DVSS.n645 DVSS.n639 0.0392324
R24703 DVSS.n2587 DVSS.n2586 0.0385184
R24704 DVSS.n61 DVSS.n58 0.036243
R24705 DVSS.n1934 DVSS.n1796 0.036243
R24706 DVSS.n753 DVSS.n745 0.036243
R24707 DVSS.n706 DVSS.n703 0.036243
R24708 DVSS.n3034 DVSS.n47 0.0333283
R24709 DVSS.n1909 DVSS.n1908 0.0333283
R24710 DVSS.n2736 DVSS.n2735 0.0333283
R24711 DVSS.n2789 DVSS.n690 0.0333283
R24712 DVSS.n3047 DVSS.n29 0.03175
R24713 DVSS.n563 DVSS.n559 0.03175
R24714 DVSS.n3048 DVSS.n3047 0.0304745
R24715 DVSS.n564 DVSS.n563 0.0304745
R24716 DVSS.n2927 DVSS.n2906 0.0303295
R24717 DVSS.n3064 DVSS.n3059 0.0302256
R24718 DVSS.n3061 DVSS 0.0302256
R24719 DVSS.n2472 DVSS.n2471 0.0299471
R24720 DVSS.n2460 DVSS.n2459 0.0299471
R24721 DVSS.n2952 DVSS.n2951 0.0298561
R24722 DVSS.n2895 DVSS.n2893 0.0296353
R24723 DVSS.n3078 DVSS.n12 0.0295179
R24724 DVSS.n3075 DVSS 0.0295179
R24725 DVSS.n1854 DVSS.n1853 0.0292559
R24726 DVSS.n1842 DVSS.n1812 0.0292559
R24727 DVSS.n2472 DVSS.n1774 0.0287452
R24728 DVSS.n2461 DVSS.n2460 0.0287452
R24729 DVSS.n2551 DVSS.n1256 0.0287258
R24730 DVSS.n2558 DVSS.n1246 0.0287258
R24731 DVSS.n181 DVSS 0.0286915
R24732 DVSS.n2054 DVSS 0.0286915
R24733 DVSS.n862 DVSS 0.0286915
R24734 DVSS.n1384 DVSS 0.0286915
R24735 DVSS.n2982 DVSS.n2981 0.0286642
R24736 DVSS.n2630 DVSS.n47 0.0282778
R24737 DVSS.n1910 DVSS.n1909 0.0282778
R24738 DVSS.n2736 DVSS.n735 0.0282778
R24739 DVSS.n690 DVSS.n689 0.0282778
R24740 DVSS.n1854 DVSS.n1818 0.0280822
R24741 DVSS.n1843 DVSS.n1842 0.0280822
R24742 DVSS.n2955 DVSS.n2898 0.0279621
R24743 DVSS.n2968 DVSS.n2967 0.0277556
R24744 DVSS.n2551 DVSS.n2550 0.0275737
R24745 DVSS.n2558 DVSS.n2556 0.0275737
R24746 DVSS.n2419 DVSS.n2416 0.0275051
R24747 DVSS.n610 DVSS.n543 0.0271646
R24748 DVSS.n2699 DVSS.n2698 0.0271646
R24749 DVSS.n1746 DVSS.n1274 0.0271646
R24750 DVSS.n3018 DVSS.n61 0.026142
R24751 DVSS.n1935 DVSS.n1934 0.026142
R24752 DVSS.n2713 DVSS.n753 0.026142
R24753 DVSS.n2774 DVSS.n706 0.026142
R24754 DVSS.n3064 DVSS.n3063 0.0256524
R24755 DVSS.n2942 DVSS.n2941 0.0250855
R24756 DVSS.n3078 DVSS.n3077 0.0250536
R24757 DVSS.n541 DVSS.n73 0.0249644
R24758 DVSS.n2414 DVSS.n1789 0.0249644
R24759 DVSS.n2702 DVSS.n757 0.0249644
R24760 DVSS.n1744 DVSS.n1277 0.0249644
R24761 DVSS.n2685 DVSS.n2684 0.0245
R24762 DVSS.n2431 DVSS.n1786 0.0245
R24763 DVSS.n2418 DVSS.n2417 0.0237334
R24764 DVSS.n74 DVSS 0.0237145
R24765 DVSS.n1790 DVSS 0.0237145
R24766 DVSS.n2704 DVSS 0.0237145
R24767 DVSS.n1278 DVSS 0.0237145
R24768 DVSS.n2864 DVSS.n2863 0.0237108
R24769 DVSS.n611 DVSS 0.0236262
R24770 DVSS.n2527 DVSS.n1266 0.0235326
R24771 DVSS DVSS.n2963 0.0232273
R24772 DVSS.n2966 DVSS 0.0230564
R24773 DVSS.n211 DVSS.n209 0.0228214
R24774 DVSS.n190 DVSS.n188 0.0228214
R24775 DVSS.n2084 DVSS.n2082 0.0228214
R24776 DVSS.n2063 DVSS.n2061 0.0228214
R24777 DVSS.n892 DVSS.n890 0.0228214
R24778 DVSS.n871 DVSS.n869 0.0228214
R24779 DVSS.n1414 DVSS.n1412 0.0228214
R24780 DVSS.n1393 DVSS.n1391 0.0228214
R24781 DVSS DVSS.n2522 0.0223216
R24782 DVSS.n2941 DVSS.n2902 0.0222446
R24783 DVSS DVSS.n2420 0.0214378
R24784 DVSS DVSS.n1223 0.0214378
R24785 DVSS.n2686 DVSS.n2685 0.02125
R24786 DVSS.n2421 DVSS.n1786 0.02125
R24787 DVSS.n609 DVSS.n608 0.0204913
R24788 DVSS.n542 DVSS.n71 0.0198972
R24789 DVSS.n2415 DVSS.n1788 0.0198972
R24790 DVSS.n2703 DVSS.n2700 0.0198972
R24791 DVSS.n1745 DVSS.n1275 0.0198972
R24792 DVSS.n222 DVSS.n203 0.0198452
R24793 DVSS.n201 DVSS.n182 0.0198452
R24794 DVSS.n2095 DVSS.n2076 0.0198452
R24795 DVSS.n2074 DVSS.n2055 0.0198452
R24796 DVSS.n903 DVSS.n884 0.0198452
R24797 DVSS.n882 DVSS.n863 0.0198452
R24798 DVSS.n1425 DVSS.n1406 0.0198452
R24799 DVSS.n1404 DVSS.n1385 0.0198452
R24800 DVSS.n585 DVSS.n583 0.0196327
R24801 DVSS.n2506 DVSS.n2505 0.0194094
R24802 DVSS.n2697 DVSS.n2696 0.0186762
R24803 DVSS.n421 DVSS.n420 0.0185851
R24804 DVSS.n425 DVSS.n421 0.0185851
R24805 DVSS.n425 DVSS.n424 0.0185851
R24806 DVSS.n424 DVSS.n423 0.0185851
R24807 DVSS.n423 DVSS.n118 0.0185851
R24808 DVSS.n437 DVSS.n118 0.0185851
R24809 DVSS.n445 DVSS.n444 0.0185851
R24810 DVSS.n440 DVSS.n439 0.0185851
R24811 DVSS.n439 DVSS.n104 0.0185851
R24812 DVSS.n459 DVSS.n104 0.0185851
R24813 DVSS.n460 DVSS.n459 0.0185851
R24814 DVSS.n465 DVSS.n102 0.0185851
R24815 DVSS.n466 DVSS.n465 0.0185851
R24816 DVSS.n493 DVSS.n466 0.0185851
R24817 DVSS.n491 DVSS.n467 0.0185851
R24818 DVSS.n467 DVSS.n86 0.0185851
R24819 DVSS.n86 DVSS.n84 0.0185851
R24820 DVSS.n531 DVSS.n84 0.0185851
R24821 DVSS.n532 DVSS.n531 0.0185851
R24822 DVSS.n533 DVSS.n532 0.0185851
R24823 DVSS.n2294 DVSS.n2293 0.0185851
R24824 DVSS.n2298 DVSS.n2294 0.0185851
R24825 DVSS.n2298 DVSS.n2297 0.0185851
R24826 DVSS.n2297 DVSS.n2296 0.0185851
R24827 DVSS.n2296 DVSS.n1991 0.0185851
R24828 DVSS.n2310 DVSS.n1991 0.0185851
R24829 DVSS.n2318 DVSS.n2317 0.0185851
R24830 DVSS.n2313 DVSS.n2312 0.0185851
R24831 DVSS.n2312 DVSS.n1977 0.0185851
R24832 DVSS.n2332 DVSS.n1977 0.0185851
R24833 DVSS.n2333 DVSS.n2332 0.0185851
R24834 DVSS.n2338 DVSS.n1975 0.0185851
R24835 DVSS.n2339 DVSS.n2338 0.0185851
R24836 DVSS.n2366 DVSS.n2339 0.0185851
R24837 DVSS.n2364 DVSS.n2340 0.0185851
R24838 DVSS.n2340 DVSS.n1959 0.0185851
R24839 DVSS.n1959 DVSS.n1957 0.0185851
R24840 DVSS.n2404 DVSS.n1957 0.0185851
R24841 DVSS.n2405 DVSS.n2404 0.0185851
R24842 DVSS.n2406 DVSS.n2405 0.0185851
R24843 DVSS.n1102 DVSS.n1101 0.0185851
R24844 DVSS.n1106 DVSS.n1102 0.0185851
R24845 DVSS.n1106 DVSS.n1105 0.0185851
R24846 DVSS.n1105 DVSS.n1104 0.0185851
R24847 DVSS.n1104 DVSS.n799 0.0185851
R24848 DVSS.n1118 DVSS.n799 0.0185851
R24849 DVSS.n1126 DVSS.n1125 0.0185851
R24850 DVSS.n1121 DVSS.n1120 0.0185851
R24851 DVSS.n1120 DVSS.n785 0.0185851
R24852 DVSS.n1140 DVSS.n785 0.0185851
R24853 DVSS.n1141 DVSS.n1140 0.0185851
R24854 DVSS.n1146 DVSS.n783 0.0185851
R24855 DVSS.n1147 DVSS.n1146 0.0185851
R24856 DVSS.n1174 DVSS.n1147 0.0185851
R24857 DVSS.n1172 DVSS.n1148 0.0185851
R24858 DVSS.n1148 DVSS.n767 0.0185851
R24859 DVSS.n767 DVSS.n765 0.0185851
R24860 DVSS.n1212 DVSS.n765 0.0185851
R24861 DVSS.n1213 DVSS.n1212 0.0185851
R24862 DVSS.n1214 DVSS.n1213 0.0185851
R24863 DVSS.n1624 DVSS.n1623 0.0185851
R24864 DVSS.n1628 DVSS.n1624 0.0185851
R24865 DVSS.n1628 DVSS.n1627 0.0185851
R24866 DVSS.n1627 DVSS.n1626 0.0185851
R24867 DVSS.n1626 DVSS.n1321 0.0185851
R24868 DVSS.n1640 DVSS.n1321 0.0185851
R24869 DVSS.n1648 DVSS.n1647 0.0185851
R24870 DVSS.n1643 DVSS.n1642 0.0185851
R24871 DVSS.n1642 DVSS.n1307 0.0185851
R24872 DVSS.n1662 DVSS.n1307 0.0185851
R24873 DVSS.n1663 DVSS.n1662 0.0185851
R24874 DVSS.n1668 DVSS.n1305 0.0185851
R24875 DVSS.n1669 DVSS.n1668 0.0185851
R24876 DVSS.n1696 DVSS.n1669 0.0185851
R24877 DVSS.n1694 DVSS.n1670 0.0185851
R24878 DVSS.n1670 DVSS.n1289 0.0185851
R24879 DVSS.n1289 DVSS.n1287 0.0185851
R24880 DVSS.n1734 DVSS.n1287 0.0185851
R24881 DVSS.n1735 DVSS.n1734 0.0185851
R24882 DVSS.n1736 DVSS.n1735 0.0185851
R24883 DVSS.n2488 DVSS.n2487 0.0185288
R24884 DVSS.n2956 DVSS.n2955 0.0184924
R24885 DVSS.n2969 DVSS.n2968 0.0183571
R24886 DVSS.n2981 DVSS.n2978 0.0183259
R24887 DVSS.n2633 DVSS.n2630 0.0181768
R24888 DVSS.n3029 DVSS.n3028 0.0181768
R24889 DVSS.n1911 DVSS.n1910 0.0181768
R24890 DVSS.n1920 DVSS.n1799 0.0181768
R24891 DVSS.n2738 DVSS.n735 0.0181768
R24892 DVSS.n2726 DVSS.n2723 0.0181768
R24893 DVSS.n689 DVSS.n683 0.0181768
R24894 DVSS.n2784 DVSS.n2783 0.0181768
R24895 DVSS.n2848 DVSS.n639 0.0181056
R24896 DVSS.n609 DVSS.n70 0.0180768
R24897 DVSS.n540 DVSS.n71 0.0179419
R24898 DVSS.n2413 DVSS.n1788 0.0179419
R24899 DVSS.n2703 DVSS.n1221 0.0179419
R24900 DVSS.n1743 DVSS.n1275 0.0179419
R24901 DVSS.n2587 DVSS.n2585 0.0177811
R24902 DVSS.n541 DVSS.n76 0.0175455
R24903 DVSS.n2414 DVSS.n1949 0.0175455
R24904 DVSS.n2705 DVSS.n757 0.0175455
R24905 DVSS.n1744 DVSS.n1279 0.0175455
R24906 DVSS.n2505 DVSS.n1747 0.0171144
R24907 DVSS.n461 DVSS.n102 0.0169894
R24908 DVSS.n2334 DVSS.n1975 0.0169894
R24909 DVSS.n1142 DVSS.n783 0.0169894
R24910 DVSS.n1664 DVSS.n1305 0.0169894
R24911 DVSS.n2956 DVSS.n2952 0.0165985
R24912 DVSS.n2969 DVSS.n2895 0.0164774
R24913 DVSS.n2697 DVSS.n1222 0.0164622
R24914 DVSS.n564 DVSS.n560 0.0164439
R24915 DVSS.n574 DVSS.n573 0.0164439
R24916 DVSS.n612 DVSS.n70 0.0164439
R24917 DVSS.n2937 DVSS.n2906 0.016125
R24918 DVSS.n2462 DVSS.n2461 0.015524
R24919 DVSS.n2476 DVSS.n1764 0.015524
R24920 DVSS.n2521 DVSS.n1747 0.015524
R24921 DVSS.n2674 DVSS.n2671 0.0152059
R24922 DVSS.n1844 DVSS.n1843 0.0151714
R24923 DVSS.n2850 DVSS.n638 0.0151714
R24924 DVSS.n3045 DVSS.n29 0.0151684
R24925 DVSS.n2417 DVSS.n659 0.0149009
R24926 DVSS.n2560 DVSS.n2556 0.0149009
R24927 DVSS.n2576 DVSS.n2575 0.0149009
R24928 DVSS.n1226 DVSS.n1222 0.0149009
R24929 DVSS.n443 DVSS.n440 0.0148617
R24930 DVSS.n2316 DVSS.n2313 0.0148617
R24931 DVSS.n1124 DVSS.n1121 0.0148617
R24932 DVSS.n1646 DVSS.n1643 0.0148617
R24933 DVSS.n2684 DVSS.n2665 0.01475
R24934 DVSS.n2433 DVSS.n2431 0.01475
R24935 DVSS DVSS.n590 0.0145306
R24936 DVSS.n2471 DVSS.n1773 0.0143221
R24937 DVSS.n2863 DVSS.n2862 0.0142814
R24938 DVSS.n2668 DVSS 0.01425
R24939 DVSS.n1785 DVSS 0.01425
R24940 DVSS.n2537 DVSS.n1266 0.0141756
R24941 DVSS.n1831 DVSS.n1830 0.0140747
R24942 DVSS.n1853 DVSS.n1817 0.0139977
R24943 DVSS.n2541 DVSS.n2540 0.0138333
R24944 DVSS.n3 DVSS.n2 0.0137979
R24945 DVSS DVSS.n1825 0.0137979
R24946 DVSS.n2553 DVSS.n1256 0.0137488
R24947 DVSS.n2512 DVSS 0.0137212
R24948 DVSS.n2526 DVSS.n2525 0.0136958
R24949 DVSS.n1265 DVSS 0.0136958
R24950 DVSS.n656 DVSS 0.0134108
R24951 DVSS.n2602 DVSS 0.0131728
R24952 DVSS.n593 DVSS.n589 0.0119796
R24953 DVSS.n73 DVSS.n72 0.0117068
R24954 DVSS.n1938 DVSS.n1789 0.0117068
R24955 DVSS.n2702 DVSS.n2701 0.0117068
R24956 DVSS.n1277 DVSS.n1276 0.0117068
R24957 DVSS.n2492 DVSS.n1759 0.0113173
R24958 DVSS.n2840 DVSS.n650 0.0110634
R24959 DVSS.n657 DVSS.n656 0.0110634
R24960 DVSS.n2592 DVSS.n2591 0.0108687
R24961 DVSS.n2418 DVSS.n658 0.0104846
R24962 DVSS.n3073 DVSS.n15 0.0104085
R24963 DVSS.n2667 DVSS.n2665 0.01025
R24964 DVSS.n2675 DVSS 0.01025
R24965 DVSS.n2433 DVSS.n2432 0.01025
R24966 DVSS.n2435 DVSS 0.01025
R24967 DVSS.n3088 DVSS.n3087 0.0101726
R24968 DVSS.n608 DVSS.n607 0.0100663
R24969 DVSS.n2862 DVSS.n2861 0.0099294
R24970 DVSS DVSS.n1827 0.0099294
R24971 DVSS.n2537 DVSS.n2536 0.00985701
R24972 DVSS DVSS.n2539 0.00985701
R24973 DVSS.n2507 DVSS.n2506 0.00951442
R24974 DVSS.n72 DVSS.n62 0.00933838
R24975 DVSS.n1939 DVSS.n1938 0.00933838
R24976 DVSS.n2701 DVSS.n754 0.00933838
R24977 DVSS.n1276 DVSS.n707 0.00933838
R24978 DVSS.n2827 DVSS.n658 0.00914055
R24979 DVSS.n2696 DVSS.n1224 0.00914055
R24980 DVSS.n612 DVSS.n611 0.00895784
R24981 DVSS.n76 DVSS.n74 0.00856303
R24982 DVSS.n1949 DVSS.n1790 0.00856303
R24983 DVSS.n2705 DVSS.n2704 0.00856303
R24984 DVSS.n1279 DVSS.n1278 0.00856303
R24985 DVSS.n2522 DVSS.n2521 0.0084995
R24986 DVSS.n2420 DVSS.n659 0.00818896
R24987 DVSS.n1226 DVSS.n1223 0.00818896
R24988 DVSS DVSS.n2667 0.008
R24989 DVSS.n2432 DVSS 0.008
R24990 DVSS.n2861 DVSS 0.00775339
R24991 DVSS.n2536 DVSS 0.0076977
R24992 DVSS.n3062 DVSS.n3061 0.00735976
R24993 DVSS.n2864 DVSS.n3 0.00726983
R24994 DVSS.n2527 DVSS.n2526 0.00721785
R24995 DVSS.n3076 DVSS.n3075 0.00719643
R24996 DVSS.n416 DVSS.n154 0.00688298
R24997 DVSS.n2289 DVSS.n2027 0.00688298
R24998 DVSS.n1097 DVSS.n835 0.00688298
R24999 DVSS.n1619 DVSS.n1357 0.00688298
R25000 DVSS DVSS.n3062 0.00659756
R25001 DVSS.n208 DVSS.n203 0.00645238
R25002 DVSS.n187 DVSS.n182 0.00645238
R25003 DVSS.n2081 DVSS.n2076 0.00645238
R25004 DVSS.n2060 DVSS.n2055 0.00645238
R25005 DVSS.n889 DVSS.n884 0.00645238
R25006 DVSS.n868 DVSS.n863 0.00645238
R25007 DVSS.n1411 DVSS.n1406 0.00645238
R25008 DVSS.n1390 DVSS.n1385 0.00645238
R25009 DVSS DVSS.n3076 0.00645238
R25010 DVSS.n411 DVSS.n202 0.00565464
R25011 DVSS.n2284 DVSS.n2075 0.00565464
R25012 DVSS.n1092 DVSS.n883 0.00565464
R25013 DVSS.n1614 DVSS.n1405 0.00565464
R25014 DVSS.n2657 DVSS.n2616 0.00491919
R25015 DVSS.n1886 DVSS.n1885 0.00491919
R25016 DVSS.n2760 DVSS.n2759 0.00491919
R25017 DVSS.n672 DVSS.n668 0.00491919
R25018 DVSS.n2928 DVSS.n2927 0.00476136
R25019 DVSS.n416 DVSS.n415 0.00475532
R25020 DVSS.n2289 DVSS.n2288 0.00475532
R25021 DVSS.n1097 DVSS.n1096 0.00475532
R25022 DVSS.n1619 DVSS.n1618 0.00475532
R25023 DVSS.n584 DVSS.n552 0.00432653
R25024 DVSS.n414 DVSS.n413 0.00423171
R25025 DVSS.n2287 DVSS.n2286 0.00423171
R25026 DVSS.n1095 DVSS.n1094 0.00423171
R25027 DVSS.n1617 DVSS.n1616 0.00423171
R25028 DVSS.n444 DVSS.n443 0.0042234
R25029 DVSS.n2317 DVSS.n2316 0.0042234
R25030 DVSS.n1125 DVSS.n1124 0.0042234
R25031 DVSS.n1647 DVSS.n1646 0.0042234
R25032 DVSS.n2494 DVSS.n2493 0.00410577
R25033 DVSS.n646 DVSS.n645 0.00402113
R25034 DVSS.n2586 DVSS.n1237 0.00395622
R25035 DVSS.n2687 DVSS.n2686 0.00375
R25036 DVSS.n2422 DVSS.n2421 0.00375
R25037 DVSS.n2 DVSS.n1 0.00364313
R25038 DVSS.n2525 DVSS.n2524 0.003619
R25039 DVSS.n212 DVSS.n211 0.00347619
R25040 DVSS.n191 DVSS.n190 0.00347619
R25041 DVSS.n2085 DVSS.n2084 0.00347619
R25042 DVSS.n2064 DVSS.n2063 0.00347619
R25043 DVSS.n893 DVSS.n892 0.00347619
R25044 DVSS.n872 DVSS.n871 0.00347619
R25045 DVSS.n1415 DVSS.n1414 0.00347619
R25046 DVSS.n1394 DVSS.n1393 0.00347619
R25047 DVSS.n3032 DVSS.n48 0.00302525
R25048 DVSS.n1930 DVSS.n1929 0.00302525
R25049 DVSS.n2727 DVSS.n744 0.00302525
R25050 DVSS.n2787 DVSS.n691 0.00302525
R25051 DVSS.n2676 DVSS.n2675 0.00275
R25052 DVSS.n2436 DVSS.n2435 0.00275
R25053 DVSS.n1827 DVSS.n1826 0.00267602
R25054 DVSS.n2539 DVSS.n1264 0.00265931
R25055 DVSS.n2676 DVSS 0.0025
R25056 DVSS.n2436 DVSS 0.0025
R25057 DVSS.n1826 DVSS 0.00243424
R25058 DVSS DVSS.n1264 0.00241939
R25059 DVSS.n3016 DVSS.n62 0.00239394
R25060 DVSS.n1940 DVSS.n1939 0.00239394
R25061 DVSS.n2711 DVSS.n754 0.00239394
R25062 DVSS.n2772 DVSS.n707 0.00239394
R25063 DVSS.n461 DVSS.n460 0.00209574
R25064 DVSS.n2334 DVSS.n2333 0.00209574
R25065 DVSS.n1142 DVSS.n1141 0.00209574
R25066 DVSS.n1664 DVSS.n1663 0.00209574
R25067 DVSS.n607 DVSS.n544 0.00177551
R25068 DVSS.n2510 DVSS.n2507 0.00170192
R25069 DVSS.n2828 DVSS.n2827 0.00165207
R25070 DVSS.n2604 DVSS.n1224 0.00165207
R25071 DVSS.n533 DVSS.n77 0.00156383
R25072 DVSS.n2406 DVSS.n1950 0.00156383
R25073 DVSS.n1214 DVSS.n758 0.00156383
R25074 DVSS.n1736 DVSS.n1280 0.00156383
R25075 DVSS.n415 DVSS.n414 0.00149989
R25076 DVSS.n2288 DVSS.n2287 0.00149989
R25077 DVSS.n1096 DVSS.n1095 0.00149989
R25078 DVSS.n1618 DVSS.n1617 0.00149989
R25079 DVSS.n2417 DVSS.n2416 0.00149701
R25080 DVSS.n2668 DVSS 0.00125
R25081 DVSS DVSS.n1785 0.00125
R25082 DVSS.n1825 DVSS 0.00122534
R25083 DVSS DVSS.n1265 0.00121977
R25084 DVSS.n571 DVSS.n558 0.00113776
R25085 DVSS.n2477 DVSS.n1769 0.00110096
R25086 DVSS.n1858 DVSS.n1813 0.00108685
R25087 DVSS.n2573 DVSS.n1244 0.00107604
R25088 DVSS.n542 DVSS.n541 0.001
R25089 DVSS.n2415 DVSS.n2414 0.001
R25090 DVSS.n2700 DVSS.n757 0.001
R25091 DVSS.n1745 DVSS.n1744 0.001
R25092 DVSS.n543 DVSS.n70 0.001
R25093 DVSS.n1747 DVSS.n1746 0.001
R25094 DVSS.n2699 DVSS.n1222 0.001
R25095 DVSS.n413 DVSS.n154 0.000500988
R25096 DVSS.n418 DVSS.n154 0.000500988
R25097 DVSS.n2286 DVSS.n2027 0.000500988
R25098 DVSS.n2291 DVSS.n2027 0.000500988
R25099 DVSS.n1094 DVSS.n835 0.000500988
R25100 DVSS.n1099 DVSS.n835 0.000500988
R25101 DVSS.n1616 DVSS.n1357 0.000500988
R25102 DVSS.n1621 DVSS.n1357 0.000500988
R25103 DVSS.n443 DVSS.n442 0.000500379
R25104 DVSS.n2316 DVSS.n2315 0.000500379
R25105 DVSS.n1124 DVSS.n1123 0.000500379
R25106 DVSS.n1646 DVSS.n1645 0.000500379
R25107 DVSS.n78 DVSS.n77 0.000500334
R25108 DVSS.n1951 DVSS.n1950 0.000500334
R25109 DVSS.n759 DVSS.n758 0.000500334
R25110 DVSS.n1281 DVSS.n1280 0.000500334
R25111 DVSS.n462 DVSS.n461 0.000500219
R25112 DVSS.n2335 DVSS.n2334 0.000500219
R25113 DVSS.n1143 DVSS.n1142 0.000500219
R25114 DVSS.n1665 DVSS.n1664 0.000500219
R25115 DVSS.n2964 DVSS.n0 0.000500012
R25116 B1.n66 B1.n65 185
R25117 B1.n64 B1.n57 185
R25118 B1.n24 B1.n15 185
R25119 B1.n23 B1.n22 185
R25120 B1.n69 B1.t0 120.037
R25121 B1.t1 B1.n14 120.037
R25122 B1.n59 B1.n57 112.831
R25123 B1.n22 B1.n21 112.831
R25124 B1.n68 B1.n67 104.172
R25125 B1.n27 B1.n26 104.172
R25126 B1.n68 B1.n56 92.5005
R25127 B1.n28 B1.n27 92.5005
R25128 B1.t0 B1.n68 66.8281
R25129 B1.n27 B1.t1 66.8281
R25130 B1.n6 B1.t4 35.2053
R25131 B1.n3 B1.t5 34.0571
R25132 B1.n67 B1.n66 29.4833
R25133 B1.n26 B1.n15 29.4833
R25134 B1.n1 B1.t2 27.6955
R25135 B1.n1 B1.t3 27.6955
R25136 B1.n45 B1.n44 19.0955
R25137 B1.n69 B1.n56 15.4558
R25138 B1.n28 B1.n14 15.4558
R25139 B1.n64 B1.n63 13.5534
R25140 B1.n23 B1.n18 13.5534
R25141 B1.n2 B1.n1 9.67857
R25142 B1.n41 B1.n34 9.30581
R25143 B1.n59 B1.n58 9.30424
R25144 B1.n21 B1.n20 9.30413
R25145 B1.n40 B1.n39 9.3005
R25146 B1.n46 B1.n45 9.3005
R25147 B1.n71 B1.n70 9.3005
R25148 B1.n55 B1.n52 9.3005
R25149 B1.n67 B1.n55 9.3005
R25150 B1.n63 B1.n62 9.3005
R25151 B1.n72 B1.n54 9.3005
R25152 B1.n29 B1.n13 9.3005
R25153 B1.n25 B1.n11 9.3005
R25154 B1.n26 B1.n25 9.3005
R25155 B1.n18 B1.n17 9.3005
R25156 B1.n31 B1.n30 9.3005
R25157 B1.n71 B1.n56 9.03579
R25158 B1.n29 B1.n28 9.03579
R25159 B1.n43 B1.n41 8.49366
R25160 B1.n43 B1.t7 8.2655
R25161 B1.n43 B1.t6 8.2655
R25162 B1.n44 B1.n43 7.97749
R25163 B1.n42 B1.n40 7.26743
R25164 B1.n43 B1.n42 6.15568
R25165 B1.n65 B1.n55 5.64756
R25166 B1.n25 B1.n24 5.64756
R25167 B1.n41 B1.n35 4.89462
R25168 B1.n60 B1.n59 4.89462
R25169 B1.n21 B1.n19 4.89462
R25170 B1.n73 B1.n55 4.51815
R25171 B1.n72 B1.n71 4.51815
R25172 B1.n25 B1.n12 4.51815
R25173 B1.n30 B1.n29 4.51815
R25174 B1.n5 B1.n4 4.5005
R25175 B1.n4 B1.n2 4.5005
R25176 B1.n51 B1.n9 4.5005
R25177 B1.n49 B1.n9 4.5005
R25178 B1.n51 B1.n50 4.5005
R25179 B1.n50 B1.n49 4.5005
R25180 B1.n74 B1.n53 4.5005
R25181 B1.n75 B1.n8 4.5005
R25182 B1.n53 B1.n8 4.5005
R25183 B1.n75 B1.n74 4.5005
R25184 B1.n48 B1.n32 4.5005
R25185 B1.n47 B1.n36 4.5005
R25186 B1.n48 B1.n47 4.5005
R25187 B1.n36 B1.n32 4.5005
R25188 B1.n38 B1.n33 4.5005
R25189 B1.n66 B1.n57 3.93153
R25190 B1.n22 B1.n15 3.93153
R25191 B1.n19 B1.n9 3.03311
R25192 B1.n50 B1.n12 3.03311
R25193 B1.n60 B1.n8 3.03311
R25194 B1.n74 B1.n73 3.03311
R25195 B1.n47 B1.n35 3.03311
R25196 B1.n3 B1.n0 2.2714
R25197 B1.n58 B1.n7 2.25261
R25198 B1.n20 B1.n10 2.25256
R25199 B1.n34 B1.n33 2.25127
R25200 B1.n37 B1.n33 2.24434
R25201 B1.n73 B1.n72 1.88285
R25202 B1.n30 B1.n12 1.88285
R25203 B1.n45 B1.n35 1.50638
R25204 B1.n63 B1.n60 1.50638
R25205 B1.n19 B1.n18 1.50638
R25206 B1.n16 B1.n10 1.49213
R25207 B1.n70 B1.n69 1.49212
R25208 B1.n61 B1.n7 1.49182
R25209 B1.n14 B1.n13 1.49166
R25210 B1.n65 B1.n64 0.753441
R25211 B1.n24 B1.n23 0.753441
R25212 B1.n44 B1.n40 0.521921
R25213 B1.n77 B1.n6 0.29767
R25214 B1.n49 B1.n48 0.238951
R25215 B1.n77 B1.n76 0.196255
R25216 B1 B1.n77 0.1855
R25217 B1.n6 B1.n5 0.149538
R25218 B1.n75 B1.n51 0.124821
R25219 B1.n42 B1.n32 0.0579027
R25220 B1.n62 B1.n61 0.0396286
R25221 B1.n17 B1.n16 0.0383668
R25222 B1.n46 B1.n37 0.0314092
R25223 B1.n5 B1.n0 0.0281442
R25224 B1.n39 B1.n37 0.0271357
R25225 B1.n61 B1.n52 0.0202788
R25226 B1.n16 B1.n11 0.0196501
R25227 B1.n51 B1.n10 0.0168043
R25228 B1.n36 B1.n33 0.016125
R25229 B1.n74 B1.n52 0.013431
R25230 B1.n70 B1.n54 0.013431
R25231 B1.n50 B1.n11 0.013
R25232 B1.n31 B1.n13 0.013
R25233 B1.n38 B1.n32 0.0122521
R25234 B1.n58 B1.n8 0.0117689
R25235 B1.n20 B1.n9 0.0114102
R25236 B1.n47 B1.n34 0.0100704
R25237 B1.n76 B1.n7 0.0100109
R25238 B1.n74 B1.n54 0.00588793
R25239 B1.n50 B1.n31 0.00570833
R25240 B1.n62 B1.n8 0.00481034
R25241 B1.n47 B1.n46 0.0047735
R25242 B1.n17 B1.n9 0.00466667
R25243 B1.n53 B1.n7 0.00457609
R25244 B1.n76 B1.n75 0.00457609
R25245 B1.n2 B1.n0 0.00410577
R25246 B1.n39 B1.n38 0.00370513
R25247 B1.n48 B1.n33 0.00253804
R25248 B1.n4 B1.n3 0.00185919
R25249 B1.n49 B1.n10 0.0018587
R25250 a_2221_8623.n79 a_2221_8623.t9 60.2505
R25251 a_2221_8623.n57 a_2221_8623.t6 60.2505
R25252 a_2221_8623.n43 a_2221_8623.t8 60.2505
R25253 a_2221_8623.n21 a_2221_8623.t7 60.2505
R25254 a_2221_8623.n0 a_2221_8623.n131 9.3005
R25255 a_2221_8623.n0 a_2221_8623.n129 9.3005
R25256 a_2221_8623.n4 a_2221_8623.n65 9.3005
R25257 a_2221_8623.n4 a_2221_8623.n66 9.3005
R25258 a_2221_8623.n4 a_2221_8623.n64 9.3005
R25259 a_2221_8623.n64 a_2221_8623.n63 9.3005
R25260 a_2221_8623.n5 a_2221_8623.n72 9.3005
R25261 a_2221_8623.n6 a_2221_8623.n89 9.3005
R25262 a_2221_8623.n5 a_2221_8623.n78 9.3005
R25263 a_2221_8623.n78 a_2221_8623.n77 9.3005
R25264 a_2221_8623.n5 a_2221_8623.n71 9.3005
R25265 a_2221_8623.n6 a_2221_8623.n87 9.3005
R25266 a_2221_8623.n87 a_2221_8623.n86 9.3005
R25267 a_2221_8623.n6 a_2221_8623.n88 9.3005
R25268 a_2221_8623.n3 a_2221_8623.n29 9.3005
R25269 a_2221_8623.n3 a_2221_8623.n30 9.3005
R25270 a_2221_8623.n3 a_2221_8623.n28 9.3005
R25271 a_2221_8623.n28 a_2221_8623.n27 9.3005
R25272 a_2221_8623.n2 a_2221_8623.n36 9.3005
R25273 a_2221_8623.n2 a_2221_8623.n42 9.3005
R25274 a_2221_8623.n42 a_2221_8623.n41 9.3005
R25275 a_2221_8623.n2 a_2221_8623.n35 9.3005
R25276 a_2221_8623.n1 a_2221_8623.n51 9.3005
R25277 a_2221_8623.n51 a_2221_8623.n50 9.3005
R25278 a_2221_8623.n1 a_2221_8623.n53 9.3005
R25279 a_2221_8623.n1 a_2221_8623.n52 9.3005
R25280 a_2221_8623.n8 a_2221_8623.n19 9.3005
R25281 a_2221_8623.n7 a_2221_8623.n14 9.3005
R25282 a_2221_8623.n162 a_2221_8623.n159 9.3005
R25283 a_2221_8623.n162 a_2221_8623.n160 9.3005
R25284 a_2221_8623.n80 a_2221_8623.n79 8.76429
R25285 a_2221_8623.n44 a_2221_8623.n43 8.76429
R25286 a_2221_8623.n85 a_2221_8623.n84 7.45411
R25287 a_2221_8623.n76 a_2221_8623.n75 7.45411
R25288 a_2221_8623.n62 a_2221_8623.n61 7.45411
R25289 a_2221_8623.n40 a_2221_8623.n39 7.45411
R25290 a_2221_8623.n49 a_2221_8623.n48 7.45411
R25291 a_2221_8623.n26 a_2221_8623.n25 7.45411
R25292 a_2221_8623.n58 a_2221_8623.n57 6.80105
R25293 a_2221_8623.n22 a_2221_8623.n21 6.80105
R25294 a_2221_8623.n83 a_2221_8623.n82 5.64756
R25295 a_2221_8623.n74 a_2221_8623.n73 5.64756
R25296 a_2221_8623.n60 a_2221_8623.n59 5.64756
R25297 a_2221_8623.n38 a_2221_8623.n37 5.64756
R25298 a_2221_8623.n47 a_2221_8623.n46 5.64756
R25299 a_2221_8623.n24 a_2221_8623.n23 5.64756
R25300 a_2221_8623.n112 a_2221_8623.t2 5.5395
R25301 a_2221_8623.n112 a_2221_8623.t1 5.5395
R25302 a_2221_8623.t3 a_2221_8623.n162 5.5395
R25303 a_2221_8623.n162 a_2221_8623.t0 5.5395
R25304 a_2221_8623.n70 a_2221_8623.n69 4.73575
R25305 a_2221_8623.n68 a_2221_8623.n67 4.73575
R25306 a_2221_8623.n34 a_2221_8623.n33 4.73575
R25307 a_2221_8623.n32 a_2221_8623.n31 4.73575
R25308 a_2221_8623.n81 a_2221_8623.n80 4.6505
R25309 a_2221_8623.n45 a_2221_8623.n44 4.6505
R25310 a_2221_8623.n135 a_2221_8623.n134 4.51815
R25311 a_2221_8623.n17 a_2221_8623.n16 4.51815
R25312 a_2221_8623.n155 a_2221_8623.n154 4.51815
R25313 a_2221_8623.n0 a_2221_8623.n128 4.5005
R25314 a_2221_8623.n124 a_2221_8623.n133 4.5005
R25315 a_2221_8623.n125 a_2221_8623.n123 4.5005
R25316 a_2221_8623.n118 a_2221_8623.n116 4.5005
R25317 a_2221_8623.n8 a_2221_8623.n12 4.5005
R25318 a_2221_8623.n7 a_2221_8623.n17 4.5005
R25319 a_2221_8623.n102 a_2221_8623.n107 4.5005
R25320 a_2221_8623.n139 a_2221_8623.n147 4.5005
R25321 a_2221_8623.n152 a_2221_8623.n151 4.5005
R25322 a_2221_8623.n138 a_2221_8623.n141 4.5005
R25323 a_2221_8623.n162 a_2221_8623.n161 4.35791
R25324 a_2221_8623.n91 a_2221_8623.n93 4.24504
R25325 a_2221_8623.n54 a_2221_8623.n56 4.24504
R25326 a_2221_8623.n12 a_2221_8623.n11 3.76521
R25327 a_2221_8623.n4 a_2221_8623.n58 3.42768
R25328 a_2221_8623.n3 a_2221_8623.n22 3.42768
R25329 a_2221_8623.n123 a_2221_8623.n119 3.38874
R25330 a_2221_8623.n147 a_2221_8623.n144 3.38874
R25331 a_2221_8623.n131 a_2221_8623.n130 3.38537
R25332 a_2221_8623.n158 a_2221_8623.n157 3.38537
R25333 a_2221_8623.n97 a_2221_8623.t4 3.3065
R25334 a_2221_8623.n97 a_2221_8623.t5 3.3065
R25335 a_2221_8623.n107 a_2221_8623.n105 3.28194
R25336 a_2221_8623.n99 a_2221_8623.n98 3.15821
R25337 a_2221_8623.n117 a_2221_8623.n135 3.03311
R25338 a_2221_8623.n153 a_2221_8623.n155 3.03311
R25339 a_2221_8623.n107 a_2221_8623.n106 3.01226
R25340 a_2221_8623.n12 a_2221_8623.n10 2.63579
R25341 a_2221_8623.n14 a_2221_8623.n13 2.61733
R25342 a_2221_8623.n0 a_2221_8623.n126 2.57914
R25343 a_2221_8623.n122 a_2221_8623.n121 2.25932
R25344 a_2221_8623.n146 a_2221_8623.n145 2.25932
R25345 a_2221_8623.n19 a_2221_8623.n18 2.24766
R25346 a_2221_8623.n116 a_2221_8623.n114 2.22452
R25347 a_2221_8623.n151 a_2221_8623.n149 2.22452
R25348 a_2221_8623.n162 a_2221_8623.n148 1.99078
R25349 a_2221_8623.n17 a_2221_8623.n15 1.88285
R25350 a_2221_8623.n113 a_2221_8623.n112 1.72048
R25351 a_2221_8623.n99 a_2221_8623.n97 1.61799
R25352 a_2221_8623.n108 a_2221_8623.n96 1.51434
R25353 a_2221_8623.n96 a_2221_8623.n8 1.51334
R25354 a_2221_8623.n128 a_2221_8623.n127 1.50638
R25355 a_2221_8623.n159 a_2221_8623.n158 1.50638
R25356 a_2221_8623.n142 a_2221_8623.n143 1.50638
R25357 a_2221_8623.n101 a_2221_8623.n100 1.12991
R25358 a_2221_8623.n95 a_2221_8623.n94 3.28829
R25359 a_2221_8623.n86 a_2221_8623.n85 0.994314
R25360 a_2221_8623.n77 a_2221_8623.n76 0.994314
R25361 a_2221_8623.n63 a_2221_8623.n62 0.994314
R25362 a_2221_8623.n41 a_2221_8623.n40 0.994314
R25363 a_2221_8623.n50 a_2221_8623.n49 0.994314
R25364 a_2221_8623.n27 a_2221_8623.n26 0.994314
R25365 a_2221_8623.n111 a_2221_8623.n156 0.829361
R25366 a_2221_8623.n133 a_2221_8623.n132 0.753441
R25367 a_2221_8623.n87 a_2221_8623.n83 0.753441
R25368 a_2221_8623.n78 a_2221_8623.n74 0.753441
R25369 a_2221_8623.n64 a_2221_8623.n60 0.753441
R25370 a_2221_8623.n42 a_2221_8623.n38 0.753441
R25371 a_2221_8623.n51 a_2221_8623.n47 0.753441
R25372 a_2221_8623.n28 a_2221_8623.n24 0.753441
R25373 a_2221_8623.n141 a_2221_8623.n140 0.753441
R25374 a_2221_8623.n137 a_2221_8623.n136 0.754708
R25375 a_2221_8623.n93 a_2221_8623.n92 0.709906
R25376 a_2221_8623.n56 a_2221_8623.n55 0.709906
R25377 a_2221_8623.n109 a_2221_8623.n137 0.678625
R25378 a_2221_8623.n70 a_2221_8623.n68 0.458354
R25379 a_2221_8623.n34 a_2221_8623.n32 0.458354
R25380 a_2221_8623.n123 a_2221_8623.n122 0.376971
R25381 a_2221_8623.n121 a_2221_8623.n120 0.376971
R25382 a_2221_8623.n104 a_2221_8623.n103 0.376971
R25383 a_2221_8623.n147 a_2221_8623.n146 0.376971
R25384 a_2221_8623.n95 a_2221_8623.n20 0.242354
R25385 a_2221_8623.n136 a_2221_8623.n113 0.225683
R25386 a_2221_8623.n108 a_2221_8623.n99 0.224119
R25387 a_2221_8623.n6 a_2221_8623.n81 0.190717
R25388 a_2221_8623.n81 a_2221_8623.n5 0.190717
R25389 a_2221_8623.n45 a_2221_8623.n2 0.190717
R25390 a_2221_8623.n1 a_2221_8623.n45 0.190717
R25391 a_2221_8623.n94 a_2221_8623.n54 0.159981
R25392 a_2221_8623.n94 a_2221_8623.n91 0.159717
R25393 a_2221_8623.n138 a_2221_8623.n142 4.63429
R25394 a_2221_8623.n105 a_2221_8623.n104 0.0902327
R25395 a_2221_8623.n117 a_2221_8623.n125 0.0900802
R25396 a_2221_8623.n136 a_2221_8623.n118 0.0608541
R25397 a_2221_8623.n111 a_2221_8623.n110 0.0528649
R25398 a_2221_8623.n156 a_2221_8623.n153 0.0511262
R25399 a_2221_8623.n156 a_2221_8623.n139 0.040511
R25400 a_2221_8623.n114 a_2221_8623.n115 0.0303633
R25401 a_2221_8623.n149 a_2221_8623.n150 0.0303633
R25402 a_2221_8623.n102 a_2221_8623.n101 4.54542
R25403 a_2221_8623.n152 a_2221_8623.n148 0.0122188
R25404 a_2221_8623.n153 a_2221_8623.n152 0.0454219
R25405 a_2221_8623.n139 a_2221_8623.n138 0.0454219
R25406 a_2221_8623.n118 a_2221_8623.n117 0.0454219
R25407 a_2221_8623.n125 a_2221_8623.n124 0.0454219
R25408 a_2221_8623.n111 a_2221_8623.n109 0.022561
R25409 a_2221_8623.n111 a_2221_8623.n20 0.847626
R25410 a_2221_8623.n108 a_2221_8623.n102 0.0883906
R25411 a_2221_8623.n96 a_2221_8623.n95 0.905839
R25412 a_2221_8623.n91 a_2221_8623.n90 0.0410417
R25413 a_2221_8623.n8 a_2221_8623.n9 2.77239
R25414 a_2221_8623.n5 a_2221_8623.n70 0.205546
R25415 a_2221_8623.n68 a_2221_8623.n4 0.205546
R25416 a_2221_8623.n32 a_2221_8623.n3 0.205546
R25417 a_2221_8623.n2 a_2221_8623.n34 0.205546
R25418 a_2221_8623.n54 a_2221_8623.n1 0.177485
R25419 a_2221_8623.n124 a_2221_8623.n0 0.171838
R25420 a_2221_8623.n8 a_2221_8623.n7 0.167464
R25421 a_2221_8623.n90 a_2221_8623.n6 0.137941
R25422 a_2093_3714.n47 a_2093_3714.n46 6.31679
R25423 a_2093_3714.n1 a_2093_3714.n19 6.12763
R25424 a_2093_3714.n3 a_2093_3714.n25 6.12763
R25425 a_2093_3714.n6 a_2093_3714.n41 6.12763
R25426 a_2093_3714.n17 a_2093_3714.t6 5.5395
R25427 a_2093_3714.n17 a_2093_3714.t9 5.5395
R25428 a_2093_3714.n23 a_2093_3714.t10 5.5395
R25429 a_2093_3714.n23 a_2093_3714.t11 5.5395
R25430 a_2093_3714.n29 a_2093_3714.t8 5.5395
R25431 a_2093_3714.n29 a_2093_3714.t4 5.5395
R25432 a_2093_3714.n34 a_2093_3714.t3 5.5395
R25433 a_2093_3714.n34 a_2093_3714.t2 5.5395
R25434 a_2093_3714.n39 a_2093_3714.t5 5.5395
R25435 a_2093_3714.n39 a_2093_3714.t7 5.5395
R25436 a_2093_3714.n48 a_2093_3714.t0 5.5395
R25437 a_2093_3714.t1 a_2093_3714.n48 5.5395
R25438 a_2093_3714.n5 a_2093_3714.n38 4.5005
R25439 a_2093_3714.n4 a_2093_3714.n33 4.5005
R25440 a_2093_3714.n2 a_2093_3714.n22 4.5005
R25441 a_2093_3714.n7 a_2093_3714.n28 4.5005
R25442 a_2093_3714.n0 a_2093_3714.n16 4.5005
R25443 a_2093_3714.n8 a_2093_3714.n43 4.5005
R25444 a_2093_3714.n9 a_2093_3714.n45 4.5005
R25445 a_2093_3714.n16 a_2093_3714.n14 3.76521
R25446 a_2093_3714.n22 a_2093_3714.n20 3.76521
R25447 a_2093_3714.n28 a_2093_3714.n26 3.76521
R25448 a_2093_3714.n33 a_2093_3714.n31 3.76521
R25449 a_2093_3714.n38 a_2093_3714.n36 3.76521
R25450 a_2093_3714.n45 a_2093_3714.n44 3.76521
R25451 a_2093_3714.n43 a_2093_3714.n42 3.01226
R25452 a_2093_3714.n16 a_2093_3714.n15 2.63579
R25453 a_2093_3714.n22 a_2093_3714.n21 2.63579
R25454 a_2093_3714.n28 a_2093_3714.n27 2.63579
R25455 a_2093_3714.n33 a_2093_3714.n32 2.63579
R25456 a_2093_3714.n38 a_2093_3714.n37 2.63579
R25457 a_2093_3714.n11 a_2093_3714.n1 2.20191
R25458 a_2093_3714.n13 a_2093_3714.n6 1.48434
R25459 a_2093_3714.n10 a_2093_3714.n4 1.74534
R25460 a_2093_3714.n11 a_2093_3714.n3 1.48434
R25461 a_2093_3714.n12 a_2093_3714.n7 1.745
R25462 a_2093_3714.n7 a_2093_3714.n30 1.4669
R25463 a_2093_3714.n0 a_2093_3714.n18 1.46689
R25464 a_2093_3714.n2 a_2093_3714.n24 1.46689
R25465 a_2093_3714.n4 a_2093_3714.n35 1.46689
R25466 a_2093_3714.n5 a_2093_3714.n40 1.46689
R25467 a_2093_3714.n47 a_2093_3714.n9 1.46687
R25468 a_2093_3714.n12 a_2093_3714.n11 0.700686
R25469 a_2093_3714.n8 a_2093_3714.n13 2.18453
R25470 a_2093_3714.n13 a_2093_3714.n10 0.735439
R25471 a_2093_3714.n10 a_2093_3714.n12 0.718062
R25472 a_2093_3714.n30 a_2093_3714.n29 0.400769
R25473 a_2093_3714.n18 a_2093_3714.n17 0.400768
R25474 a_2093_3714.n24 a_2093_3714.n23 0.400768
R25475 a_2093_3714.n35 a_2093_3714.n34 0.400768
R25476 a_2093_3714.n40 a_2093_3714.n39 0.400768
R25477 a_2093_3714.n48 a_2093_3714.n47 0.40076
R25478 a_2093_3714.n1 a_2093_3714.n0 0.261498
R25479 a_2093_3714.n6 a_2093_3714.n5 0.261477
R25480 a_2093_3714.n3 a_2093_3714.n2 0.261477
R25481 a_2093_3714.n9 a_2093_3714.n8 0.261136
R25482 a_2151_594.n7 a_2151_594.t0 60.2505
R25483 a_2151_594.n64 a_2151_594.t2 60.2505
R25484 a_2151_594.n21 a_2151_594.t9 60.2505
R25485 a_2151_594.n42 a_2151_594.t8 60.2505
R25486 a_2151_594.n4 a_2151_594.n73 9.3005
R25487 a_2151_594.n3 a_2151_594.n57 9.3005
R25488 a_2151_594.n2 a_2151_594.n51 9.3005
R25489 a_2151_594.n1 a_2151_594.n35 9.3005
R25490 a_2151_594.n1 a_2151_594.n34 9.3005
R25491 a_2151_594.n2 a_2151_594.n52 9.3005
R25492 a_2151_594.n2 a_2151_594.n50 9.3005
R25493 a_2151_594.n50 a_2151_594.n49 9.3005
R25494 a_2151_594.n1 a_2151_594.n41 9.3005
R25495 a_2151_594.n41 a_2151_594.n40 9.3005
R25496 a_2151_594.n0 a_2151_594.n29 9.3005
R25497 a_2151_594.n0 a_2151_594.n30 9.3005
R25498 a_2151_594.n0 a_2151_594.n28 9.3005
R25499 a_2151_594.n28 a_2151_594.n27 9.3005
R25500 a_2151_594.n4 a_2151_594.n74 9.3005
R25501 a_2151_594.n4 a_2151_594.n72 9.3005
R25502 a_2151_594.n72 a_2151_594.n71 9.3005
R25503 a_2151_594.n3 a_2151_594.n63 9.3005
R25504 a_2151_594.n63 a_2151_594.n62 9.3005
R25505 a_2151_594.n3 a_2151_594.n56 9.3005
R25506 a_2151_594.n5 a_2151_594.n14 9.3005
R25507 a_2151_594.n14 a_2151_594.n13 9.3005
R25508 a_2151_594.n5 a_2151_594.n16 9.3005
R25509 a_2151_594.n5 a_2151_594.n15 9.3005
R25510 a_2151_594.n43 a_2151_594.n42 8.76429
R25511 a_2151_594.n65 a_2151_594.n64 8.76429
R25512 a_2151_594.n26 a_2151_594.n25 8.21641
R25513 a_2151_594.n48 a_2151_594.n47 8.21641
R25514 a_2151_594.n39 a_2151_594.n38 8.21641
R25515 a_2151_594.n70 a_2151_594.n69 8.21641
R25516 a_2151_594.n61 a_2151_594.n60 8.21641
R25517 a_2151_594.n12 a_2151_594.n11 8.21641
R25518 a_2151_594.n22 a_2151_594.n21 6.92011
R25519 a_2151_594.n8 a_2151_594.n7 6.92007
R25520 a_2151_594.n24 a_2151_594.n23 5.64756
R25521 a_2151_594.n46 a_2151_594.n45 5.64756
R25522 a_2151_594.n37 a_2151_594.n36 5.64756
R25523 a_2151_594.n68 a_2151_594.n67 5.64756
R25524 a_2151_594.n59 a_2151_594.n58 5.64756
R25525 a_2151_594.n10 a_2151_594.n9 5.64756
R25526 a_2151_594.n97 a_2151_594.t6 5.5395
R25527 a_2151_594.n97 a_2151_594.t5 5.5395
R25528 a_2151_594.n115 a_2151_594.t4 5.5395
R25529 a_2151_594.t7 a_2151_594.n115 5.5395
R25530 a_2151_594.n78 a_2151_594.n77 5.27461
R25531 a_2151_594.n31 a_2151_594.n20 4.76425
R25532 a_2151_594.n53 a_2151_594.n19 4.76425
R25533 a_2151_594.n33 a_2151_594.n32 4.76425
R25534 a_2151_594.n75 a_2151_594.n18 4.76425
R25535 a_2151_594.n55 a_2151_594.n54 4.76425
R25536 a_2151_594.n17 a_2151_594.n6 4.76425
R25537 a_2151_594.n44 a_2151_594.n43 4.6505
R25538 a_2151_594.n66 a_2151_594.n65 4.6505
R25539 a_2151_594.n104 a_2151_594.n103 4.51815
R25540 a_2151_594.n109 a_2151_594.n108 4.51815
R25541 a_2151_594.n79 a_2151_594.n90 6.0005
R25542 a_2151_594.n80 a_2151_594.n82 4.5005
R25543 a_2151_594.n96 a_2151_594.n101 4.5005
R25544 a_2151_594.n92 a_2151_594.n112 4.5005
R25545 a_2151_594.n5 a_2151_594.n8 3.47842
R25546 a_2151_594.n0 a_2151_594.n22 3.47753
R25547 a_2151_594.n90 a_2151_594.n89 3.38238
R25548 a_2151_594.n95 a_2151_594.t1 3.3065
R25549 a_2151_594.n95 a_2151_594.t3 3.3065
R25550 a_2151_594.n84 a_2151_594.n95 3.21134
R25551 a_2151_594.n102 a_2151_594.n104 3.03311
R25552 a_2151_594.n93 a_2151_594.n109 3.03311
R25553 a_2151_594.n115 a_2151_594.n91 2.85325
R25554 a_2151_594.n94 a_2151_594.n84 2.63601
R25555 a_2151_594.n100 a_2151_594.n99 2.25932
R25556 a_2151_594.n111 a_2151_594.n110 2.25932
R25557 a_2151_594.n90 a_2151_594.n88 1.88285
R25558 a_2151_594.n115 a_2151_594.n114 1.64452
R25559 a_2151_594.n98 a_2151_594.n97 1.64446
R25560 a_2151_594.n94 a_2151_594.n106 1.62064
R25561 a_2151_594.n83 a_2151_594.n86 6.0005
R25562 a_2151_594.n86 a_2151_594.n85 1.12991
R25563 a_2151_594.n27 a_2151_594.n26 1.09595
R25564 a_2151_594.n49 a_2151_594.n48 1.09595
R25565 a_2151_594.n40 a_2151_594.n39 1.09595
R25566 a_2151_594.n71 a_2151_594.n70 1.09595
R25567 a_2151_594.n62 a_2151_594.n61 1.09595
R25568 a_2151_594.n13 a_2151_594.n12 1.09595
R25569 a_2151_594.n101 a_2151_594.n100 0.753441
R25570 a_2151_594.n28 a_2151_594.n24 0.753441
R25571 a_2151_594.n50 a_2151_594.n46 0.753441
R25572 a_2151_594.n41 a_2151_594.n37 0.753441
R25573 a_2151_594.n72 a_2151_594.n68 0.753441
R25574 a_2151_594.n63 a_2151_594.n59 0.753441
R25575 a_2151_594.n14 a_2151_594.n10 0.753441
R25576 a_2151_594.n88 a_2151_594.n87 0.753441
R25577 a_2151_594.n112 a_2151_594.n111 0.753441
R25578 a_2151_594.n107 a_2151_594.n94 0.599869
R25579 a_2151_594.n106 a_2151_594.n105 0.561382
R25580 a_2151_594.n114 a_2151_594.n113 0.462706
R25581 a_2151_594.n55 a_2151_594.n53 0.458354
R25582 a_2151_594.n33 a_2151_594.n31 0.458354
R25583 a_2151_594.n82 a_2151_594.n81 0.376971
R25584 a_2151_594.n76 a_2151_594.n17 0.229427
R25585 a_2151_594.n76 a_2151_594.n75 0.229427
R25586 a_2151_594.n78 a_2151_594.n76 0.191391
R25587 a_2151_594.n4 a_2151_594.n66 0.190717
R25588 a_2151_594.n66 a_2151_594.n3 0.190717
R25589 a_2151_594.n2 a_2151_594.n44 0.190717
R25590 a_2151_594.n44 a_2151_594.n1 0.190717
R25591 a_2151_594.n83 a_2151_594.n84 0.0960207
R25592 a_2151_594.n102 a_2151_594.n96 0.135435
R25593 a_2151_594.n92 a_2151_594.n93 0.134305
R25594 a_2151_594.n79 a_2151_594.n83 0.0765135
R25595 a_2151_594.n80 a_2151_594.n78 0.125375
R25596 a_2151_594.n106 a_2151_594.n102 0.0711242
R25597 a_2151_594.n93 a_2151_594.n107 0.0536188
R25598 a_2151_594.n113 a_2151_594.n92 0.0954783
R25599 a_2151_594.n96 a_2151_594.n98 0.55664
R25600 a_2151_594.n80 a_2151_594.n79 1.53935
R25601 a_2151_594.n17 a_2151_594.n5 0.205546
R25602 a_2151_594.n75 a_2151_594.n4 0.205546
R25603 a_2151_594.n3 a_2151_594.n55 0.205546
R25604 a_2151_594.n53 a_2151_594.n2 0.205546
R25605 a_2151_594.n1 a_2151_594.n33 0.205546
R25606 a_2151_594.n31 a_2151_594.n0 0.205546
R25607 a_2551_620.n27 a_2551_620.t6 60.2505
R25608 a_2551_620.n48 a_2551_620.t7 60.2505
R25609 a_2551_620.n70 a_2551_620.t4 60.2505
R25610 a_2551_620.n82 a_2551_620.t2 60.2505
R25611 a_2551_620.n1 a_2551_620.n90 9.3005
R25612 a_2551_620.n1 a_2551_620.n91 9.3005
R25613 a_2551_620.n1 a_2551_620.n89 9.3005
R25614 a_2551_620.n89 a_2551_620.n88 9.3005
R25615 a_2551_620.n2 a_2551_620.n79 9.3005
R25616 a_2551_620.n3 a_2551_620.n63 9.3005
R25617 a_2551_620.n3 a_2551_620.n62 9.3005
R25618 a_2551_620.n3 a_2551_620.n69 9.3005
R25619 a_2551_620.n69 a_2551_620.n68 9.3005
R25620 a_2551_620.n2 a_2551_620.n78 9.3005
R25621 a_2551_620.n78 a_2551_620.n77 9.3005
R25622 a_2551_620.n2 a_2551_620.n80 9.3005
R25623 a_2551_620.n4 a_2551_620.n57 9.3005
R25624 a_2551_620.n5 a_2551_620.n41 9.3005
R25625 a_2551_620.n5 a_2551_620.n40 9.3005
R25626 a_2551_620.n5 a_2551_620.n47 9.3005
R25627 a_2551_620.n47 a_2551_620.n46 9.3005
R25628 a_2551_620.n4 a_2551_620.n56 9.3005
R25629 a_2551_620.n56 a_2551_620.n55 9.3005
R25630 a_2551_620.n4 a_2551_620.n58 9.3005
R25631 a_2551_620.n6 a_2551_620.n35 9.3005
R25632 a_2551_620.n6 a_2551_620.n34 9.3005
R25633 a_2551_620.n34 a_2551_620.n33 9.3005
R25634 a_2551_620.n6 a_2551_620.n36 9.3005
R25635 a_2551_620.n7 a_2551_620.n98 9.3005
R25636 a_2551_620.n7 a_2551_620.n97 9.3005
R25637 a_2551_620.n100 a_2551_620.n99 9.3005
R25638 a_2551_620.n102 a_2551_620.n101 9.3005
R25639 a_2551_620.n104 a_2551_620.n103 9.3005
R25640 a_2551_620.n0 a_2551_620.n105 9.3005
R25641 a_2551_620.n125 a_2551_620.n112 9.909
R25642 a_2551_620.n125 a_2551_620.n113 11.0386
R25643 a_2551_620.n125 a_2551_620.n124 8.89115
R25644 a_2551_620.n125 a_2551_620.n121 8.88036
R25645 a_2551_620.n125 a_2551_620.n118 8.86963
R25646 a_2551_620.n125 a_2551_620.n115 8.85895
R25647 a_2551_620.n71 a_2551_620.n70 8.76429
R25648 a_2551_620.n49 a_2551_620.n48 8.76429
R25649 a_2551_620.n32 a_2551_620.n31 7.45411
R25650 a_2551_620.n45 a_2551_620.n44 7.45411
R25651 a_2551_620.n54 a_2551_620.n53 7.45411
R25652 a_2551_620.n67 a_2551_620.n66 7.45411
R25653 a_2551_620.n76 a_2551_620.n75 7.45411
R25654 a_2551_620.n87 a_2551_620.n86 7.45411
R25655 a_2551_620.n20 a_2551_620.n19 7.45281
R25656 a_2551_620.n28 a_2551_620.n27 6.80105
R25657 a_2551_620.n83 a_2551_620.n82 6.80105
R25658 a_2551_620.n0 a_2551_620.n11 6.29716
R25659 a_2551_620.n30 a_2551_620.n29 5.64756
R25660 a_2551_620.n43 a_2551_620.n42 5.64756
R25661 a_2551_620.n52 a_2551_620.n51 5.64756
R25662 a_2551_620.n65 a_2551_620.n64 5.64756
R25663 a_2551_620.n74 a_2551_620.n73 5.64756
R25664 a_2551_620.n85 a_2551_620.n84 5.64756
R25665 a_2551_620.n125 a_2551_620.t5 5.5395
R25666 a_2551_620.t3 a_2551_620.n125 5.5395
R25667 a_2551_620.n96 a_2551_620.n95 4.95534
R25668 a_2551_620.n37 a_2551_620.n26 4.73575
R25669 a_2551_620.n39 a_2551_620.n38 4.73575
R25670 a_2551_620.n59 a_2551_620.n25 4.73575
R25671 a_2551_620.n61 a_2551_620.n60 4.73575
R25672 a_2551_620.n81 a_2551_620.n24 4.73575
R25673 a_2551_620.n93 a_2551_620.n92 4.73575
R25674 a_2551_620.n72 a_2551_620.n71 4.6505
R25675 a_2551_620.n50 a_2551_620.n49 4.6505
R25676 a_2551_620.n8 a_2551_620.n21 4.5005
R25677 a_2551_620.n9 a_2551_620.n20 4.5005
R25678 a_2551_620.n8 a_2551_620.n108 4.5005
R25679 a_2551_620.n0 a_2551_620.n23 4.5005
R25680 a_2551_620.n9 a_2551_620.n110 4.5005
R25681 a_2551_620.n6 a_2551_620.n28 3.42768
R25682 a_2551_620.n1 a_2551_620.n83 3.42768
R25683 a_2551_620.n110 a_2551_620.n109 3.38874
R25684 a_2551_620.n117 a_2551_620.n116 3.38874
R25685 a_2551_620.n17 a_2551_620.n16 3.38238
R25686 a_2551_620.n106 a_2551_620.t1 3.3065
R25687 a_2551_620.n106 a_2551_620.t0 3.3065
R25688 a_2551_620.n11 a_2551_620.n106 3.21133
R25689 a_2551_620.n20 a_2551_620.n18 2.63579
R25690 a_2551_620.n120 a_2551_620.n119 2.63579
R25691 a_2551_620.n17 a_2551_620.n15 1.88285
R25692 a_2551_620.n23 a_2551_620.n22 1.88285
R25693 a_2551_620.n123 a_2551_620.n122 1.88285
R25694 a_2551_620.n125 a_2551_620.n111 1.67004
R25695 a_2551_620.n108 a_2551_620.n107 1.50638
R25696 a_2551_620.n10 a_2551_620.n13 6.0005
R25697 a_2551_620.n13 a_2551_620.n12 1.12991
R25698 a_2551_620.n33 a_2551_620.n32 0.994314
R25699 a_2551_620.n46 a_2551_620.n45 0.994314
R25700 a_2551_620.n55 a_2551_620.n54 0.994314
R25701 a_2551_620.n68 a_2551_620.n67 0.994314
R25702 a_2551_620.n77 a_2551_620.n76 0.994314
R25703 a_2551_620.n88 a_2551_620.n87 0.994314
R25704 a_2551_620.n111 a_2551_620.n9 0.944917
R25705 a_2551_620.n15 a_2551_620.n14 0.753441
R25706 a_2551_620.n34 a_2551_620.n30 0.753441
R25707 a_2551_620.n47 a_2551_620.n43 0.753441
R25708 a_2551_620.n56 a_2551_620.n52 0.753441
R25709 a_2551_620.n69 a_2551_620.n65 0.753441
R25710 a_2551_620.n78 a_2551_620.n74 0.753441
R25711 a_2551_620.n89 a_2551_620.n85 0.753441
R25712 a_2551_620.n39 a_2551_620.n37 0.458354
R25713 a_2551_620.n61 a_2551_620.n59 0.458354
R25714 a_2551_620.n94 a_2551_620.n81 0.229427
R25715 a_2551_620.n94 a_2551_620.n93 0.229427
R25716 a_2551_620.n96 a_2551_620.n94 0.215848
R25717 a_2551_620.n104 a_2551_620.n102 0.190717
R25718 a_2551_620.n50 a_2551_620.n5 0.190717
R25719 a_2551_620.n4 a_2551_620.n50 0.190717
R25720 a_2551_620.n72 a_2551_620.n3 0.190717
R25721 a_2551_620.n2 a_2551_620.n72 0.190717
R25722 a_2551_620.n0 a_2551_620.n104 0.190717
R25723 a_2551_620.n102 a_2551_620.n100 0.190717
R25724 a_2551_620.n7 a_2551_620.n96 0.164777
R25725 a_2551_620.n115 a_2551_620.n114 0.160869
R25726 a_2551_620.n118 a_2551_620.n117 0.14967
R25727 a_2551_620.n121 a_2551_620.n120 0.138414
R25728 a_2551_620.n124 a_2551_620.n123 0.127101
R25729 a_2551_620.n10 a_2551_620.n11 0.0960207
R25730 a_2551_620.n17 a_2551_620.n10 6.07651
R25731 a_2551_620.n8 a_2551_620.n0 0.208476
R25732 a_2551_620.n37 a_2551_620.n6 0.205546
R25733 a_2551_620.n5 a_2551_620.n39 0.205546
R25734 a_2551_620.n59 a_2551_620.n4 0.205546
R25735 a_2551_620.n3 a_2551_620.n61 0.205546
R25736 a_2551_620.n81 a_2551_620.n2 0.205546
R25737 a_2551_620.n93 a_2551_620.n1 0.205546
R25738 a_2551_620.n100 a_2551_620.n7 0.190717
R25739 a_2551_620.n9 a_2551_620.n8 0.135431
R25740 a_5299_3714.n53 a_5299_3714.t2 60.2505
R25741 a_5299_3714.n31 a_5299_3714.t9 60.2505
R25742 a_5299_3714.n9 a_5299_3714.t8 60.2505
R25743 a_5299_3714.n66 a_5299_3714.t0 60.2505
R25744 a_5299_3714.n0 a_5299_3714.n74 9.3005
R25745 a_5299_3714.n0 a_5299_3714.n75 9.3005
R25746 a_5299_3714.n0 a_5299_3714.n73 9.3005
R25747 a_5299_3714.n73 a_5299_3714.n72 9.3005
R25748 a_5299_3714.n3 a_5299_3714.n41 9.3005
R25749 a_5299_3714.n4 a_5299_3714.n23 9.3005
R25750 a_5299_3714.n5 a_5299_3714.n18 9.3005
R25751 a_5299_3714.n5 a_5299_3714.n17 9.3005
R25752 a_5299_3714.n5 a_5299_3714.n16 9.3005
R25753 a_5299_3714.n16 a_5299_3714.n15 9.3005
R25754 a_5299_3714.n4 a_5299_3714.n24 9.3005
R25755 a_5299_3714.n4 a_5299_3714.n30 9.3005
R25756 a_5299_3714.n30 a_5299_3714.n29 9.3005
R25757 a_5299_3714.n3 a_5299_3714.n40 9.3005
R25758 a_5299_3714.n3 a_5299_3714.n39 9.3005
R25759 a_5299_3714.n39 a_5299_3714.n38 9.3005
R25760 a_5299_3714.n2 a_5299_3714.n45 9.3005
R25761 a_5299_3714.n2 a_5299_3714.n52 9.3005
R25762 a_5299_3714.n52 a_5299_3714.n51 9.3005
R25763 a_5299_3714.n2 a_5299_3714.n46 9.3005
R25764 a_5299_3714.n1 a_5299_3714.n61 9.3005
R25765 a_5299_3714.n61 a_5299_3714.n60 9.3005
R25766 a_5299_3714.n1 a_5299_3714.n63 9.3005
R25767 a_5299_3714.n1 a_5299_3714.n62 9.3005
R25768 a_5299_3714.n32 a_5299_3714.n31 8.76429
R25769 a_5299_3714.n54 a_5299_3714.n53 8.76429
R25770 a_5299_3714.n14 a_5299_3714.n13 8.21641
R25771 a_5299_3714.n28 a_5299_3714.n27 8.21641
R25772 a_5299_3714.n37 a_5299_3714.n36 8.21641
R25773 a_5299_3714.n71 a_5299_3714.n70 8.21641
R25774 a_5299_3714.n50 a_5299_3714.n49 8.21641
R25775 a_5299_3714.n59 a_5299_3714.n58 8.21641
R25776 a_5299_3714.n10 a_5299_3714.n9 6.92242
R25777 a_5299_3714.n67 a_5299_3714.n66 6.92012
R25778 a_5299_3714.n12 a_5299_3714.n11 5.64756
R25779 a_5299_3714.n26 a_5299_3714.n25 5.64756
R25780 a_5299_3714.n35 a_5299_3714.n34 5.64756
R25781 a_5299_3714.n69 a_5299_3714.n68 5.64756
R25782 a_5299_3714.n48 a_5299_3714.n47 5.64756
R25783 a_5299_3714.n57 a_5299_3714.n56 5.64756
R25784 a_5299_3714.n98 a_5299_3714.t5 5.5395
R25785 a_5299_3714.n98 a_5299_3714.t4 5.5395
R25786 a_5299_3714.n115 a_5299_3714.t6 5.5395
R25787 a_5299_3714.t7 a_5299_3714.n115 5.5395
R25788 a_5299_3714.n79 a_5299_3714.n78 5.27461
R25789 a_5299_3714.n20 a_5299_3714.n19 4.76425
R25790 a_5299_3714.n22 a_5299_3714.n21 4.76425
R25791 a_5299_3714.n43 a_5299_3714.n42 4.76425
R25792 a_5299_3714.n76 a_5299_3714.n65 4.76425
R25793 a_5299_3714.n44 a_5299_3714.n8 4.76425
R25794 a_5299_3714.n64 a_5299_3714.n7 4.76425
R25795 a_5299_3714.n33 a_5299_3714.n32 4.6505
R25796 a_5299_3714.n55 a_5299_3714.n54 4.6505
R25797 a_5299_3714.n105 a_5299_3714.n104 4.51815
R25798 a_5299_3714.n110 a_5299_3714.n109 4.51815
R25799 a_5299_3714.n80 a_5299_3714.n91 6.0005
R25800 a_5299_3714.n81 a_5299_3714.n83 4.5005
R25801 a_5299_3714.n97 a_5299_3714.n102 4.5005
R25802 a_5299_3714.n93 a_5299_3714.n113 4.5005
R25803 a_5299_3714.n0 a_5299_3714.n67 3.47756
R25804 a_5299_3714.n5 a_5299_3714.n10 3.4767
R25805 a_5299_3714.n91 a_5299_3714.n90 3.38238
R25806 a_5299_3714.n95 a_5299_3714.t3 3.3065
R25807 a_5299_3714.n95 a_5299_3714.t1 3.3065
R25808 a_5299_3714.n85 a_5299_3714.n95 3.21134
R25809 a_5299_3714.n103 a_5299_3714.n105 3.03311
R25810 a_5299_3714.n94 a_5299_3714.n110 3.03311
R25811 a_5299_3714.n115 a_5299_3714.n92 2.85325
R25812 a_5299_3714.n6 a_5299_3714.n85 2.81636
R25813 a_5299_3714.n101 a_5299_3714.n100 2.25932
R25814 a_5299_3714.n112 a_5299_3714.n111 2.25932
R25815 a_5299_3714.n91 a_5299_3714.n89 1.88285
R25816 a_5299_3714.n99 a_5299_3714.n98 1.64453
R25817 a_5299_3714.n115 a_5299_3714.n114 1.64449
R25818 a_5299_3714.n84 a_5299_3714.n87 6.0005
R25819 a_5299_3714.n87 a_5299_3714.n86 1.12991
R25820 a_5299_3714.n15 a_5299_3714.n14 1.09595
R25821 a_5299_3714.n29 a_5299_3714.n28 1.09595
R25822 a_5299_3714.n38 a_5299_3714.n37 1.09595
R25823 a_5299_3714.n72 a_5299_3714.n71 1.09595
R25824 a_5299_3714.n51 a_5299_3714.n50 1.09595
R25825 a_5299_3714.n60 a_5299_3714.n59 1.09595
R25826 a_5299_3714.n107 a_5299_3714.n106 0.760382
R25827 a_5299_3714.n16 a_5299_3714.n12 0.753441
R25828 a_5299_3714.n30 a_5299_3714.n26 0.753441
R25829 a_5299_3714.n39 a_5299_3714.n35 0.753441
R25830 a_5299_3714.n73 a_5299_3714.n69 0.753441
R25831 a_5299_3714.n52 a_5299_3714.n48 0.753441
R25832 a_5299_3714.n61 a_5299_3714.n57 0.753441
R25833 a_5299_3714.n89 a_5299_3714.n88 0.753441
R25834 a_5299_3714.n102 a_5299_3714.n101 0.753441
R25835 a_5299_3714.n113 a_5299_3714.n112 0.753441
R25836 a_5299_3714.n6 a_5299_3714.n107 0.678625
R25837 a_5299_3714.n106 a_5299_3714.n96 0.573452
R25838 a_5299_3714.n22 a_5299_3714.n20 0.458354
R25839 a_5299_3714.n44 a_5299_3714.n43 0.458354
R25840 a_5299_3714.n83 a_5299_3714.n82 0.376971
R25841 a_5299_3714.n77 a_5299_3714.n64 0.229427
R25842 a_5299_3714.n77 a_5299_3714.n76 0.229427
R25843 a_5299_3714.n79 a_5299_3714.n77 0.191391
R25844 a_5299_3714.n33 a_5299_3714.n4 0.190717
R25845 a_5299_3714.n3 a_5299_3714.n33 0.190717
R25846 a_5299_3714.n55 a_5299_3714.n2 0.190717
R25847 a_5299_3714.n1 a_5299_3714.n55 0.190717
R25848 a_5299_3714.n84 a_5299_3714.n85 0.0960207
R25849 a_5299_3714.n93 a_5299_3714.n94 0.135434
R25850 a_5299_3714.n103 a_5299_3714.n97 0.13503
R25851 a_5299_3714.n80 a_5299_3714.n84 0.0765135
R25852 a_5299_3714.n81 a_5299_3714.n79 0.125375
R25853 a_5299_3714.n106 a_5299_3714.n103 0.0591603
R25854 a_5299_3714.n94 a_5299_3714.n108 0.0540944
R25855 a_5299_3714.n114 a_5299_3714.n93 0.556715
R25856 a_5299_3714.n97 a_5299_3714.n99 0.556623
R25857 a_5299_3714.n81 a_5299_3714.n80 1.53935
R25858 a_5299_3714.n108 a_5299_3714.n6 0.620875
R25859 a_5299_3714.n20 a_5299_3714.n5 0.205546
R25860 a_5299_3714.n4 a_5299_3714.n22 0.205546
R25861 a_5299_3714.n43 a_5299_3714.n3 0.205546
R25862 a_5299_3714.n2 a_5299_3714.n44 0.205546
R25863 a_5299_3714.n64 a_5299_3714.n1 0.205546
R25864 a_5299_3714.n76 a_5299_3714.n0 0.205546
R25865 a_2093_1782.n88 a_2093_1782.n22 8.05594
R25866 a_2093_1782.n88 a_2093_1782.n20 8.02924
R25867 a_2093_1782.n87 a_2093_1782.n86 6.13632
R25868 a_2093_1782.n83 a_2093_1782.n82 5.61043
R25869 a_2093_1782.n48 a_2093_1782.n47 5.61041
R25870 a_2093_1782.n51 a_2093_1782.n50 5.61041
R25871 a_2093_1782.n28 a_2093_1782.n27 5.61037
R25872 a_2093_1782.n62 a_2093_1782.n61 5.61037
R25873 a_2093_1782.n81 a_2093_1782.n80 5.61037
R25874 a_2093_1782.n8 a_2093_1782.n78 4.5005
R25875 a_2093_1782.n15 a_2093_1782.n70 4.5005
R25876 a_2093_1782.n6 a_2093_1782.n66 4.5005
R25877 a_2093_1782.n4 a_2093_1782.n59 4.5005
R25878 a_2093_1782.n14 a_2093_1782.n55 4.5005
R25879 a_2093_1782.n38 a_2093_1782.n41 4.5005
R25880 a_2093_1782.n13 a_2093_1782.n36 4.5005
R25881 a_2093_1782.n0 a_2093_1782.n32 4.5005
R25882 a_2093_1782.n2 a_2093_1782.n45 4.5005
R25883 a_2093_1782.n16 a_2093_1782.n74 4.5005
R25884 a_2093_1782.n25 a_2093_1782.n24 4.5005
R25885 a_2093_1782.n17 a_2093_1782.n85 4.5005
R25886 a_2093_1782.n36 a_2093_1782.n35 3.76521
R25887 a_2093_1782.n41 a_2093_1782.n40 3.76521
R25888 a_2093_1782.n55 a_2093_1782.n54 3.76521
R25889 a_2093_1782.n70 a_2093_1782.n69 3.76521
R25890 a_2093_1782.n74 a_2093_1782.n73 3.76521
R25891 a_2093_1782.n24 a_2093_1782.n23 3.76521
R25892 a_2093_1782.n32 a_2093_1782.n30 3.38874
R25893 a_2093_1782.n45 a_2093_1782.n43 3.38874
R25894 a_2093_1782.n59 a_2093_1782.n57 3.38874
R25895 a_2093_1782.n66 a_2093_1782.n64 3.38874
R25896 a_2093_1782.n78 a_2093_1782.n76 3.38874
R25897 a_2093_1782.n33 a_2093_1782.t6 3.3065
R25898 a_2093_1782.n33 a_2093_1782.t8 3.3065
R25899 a_2093_1782.n37 a_2093_1782.t9 3.3065
R25900 a_2093_1782.n37 a_2093_1782.t11 3.3065
R25901 a_2093_1782.n52 a_2093_1782.t10 3.3065
R25902 a_2093_1782.n52 a_2093_1782.t4 3.3065
R25903 a_2093_1782.n67 a_2093_1782.t3 3.3065
R25904 a_2093_1782.n67 a_2093_1782.t2 3.3065
R25905 a_2093_1782.n71 a_2093_1782.t1 3.3065
R25906 a_2093_1782.n71 a_2093_1782.t0 3.3065
R25907 a_2093_1782.t5 a_2093_1782.n88 3.3065
R25908 a_2093_1782.n88 a_2093_1782.t7 3.3065
R25909 a_2093_1782.n32 a_2093_1782.n31 3.01226
R25910 a_2093_1782.n45 a_2093_1782.n44 3.01226
R25911 a_2093_1782.n59 a_2093_1782.n58 3.01226
R25912 a_2093_1782.n66 a_2093_1782.n65 3.01226
R25913 a_2093_1782.n78 a_2093_1782.n77 3.01226
R25914 a_2093_1782.n85 a_2093_1782.n84 3.01226
R25915 a_2093_1782.n36 a_2093_1782.n34 2.63579
R25916 a_2093_1782.n41 a_2093_1782.n39 2.63579
R25917 a_2093_1782.n55 a_2093_1782.n53 2.63579
R25918 a_2093_1782.n70 a_2093_1782.n68 2.63579
R25919 a_2093_1782.n74 a_2093_1782.n72 2.63579
R25920 a_2093_1782.n11 a_2093_1782.n9 2.18375
R25921 a_2093_1782.n18 a_2093_1782.n1 2.18356
R25922 a_2093_1782.n38 a_2093_1782.n37 1.85087
R25923 a_2093_1782.n13 a_2093_1782.n33 1.85087
R25924 a_2093_1782.n14 a_2093_1782.n52 1.85087
R25925 a_2093_1782.n15 a_2093_1782.n67 1.85087
R25926 a_2093_1782.n16 a_2093_1782.n71 1.85087
R25927 a_2093_1782.n87 a_2093_1782.n25 1.48737
R25928 a_2093_1782.n12 a_2093_1782.n5 1.48434
R25929 a_2093_1782.n18 a_2093_1782.n3 1.48434
R25930 a_2093_1782.n19 a_2093_1782.n7 1.48434
R25931 a_2093_1782.n10 a_2093_1782.n11 1.48434
R25932 a_2093_1782.n11 a_2093_1782.n19 0.736217
R25933 a_2093_1782.n19 a_2093_1782.n12 0.735439
R25934 a_2093_1782.n12 a_2093_1782.n18 0.718062
R25935 a_2093_1782.n27 a_2093_1782.n26 0.461175
R25936 a_2093_1782.n47 a_2093_1782.n46 0.461175
R25937 a_2093_1782.n50 a_2093_1782.n49 0.461175
R25938 a_2093_1782.n61 a_2093_1782.n60 0.461175
R25939 a_2093_1782.n80 a_2093_1782.n79 0.461175
R25940 a_2093_1782.n30 a_2093_1782.n29 0.430121
R25941 a_2093_1782.n43 a_2093_1782.n42 0.430121
R25942 a_2093_1782.n57 a_2093_1782.n56 0.430121
R25943 a_2093_1782.n64 a_2093_1782.n63 0.430121
R25944 a_2093_1782.n76 a_2093_1782.n75 0.430121
R25945 a_2093_1782.n22 a_2093_1782.n21 0.429625
R25946 a_2093_1782.n88 a_2093_1782.n87 0.363993
R25947 a_2093_1782.n9 a_2093_1782.n81 0.297864
R25948 a_2093_1782.n1 a_2093_1782.n28 0.297864
R25949 a_2093_1782.n7 a_2093_1782.n62 0.297864
R25950 a_2093_1782.n3 a_2093_1782.n48 0.297822
R25951 a_2093_1782.n5 a_2093_1782.n51 0.297822
R25952 a_2093_1782.n10 a_2093_1782.n83 0.297796
R25953 a_2093_1782.n17 a_2093_1782.n10 0.155159
R25954 a_2093_1782.n0 a_2093_1782.n13 0.14384
R25955 a_2093_1782.n2 a_2093_1782.n38 0.142841
R25956 a_2093_1782.n6 a_2093_1782.n15 0.142841
R25957 a_2093_1782.n4 a_2093_1782.n14 0.142841
R25958 a_2093_1782.n8 a_2093_1782.n16 0.141862
R25959 a_2093_1782.n9 a_2093_1782.n8 0.136602
R25960 a_2093_1782.n7 a_2093_1782.n6 0.136602
R25961 a_2093_1782.n5 a_2093_1782.n4 0.136602
R25962 a_2093_1782.n3 a_2093_1782.n2 0.136602
R25963 a_2093_1782.n1 a_2093_1782.n0 0.136602
R25964 a_2093_1782.n25 a_2093_1782.n17 0.124283
R25965 VO.n7 VO.n6 585
R25966 VO.n3 VO.n2 291.406
R25967 VO.n12 VO.t0 194.387
R25968 VO.n5 VO.n4 148.663
R25969 VO.t0 VO.n11 122.728
R25970 VO.n3 VO.t1 22.4191
R25971 VO.n7 VO.n4 10.5541
R25972 VO VO.n5 9.62836
R25973 VO.n18 VO.n17 9.3005
R25974 VO.n15 VO.n14 9.3005
R25975 VO.n8 VO.n7 9.3005
R25976 VO VO.n10 7.00682
R25977 VO VO.n9 6.32867
R25978 VO.n13 VO.n12 5.92892
R25979 VO.n14 VO.n13 4.72813
R25980 VO VO.n11 4.69453
R25981 VO.n10 VO.n0 4.6505
R25982 VO.n16 VO.n1 4.6505
R25983 VO.n10 VO 2.96471
R25984 VO VO.n19 2.51698
R25985 VO.n13 VO 2.42576
R25986 VO.n4 VO.n3 2.19143
R25987 VO.n17 VO 2.15629
R25988 VO.n9 VO.n0 2.04091
R25989 VO.n16 VO.n15 1.75208
R25990 VO.n6 VO.n2 1.61734
R25991 VO.n12 VO 1.61734
R25992 VO.n9 VO.n8 0.816947
R25993 VO.n15 VO.n11 0.795743
R25994 VO.n8 VO.n2 0.674184
R25995 VO.n17 VO.n16 0.539447
R25996 VO.n5 VO 0.343399
R25997 VO.n6 VO 0.269974
R25998 VO.n19 VO.n18 0.0807632
R25999 VO.n14 VO.n1 0.0176053
R26000 VO.n19 VO.n0 0.00971053
R26001 VO.n18 VO.n1 0.00576316
R26002 SELA.n6 SELA.t2 186.374
R26003 SELA.n6 SELA.t3 170.308
R26004 SELA.n7 SELA.n6 139.876
R26005 SELA.n0 SELA.t4 84.8325
R26006 SELA.n1 SELA.t0 84.8325
R26007 SELA.n1 SELA.n0 60.1541
R26008 SELA.n2 SELA.n1 50.1642
R26009 SELA.n0 SELA.t5 48.6825
R26010 SELA.n1 SELA.t1 48.6825
R26011 SELA.n5 SELA 42.9181
R26012 SELA.n4 SELA 17.169
R26013 SELA.n3 SELA.n2 15.2731
R26014 SELA.n11 SELA.n9 14.3125
R26015 SELA.n5 SELA 12.8005
R26016 SELA.n4 SELA.n3 4.77356
R26017 SELA.n8 SELA 2.73914
R26018 SELA SELA.n3 2.13383
R26019 SELA SELA.n7 1.61978
R26020 SELA.n9 SELA.n8 1.31185
R26021 SELA.n2 SELA 1.1768
R26022 SELA SELA.n13 0.979433
R26023 SELA.n7 SELA.n5 0.925801
R26024 SELA.n13 SELA.n12 0.675199
R26025 SELA.n10 SELA 0.34425
R26026 SELA.n13 SELA 0.321549
R26027 SELA SELA.n11 0.0255
R26028 SELA.n11 SELA.n10 0.0194024
R26029 SELA SELA.n4 0.0180439
R26030 SELA.n12 SELA 0.0151341
R26031 SELA.n8 SELA 0.00770734
R26032 SELA.n12 SELA 0.00415854
R26033 SELA.n10 SELA 0.00171951
R26034 SELA.n12 SELA.n9 0.000502048
R26035 DVDD.n4 DVDD.t13 591.327
R26036 DVDD.n6 DVDD.t8 591.327
R26037 DVDD.n15 DVDD.n14 585
R26038 DVDD.n194 DVDD.n181 321.882
R26039 DVDD.n228 DVDD.n181 321.882
R26040 DVDD.n228 DVDD.n179 321.882
R26041 DVDD.n54 DVDD.n41 321.882
R26042 DVDD.n88 DVDD.n41 321.882
R26043 DVDD.n88 DVDD.n39 321.882
R26044 DVDD.n229 DVDD.n180 175.386
R26045 DVDD.n89 DVDD.n40 175.386
R26046 DVDD.n194 DVDD.t2 171.452
R26047 DVDD.n54 DVDD.t27 171.452
R26048 DVDD.n310 DVDD.n309 161.37
R26049 DVDD.n110 DVDD.n103 161.37
R26050 DVDD.n257 DVDD.n256 161.37
R26051 DVDD.n158 DVDD.n157 161.37
R26052 DVDD.n201 DVDD.t3 160.743
R26053 DVDD.n61 DVDD.t28 160.743
R26054 DVDD.n213 DVDD.t7 158.225
R26055 DVDD.n73 DVDD.t20 158.225
R26056 DVDD.n9 DVDD.t14 148.294
R26057 DVDD.t23 DVDD.n305 129.546
R26058 DVDD.t11 DVDD.n105 129.546
R26059 DVDD.t21 DVDD.n252 129.546
R26060 DVDD.t25 DVDD.n153 129.546
R26061 DVDD.n231 DVDD.n230 124.013
R26062 DVDD.n91 DVDD.n90 124.013
R26063 DVDD.n13 DVDD.n10 107.746
R26064 DVDD.n306 DVDD.t23 100.874
R26065 DVDD.n106 DVDD.t11 100.874
R26066 DVDD.n253 DVDD.t21 100.874
R26067 DVDD.n154 DVDD.t25 100.874
R26068 DVDD.t6 DVDD.n229 96.8274
R26069 DVDD.t19 DVDD.n89 96.8274
R26070 DVDD.n307 DVDD.n305 92.5005
R26071 DVDD.n305 DVDD.n304 92.5005
R26072 DVDD.n107 DVDD.n105 92.5005
R26073 DVDD.n105 DVDD.n104 92.5005
R26074 DVDD.n254 DVDD.n252 92.5005
R26075 DVDD.n252 DVDD.n251 92.5005
R26076 DVDD.n155 DVDD.n153 92.5005
R26077 DVDD.n153 DVDD.n152 92.5005
R26078 DVDD.n6 DVDD.n1 92.5005
R26079 DVDD.n6 DVDD.n5 81.7536
R26080 DVDD.n230 DVDD.t6 81.7266
R26081 DVDD.n90 DVDD.t19 81.7266
R26082 DVDD.n308 DVDD.n304 55.3934
R26083 DVDD.n108 DVDD.n104 55.3934
R26084 DVDD.n255 DVDD.n251 55.3934
R26085 DVDD.n156 DVDD.n152 55.3934
R26086 DVDD.n9 DVDD.n2 52.9371
R26087 DVDD.n16 DVDD.n1 49.5938
R26088 DVDD.n7 DVDD.n6 47.5553
R26089 DVDD.n305 DVDD.t15 47.2949
R26090 DVDD.n105 DVDD.t0 47.2949
R26091 DVDD.n252 DVDD.t17 47.2949
R26092 DVDD.n153 DVDD.t4 47.2949
R26093 DVDD.n308 DVDD.n307 46.2505
R26094 DVDD.n108 DVDD.n107 46.2505
R26095 DVDD.n255 DVDD.n254 46.2505
R26096 DVDD.n156 DVDD.n155 46.2505
R26097 DVDD.n9 DVDD.n8 46.2505
R26098 DVDD.n7 DVDD.n2 42.3392
R26099 DVDD.n5 DVDD.n4 40.8773
R26100 DVDD.n195 DVDD.n182 36.1417
R26101 DVDD.n227 DVDD.n182 36.1417
R26102 DVDD.n227 DVDD.n178 36.1417
R26103 DVDD.n231 DVDD.n178 36.1417
R26104 DVDD.n55 DVDD.n42 36.1417
R26105 DVDD.n87 DVDD.n42 36.1417
R26106 DVDD.n87 DVDD.n38 36.1417
R26107 DVDD.n91 DVDD.n38 36.1417
R26108 DVDD.n5 DVDD.n2 34.4168
R26109 DVDD.n309 DVDD.t24 32.8338
R26110 DVDD.n309 DVDD.t16 32.8338
R26111 DVDD.n103 DVDD.t12 32.8338
R26112 DVDD.n103 DVDD.t1 32.8338
R26113 DVDD.n256 DVDD.t22 32.8338
R26114 DVDD.n256 DVDD.t18 32.8338
R26115 DVDD.n157 DVDD.t26 32.8338
R26116 DVDD.n157 DVDD.t5 32.8338
R26117 DVDD.n4 DVDD.n3 32.0046
R26118 DVDD.n8 DVDD.n3 28.4938
R26119 DVDD.n3 DVDD.n1 28.4938
R26120 DVDD.n306 DVDD.n304 26.4697
R26121 DVDD.n307 DVDD.n306 26.4697
R26122 DVDD.n106 DVDD.n104 26.4697
R26123 DVDD.n107 DVDD.n106 26.4697
R26124 DVDD.n253 DVDD.n251 26.4697
R26125 DVDD.n254 DVDD.n253 26.4697
R26126 DVDD.n154 DVDD.n152 26.4697
R26127 DVDD.n155 DVDD.n154 26.4697
R26128 DVDD.n12 DVDD.t9 22.8666
R26129 DVDD.n8 DVDD.n7 21.17
R26130 DVDD.n312 DVDD.n311 17.8772
R26131 DVDD.n109 DVDD.n102 17.8772
R26132 DVDD.n259 DVDD.n258 17.8772
R26133 DVDD.n160 DVDD.n159 17.8772
R26134 DVDD.n311 DVDD.n310 17.4938
R26135 DVDD.n110 DVDD.n109 17.4938
R26136 DVDD.n258 DVDD.n257 17.4938
R26137 DVDD.n159 DVDD.n158 17.4938
R26138 DVDD.n14 DVDD.n13 13.514
R26139 DVDD.t2 DVDD.n180 12.789
R26140 DVDD.t27 DVDD.n40 12.789
R26141 DVDD.n14 DVDD.t10 11.4335
R26142 DVDD.n17 DVDD.n16 10.8623
R26143 DVDD.n201 DVDD.n200 9.3005
R26144 DVDD.n201 DVDD.n190 9.3005
R26145 DVDD.n201 DVDD.n189 9.3005
R26146 DVDD.n61 DVDD.n60 9.3005
R26147 DVDD.n61 DVDD.n50 9.3005
R26148 DVDD.n61 DVDD.n49 9.3005
R26149 DVDD.n12 DVDD.n11 9.3005
R26150 DVDD.n195 DVDD.n194 8.85536
R26151 DVDD.n182 DVDD.n181 8.85536
R26152 DVDD.n181 DVDD.n180 8.85536
R26153 DVDD.n228 DVDD.n227 8.85536
R26154 DVDD.n229 DVDD.n228 8.85536
R26155 DVDD.n179 DVDD.n178 8.85536
R26156 DVDD.n55 DVDD.n54 8.85536
R26157 DVDD.n42 DVDD.n41 8.85536
R26158 DVDD.n41 DVDD.n40 8.85536
R26159 DVDD.n88 DVDD.n87 8.85536
R26160 DVDD.n89 DVDD.n88 8.85536
R26161 DVDD.n39 DVDD.n38 8.85536
R26162 DVDD.n230 DVDD.n179 5.53567
R26163 DVDD.n90 DVDD.n39 5.53567
R26164 DVDD.n310 DVDD.n303 4.6505
R26165 DVDD.n111 DVDD.n110 4.6505
R26166 DVDD.n257 DVDD.n250 4.6505
R26167 DVDD.n158 DVDD.n151 4.6505
R26168 DVDD.n213 DVDD.n177 4.6505
R26169 DVDD.n220 DVDD.n213 4.6505
R26170 DVDD.n202 DVDD.n201 4.6505
R26171 DVDD.n73 DVDD.n37 4.6505
R26172 DVDD.n80 DVDD.n73 4.6505
R26173 DVDD.n62 DVDD.n61 4.6505
R26174 DVDD.n292 DVDD.n26 4.5005
R26175 DVDD.n23 DVDD.n22 4.5005
R26176 DVDD.n284 DVDD.n98 4.5005
R26177 DVDD.n268 DVDD.n116 4.5005
R26178 DVDD.n279 DVDD.n278 4.5005
R26179 DVDD.n263 DVDD.n262 4.5005
R26180 DVDD.n121 DVDD.n120 4.5005
R26181 DVDD.n240 DVDD.n239 4.5005
R26182 DVDD.n164 DVDD.n163 4.5005
R26183 DVDD.n132 DVDD.n131 4.5005
R26184 DVDD.n140 DVDD.n136 4.5005
R26185 DVDD.n197 DVDD.n196 4.5005
R26186 DVDD.n199 DVDD.n198 4.5005
R26187 DVDD.n204 DVDD.n203 4.5005
R26188 DVDD.n207 DVDD.n206 4.5005
R26189 DVDD.n210 DVDD.n209 4.5005
R26190 DVDD.n226 DVDD.n225 4.5005
R26191 DVDD.n223 DVDD.n222 4.5005
R26192 DVDD.n218 DVDD.n217 4.5005
R26193 DVDD.n174 DVDD.n172 4.5005
R26194 DVDD DVDD.n173 4.5005
R26195 DVDD.n205 DVDD.n186 4.5005
R26196 DVDD.n211 DVDD.n183 4.5005
R26197 DVDD.n221 DVDD.n212 4.5005
R26198 DVDD.n216 DVDD.n215 4.5005
R26199 DVDD.n176 DVDD.n175 4.5005
R26200 DVDD.n57 DVDD.n56 4.5005
R26201 DVDD.n59 DVDD.n58 4.5005
R26202 DVDD.n64 DVDD.n63 4.5005
R26203 DVDD.n67 DVDD.n66 4.5005
R26204 DVDD.n70 DVDD.n69 4.5005
R26205 DVDD.n86 DVDD.n85 4.5005
R26206 DVDD.n83 DVDD.n82 4.5005
R26207 DVDD.n78 DVDD.n77 4.5005
R26208 DVDD.n34 DVDD.n32 4.5005
R26209 DVDD DVDD.n33 4.5005
R26210 DVDD.n65 DVDD.n46 4.5005
R26211 DVDD.n71 DVDD.n43 4.5005
R26212 DVDD.n81 DVDD.n72 4.5005
R26213 DVDD.n76 DVDD.n75 4.5005
R26214 DVDD.n36 DVDD.n35 4.5005
R26215 DVDD.n311 DVDD.n308 4.32258
R26216 DVDD.n109 DVDD.n108 4.32258
R26217 DVDD.n258 DVDD.n255 4.32258
R26218 DVDD.n159 DVDD.n156 4.32258
R26219 DVDD.n16 DVDD.n15 3.76521
R26220 DVDD.n16 DVDD.n9 3.34378
R26221 DVDD.n322 DVDD.n321 3.15264
R26222 DVDD.n214 DVDD.n213 3.09891
R26223 DVDD.n74 DVDD.n73 3.09891
R26224 DVDD.n199 DVDD.n195 3.03311
R26225 DVDD.n207 DVDD.n182 3.03311
R26226 DVDD.n227 DVDD.n226 3.03311
R26227 DVDD.n218 DVDD.n178 3.03311
R26228 DVDD DVDD.n231 3.03311
R26229 DVDD.n59 DVDD.n55 3.03311
R26230 DVDD.n67 DVDD.n42 3.03311
R26231 DVDD.n87 DVDD.n86 3.03311
R26232 DVDD.n78 DVDD.n38 3.03311
R26233 DVDD DVDD.n91 3.03311
R26234 DVDD.n15 DVDD.n10 2.82403
R26235 DVDD DVDD.n17 2.78431
R26236 DVDD.n11 DVDD.n0 2.54327
R26237 DVDD.n313 DVDD 1.93032
R26238 DVDD DVDD.n101 1.93032
R26239 DVDD.n260 DVDD 1.93032
R26240 DVDD.n161 DVDD 1.93032
R26241 DVDD.n0 DVDD 1.8288
R26242 DVDD DVDD.n169 1.75727
R26243 DVDD DVDD.n29 1.75727
R26244 DVDD.n313 DVDD 1.61911
R26245 DVDD.n101 DVDD 1.61911
R26246 DVDD.n260 DVDD 1.61911
R26247 DVDD.n161 DVDD 1.61911
R26248 DVDD.n13 DVDD.n12 1.43457
R26249 DVDD.n302 DVDD 1.11892
R26250 DVDD.n112 DVDD 1.11892
R26251 DVDD.n249 DVDD 1.11892
R26252 DVDD.n150 DVDD 1.11892
R26253 DVDD.n272 DVDD.n267 0.433917
R26254 DVDD.n321 DVDD.n320 0.432745
R26255 DVDD.n303 DVDD.n302 0.417167
R26256 DVDD.n112 DVDD.n111 0.417167
R26257 DVDD.n250 DVDD.n249 0.417167
R26258 DVDD.n151 DVDD.n150 0.417167
R26259 DVDD.n27 DVDD 0.377693
R26260 DVDD.n269 DVDD 0.377693
R26261 DVDD.n126 DVDD 0.377693
R26262 DVDD.n137 DVDD 0.377693
R26263 DVDD.n11 DVDD.n10 0.376971
R26264 DVDD.n289 DVDD.n288 0.312991
R26265 DVDD.n236 DVDD.n168 0.296735
R26266 DVDD DVDD.n122 0.272089
R26267 DVDD DVDD.n312 0.268044
R26268 DVDD.n102 DVDD 0.268044
R26269 DVDD DVDD.n259 0.268044
R26270 DVDD DVDD.n160 0.268044
R26271 DVDD DVDD.n133 0.243821
R26272 DVDD DVDD.n18 0.238894
R26273 DVDD.n321 DVDD 0.235903
R26274 DVDD.n282 DVDD 0.234986
R26275 DVDD DVDD.n235 0.206256
R26276 DVDD.n289 DVDD.n95 0.185367
R26277 DVDD.n17 DVDD.n0 0.163151
R26278 DVDD.n312 DVDD.n303 0.158395
R26279 DVDD.n111 DVDD.n102 0.158395
R26280 DVDD.n259 DVDD.n250 0.158395
R26281 DVDD.n160 DVDD.n151 0.158395
R26282 DVDD.n27 DVDD 0.15085
R26283 DVDD.n269 DVDD 0.15085
R26284 DVDD.n126 DVDD 0.15085
R26285 DVDD.n137 DVDD 0.15085
R26286 DVDD.n147 DVDD 0.14163
R26287 DVDD.n246 DVDD 0.14163
R26288 DVDD.n299 DVDD 0.124528
R26289 DVDD DVDD.n281 0.12237
R26290 DVDD.n290 DVDD 0.112517
R26291 DVDD.n237 DVDD.n236 0.110693
R26292 DVDD.n314 DVDD.n313 0.0728282
R26293 DVDD.n101 DVDD.n99 0.0728282
R26294 DVDD.n261 DVDD.n260 0.0728282
R26295 DVDD.n162 DVDD.n161 0.0728282
R26296 DVDD.n28 DVDD.n27 0.0471653
R26297 DVDD.n270 DVDD.n269 0.0471653
R26298 DVDD.n127 DVDD.n126 0.0471653
R26299 DVDD.n138 DVDD.n137 0.0471653
R26300 DVDD.n302 DVDD.n301 0.0401723
R26301 DVDD.n113 DVDD.n112 0.0401723
R26302 DVDD.n249 DVDD.n248 0.0401723
R26303 DVDD.n150 DVDD.n149 0.0401723
R26304 DVDD.n288 DVDD.n287 0.0390074
R26305 DVDD.n267 DVDD.n266 0.0390074
R26306 DVDD.n168 DVDD.n167 0.0390074
R26307 DVDD.n284 DVDD.n283 0.0378134
R26308 DVDD.n263 DVDD.n119 0.0378134
R26309 DVDD.n164 DVDD.n130 0.0378134
R26310 DVDD.n301 DVDD.n22 0.0359671
R26311 DVDD.n28 DVDD.n26 0.0359671
R26312 DVDD.n278 DVDD.n113 0.0359671
R26313 DVDD.n270 DVDD.n268 0.0359671
R26314 DVDD.n248 DVDD.n120 0.0359671
R26315 DVDD.n240 DVDD.n127 0.0359671
R26316 DVDD.n149 DVDD.n131 0.0359671
R26317 DVDD.n138 DVDD.n136 0.0359671
R26318 DVDD.n300 DVDD.n23 0.0357113
R26319 DVDD.n297 DVDD.n23 0.0357113
R26320 DVDD.n297 DVDD.n25 0.0357113
R26321 DVDD.n293 DVDD.n25 0.0357113
R26322 DVDD.n293 DVDD.n292 0.0357113
R26323 DVDD.n292 DVDD.n291 0.0357113
R26324 DVDD.n280 DVDD.n279 0.0357113
R26325 DVDD.n279 DVDD.n114 0.0357113
R26326 DVDD.n275 DVDD.n114 0.0357113
R26327 DVDD.n275 DVDD.n274 0.0357113
R26328 DVDD.n274 DVDD.n116 0.0357113
R26329 DVDD.n271 DVDD.n116 0.0357113
R26330 DVDD.n247 DVDD.n121 0.0357113
R26331 DVDD.n244 DVDD.n121 0.0357113
R26332 DVDD.n244 DVDD.n243 0.0357113
R26333 DVDD.n243 DVDD.n125 0.0357113
R26334 DVDD.n239 DVDD.n125 0.0357113
R26335 DVDD.n239 DVDD.n238 0.0357113
R26336 DVDD.n148 DVDD.n132 0.0357113
R26337 DVDD.n145 DVDD.n132 0.0357113
R26338 DVDD.n145 DVDD.n135 0.0357113
R26339 DVDD.n141 DVDD.n135 0.0357113
R26340 DVDD.n141 DVDD.n140 0.0357113
R26341 DVDD.n140 DVDD.n139 0.0357113
R26342 DVDD.n296 DVDD.n22 0.035465
R26343 DVDD.n296 DVDD.n295 0.035465
R26344 DVDD.n295 DVDD.n294 0.035465
R26345 DVDD.n294 DVDD.n26 0.035465
R26346 DVDD.n278 DVDD.n277 0.035465
R26347 DVDD.n277 DVDD.n276 0.035465
R26348 DVDD.n276 DVDD.n115 0.035465
R26349 DVDD.n268 DVDD.n115 0.035465
R26350 DVDD.n124 DVDD.n120 0.035465
R26351 DVDD.n242 DVDD.n124 0.035465
R26352 DVDD.n242 DVDD.n241 0.035465
R26353 DVDD.n241 DVDD.n240 0.035465
R26354 DVDD.n144 DVDD.n131 0.035465
R26355 DVDD.n144 DVDD.n143 0.035465
R26356 DVDD.n143 DVDD.n142 0.035465
R26357 DVDD.n142 DVDD.n136 0.035465
R26358 DVDD.n317 DVDD.n20 0.0340821
R26359 DVDD.n285 DVDD.n284 0.0340821
R26360 DVDD.n264 DVDD.n263 0.0340821
R26361 DVDD.n165 DVDD.n164 0.0340821
R26362 DVDD.n197 DVDD.n187 0.0333947
R26363 DVDD.n212 DVDD.n171 0.0333947
R26364 DVDD.n175 DVDD.n169 0.0333947
R26365 DVDD.n57 DVDD.n47 0.0333947
R26366 DVDD.n72 DVDD.n31 0.0333947
R26367 DVDD.n35 DVDD.n29 0.0333947
R26368 DVDD.n316 DVDD.n315 0.0333467
R26369 DVDD.n286 DVDD.n98 0.0333467
R26370 DVDD.n262 DVDD.n118 0.0333467
R26371 DVDD.n163 DVDD.n129 0.0333467
R26372 DVDD.n198 DVDD.n193 0.03175
R26373 DVDD.n224 DVDD.n223 0.03175
R26374 DVDD.n58 DVDD.n53 0.03175
R26375 DVDD.n84 DVDD.n83 0.03175
R26376 DVDD.n205 DVDD.n204 0.0284605
R26377 DVDD.n217 DVDD.n216 0.0284605
R26378 DVDD.n65 DVDD.n64 0.0284605
R26379 DVDD.n77 DVDD.n76 0.0284605
R26380 DVDD DVDD.n314 0.0274625
R26381 DVDD.n99 DVDD 0.0274625
R26382 DVDD DVDD.n261 0.0274625
R26383 DVDD DVDD.n162 0.0274625
R26384 DVDD.n322 DVDD 0.0264901
R26385 DVDD DVDD.n322 0.0262353
R26386 DVDD.n193 DVDD.n192 0.0255919
R26387 DVDD.n53 DVDD.n52 0.0255919
R26388 DVDD.n192 DVDD.n191 0.0252368
R26389 DVDD.n191 DVDD.n170 0.0252368
R26390 DVDD.n52 DVDD.n51 0.0252368
R26391 DVDD.n51 DVDD.n30 0.0252368
R26392 DVDD.n225 DVDD.n211 0.0251711
R26393 DVDD.n85 DVDD.n71 0.0251711
R26394 DVDD.n139 DVDD.n134 0.024355
R26395 DVDD.n267 DVDD.n117 0.0242975
R26396 DVDD.n122 DVDD.n117 0.0242975
R26397 DVDD.n147 DVDD.n146 0.024
R26398 DVDD.n146 DVDD.n134 0.024
R26399 DVDD.n246 DVDD.n245 0.024
R26400 DVDD.n245 DVDD.n123 0.024
R26401 DVDD.n237 DVDD.n123 0.024
R26402 DVDD.n220 DVDD.n219 0.0232804
R26403 DVDD.n80 DVDD.n79 0.0232804
R26404 DVDD.n222 DVDD.n184 0.0226963
R26405 DVDD.n82 DVDD.n44 0.0226963
R26406 DVDD.n206 DVDD.n185 0.0218816
R26407 DVDD.n233 DVDD.n172 0.0218816
R26408 DVDD.n66 DVDD.n45 0.0218816
R26409 DVDD.n93 DVDD.n32 0.0218816
R26410 DVDD.n190 DVDD.n188 0.021528
R26411 DVDD.n50 DVDD.n48 0.021528
R26412 DVDD.n168 DVDD.n128 0.0215056
R26413 DVDD.n133 DVDD.n128 0.0215056
R26414 DVDD.n320 DVDD.n319 0.0213889
R26415 DVDD.n319 DVDD.n18 0.0213889
R26416 DVDD.n299 DVDD.n298 0.0213889
R26417 DVDD.n298 DVDD.n24 0.0213889
R26418 DVDD.n290 DVDD.n24 0.0213889
R26419 DVDD.n288 DVDD.n96 0.0210464
R26420 DVDD.n282 DVDD.n96 0.0210464
R26421 DVDD.n281 DVDD.n100 0.0208243
R26422 DVDD.n273 DVDD.n100 0.0208243
R26423 DVDD.n273 DVDD.n272 0.0208243
R26424 DVDD.n210 DVDD.n185 0.0185921
R26425 DVDD.n233 DVDD.n173 0.0185921
R26426 DVDD.n70 DVDD.n45 0.0185921
R26427 DVDD.n93 DVDD.n33 0.0185921
R26428 DVDD.n226 DVDD.n183 0.0180234
R26429 DVDD.n176 DVDD 0.0180234
R26430 DVDD.n86 DVDD.n43 0.0180234
R26431 DVDD.n36 DVDD 0.0180234
R26432 DVDD.n200 DVDD.n193 0.016626
R26433 DVDD.n60 DVDD.n53 0.016626
R26434 DVDD.n208 DVDD.n207 0.0156869
R26435 DVDD.n232 DVDD.n174 0.0156869
R26436 DVDD.n68 DVDD.n67 0.0156869
R26437 DVDD.n92 DVDD.n34 0.0156869
R26438 DVDD.n218 DVDD.n214 0.0153479
R26439 DVDD.n78 DVDD.n74 0.0153479
R26440 DVDD.n211 DVDD.n210 0.0153026
R26441 DVDD.n175 DVDD.n173 0.0153026
R26442 DVDD.n71 DVDD.n70 0.0153026
R26443 DVDD.n35 DVDD.n33 0.0153026
R26444 DVDD.n203 DVDD.n202 0.0151028
R26445 DVDD.n63 DVDD.n62 0.0151028
R26446 DVDD.n209 DVDD.n208 0.0133505
R26447 DVDD.n232 DVDD 0.0133505
R26448 DVDD.n69 DVDD.n68 0.0133505
R26449 DVDD.n92 DVDD 0.0133505
R26450 DVDD.n206 DVDD.n205 0.0120132
R26451 DVDD.n216 DVDD.n172 0.0120132
R26452 DVDD.n66 DVDD.n65 0.0120132
R26453 DVDD.n76 DVDD.n32 0.0120132
R26454 DVDD.n209 DVDD.n183 0.011014
R26455 DVDD.n69 DVDD.n43 0.011014
R26456 DVDD.n315 DVDD 0.0105365
R26457 DVDD DVDD.n98 0.0105365
R26458 DVDD.n262 DVDD 0.0105365
R26459 DVDD.n163 DVDD 0.0105365
R26460 DVDD.n235 DVDD.n170 0.0103947
R26461 DVDD.n95 DVDD.n30 0.0103947
R26462 DVDD.n235 DVDD.n169 0.00951292
R26463 DVDD.n95 DVDD.n29 0.00951292
R26464 DVDD.n177 DVDD.n176 0.00926168
R26465 DVDD.n37 DVDD.n36 0.00926168
R26466 DVDD DVDD.n289 0.00885556
R26467 DVDD.n225 DVDD.n224 0.00872368
R26468 DVDD.n85 DVDD.n84 0.00872368
R26469 DVDD.n207 DVDD.n186 0.00867757
R26470 DVDD.n215 DVDD.n174 0.00867757
R26471 DVDD.n67 DVDD.n46 0.00867757
R26472 DVDD.n75 DVDD.n34 0.00867757
R26473 DVDD.n215 DVDD.n214 0.00750551
R26474 DVDD.n75 DVDD.n74 0.00750551
R26475 DVDD.n200 DVDD.n199 0.00692523
R26476 DVDD.n60 DVDD.n59 0.00692523
R26477 DVDD.n226 DVDD.n184 0.00634112
R26478 DVDD.n86 DVDD.n44 0.00634112
R26479 DVDD.n202 DVDD.n186 0.00575701
R26480 DVDD.n62 DVDD.n46 0.00575701
R26481 DVDD.n204 DVDD.n187 0.00543421
R26482 DVDD.n217 DVDD.n171 0.00543421
R26483 DVDD.n64 DVDD.n47 0.00543421
R26484 DVDD.n77 DVDD.n31 0.00543421
R26485 DVDD.n236 DVDD 0.00493889
R26486 DVDD.n287 DVDD.n286 0.00482522
R26487 DVDD.n266 DVDD.n118 0.00482522
R26488 DVDD.n167 DVDD.n129 0.00482522
R26489 DVDD.n318 DVDD.n317 0.00423134
R26490 DVDD.n285 DVDD.n97 0.00423134
R26491 DVDD.n265 DVDD.n264 0.00423134
R26492 DVDD.n166 DVDD.n165 0.00423134
R26493 DVDD.n203 DVDD.n188 0.00400467
R26494 DVDD.n219 DVDD.n218 0.00400467
R26495 DVDD.n63 DVDD.n48 0.00400467
R26496 DVDD.n79 DVDD.n78 0.00400467
R26497 DVDD.n196 DVDD.n190 0.00283645
R26498 DVDD.n56 DVDD.n50 0.00283645
R26499 DVDD.n235 DVDD.n234 0.00258889
R26500 DVDD.n95 DVDD.n94 0.00258889
R26501 DVDD DVDD.n177 0.00225234
R26502 DVDD DVDD.n37 0.00225234
R26503 DVDD.n198 DVDD.n197 0.00214474
R26504 DVDD.n223 DVDD.n212 0.00214474
R26505 DVDD.n58 DVDD.n57 0.00214474
R26506 DVDD.n83 DVDD.n72 0.00214474
R26507 DVDD.n222 DVDD.n221 0.00166822
R26508 DVDD.n82 DVDD.n81 0.00166822
R26509 DVDD.n301 DVDD.n300 0.00135292
R26510 DVDD.n291 DVDD.n28 0.00135292
R26511 DVDD.n280 DVDD.n113 0.00135292
R26512 DVDD.n271 DVDD.n270 0.00135292
R26513 DVDD.n248 DVDD.n247 0.00135292
R26514 DVDD.n238 DVDD.n127 0.00135292
R26515 DVDD.n149 DVDD.n148 0.00135292
R26516 DVDD.n139 DVDD.n138 0.00135292
R26517 DVDD.n314 DVDD.n21 0.00135241
R26518 DVDD.n283 DVDD.n99 0.00135241
R26519 DVDD.n261 DVDD.n119 0.00135241
R26520 DVDD.n162 DVDD.n130 0.00135241
R26521 DVDD.n266 DVDD.n265 0.00117863
R26522 DVDD.n167 DVDD.n166 0.00117863
R26523 DVDD.n287 DVDD.n97 0.00117863
R26524 DVDD.n318 DVDD.n19 0.00117863
R26525 DVDD.n199 DVDD.n189 0.00108411
R26526 DVDD.n196 DVDD.n189 0.00108411
R26527 DVDD.n221 DVDD.n220 0.00108411
R26528 DVDD.n59 DVDD.n49 0.00108411
R26529 DVDD.n56 DVDD.n49 0.00108411
R26530 DVDD.n81 DVDD.n80 0.00108411
R26531 DVDD.n145 DVDD.n144 0.00085506
R26532 DVDD.n142 DVDD.n141 0.00085506
R26533 DVDD.n188 DVDD.n187 0.00085506
R26534 DVDD.n208 DVDD.n185 0.00085506
R26535 DVDD.n219 DVDD.n171 0.00085506
R26536 DVDD.n233 DVDD.n232 0.00085506
R26537 DVDD.n244 DVDD.n124 0.00085506
R26538 DVDD.n241 DVDD.n125 0.00085506
R26539 DVDD.n274 DVDD.n115 0.00085506
R26540 DVDD.n277 DVDD.n114 0.00085506
R26541 DVDD.n48 DVDD.n47 0.00085506
R26542 DVDD.n68 DVDD.n45 0.00085506
R26543 DVDD.n79 DVDD.n31 0.00085506
R26544 DVDD.n93 DVDD.n92 0.00085506
R26545 DVDD.n294 DVDD.n293 0.00085506
R26546 DVDD.n297 DVDD.n296 0.00085506
R26547 DVDD.n148 DVDD.n147 0.000855023
R26548 DVDD.n146 DVDD.n145 0.000855023
R26549 DVDD.n141 DVDD.n134 0.000855023
R26550 DVDD.n166 DVDD.n128 0.000855023
R26551 DVDD.n133 DVDD.n130 0.000855023
R26552 DVDD.n192 DVDD.n187 0.000855023
R26553 DVDD.n191 DVDD.n185 0.000855023
R26554 DVDD.n224 DVDD.n170 0.000855023
R26555 DVDD.n234 DVDD.n171 0.000855023
R26556 DVDD.n234 DVDD.n233 0.000855023
R26557 DVDD.n247 DVDD.n246 0.000855023
R26558 DVDD.n245 DVDD.n244 0.000855023
R26559 DVDD.n125 DVDD.n123 0.000855023
R26560 DVDD.n238 DVDD.n237 0.000855023
R26561 DVDD.n265 DVDD.n117 0.000855023
R26562 DVDD.n122 DVDD.n119 0.000855023
R26563 DVDD.n274 DVDD.n273 0.000855023
R26564 DVDD.n114 DVDD.n100 0.000855023
R26565 DVDD.n281 DVDD.n280 0.000855023
R26566 DVDD.n272 DVDD.n271 0.000855023
R26567 DVDD.n97 DVDD.n96 0.000855023
R26568 DVDD.n283 DVDD.n282 0.000855023
R26569 DVDD.n52 DVDD.n47 0.000855023
R26570 DVDD.n51 DVDD.n45 0.000855023
R26571 DVDD.n84 DVDD.n30 0.000855023
R26572 DVDD.n94 DVDD.n31 0.000855023
R26573 DVDD.n94 DVDD.n93 0.000855023
R26574 DVDD.n293 DVDD.n24 0.000855023
R26575 DVDD.n298 DVDD.n297 0.000855023
R26576 DVDD.n300 DVDD.n299 0.000855023
R26577 DVDD.n319 DVDD.n318 0.000855023
R26578 DVDD.n21 DVDD.n18 0.000855023
R26579 DVDD.n291 DVDD.n290 0.000855023
R26580 DVDD.n224 DVDD.n184 0.000854948
R26581 DVDD.n84 DVDD.n44 0.000854948
R26582 DVDD.n264 DVDD.n118 0.000500614
R26583 DVDD.n165 DVDD.n129 0.000500614
R26584 DVDD.n317 DVDD.n316 0.000500614
R26585 DVDD.n286 DVDD.n285 0.000500614
R26586 DVDD.n243 DVDD.n242 0.000500461
R26587 DVDD.n143 DVDD.n135 0.000500461
R26588 DVDD.n295 DVDD.n25 0.000500461
R26589 DVDD.n276 DVDD.n275 0.000500461
R26590 a_5299_620.n27 a_5299_620.t9 129.037
R26591 a_5299_620.n27 a_5299_620.t8 68.9672
R26592 a_5299_620.n42 a_5299_620.n40 8.0439
R26593 a_5299_620.n3 a_5299_620.n20 7.45281
R26594 a_5299_620.n35 a_5299_620.n33 5.63
R26595 a_5299_620.n36 a_5299_620.t4 5.5395
R26596 a_5299_620.n36 a_5299_620.t5 5.5395
R26597 a_5299_620.n24 a_5299_620.t7 5.5395
R26598 a_5299_620.n24 a_5299_620.t6 5.5395
R26599 a_5299_620.n2 a_5299_620.n1 4.54542
R26600 a_5299_620.n6 a_5299_620.n39 4.5005
R26601 a_5299_620.n5 a_5299_620.n31 4.5005
R26602 a_5299_620.n0 a_5299_620.n42 4.5005
R26603 a_5299_620.n0 a_5299_620.n46 4.5005
R26604 a_5299_620.n4 a_5299_620.n23 4.5005
R26605 a_5299_620.n2 a_5299_620.n17 4.5005
R26606 a_5299_620.n2 a_5299_620.n12 4.5005
R26607 a_5299_620.n2 a_5299_620.n14 4.5005
R26608 a_5299_620.n47 a_5299_620.n0 4.3695
R26609 a_5299_620.n23 a_5299_620.n21 4.14168
R26610 a_5299_620.n7 a_5299_620.n26 3.82535
R26611 a_5299_620.n39 a_5299_620.n38 3.76521
R26612 a_5299_620.n46 a_5299_620.n45 3.76521
R26613 a_5299_620.n31 a_5299_620.n28 3.38874
R26614 a_5299_620.n42 a_5299_620.n41 3.38874
R26615 a_5299_620.n12 a_5299_620.n11 3.38238
R26616 a_5299_620.n44 a_5299_620.t3 3.3065
R26617 a_5299_620.n44 a_5299_620.t2 3.3065
R26618 a_5299_620.t1 a_5299_620.n50 3.3065
R26619 a_5299_620.n50 a_5299_620.t0 3.3065
R26620 a_5299_620.n31 a_5299_620.n30 3.01226
R26621 a_5299_620.n16 a_5299_620.n15 3.01226
R26622 a_5299_620.n39 a_5299_620.n37 2.63579
R26623 a_5299_620.n3 a_5299_620.n19 2.63579
R26624 a_5299_620.n7 a_5299_620.n27 2.423
R26625 a_5299_620.n18 a_5299_620.n48 2.2208
R26626 a_5299_620.n25 a_5299_620.n24 2.12431
R26627 a_5299_620.n47 a_5299_620.n6 3.11985
R26628 a_5299_620.n6 a_5299_620.n36 1.90815
R26629 a_5299_620.n12 a_5299_620.n10 1.88285
R26630 a_5299_620.n0 a_5299_620.n44 2.5496
R26631 a_5299_620.n23 a_5299_620.n22 1.50638
R26632 a_5299_620.n50 a_5299_620.n49 1.33804
R26633 a_5299_620.n14 a_5299_620.n13 1.12991
R26634 a_5299_620.n17 a_5299_620.n16 1.12991
R26635 a_5299_620.n26 a_5299_620.n4 0.922158
R26636 a_5299_620.n48 a_5299_620.n7 0.824928
R26637 a_5299_620.n10 a_5299_620.n9 0.753441
R26638 a_5299_620.n7 a_5299_620.n47 0.504252
R26639 a_5299_620.n1 a_5299_620.n8 0.376971
R26640 a_5299_620.n49 a_5299_620.n18 0.352626
R26641 a_5299_620.n32 a_5299_620.n35 0.278788
R26642 a_5299_620.n33 a_5299_620.n34 0.161367
R26643 a_5299_620.n28 a_5299_620.n29 0.150167
R26644 a_5299_620.n6 a_5299_620.n5 0.143833
R26645 a_5299_620.n5 a_5299_620.n32 0.1366
R26646 a_5299_620.n4 a_5299_620.n3 4.63501
R26647 a_5299_620.n0 a_5299_620.n43 1.11727
R26648 a_5299_620.n4 a_5299_620.n25 0.422157
R26649 a_5299_620.n18 a_5299_620.n2 0.221203
R26650 A1.n66 A1.n65 185
R26651 A1.n64 A1.n57 185
R26652 A1.n24 A1.n15 185
R26653 A1.n23 A1.n22 185
R26654 A1.n69 A1.t4 120.037
R26655 A1.t5 A1.n14 120.037
R26656 A1.n59 A1.n57 112.831
R26657 A1.n22 A1.n21 112.831
R26658 A1.n68 A1.n67 104.172
R26659 A1.n27 A1.n26 104.172
R26660 A1.n68 A1.n56 92.5005
R26661 A1.n28 A1.n27 92.5005
R26662 A1.t4 A1.n68 66.8281
R26663 A1.n27 A1.t5 66.8281
R26664 A1.n6 A1.t0 35.2053
R26665 A1.n3 A1.t1 34.0571
R26666 A1.n67 A1.n66 29.4833
R26667 A1.n26 A1.n15 29.4833
R26668 A1.n1 A1.t6 27.6955
R26669 A1.n1 A1.t7 27.6955
R26670 A1.n45 A1.n44 19.0955
R26671 A1.n69 A1.n56 15.4558
R26672 A1.n28 A1.n14 15.4558
R26673 A1.n64 A1.n63 13.5534
R26674 A1.n23 A1.n18 13.5534
R26675 A1.n2 A1.n1 9.67857
R26676 A1.n41 A1.n34 9.30581
R26677 A1.n59 A1.n58 9.30424
R26678 A1.n21 A1.n20 9.30413
R26679 A1.n40 A1.n39 9.3005
R26680 A1.n46 A1.n45 9.3005
R26681 A1.n71 A1.n70 9.3005
R26682 A1.n55 A1.n52 9.3005
R26683 A1.n67 A1.n55 9.3005
R26684 A1.n63 A1.n62 9.3005
R26685 A1.n72 A1.n54 9.3005
R26686 A1.n29 A1.n13 9.3005
R26687 A1.n25 A1.n11 9.3005
R26688 A1.n26 A1.n25 9.3005
R26689 A1.n18 A1.n17 9.3005
R26690 A1.n31 A1.n30 9.3005
R26691 A1.n71 A1.n56 9.03579
R26692 A1.n29 A1.n28 9.03579
R26693 A1.n43 A1.n41 8.49366
R26694 A1.n43 A1.t2 8.2655
R26695 A1.n43 A1.t3 8.2655
R26696 A1.n44 A1.n43 7.97749
R26697 A1.n42 A1.n40 7.26743
R26698 A1.n43 A1.n42 6.15568
R26699 A1.n65 A1.n55 5.64756
R26700 A1.n25 A1.n24 5.64756
R26701 A1.n41 A1.n35 4.89462
R26702 A1.n60 A1.n59 4.89462
R26703 A1.n21 A1.n19 4.89462
R26704 A1.n73 A1.n55 4.51815
R26705 A1.n72 A1.n71 4.51815
R26706 A1.n25 A1.n12 4.51815
R26707 A1.n30 A1.n29 4.51815
R26708 A1.n5 A1.n4 4.5005
R26709 A1.n4 A1.n2 4.5005
R26710 A1.n51 A1.n9 4.5005
R26711 A1.n49 A1.n9 4.5005
R26712 A1.n51 A1.n50 4.5005
R26713 A1.n50 A1.n49 4.5005
R26714 A1.n74 A1.n53 4.5005
R26715 A1.n75 A1.n8 4.5005
R26716 A1.n53 A1.n8 4.5005
R26717 A1.n75 A1.n74 4.5005
R26718 A1.n48 A1.n32 4.5005
R26719 A1.n47 A1.n36 4.5005
R26720 A1.n48 A1.n47 4.5005
R26721 A1.n36 A1.n32 4.5005
R26722 A1.n38 A1.n33 4.5005
R26723 A1.n66 A1.n57 3.93153
R26724 A1.n22 A1.n15 3.93153
R26725 A1.n19 A1.n9 3.03311
R26726 A1.n50 A1.n12 3.03311
R26727 A1.n60 A1.n8 3.03311
R26728 A1.n74 A1.n73 3.03311
R26729 A1.n47 A1.n35 3.03311
R26730 A1.n3 A1.n0 2.2714
R26731 A1.n58 A1.n7 2.25261
R26732 A1.n20 A1.n10 2.25256
R26733 A1.n34 A1.n33 2.25127
R26734 A1.n37 A1.n33 2.24434
R26735 A1.n73 A1.n72 1.88285
R26736 A1.n30 A1.n12 1.88285
R26737 A1.n45 A1.n35 1.50638
R26738 A1.n63 A1.n60 1.50638
R26739 A1.n19 A1.n18 1.50638
R26740 A1.n16 A1.n10 1.49213
R26741 A1.n70 A1.n69 1.49212
R26742 A1.n61 A1.n7 1.49182
R26743 A1.n14 A1.n13 1.49166
R26744 A1.n65 A1.n64 0.753441
R26745 A1.n24 A1.n23 0.753441
R26746 A1.n44 A1.n40 0.521921
R26747 A1.n77 A1.n6 0.29767
R26748 A1.n49 A1.n48 0.238951
R26749 A1.n77 A1.n76 0.196255
R26750 A1 A1.n77 0.1855
R26751 A1.n6 A1.n5 0.149538
R26752 A1.n75 A1.n51 0.124821
R26753 A1.n42 A1.n32 0.0579027
R26754 A1.n78 A1 0.0523868
R26755 A1.n62 A1.n61 0.0396286
R26756 A1.n17 A1.n16 0.0383668
R26757 A1.n46 A1.n37 0.0314092
R26758 A1.n5 A1.n0 0.0281442
R26759 A1.n39 A1.n37 0.0271357
R26760 A1.n61 A1.n52 0.0202788
R26761 A1.n16 A1.n11 0.0196501
R26762 A1.n51 A1.n10 0.0168043
R26763 A1.n36 A1.n33 0.016125
R26764 A1 A1.n78 0.0137212
R26765 A1.n78 A1 0.0134717
R26766 A1.n74 A1.n52 0.013431
R26767 A1.n70 A1.n54 0.013431
R26768 A1.n50 A1.n11 0.013
R26769 A1.n31 A1.n13 0.013
R26770 A1.n38 A1.n32 0.0122521
R26771 A1.n58 A1.n8 0.0117689
R26772 A1.n20 A1.n9 0.0114102
R26773 A1.n47 A1.n34 0.0100704
R26774 A1.n76 A1.n7 0.0100109
R26775 A1.n74 A1.n54 0.00588793
R26776 A1.n50 A1.n31 0.00570833
R26777 A1.n62 A1.n8 0.00481034
R26778 A1.n47 A1.n46 0.0047735
R26779 A1.n17 A1.n9 0.00466667
R26780 A1.n53 A1.n7 0.00457609
R26781 A1.n76 A1.n75 0.00457609
R26782 A1.n2 A1.n0 0.00410577
R26783 A1.n39 A1.n38 0.00370513
R26784 A1.n48 A1.n33 0.00253804
R26785 A1.n4 A1.n3 0.00185919
R26786 A1.n49 A1.n10 0.0018587
R26787 a_5299_1782.n21 a_5299_1782.t8 60.2505
R26788 a_5299_1782.n42 a_5299_1782.t9 60.2505
R26789 a_5299_1782.n64 a_5299_1782.t0 60.2505
R26790 a_5299_1782.n76 a_5299_1782.t2 60.2505
R26791 a_5299_1782.n2 a_5299_1782.n84 9.3005
R26792 a_5299_1782.n2 a_5299_1782.n85 9.3005
R26793 a_5299_1782.n2 a_5299_1782.n83 9.3005
R26794 a_5299_1782.n83 a_5299_1782.n82 9.3005
R26795 a_5299_1782.n3 a_5299_1782.n73 9.3005
R26796 a_5299_1782.n4 a_5299_1782.n57 9.3005
R26797 a_5299_1782.n4 a_5299_1782.n56 9.3005
R26798 a_5299_1782.n4 a_5299_1782.n63 9.3005
R26799 a_5299_1782.n63 a_5299_1782.n62 9.3005
R26800 a_5299_1782.n3 a_5299_1782.n72 9.3005
R26801 a_5299_1782.n72 a_5299_1782.n71 9.3005
R26802 a_5299_1782.n3 a_5299_1782.n74 9.3005
R26803 a_5299_1782.n5 a_5299_1782.n51 9.3005
R26804 a_5299_1782.n6 a_5299_1782.n35 9.3005
R26805 a_5299_1782.n6 a_5299_1782.n34 9.3005
R26806 a_5299_1782.n6 a_5299_1782.n41 9.3005
R26807 a_5299_1782.n41 a_5299_1782.n40 9.3005
R26808 a_5299_1782.n5 a_5299_1782.n50 9.3005
R26809 a_5299_1782.n50 a_5299_1782.n49 9.3005
R26810 a_5299_1782.n5 a_5299_1782.n52 9.3005
R26811 a_5299_1782.n7 a_5299_1782.n29 9.3005
R26812 a_5299_1782.n7 a_5299_1782.n28 9.3005
R26813 a_5299_1782.n28 a_5299_1782.n27 9.3005
R26814 a_5299_1782.n7 a_5299_1782.n30 9.3005
R26815 a_5299_1782.n1 a_5299_1782.n91 9.3005
R26816 a_5299_1782.n119 a_5299_1782.n118 10.743
R26817 a_5299_1782.n65 a_5299_1782.n64 8.76429
R26818 a_5299_1782.n43 a_5299_1782.n42 8.76429
R26819 a_5299_1782.n26 a_5299_1782.n25 7.45411
R26820 a_5299_1782.n39 a_5299_1782.n38 7.45411
R26821 a_5299_1782.n48 a_5299_1782.n47 7.45411
R26822 a_5299_1782.n61 a_5299_1782.n60 7.45411
R26823 a_5299_1782.n70 a_5299_1782.n69 7.45411
R26824 a_5299_1782.n81 a_5299_1782.n80 7.45411
R26825 a_5299_1782.n22 a_5299_1782.n21 6.80105
R26826 a_5299_1782.n77 a_5299_1782.n76 6.80105
R26827 a_5299_1782.n24 a_5299_1782.n23 5.64756
R26828 a_5299_1782.n37 a_5299_1782.n36 5.64756
R26829 a_5299_1782.n46 a_5299_1782.n45 5.64756
R26830 a_5299_1782.n59 a_5299_1782.n58 5.64756
R26831 a_5299_1782.n68 a_5299_1782.n67 5.64756
R26832 a_5299_1782.n79 a_5299_1782.n78 5.64756
R26833 a_5299_1782.n96 a_5299_1782.t1 5.5395
R26834 a_5299_1782.n96 a_5299_1782.t3 5.5395
R26835 a_5299_1782.n90 a_5299_1782.n89 4.95584
R26836 a_5299_1782.n31 a_5299_1782.n20 4.73575
R26837 a_5299_1782.n33 a_5299_1782.n32 4.73575
R26838 a_5299_1782.n53 a_5299_1782.n19 4.73575
R26839 a_5299_1782.n55 a_5299_1782.n54 4.73575
R26840 a_5299_1782.n75 a_5299_1782.n18 4.73575
R26841 a_5299_1782.n87 a_5299_1782.n86 4.73575
R26842 a_5299_1782.n11 a_5299_1782.n13 4.66695
R26843 a_5299_1782.n66 a_5299_1782.n65 4.6505
R26844 a_5299_1782.n44 a_5299_1782.n43 4.6505
R26845 a_5299_1782.n1 a_5299_1782.n17 4.5005
R26846 a_5299_1782.n13 a_5299_1782.n99 4.5005
R26847 a_5299_1782.n12 a_5299_1782.n95 4.5005
R26848 a_5299_1782.n0 a_5299_1782.n110 4.5005
R26849 a_5299_1782.n0 a_5299_1782.n105 4.5005
R26850 a_5299_1782.n10 a_5299_1782.n117 4.5005
R26851 a_5299_1782.n9 a_5299_1782.n114 4.5005
R26852 a_5299_1782.n9 a_5299_1782.n112 4.5005
R26853 a_5299_1782.n110 a_5299_1782.n109 4.14168
R26854 a_5299_1782.n99 a_5299_1782.n98 3.76521
R26855 a_5299_1782.n114 a_5299_1782.n113 3.76521
R26856 a_5299_1782.n7 a_5299_1782.n22 3.42768
R26857 a_5299_1782.n2 a_5299_1782.n77 3.42768
R26858 a_5299_1782.n95 a_5299_1782.n93 3.38874
R26859 a_5299_1782.n17 a_5299_1782.n16 3.38874
R26860 a_5299_1782.n106 a_5299_1782.t5 3.3065
R26861 a_5299_1782.n106 a_5299_1782.t4 3.3065
R26862 a_5299_1782.n119 a_5299_1782.t6 3.3065
R26863 a_5299_1782.t7 a_5299_1782.n119 3.3065
R26864 a_5299_1782.n95 a_5299_1782.n94 3.01226
R26865 a_5299_1782.n17 a_5299_1782.n15 3.01226
R26866 a_5299_1782.n119 a_5299_1782.n100 2.66355
R26867 a_5299_1782.n99 a_5299_1782.n97 2.63579
R26868 a_5299_1782.n104 a_5299_1782.n103 2.25932
R26869 a_5299_1782.n116 a_5299_1782.n115 2.25932
R26870 a_5299_1782.n9 a_5299_1782.n11 1.68471
R26871 a_5299_1782.n107 a_5299_1782.n106 1.46875
R26872 a_5299_1782.n27 a_5299_1782.n26 0.994314
R26873 a_5299_1782.n40 a_5299_1782.n39 0.994314
R26874 a_5299_1782.n49 a_5299_1782.n48 0.994314
R26875 a_5299_1782.n62 a_5299_1782.n61 0.994314
R26876 a_5299_1782.n71 a_5299_1782.n70 0.994314
R26877 a_5299_1782.n82 a_5299_1782.n81 0.994314
R26878 a_5299_1782.n28 a_5299_1782.n24 0.753441
R26879 a_5299_1782.n41 a_5299_1782.n37 0.753441
R26880 a_5299_1782.n50 a_5299_1782.n46 0.753441
R26881 a_5299_1782.n63 a_5299_1782.n59 0.753441
R26882 a_5299_1782.n72 a_5299_1782.n68 0.753441
R26883 a_5299_1782.n83 a_5299_1782.n79 0.753441
R26884 a_5299_1782.n102 a_5299_1782.n101 0.603501
R26885 a_5299_1782.n119 a_5299_1782.n10 2.11613
R26886 a_5299_1782.n8 a_5299_1782.n107 0.555049
R26887 a_5299_1782.n33 a_5299_1782.n31 0.458354
R26888 a_5299_1782.n55 a_5299_1782.n53 0.458354
R26889 a_5299_1782.n13 a_5299_1782.n96 1.90913
R26890 a_5299_1782.n11 a_5299_1782.n102 0.710352
R26891 a_5299_1782.n110 a_5299_1782.n108 0.376971
R26892 a_5299_1782.n105 a_5299_1782.n104 0.376971
R26893 a_5299_1782.n112 a_5299_1782.n111 0.376971
R26894 a_5299_1782.n117 a_5299_1782.n116 0.376971
R26895 a_5299_1782.n88 a_5299_1782.n75 0.229427
R26896 a_5299_1782.n88 a_5299_1782.n87 0.229427
R26897 a_5299_1782.n90 a_5299_1782.n88 0.215848
R26898 a_5299_1782.n31 a_5299_1782.n7 0.205546
R26899 a_5299_1782.n6 a_5299_1782.n33 0.205546
R26900 a_5299_1782.n53 a_5299_1782.n5 0.205546
R26901 a_5299_1782.n4 a_5299_1782.n55 0.205546
R26902 a_5299_1782.n75 a_5299_1782.n3 0.205546
R26903 a_5299_1782.n87 a_5299_1782.n2 0.205546
R26904 a_5299_1782.n44 a_5299_1782.n6 0.190717
R26905 a_5299_1782.n5 a_5299_1782.n44 0.190717
R26906 a_5299_1782.n66 a_5299_1782.n4 0.190717
R26907 a_5299_1782.n3 a_5299_1782.n66 0.190717
R26908 a_5299_1782.n0 a_5299_1782.n8 0.183965
R26909 a_5299_1782.n12 a_5299_1782.n1 0.169804
R26910 a_5299_1782.n15 a_5299_1782.n14 0.161367
R26911 a_5299_1782.n93 a_5299_1782.n92 0.150167
R26912 a_5299_1782.n1 a_5299_1782.n90 0.140745
R26913 a_5299_1782.n13 a_5299_1782.n12 0.14187
R26914 a_5299_1782.n10 a_5299_1782.n9 0.135427
R26915 a_5299_1782.n102 a_5299_1782.n0 0.107619
R26916 B2.n66 B2.n65 185
R26917 B2.n64 B2.n57 185
R26918 B2.n24 B2.n15 185
R26919 B2.n23 B2.n22 185
R26920 B2.n69 B2.t4 120.037
R26921 B2.t5 B2.n14 120.037
R26922 B2.n59 B2.n57 112.831
R26923 B2.n22 B2.n21 112.831
R26924 B2.n68 B2.n67 104.172
R26925 B2.n27 B2.n26 104.172
R26926 B2.n68 B2.n56 92.5005
R26927 B2.n28 B2.n27 92.5005
R26928 B2.t4 B2.n68 66.8281
R26929 B2.n27 B2.t5 66.8281
R26930 B2.n6 B2.t0 35.2053
R26931 B2.n3 B2.t1 34.0571
R26932 B2.n67 B2.n66 29.4833
R26933 B2.n26 B2.n15 29.4833
R26934 B2.n1 B2.t7 27.6955
R26935 B2.n1 B2.t6 27.6955
R26936 B2.n45 B2.n44 19.0955
R26937 B2.n69 B2.n56 15.4558
R26938 B2.n28 B2.n14 15.4558
R26939 B2.n64 B2.n63 13.5534
R26940 B2.n23 B2.n18 13.5534
R26941 B2.n2 B2.n1 9.67857
R26942 B2.n41 B2.n34 9.30581
R26943 B2.n59 B2.n58 9.30424
R26944 B2.n21 B2.n20 9.30413
R26945 B2.n40 B2.n39 9.3005
R26946 B2.n46 B2.n45 9.3005
R26947 B2.n71 B2.n70 9.3005
R26948 B2.n55 B2.n52 9.3005
R26949 B2.n67 B2.n55 9.3005
R26950 B2.n63 B2.n62 9.3005
R26951 B2.n72 B2.n54 9.3005
R26952 B2.n29 B2.n13 9.3005
R26953 B2.n25 B2.n11 9.3005
R26954 B2.n26 B2.n25 9.3005
R26955 B2.n18 B2.n17 9.3005
R26956 B2.n31 B2.n30 9.3005
R26957 B2.n71 B2.n56 9.03579
R26958 B2.n29 B2.n28 9.03579
R26959 B2.n43 B2.n41 8.49366
R26960 B2.n43 B2.t3 8.2655
R26961 B2.n43 B2.t2 8.2655
R26962 B2.n44 B2.n43 7.97749
R26963 B2.n42 B2.n40 7.26743
R26964 B2.n43 B2.n42 6.15568
R26965 B2.n65 B2.n55 5.64756
R26966 B2.n25 B2.n24 5.64756
R26967 B2.n41 B2.n35 4.89462
R26968 B2.n60 B2.n59 4.89462
R26969 B2.n21 B2.n19 4.89462
R26970 B2.n73 B2.n55 4.51815
R26971 B2.n72 B2.n71 4.51815
R26972 B2.n25 B2.n12 4.51815
R26973 B2.n30 B2.n29 4.51815
R26974 B2.n5 B2.n4 4.5005
R26975 B2.n4 B2.n2 4.5005
R26976 B2.n51 B2.n9 4.5005
R26977 B2.n49 B2.n9 4.5005
R26978 B2.n51 B2.n50 4.5005
R26979 B2.n50 B2.n49 4.5005
R26980 B2.n74 B2.n53 4.5005
R26981 B2.n75 B2.n8 4.5005
R26982 B2.n53 B2.n8 4.5005
R26983 B2.n75 B2.n74 4.5005
R26984 B2.n48 B2.n32 4.5005
R26985 B2.n47 B2.n36 4.5005
R26986 B2.n48 B2.n47 4.5005
R26987 B2.n36 B2.n32 4.5005
R26988 B2.n38 B2.n33 4.5005
R26989 B2.n66 B2.n57 3.93153
R26990 B2.n22 B2.n15 3.93153
R26991 B2.n19 B2.n9 3.03311
R26992 B2.n50 B2.n12 3.03311
R26993 B2.n60 B2.n8 3.03311
R26994 B2.n74 B2.n73 3.03311
R26995 B2.n47 B2.n35 3.03311
R26996 B2.n3 B2.n0 2.2714
R26997 B2.n58 B2.n7 2.25261
R26998 B2.n20 B2.n10 2.25256
R26999 B2.n34 B2.n33 2.25127
R27000 B2.n37 B2.n33 2.24434
R27001 B2.n73 B2.n72 1.88285
R27002 B2.n30 B2.n12 1.88285
R27003 B2.n45 B2.n35 1.50638
R27004 B2.n63 B2.n60 1.50638
R27005 B2.n19 B2.n18 1.50638
R27006 B2.n16 B2.n10 1.49213
R27007 B2.n70 B2.n69 1.49212
R27008 B2.n61 B2.n7 1.49182
R27009 B2.n14 B2.n13 1.49166
R27010 B2.n65 B2.n64 0.753441
R27011 B2.n24 B2.n23 0.753441
R27012 B2.n44 B2.n40 0.521921
R27013 B2.n77 B2.n6 0.29767
R27014 B2.n49 B2.n48 0.238951
R27015 B2.n77 B2.n76 0.196255
R27016 B2 B2.n77 0.1855
R27017 B2.n6 B2.n5 0.149538
R27018 B2.n75 B2.n51 0.124821
R27019 B2.n42 B2.n32 0.0579027
R27020 B2.n62 B2.n61 0.0396286
R27021 B2.n17 B2.n16 0.0383668
R27022 B2.n46 B2.n37 0.0314092
R27023 B2.n5 B2.n0 0.0281442
R27024 B2.n39 B2.n37 0.0271357
R27025 B2.n61 B2.n52 0.0202788
R27026 B2.n16 B2.n11 0.0196501
R27027 B2.n51 B2.n10 0.0168043
R27028 B2.n36 B2.n33 0.016125
R27029 B2.n74 B2.n52 0.013431
R27030 B2.n70 B2.n54 0.013431
R27031 B2.n50 B2.n11 0.013
R27032 B2.n31 B2.n13 0.013
R27033 B2.n38 B2.n32 0.0122521
R27034 B2.n58 B2.n8 0.0117689
R27035 B2.n20 B2.n9 0.0114102
R27036 B2.n47 B2.n34 0.0100704
R27037 B2.n76 B2.n7 0.0100109
R27038 B2.n74 B2.n54 0.00588793
R27039 B2.n50 B2.n31 0.00570833
R27040 B2.n62 B2.n8 0.00481034
R27041 B2.n47 B2.n46 0.0047735
R27042 B2.n17 B2.n9 0.00466667
R27043 B2.n53 B2.n7 0.00457609
R27044 B2.n76 B2.n75 0.00457609
R27045 B2.n2 B2.n0 0.00410577
R27046 B2.n39 B2.n38 0.00370513
R27047 B2.n48 B2.n33 0.00253804
R27048 B2.n4 B2.n3 0.00185919
R27049 B2.n49 B2.n10 0.0018587
R27050 SELB.n6 SELB.t4 186.374
R27051 SELB.n6 SELB.t5 170.308
R27052 SELB.n7 SELB.n6 139.876
R27053 SELB.n0 SELB.t1 84.8325
R27054 SELB.n1 SELB.t0 84.8325
R27055 SELB.n1 SELB.n0 60.1541
R27056 SELB.n2 SELB.n1 50.1642
R27057 SELB.n0 SELB.t3 48.6825
R27058 SELB.n1 SELB.t2 48.6825
R27059 SELB.n5 SELB 42.9181
R27060 SELB.n4 SELB 17.169
R27061 SELB.n3 SELB.n2 15.2731
R27062 SELB.n11 SELB.n9 14.3125
R27063 SELB.n5 SELB 12.8005
R27064 SELB.n4 SELB.n3 4.77356
R27065 SELB.n8 SELB 2.73914
R27066 SELB SELB.n3 2.13383
R27067 SELB SELB.n7 1.61978
R27068 SELB.n9 SELB.n8 1.31185
R27069 SELB SELB.n13 1.25831
R27070 SELB.n2 SELB 1.1768
R27071 SELB.n7 SELB.n5 0.925801
R27072 SELB.n13 SELB.n12 0.675199
R27073 SELB.n10 SELB 0.34425
R27074 SELB.n13 SELB 0.321549
R27075 SELB SELB.n11 0.0255
R27076 SELB.n11 SELB.n10 0.0194024
R27077 SELB SELB.n4 0.0180439
R27078 SELB.n12 SELB 0.0151341
R27079 SELB.n8 SELB 0.00770734
R27080 SELB.n12 SELB 0.00415854
R27081 SELB.n10 SELB 0.00171951
R27082 SELB.n12 SELB.n9 0.000502048
R27083 A2.n66 A2.n65 185
R27084 A2.n64 A2.n57 185
R27085 A2.n24 A2.n15 185
R27086 A2.n23 A2.n22 185
R27087 A2.n69 A2.t0 120.037
R27088 A2.t1 A2.n14 120.037
R27089 A2.n59 A2.n57 112.831
R27090 A2.n22 A2.n21 112.831
R27091 A2.n68 A2.n67 104.172
R27092 A2.n27 A2.n26 104.172
R27093 A2.n68 A2.n56 92.5005
R27094 A2.n28 A2.n27 92.5005
R27095 A2.t0 A2.n68 66.8281
R27096 A2.n27 A2.t1 66.8281
R27097 A2.n6 A2.t4 35.2053
R27098 A2.n3 A2.t5 34.0571
R27099 A2.n67 A2.n66 29.4833
R27100 A2.n26 A2.n15 29.4833
R27101 A2.n1 A2.t2 27.6955
R27102 A2.n1 A2.t3 27.6955
R27103 A2.n45 A2.n44 19.0955
R27104 A2.n69 A2.n56 15.4558
R27105 A2.n28 A2.n14 15.4558
R27106 A2.n64 A2.n63 13.5534
R27107 A2.n23 A2.n18 13.5534
R27108 A2.n2 A2.n1 9.67857
R27109 A2.n41 A2.n34 9.30581
R27110 A2.n59 A2.n58 9.30424
R27111 A2.n21 A2.n20 9.30413
R27112 A2.n40 A2.n39 9.3005
R27113 A2.n46 A2.n45 9.3005
R27114 A2.n71 A2.n70 9.3005
R27115 A2.n55 A2.n52 9.3005
R27116 A2.n67 A2.n55 9.3005
R27117 A2.n63 A2.n62 9.3005
R27118 A2.n72 A2.n54 9.3005
R27119 A2.n29 A2.n13 9.3005
R27120 A2.n25 A2.n11 9.3005
R27121 A2.n26 A2.n25 9.3005
R27122 A2.n18 A2.n17 9.3005
R27123 A2.n31 A2.n30 9.3005
R27124 A2.n71 A2.n56 9.03579
R27125 A2.n29 A2.n28 9.03579
R27126 A2.n43 A2.n41 8.49366
R27127 A2.n43 A2.t6 8.2655
R27128 A2.n43 A2.t7 8.2655
R27129 A2.n44 A2.n43 7.97749
R27130 A2.n42 A2.n40 7.26743
R27131 A2.n43 A2.n42 6.15568
R27132 A2.n65 A2.n55 5.64756
R27133 A2.n25 A2.n24 5.64756
R27134 A2.n41 A2.n35 4.89462
R27135 A2.n60 A2.n59 4.89462
R27136 A2.n21 A2.n19 4.89462
R27137 A2.n73 A2.n55 4.51815
R27138 A2.n72 A2.n71 4.51815
R27139 A2.n25 A2.n12 4.51815
R27140 A2.n30 A2.n29 4.51815
R27141 A2.n5 A2.n4 4.5005
R27142 A2.n4 A2.n2 4.5005
R27143 A2.n51 A2.n9 4.5005
R27144 A2.n49 A2.n9 4.5005
R27145 A2.n51 A2.n50 4.5005
R27146 A2.n50 A2.n49 4.5005
R27147 A2.n74 A2.n53 4.5005
R27148 A2.n75 A2.n8 4.5005
R27149 A2.n53 A2.n8 4.5005
R27150 A2.n75 A2.n74 4.5005
R27151 A2.n48 A2.n32 4.5005
R27152 A2.n47 A2.n36 4.5005
R27153 A2.n48 A2.n47 4.5005
R27154 A2.n36 A2.n32 4.5005
R27155 A2.n38 A2.n33 4.5005
R27156 A2.n66 A2.n57 3.93153
R27157 A2.n22 A2.n15 3.93153
R27158 A2.n19 A2.n9 3.03311
R27159 A2.n50 A2.n12 3.03311
R27160 A2.n60 A2.n8 3.03311
R27161 A2.n74 A2.n73 3.03311
R27162 A2.n47 A2.n35 3.03311
R27163 A2.n3 A2.n0 2.2714
R27164 A2.n58 A2.n7 2.25261
R27165 A2.n20 A2.n10 2.25256
R27166 A2.n34 A2.n33 2.25127
R27167 A2.n37 A2.n33 2.24434
R27168 A2.n73 A2.n72 1.88285
R27169 A2.n30 A2.n12 1.88285
R27170 A2.n45 A2.n35 1.50638
R27171 A2.n63 A2.n60 1.50638
R27172 A2.n19 A2.n18 1.50638
R27173 A2.n16 A2.n10 1.49213
R27174 A2.n70 A2.n69 1.49212
R27175 A2.n61 A2.n7 1.49182
R27176 A2.n14 A2.n13 1.49166
R27177 A2.n65 A2.n64 0.753441
R27178 A2.n24 A2.n23 0.753441
R27179 A2.n44 A2.n40 0.521921
R27180 A2.n77 A2.n6 0.29767
R27181 A2.n49 A2.n48 0.238951
R27182 A2.n77 A2.n76 0.196255
R27183 A2 A2.n77 0.1855
R27184 A2.n6 A2.n5 0.149538
R27185 A2.n78 A2 0.13698
R27186 A2.n75 A2.n51 0.124821
R27187 A2.n42 A2.n32 0.0579027
R27188 A2 A2.n78 0.0486771
R27189 A2.n78 A2 0.0476939
R27190 A2.n62 A2.n61 0.0396286
R27191 A2.n17 A2.n16 0.0383668
R27192 A2.n46 A2.n37 0.0314092
R27193 A2.n5 A2.n0 0.0281442
R27194 A2.n39 A2.n37 0.0271357
R27195 A2.n61 A2.n52 0.0202788
R27196 A2.n16 A2.n11 0.0196501
R27197 A2.n51 A2.n10 0.0168043
R27198 A2.n36 A2.n33 0.016125
R27199 A2.n74 A2.n52 0.013431
R27200 A2.n70 A2.n54 0.013431
R27201 A2.n50 A2.n11 0.013
R27202 A2.n31 A2.n13 0.013
R27203 A2.n38 A2.n32 0.0122521
R27204 A2.n58 A2.n8 0.0117689
R27205 A2.n20 A2.n9 0.0114102
R27206 A2.n47 A2.n34 0.0100704
R27207 A2.n76 A2.n7 0.0100109
R27208 A2.n74 A2.n54 0.00588793
R27209 A2.n50 A2.n31 0.00570833
R27210 A2.n62 A2.n8 0.00481034
R27211 A2.n47 A2.n46 0.0047735
R27212 A2.n17 A2.n9 0.00466667
R27213 A2.n53 A2.n7 0.00457609
R27214 A2.n76 A2.n75 0.00457609
R27215 A2.n2 A2.n0 0.00410577
R27216 A2.n39 A2.n38 0.00370513
R27217 A2.n48 A2.n33 0.00253804
R27218 A2.n4 A2.n3 0.00185919
R27219 A2.n49 A2.n10 0.0018587
C0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_7464_n6798# 7.03e-19
C1 a_11235_n6821# DVDD 0.19f
C2 a_6351_6657# VSS 0.0236f
C3 DVDD VO 0.466f
C4 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.34f
C5 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 5.32e-19
C6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_1.invm_0.Y 8.17e-19
C7 a_8403_n6064# DVDD 0.0139f
C8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 A2 0.518f
C9 a_11235_n6821# a_10810_n6777# 0.461f
C10 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 a_11235_n6821# 3.13e-19
C11 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.124f
C12 a_7196_n5728# a_7889_n6842# 0.265f
C13 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.00181f
C14 a_3916_n5703# a_5123_n6039# 0.289f
C15 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 5.32e-19
C16 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 2.72e-19
C17 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 0.0365f
C18 a_1263_n6838# SELA 0.00469f
C19 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.683f
C20 a_1263_n6838# VDD 0.607f
C21 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.00152f
C22 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 0.839f
C23 comparator_top_0.comparator_0.VBN comparator_top_0.VINM 0.494f
C24 a_3916_n5703# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.0154f
C25 a_10975_4108# VO 0.169f
C26 EF_AMUX21m_2.invm_0.Y DVDD 0.958f
C27 a_10542_n5707# DVDD 0.116f
C28 DVDD A1 0.00246f
C29 a_4609_n6817# VDD 0.607f
C30 EF_AMUX21m_2.invm_0.Y a_10810_n6777# 0.0217f
C31 a_7889_n6842# a_7464_n6798# 0.461f
C32 a_470_n5812# VSS 0.00701f
C33 a_10542_n5707# a_10810_n6777# 0.0272f
C34 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.07f
C35 DVDD B1 0.00248f
C36 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 a_10542_n5707# 6.2e-19
C37 a_3916_n5703# a_4184_n6773# 0.0272f
C38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X B2 8.92e-19
C39 DVDD SELA 0.92f
C40 a_570_n5724# A1 4.37e-19
C41 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_7096_n5816# 0.00188f
C42 VDD DVDD 11.6f
C43 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD 3.43f
C44 comparator_top_0.comparator_0.VOUT VO 0.0406f
C45 a_838_n6794# SELA 0.0224f
C46 a_11749_n6043# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.145f
C47 a_10810_n6777# VDD 0.154f
C48 a_838_n6794# VDD 0.154f
C49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 VDD 2.05f
C50 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X SELB 5.01e-19
C51 a_570_n5724# SELA 0.00244f
C52 a_10965_3602# VO 0.0178f
C53 a_570_n5724# VDD 1.12f
C54 comparator_top_0.comparator_0.VBP VSS 2.22f
C55 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 SELB 1.27e-19
C56 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_7096_n5816# 5.3e-19
C57 a_1263_n6838# DVDD 0.189f
C58 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_10542_n5707# 4.56e-19
C59 comparator_top_0.comparator_0.VBN VDD 9.88f
C60 a_1263_n6838# a_838_n6794# 0.461f
C61 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp B1 1.5e-19
C62 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_4184_n6773# 4.53e-21
C63 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VSS 3.09e-19
C64 a_10975_4108# VDD 0.248f
C65 a_7196_n5728# SELB 0.00244f
C66 a_570_n5724# a_1263_n6838# 0.265f
C67 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_8403_n6064# 0.00108f
C68 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp VDD 2.65f
C69 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.34f
C70 EF_AMUX21m_1.invm_0.Y SELA 0.241f
C71 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.08f
C72 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb B2 1.01f
C73 a_7096_n5816# a_7196_n5728# 0.405f
C74 a_4609_n6817# DVDD 0.186f
C75 EF_AMUX21m_1.invm_0.Y VDD 0.0233f
C76 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_4609_n6817# 7.05e-21
C77 comparator_top_0.VINP A2 2.81f
C78 comparator_top_0.VINP VSS 4.62f
C79 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.07f
C80 a_3816_n5791# VDD 0.335f
C81 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 A2 1.85e-19
C82 a_3916_n5703# A2 4.37e-19
C83 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 VSS 9.51e-19
C84 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00684f
C85 comparator_top_0.comparator_0.VOUT VDD 2.93f
C86 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 1.54e-19
C87 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 a_8403_n6064# 0.00121f
C88 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_3916_n5703# 4.56e-19
C89 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_7889_n6842# 0.00288f
C90 a_10810_n6777# DVDD 0.243f
C91 a_838_n6794# DVDD 0.238f
C92 a_6349_9307# VDD 0.701f
C93 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 DVDD 0.147f
C94 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 0.839f
C95 a_7464_n6798# SELB 0.0221f
C96 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 0.301f
C97 a_10965_3602# VDD 0.0939f
C98 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 a_10810_n6777# 1.09e-19
C99 a_570_n5724# DVDD 0.116f
C100 a_7096_n5816# a_7464_n6798# 0.139f
C101 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 0.0365f
C102 a_7196_n5728# a_8403_n6064# 0.289f
C103 a_570_n5724# a_838_n6794# 0.0272f
C104 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp B1 1.5f
C105 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_7196_n5728# 0.00139f
C106 comparator_top_0.VINM a_7196_n5728# 0.0032f
C107 a_4609_n6817# EF_AMUX21m_1.invm_0.Y 0.00503f
C108 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 2.6e-19
C109 a_470_n5812# a_1777_n6060# 3.88e-20
C110 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 a_3916_n5703# 6.2e-19
C111 a_5123_n6039# VDD 0.489f
C112 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VDD 2.65f
C113 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb A1 1.01f
C114 a_10975_4108# DVDD 0.466f
C115 a_3816_n5791# a_4609_n6817# 8.36e-19
C116 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.invm_0.Y 1.69e-19
C117 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_470_n5812# 0.00188f
C118 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 a_10542_n5707# 0.00162f
C119 EF_AMUX21m_1.invm_0.Y DVDD 0.946f
C120 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.124f
C121 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 B1 0.525f
C122 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD 3.42f
C123 a_3816_n5791# DVDD 0.435f
C124 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD 1.21f
C125 comparator_top_0.VINP a_470_n5812# 0.00115f
C126 a_8403_n6064# a_7464_n6798# 6.24e-19
C127 a_10442_n5795# a_11235_n6821# 8.36e-19
C128 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 VDD 2.17f
C129 comparator_top_0.comparator_0.VOUT DVDD 0.0256f
C130 comparator_top_0.VINM a_10442_n5795# 0.00115f
C131 a_7196_n5728# B1 4.37e-19
C132 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 SELB 1.12e-20
C133 a_11271_4224# a_11031_3400# 0.25f
C134 a_4184_n6773# VDD 0.154f
C135 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_1263_n6838# 7.05e-21
C136 a_10965_3602# DVDD 0.033f
C137 a_5123_n6039# a_4609_n6817# 2.63e-19
C138 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 a_7096_n5816# 0.00935f
C139 a_7196_n5728# VDD 1.12f
C140 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_1777_n6060# 0.00108f
C141 a_6351_7717# VDD 0.522f
C142 comparator_top_0.comparator_0.VBP comparator_top_0.VINP 0.355f
C143 comparator_top_0.VINM A2 0.00278f
C144 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X SELB 3.51e-19
C145 a_5123_n6039# DVDD 0.0134f
C146 comparator_top_0.VINP a_1777_n6060# 0.00136f
C147 a_11749_n6043# a_11235_n6821# 2.63e-19
C148 comparator_top_0.VINM VSS 4.14f
C149 a_10442_n5795# EF_AMUX21m_2.invm_0.Y 0.235f
C150 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 3.05e-19
C151 comparator_top_0.VINM B2 2.81f
C152 a_7096_n5816# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.00152f
C153 comparator_top_0.comparator_0.VOUT a_10975_4108# 0.0135f
C154 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_4609_n6817# 0.00288f
C155 a_10442_n5795# a_10542_n5707# 0.405f
C156 a_3816_n5791# EF_AMUX21m_1.invm_0.Y 0.235f
C157 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.08f
C158 comparator_top_0.VINM a_11749_n6043# 0.00136f
C159 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 a_1777_n6060# 0.00121f
C160 a_470_n5812# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.00152f
C161 a_10975_4108# a_10965_3602# 0.249f
C162 a_7464_n6798# VDD 0.153f
C163 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.124f
C164 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVDD 0.0946f
C165 a_10442_n5795# VDD 0.335f
C166 a_4609_n6817# a_4184_n6773# 0.461f
C167 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 DVDD 0.126f
C168 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 3.37e-19
C169 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 0.207f
C170 VSS A1 9e-20
C171 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp A1 1.48e-19
C172 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_570_n5724# 0.00139f
C173 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 2.6e-19
C174 a_10542_n5707# B2 4.37e-19
C175 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 0.303f
C176 comparator_top_0.VINP a_3916_n5703# 0.0032f
C177 a_4184_n6773# DVDD 0.24f
C178 a_7889_n6842# SELB 0.0046f
C179 a_8403_n6064# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.145f
C180 a_10542_n5707# a_11749_n6043# 0.289f
C181 comparator_top_0.comparator_0.VOUT a_10965_3602# 0.0309f
C182 a_7196_n5728# DVDD 0.117f
C183 VDD A2 1.89f
C184 VSS SELA 0.0267f
C185 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 a_3916_n5703# 0.00162f
C186 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp VDD 2.65f
C187 VDD VSS 0.151p
C188 a_7096_n5816# a_7889_n6842# 8.36e-19
C189 a_3816_n5791# a_5123_n6039# 3.88e-20
C190 a_1777_n6060# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.145f
C191 VDD B2 1.89f
C192 a_11749_n6043# VDD 0.489f
C193 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_11235_n6821# 0.00288f
C194 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00684f
C195 a_6351_6657# VDD 0.684f
C196 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 B1 2.1e-19
C197 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.00152f
C198 a_11271_4224# VO 0.0547f
C199 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 VDD 2.18f
C200 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X EF_AMUX21m_2.invm_0.Y 8.17e-19
C201 a_7464_n6798# DVDD 0.236f
C202 a_10809_9307# a_10811_8247# 0.139f
C203 a_10442_n5795# DVDD 0.437f
C204 EF_AMUX21m_1.invm_0.Y a_4184_n6773# 0.0217f
C205 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.282f
C206 a_10442_n5795# a_10810_n6777# 0.139f
C207 a_8403_n6064# a_7889_n6842# 2.63e-19
C208 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X B1 8.92e-19
C209 a_3816_n5791# a_4184_n6773# 0.139f
C210 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_7889_n6842# 7.05e-21
C211 comparator_top_0.comparator_0.VBP comparator_top_0.VINM 0.0131f
C212 a_470_n5812# A1 3.15e-19
C213 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD 1.2f
C214 a_10542_n5707# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.0154f
C215 DVDD A2 0.00231f
C216 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb A2 1.01f
C217 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_11235_n6821# 7.05e-21
C218 VSS DVDD 0.00708f
C219 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.34f
C220 DVDD B2 0.00233f
C221 a_470_n5812# SELA 0.235f
C222 a_5123_n6039# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.145f
C223 a_11031_3400# VO 0.0102f
C224 a_470_n5812# VDD 0.326f
C225 a_838_n6794# VSS 0.0013f
C226 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.124f
C227 a_6349_9307# a_6351_7717# 0.14f
C228 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.668f
C229 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 B2 0.518f
C230 a_11749_n6043# DVDD 0.0136f
C231 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_10442_n5795# 0.00188f
C232 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 a_4609_n6817# 3.13e-19
C233 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X VDD 1.2f
C234 a_570_n5724# VSS 0.00169f
C235 a_11749_n6043# a_10810_n6777# 6.24e-19
C236 comparator_top_0.VINM comparator_top_0.VINP 3.44f
C237 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 a_11749_n6043# 0.00121f
C238 a_5123_n6039# a_4184_n6773# 6.24e-19
C239 comparator_top_0.comparator_0.VBN VSS 11.2f
C240 a_11271_4224# VDD 0.17f
C241 a_7096_n5816# SELB 0.235f
C242 a_1777_n6060# A1 3.4e-19
C243 a_470_n5812# a_1263_n6838# 8.36e-19
C244 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_7196_n5728# 4.56e-19
C245 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 DVDD 0.11f
C246 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 0.839f
C247 comparator_top_0.VINM EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 1.54e-19
C248 a_7889_n6842# VDD 0.607f
C249 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp A1 1.5f
C250 comparator_top_0.comparator_0.VBP VDD 10.8f
C251 a_1777_n6060# SELA 5.58e-20
C252 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp B2 1.5f
C253 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_10542_n5707# 0.00139f
C254 a_1777_n6060# VDD 0.489f
C255 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_4184_n6773# 7.03e-19
C256 a_10809_9307# a_10811_7187# 4.42e-21
C257 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_11749_n6043# 0.00108f
C258 a_3816_n5791# A2 3.15e-19
C259 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVDD 0.102f
C260 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_7196_n5728# 8.72e-21
C261 comparator_top_0.VINP A1 2.82f
C262 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp VDD 2.64f
C263 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 a_7196_n5728# 6.2e-19
C264 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_3816_n5791# 0.00188f
C265 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_10810_n6777# 4.53e-21
C266 a_10809_9307# VDD 0.697f
C267 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb VDD 3.43f
C268 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 A1 0.523f
C269 comparator_top_0.comparator_0.VOUT VSS 0.872f
C270 a_8403_n6064# SELB 5.62e-20
C271 a_11031_3400# VDD 0.51f
C272 a_1777_n6060# a_1263_n6838# 2.63e-19
C273 a_470_n5812# DVDD 0.428f
C274 comparator_top_0.VINP VDD 12.7f
C275 a_6349_9307# VSS 3.54e-19
C276 a_7096_n5816# a_8403_n6064# 3.88e-20
C277 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X DVDD 0.0982f
C278 a_470_n5812# a_838_n6794# 0.139f
C279 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 SELA 1.27e-19
C280 comparator_top_0.VINM a_7096_n5816# 0.00115f
C281 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_10810_n6777# 7.03e-19
C282 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 VDD 2.16f
C283 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.282f
C284 a_470_n5812# a_570_n5724# 0.405f
C285 a_3916_n5703# VDD 1.12f
C286 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X a_7464_n6798# 1.96e-19
C287 a_11271_4224# DVDD 0.449f
C288 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 a_7464_n6798# 1.09e-19
C289 a_5123_n6039# A2 3.4e-19
C290 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp A2 1.85e-19
C291 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 a_10442_n5795# 0.0085f
C292 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_5123_n6039# 0.00108f
C293 a_7889_n6842# DVDD 0.188f
C294 EF_AMUX21m_2.invm_0.Y SELB 0.241f
C295 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 a_1263_n6838# 3.13e-19
C296 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X A1 8.93e-19
C297 a_1777_n6060# DVDD 0.0139f
C298 a_7196_n5728# a_7464_n6798# 0.0272f
C299 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X A2 8.92e-19
C300 a_1777_n6060# a_838_n6794# 6.24e-19
C301 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VSS 8.77e-20
C302 comparator_top_0.VINM a_8403_n6064# 0.00136f
C303 comparator_top_0.comparator_0.VBN comparator_top_0.comparator_0.VBP 1.78f
C304 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X SELA 3.51e-19
C305 a_7096_n5816# B1 3.15e-19
C306 VDD SELB 0.0248f
C307 a_570_n5724# a_1777_n6060# 0.289f
C308 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 a_5123_n6039# 0.00121f
C309 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X VDD 1.2f
C310 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.00724f
C311 comparator_top_0.VINM EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.682f
C312 a_11271_4224# a_10975_4108# 0.136f
C313 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 B2 1.85e-19
C314 a_11031_3400# DVDD 0.0693f
C315 a_10811_8247# a_10811_7187# 0.14f
C316 a_3916_n5703# a_4609_n6817# 0.265f
C317 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.h0 0.839f
C318 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_570_n5724# 4.56e-19
C319 a_7096_n5816# VDD 0.336f
C320 comparator_top_0.VINP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.668f
C321 a_10811_8247# VDD 0.508f
C322 a_11235_n6821# EF_AMUX21m_2.invm_0.Y 0.00503f
C323 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 DVDD 0.124f
C324 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 2.72e-19
C325 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_1263_n6838# 0.00288f
C326 a_3916_n5703# DVDD 0.115f
C327 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.X 0.282f
C328 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_3916_n5703# 0.00139f
C329 comparator_top_0.VINP a_570_n5724# 0.0032f
C330 a_10542_n5707# a_11235_n6821# 0.265f
C331 a_6351_7717# VSS 3.36e-19
C332 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 a_838_n6794# 1.09e-19
C333 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 3.11e-19
C334 comparator_top_0.comparator_0.VOUT a_11271_4224# 0.00564f
C335 comparator_top_0.comparator_0.VBN comparator_top_0.VINP 0.09f
C336 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 a_570_n5724# 6.2e-19
C337 comparator_top_0.VINM a_10542_n5707# 0.0032f
C338 a_8403_n6064# B1 3.4e-19
C339 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.34f
C340 a_10975_4108# a_11031_3400# 0.166f
C341 a_11271_4224# a_10965_3602# 7.97e-19
C342 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 a_4184_n6773# 1.09e-19
C343 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb B1 1.01f
C344 a_11235_n6821# VDD 0.607f
C345 comparator_top_0.VINM B1 2.82f
C346 VDD VO 0.268f
C347 a_6351_7717# a_6351_6657# 0.14f
C348 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.h0 a_7196_n5728# 0.00196f
C349 a_8403_n6064# VDD 0.489f
C350 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.282f
C351 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb VDD 3.43f
C352 comparator_top_0.VINM VDD 14.1f
C353 DVDD SELB 0.921f
C354 a_10442_n5795# B2 3.15e-19
C355 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X DVDD 0.101f
C356 comparator_top_0.VINP a_3816_n5791# 0.00115f
C357 a_10542_n5707# EF_AMUX21m_2.invm_0.Y 0.00242f
C358 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 EF_AMUX21m_1.invm_0.Y 1.69e-19
C359 comparator_top_0.comparator_0.VOUT a_11031_3400# 0.225f
C360 a_10442_n5795# a_11749_n6043# 3.88e-20
C361 a_3916_n5703# EF_AMUX21m_1.invm_0.Y 0.00242f
C362 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X a_838_n6794# 7.03e-19
C363 a_7196_n5728# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.0154f
C364 a_7096_n5816# DVDD 0.431f
C365 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.h0 a_3816_n5791# 0.0085f
C366 a_3816_n5791# a_3916_n5703# 0.405f
C367 a_570_n5724# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.X 0.0154f
C368 a_11031_3400# a_10965_3602# 0.17f
C369 EF_AMUX21m_2.invm_0.Y VDD 0.0233f
C370 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp A2 1.5f
C371 a_10542_n5707# VDD 1.12f
C372 VDD A1 1.9f
C373 a_10811_7187# VDD 0.512f
C374 VDD B1 1.89f
C375 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.h0 a_7889_n6842# 3.13e-19
C376 a_11749_n6043# B2 3.4e-19
C377 VDD SELA 0.0292f
C378 comparator_top_0.VINP a_5123_n6039# 0.00136f
.ends

