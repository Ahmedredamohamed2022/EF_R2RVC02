* NGSPICE file created from EF_R2RVC02.ext - technology: sky130A

.subckt EF_R2RVC02 VSS A1 A2 SELB VO B2 B1 SELA VDD DVSS DVDD EN
X0 a_4503_4914.t3 EF_AMUX2to1ISO_0.VO a_1297_4914.t1 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X1 VSS.t8 EF_R2RVCE_0.comparator_0.VBN.t9 a_1297_2982.t0 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X2 VSS.t18 a_1355_1794.t8 a_1755_1820.t5 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X3 a_6639_n11591# a_6271_n10609# DVDD.t1 DVDD.t0 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X4 DVSS.t6 a_10169_4802# a_10179_5308# DVSS.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X5 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10204_n8486.t3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t173 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.03 ps=18.1 w=1 l=0.5
X6 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t7 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A DVSS.t266 DVSS.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X7 VDD.t123 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6804_n8486.t1 VDD.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL SELB.t0 DVSS.t60 DVSS.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X9 DVSS.t173 a_10179_5308# VO.t1 DVSS.t172 sky130_fd_pr__nfet_01v8 ad=0.196 pd=2.01 as=0.196 ps=2.01 w=0.74 l=0.15
X10 VDD.t99 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3606_n8490.t1 VDD.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X11 DVSS.t94 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t2 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB DVSS.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X12 a_10235_4600# EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A VDD.t207 VDD.t206 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X13 VSS.t55 VSS.t54 VSS.t55 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X14 a_4503_4914.t7 a_4503_4914.t6 VSS.t22 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X15 a_10914_2086# a_10618_2709# DVSS.t253 DVSS.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t3 a_6804_n3484.t3 EF_AMUX2to1ISO_1.VO DVSS.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X17 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t2 DVSS.t197 DVSS.t196 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X18 VDD.t175 a_10204_n8486.t4 a_10209_n9511.t1 VDD.t174 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X19 VDD.t205 a_n227_n10525# a_466_n11639# VDD.t204 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X20 a_10464_n11635# a_10039_n11591# DVSS.t36 DVSS.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X21 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3606_n3488.t3 EF_AMUX2to1ISO_0.VO DVSS.t38 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X22 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3611_n4513# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.2 ps=33.6 w=2 l=0.5
X23 DVDD.t11 SELA.t0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL DVDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X24 VSS.t53 VSS.t51 EF_R2RVCE_0.comparator_0.VBN.t4 VSS.t52 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X25 EF_AMUX2to1ISO_0.VO a_206_n3488.t3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN DVSS.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X26 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3611_n9515.t3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X27 a_10204_n8486.t1 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD.t108 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X28 a_1297_4914.t0 EF_AMUX2to1ISO_0.VO a_4503_4914.t2 VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X29 EF_AMUX2to1ISO_0.VO a_211_n4513# EF_AMUX2to1ISO_0.VO DVSS.t148 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=0.5
X30 DVSS.t188 a_10204_n8486.t5 a_10209_n9511.t2 DVSS.t187 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X31 a_1355_1794.t7 a_1355_1794.t6 VSS.t14 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X32 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t3 DVSS.t115 DVSS.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X33 DVSS.t144 a_9671_n10609# a_9771_n10521# DVSS.t143 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X34 DVSS.t80 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_206_n8490.t2 DVSS.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X35 a_6639_n11591# a_6271_n10609# DVSS.t18 DVSS.t17 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X36 B1.t7 a_6804_n8486.t3 B1.t6 VDD.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X37 DVDD.t38 a_10180_3343# a_10136_2294# DVDD.t37 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X38 EF_AMUX2to1ISO_1.VO a_10204_n3484.t3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X39 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL SELA.t1 DVSS.t255 DVSS.t254 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X40 VDD.t22 a_10464_n11635# a_9771_n10521# VDD.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X41 VDD.t189 a_9771_n10521# a_10978_n10857# VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X42 EF_R2RVCE_0.comparator_0.VBN.t5 a_1425_9823.t6 EF_R2RVCE_0.comparator_bias_0.down VDD.t182 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
D0 DVSS.t86 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X43 B2.t7 a_10209_n9511.t3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X44 DVSS.t50 a_3441_n11595# a_3866_n11639# DVSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X45 a_9771_n10521# a_9671_n10609# DVSS.t142 DVSS.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X46 a_9771_n10521# a_9671_n10609# DVSS.t140 DVSS.t139 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X47 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t0 a_4380_n10861# VDD.t200 VDD.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X48 a_1425_9823.t4 EF_R2RVCE_0.comparator_bias_0.down VDD.t155 VDD.t154 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X49 VDD.t60 VDD.t59 VDD.t60 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X50 DVSS.t252 a_10136_2294# a_10162_2241# DVSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X51 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_8085_2982.t2 VSS.t13 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X52 DVSS.t85 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3606_n3488.t2 DVSS.t84 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X53 EF_AMUX2to1ISO_1.VO a_6809_n4509# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t7 VDD.t125 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X54 DVSS.t195 SELA.t2 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL DVSS.t194 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X55 VDD.t74 a_6371_n10521# a_7064_n11635# VDD.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X56 DVDD.t30 SELA.t3 a_n327_n10613# DVDD.t29 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X57 VSS.t7 EF_R2RVCE_0.comparator_0.VBN.t10 EF_R2RVCE_0.comparator_0.VBP.t0 VSS.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X58 DVDD.t40 a_10475_5424# a_10179_5308# DVDD.t39 sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.297 ps=2.77 w=1.12 l=0.15
X59 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3611_n4513# EF_AMUX2to1ISO_0.VO VDD.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X60 DVSS.t4 a_10169_4802# a_10179_5308# DVSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X61 EF_AMUX2to1ISO_0.VO a_3606_n3488.t4 EF_AMUX2to1ISO_0.VO VDD.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.32 ps=20.6 w=1 l=0.5
X62 DVSS.t70 a_6371_n10521# a_7578_n10857# DVSS.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X63 a_1297_4914.t7 EF_AMUX2to1ISO_1.VO a_1355_1794.t3 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X64 a_10162_2241# a_10136_2294# DVSS.t251 DVSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X65 a_3611_n4513# a_3606_n3488.t5 VDD.t19 VDD.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X66 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_206_n8490.t3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN VDD.t71 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.03 ps=18.1 w=1 l=0.5
X67 A1.t3 a_206_n8490.t4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN DVSS.t162 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X68 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t1 a_980_n10861# DVSS.t64 DVSS.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X69 a_10475_5424# a_10179_5308# DVDD.t24 DVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.297 pd=2.77 as=0.157 ps=1.4 w=1.12 l=0.15
X70 DVSS.t106 a_41_n11595# a_466_n11639# DVSS.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X71 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t1 a_10978_n10857# DVSS.t26 DVSS.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X72 EF_R2RVCE_0.comparator_0.VOUTANALOG.t2 a_1755_1820.t6 VDD.t124 VDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X73 EF_AMUX2to1ISO_0.VO a_3611_n4513# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X74 a_4503_2982.t3 EF_AMUX2to1ISO_0.VO a_1297_2982.t3 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X75 a_10162_2241# a_10618_2709# VDD.t196 VDD.t195 sky130_fd_pr__pfet_g5v0d10v5 ad=0.137 pd=1.49 as=0.111 ps=1.37 w=0.42 l=1
X76 VDD.t121 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6804_n3484.t1 VDD.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X77 DVSS.t3 a_10169_4802# a_10179_5308# DVSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X78 DVSS.t184 a_6639_n11591# a_7064_n11635# DVSS.t183 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X79 DVSS.t229 SELA.t4 a_n327_n10613# DVSS.t228 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X80 a_1425_9823.t5 VSS.t48 VSS.t50 VSS.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X81 VDD.t159 a_10204_n3484.t4 a_10209_n4509# VDD.t158 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X82 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10204_n3484.t5 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X83 a_10180_3343# EN.t0 DVSS.t150 DVSS.t149 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X84 a_5555_8917# a_10015_8387# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X85 a_10204_n3484.t1 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD.t107 VDD.t61 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X86 EF_R2RVCE_0.comparator_bias_0.down a_1425_9823.t7 EF_R2RVCE_0.comparator_0.VBN.t6 VDD.t183 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X87 VDD.t192 a_4503_2982.t6 a_4503_2982.t7 VDD.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X88 DVSS.t231 a_10204_n3484.t6 a_10209_n4509# DVSS.t230 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X89 a_1297_4914.t9 VDD.t57 VDD.t58 VDD.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X90 VDD.t133 a_10914_2086# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A VDD.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X91 VDD.t181 a_6804_n8486.t4 a_6809_n9511.t1 VDD.t180 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X92 DVSS.t221 a_n327_n10613# a_n227_n10525# DVSS.t220 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X93 a_3173_n10525# a_3073_n10613# DVSS.t209 DVSS.t208 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X94 a_1297_2982.t2 EF_AMUX2to1ISO_0.VO a_4503_2982.t2 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X95 EF_R2RVCE_0.comparator_0.VOUTANALOG.t5 a_4503_4914.t8 VSS.t21 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X96 A1.t4 a_211_n9515.t3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X97 VSS.t47 VSS.t45 VSS.t46 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X98 a_10618_2709# a_10180_3343# DVSS.t242 DVSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X99 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t5 a_6809_n4509# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t4 DVSS.t130 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X100 a_211_n9515.t1 a_206_n8490.t5 VDD.t64 VDD.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X101 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL SELA.t5 DVDD.t21 DVDD.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X102 DVSS.t224 a_6804_n8486.t5 a_6809_n9511.t2 DVSS.t223 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X103 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t10 a_6809_n9511.t3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t9 DVSS.t193 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X104 DVSS.t113 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10204_n8486.t2 DVSS.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X105 DVDD.t9 SELB.t1 a_6271_n10609# DVDD.t8 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X106 DVDD.t23 a_10179_5308# VO.t0 DVDD.t22 sky130_fd_pr__pfet_01v8_hvt ad=0.157 pd=1.4 as=0.297 ps=2.77 w=1.12 l=0.15
X107 B2.t3 a_10204_n8486.t6 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t67 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X108 a_7064_n11635# a_6639_n11591# DVSS.t182 DVSS.t181 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X109 a_3866_n11639# a_3441_n11595# DVSS.t48 DVSS.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X110 VDD.t72 a_6371_n10521# a_7578_n10857# VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X111 a_1297_4914.t10 EF_R2RVCE_0.comparator_0.VBP.t4 VDD.t190 VDD.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X112 VSS.t16 a_1355_1794.t4 a_1355_1794.t5 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
D1 DVSS.t123 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X113 a_4503_4914.t1 EF_AMUX2to1ISO_0.VO a_1297_4914.t3 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X114 a_6371_n10521# a_6271_n10609# DVSS.t16 DVSS.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X115 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_206_n3488.t4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X116 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_211_n9515.t4 A1.t7 VDD.t172 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X117 a_10464_n11635# a_10039_n11591# DVSS.t34 DVSS.t33 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X118 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t0 a_10978_n10857# VDD.t15 VDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X119 VDD.t56 VDD.t54 VDD.t56 VDD.t55 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X120 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t6 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A DVSS.t265 DVSS.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X121 EF_AMUX2to1ISO_1.VO a_6804_n3484.t4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t2 DVSS.t22 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X122 a_n227_n10525# a_n327_n10613# DVSS.t219 DVSS.t218 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X123 VDD.t168 a_3866_n11639# a_3173_n10525# VDD.t167 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X124 a_206_n3488.t1 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD.t91 VDD.t90 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X125 VSS.t44 VSS.t43 VSS.t44 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X126 B1.t0 a_6809_n9511.t4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t11 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X127 a_n227_n10525# a_n327_n10613# DVSS.t217 DVSS.t216 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X128 a_1355_1794.t2 EF_AMUX2to1ISO_1.VO a_1297_4914.t5 VDD.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X129 DVSS.t261 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10235_4600# DVSS.t260 sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X130 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t14 a_6804_n8486.t6 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t13 VDD.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X131 VDD.t161 a_1755_1820.t2 a_1755_1820.t3 VDD.t160 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X132 VSS.t20 a_4503_4914.t9 EF_R2RVCE_0.comparator_0.VOUTANALOG.t4 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X133 a_5553_10507# a_10013_10507# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X134 a_5555_7857# EF_R2RVCE_0.comparator_bias_0.up DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X135 a_5553_10507# a_10015_9447# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X136 a_1297_2982.t10 EF_AMUX2to1ISO_1.VO a_1355_5983.t7 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X137 DVSS.t264 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t5 DVSS.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X138 DVSS.t192 SELB.t2 a_6271_n10609# DVSS.t191 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X139 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t1 a_7578_n10857# DVSS.t24 DVSS.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X140 EF_R2RVCE_0.comparator_0.VOUTANALOG.t0 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t8 VSS.t10 VSS.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=2
X141 VDD.t203 a_n227_n10525# a_980_n10861# VDD.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X142 DVSS.t161 a_10235_4600# a_10475_5424# DVSS.t160 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.199 ps=2.03 w=0.75 l=0.5
X143 a_1755_6080.t3 a_1755_6080.t2 VSS.t56 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X144 VDD.t178 a_3606_n8490.t3 a_3611_n9515.t1 VDD.t177 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X145 A2.t3 a_3606_n8490.t4 A2.t2 VDD.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X146 DVSS.t215 a_n327_n10613# a_n227_n10525# DVSS.t214 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X147 VDD.t157 a_206_n3488.t5 a_211_n4513# VDD.t156 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X148 a_6804_n8486.t0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD.t119 VDD.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X149 DVSS.t164 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB DVSS.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X150 a_10475_5424# a_10235_4600# DVSS.t159 DVSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X151 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t3 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A VDD.t212 VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X152 a_3606_n8490.t0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD.t97 VDD.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X153 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10209_n9511.t4 B2.t6 VDD.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X154 VDD.t110 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD.t109 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X155 DVSS.t186 a_3606_n8490.t5 a_3611_n9515.t2 DVSS.t185 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X156 VSS.t42 VSS.t41 VSS.t42 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X157 DVSS.t146 a_10914_2086# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A DVSS.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X158 DVSS.t152 a_206_n3488.t6 a_211_n4513# DVSS.t151 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X159 a_10209_n9511.t0 a_10204_n8486.t7 VDD.t70 VDD.t69 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X160 VDD.t68 EF_R2RVCE_0.comparator_0.VOUTANALOG.t9 a_8085_2982.t0 VDD.t67 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.3 as=2.9 ps=20.6 w=10 l=2
X161 EF_AMUX2to1ISO_0.VO a_3606_n3488.t6 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t96 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X162 B2.t5 a_10209_n9511.t5 B2.t4 DVSS.t95 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X163 a_41_n11595# a_n327_n10613# DVDD.t34 DVDD.t33 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X164 a_10180_3343# EN.t1 DVDD.t28 DVDD.t27 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X165 EF_AMUX2to1ISO_1.VO a_10209_n4509# EF_AMUX2to1ISO_1.VO DVSS.t168 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.64 ps=36.6 w=2 l=0.5
X166 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t2 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A VDD.t211 VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
D2 DVSS.t111 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X167 VDD.t89 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_206_n8490.t1 VDD.t88 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X168 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t4 DVSS.t166 DVSS.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X169 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t5 VDD.t112 VDD.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X170 VSS.t15 a_1755_6080.t6 EF_R2RVCE_0.comparator_0.VOUTANALOG.t3 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X171 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t6 DVSS.t190 DVSS.t189 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X172 VSS.t5 EF_R2RVCE_0.comparator_0.VBN.t11 a_1425_9823.t0 VSS.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X173 VDD.t2 a_1355_5983.t8 a_1755_6080.t5 VDD.t1 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X174 DVSS.t250 a_10136_2294# a_10162_2241# DVSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X175 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_211_n4513# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN DVSS.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.2 ps=33.6 w=2 l=0.5
X176 VDD.t8 a_6804_n3484.t5 a_6809_n4509# VDD.t7 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X177 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t2 DVSS.t244 DVSS.t243 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X178 DVSS.t171 a_3173_n10525# a_4380_n10861# DVSS.t170 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X179 DVSS.t241 a_10180_3343# a_10618_2709# DVSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X180 a_9771_n10521# a_9671_n10609# DVSS.t138 DVSS.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X181 a_1297_2982.t11 VSS.t39 VSS.t40 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X182 DVSS.t110 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10204_n3484.t2 DVSS.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
D3 DVSS.t78 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X183 a_1755_1820.t4 a_1355_1794.t9 VSS.t12 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X184 DVSS.t62 a_6804_n3484.t6 a_6809_n4509# DVSS.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X185 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL SELB.t3 DVDD.t26 DVDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X186 VDD.t210 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t1 VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X187 EF_AMUX2to1ISO_1.VO a_10204_n3484.t7 EF_AMUX2to1ISO_1.VO VDD.t193 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.32 ps=20.6 w=1 l=0.5
X188 DVSS.t88 SELA.t6 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL DVSS.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X189 VDD.t53 VDD.t51 VDD.t53 VDD.t52 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X190 a_4503_2982.t5 a_4503_2982.t4 VDD.t166 VDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X191 a_41_n11595# a_n327_n10613# DVSS.t213 DVSS.t212 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X192 VDD.t95 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3606_n3488.t1 VDD.t94 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X193 a_7064_n11635# a_6639_n11591# DVSS.t180 DVSS.t179 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X194 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t0 a_7578_n10857# VDD.t13 VDD.t12 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X195 a_1297_2982.t1 EF_R2RVCE_0.comparator_0.VBN.t12 VSS.t3 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X196 VDD.t188 a_9771_n10521# a_10464_n11635# VDD.t187 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X197 a_4503_2982.t1 EF_AMUX2to1ISO_0.VO a_1297_2982.t5 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X198 B1.t5 a_6804_n8486.t7 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t16 DVSS.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X199 a_466_n11639# a_41_n11595# DVSS.t104 DVSS.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X200 A2.t1 a_3606_n8490.t6 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t222 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X201 A2.t7 a_3611_n9515.t4 A2.t6 DVSS.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X202 EF_R2RVCE_0.comparator_bias_0.down EF_R2RVCE_0.comparator_0.VBN.t0 EF_R2RVCE_0.comparator_0.VBN.t1 VDD.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=15
X203 EF_R2RVCE_0.comparator_0.VBN.t3 EF_R2RVCE_0.comparator_0.VBN.t2 VSS.t1 VSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X204 a_1355_5983.t3 a_1355_5983.t2 VDD.t135 VDD.t134 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X205 VDD.t50 VDD.t48 a_1297_4914.t8 VDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X206 EF_AMUX2to1ISO_0.VO a_3611_n4513# EF_AMUX2to1ISO_0.VO DVSS.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X207 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_206_n8490.t6 A1.t2 DVSS.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X208 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_211_n9515.t5 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN DVSS.t234 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X209 DVSS.t207 a_3073_n10613# a_3173_n10525# DVSS.t206 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X210 DVDD.t15 SELB.t4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL DVDD.t14 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X211 DVSS.t14 a_6271_n10609# a_6371_n10521# DVSS.t13 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X212 VDD.t47 VDD.t45 VDD.t46 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X213 a_1355_5983.t6 EF_AMUX2to1ISO_1.VO a_1297_2982.t9 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X214 DVSS.t77 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_206_n3488.t2 DVSS.t76 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X215 DVSS.t158 a_10235_4600# a_10169_4802# DVSS.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0.179 pd=1.26 as=0.12 ps=1.41 w=0.42 l=0.5
X216 DVSS.t263 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t4 DVSS.t262 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X217 a_466_n11639# a_41_n11595# DVSS.t102 DVSS.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X218 a_1297_4914.t6 EF_AMUX2to1ISO_1.VO a_1355_1794.t1 VDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X219 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t1 a_6804_n3484.t7 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t0 VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X220 DVSS.t178 a_6639_n11591# a_7064_n11635# DVSS.t177 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X221 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10204_n8486.t8 B2.t2 DVSS.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X222 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t0 a_980_n10861# VDD.t31 VDD.t30 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X223 DVSS.t156 a_10235_4600# a_10475_5424# DVSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X224 a_6804_n3484.t0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD.t117 VDD.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X225 a_3866_n11639# a_3441_n11595# DVSS.t46 DVSS.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X226 DVDD.t13 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL a_3073_n10613# DVDD.t12 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X227 a_6371_n10521# a_6271_n10609# DVSS.t12 DVSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X228 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10209_n4509# EF_AMUX2to1ISO_1.VO VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
D4 DVSS.t83 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X229 DVSS.t32 a_10039_n11591# a_10464_n11635# DVSS.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X230 VDD.t131 a_466_n11639# a_n227_n10525# VDD.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X231 a_3173_n10525# a_3073_n10613# DVSS.t205 DVSS.t204 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X232 VDD.t153 EF_R2RVCE_0.comparator_bias_0.down a_1425_9823.t3 VDD.t152 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X233 a_10209_n4509# a_10204_n3484.t8 VDD.t197 VDD.t147 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X234 DVSS.t246 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB DVSS.t245 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X235 VDD.t44 VDD.t42 VDD.t44 VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X236 DVSS.t125 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6804_n8486.t2 DVSS.t124 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X237 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL SELA.t7 DVDD.t7 DVDD.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X238 DVSS.t82 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3606_n8490.t2 DVSS.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X239 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t12 a_6809_n9511.t5 B1.t3 VDD.t186 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X240 a_3441_n11595# a_3073_n10613# DVDD.t32 DVDD.t31 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X241 VSS.t17 EF_R2RVCE_0.comparator_0.VOUTANALOG.t10 a_8085_2982.t1 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X242 A2.t5 a_3611_n9515.t5 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X243 a_7064_n11635# a_6639_n11591# DVSS.t176 DVSS.t175 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X244 EF_R2RVCE_0.comparator_0.VBP.t1 VSS.t36 VSS.t38 VSS.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X245 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_206_n3488.t7 EF_AMUX2to1ISO_0.VO DVSS.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X246 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3606_n8490.t7 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t179 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=2.03 ps=18.1 w=1 l=0.5
X247 a_6809_n9511.t0 a_6804_n8486.t8 VDD.t81 VDD.t80 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X248 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL SELB.t5 DVSS.t90 DVSS.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X249 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t9 EF_R2RVCE_0.comparator_bias_0.down VDD.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=5.8 pd=40.6 as=5.8 ps=40.6 w=20 l=2
X250 EF_AMUX2to1ISO_0.VO a_206_n3488.t8 EF_AMUX2to1ISO_0.VO VDD.t201 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X251 a_3611_n9515.t0 a_3606_n8490.t8 VDD.t62 VDD.t32 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X252 VDD.t106 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10204_n8486.t0 VDD.t105 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X253 a_1355_1794.t0 EF_AMUX2to1ISO_1.VO a_1297_4914.t4 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X254 DVSS.t249 a_10136_2294# a_10162_2241# DVSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X255 a_10464_n11635# a_10039_n11591# DVSS.t30 DVSS.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X256 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t4 DVSS.t54 DVSS.t53 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X257 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t1 a_4380_n10861# DVSS.t257 DVSS.t256 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.122 ps=1.08 w=0.75 l=0.5
X258 DVDD.t36 SELB.t6 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL DVDD.t35 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X259 DVDD.t3 SELA.t8 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL DVDD.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X260 DVSS.t72 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL a_3073_n10613# DVSS.t71 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X261 DVSS.t56 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t2 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB DVSS.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X262 EF_R2RVCE_0.comparator_0.VBN.t7 a_1425_9823.t8 EF_R2RVCE_0.comparator_bias_0.down VDD.t184 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X263 a_10169_4802# a_10235_4600# VDD.t143 VDD.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.12 ps=1.41 w=0.42 l=0.5
X264 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3611_n9515.t6 A2.t4 VDD.t82 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X265 VDD.t41 VDD.t40 VDD.t41 VDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X266 VDD.t209 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t0 VDD.t208 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X267 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t3 DVSS.t58 DVSS.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0.145 pd=1.58 as=0.145 ps=1.58 w=0.5 l=8
X268 VDD.t24 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t5 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X269 DVSS.t136 a_9671_n10609# a_9771_n10521# DVSS.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X270 EF_R2RVCE_0.comparator_0.VOUTANALOG.t6 a_1755_6080.t7 VSS.t24 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X271 a_10162_2241# a_10136_2294# DVSS.t248 DVSS.t247 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X272 DVSS.t227 SELB.t7 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL DVSS.t226 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.105 ps=1.03 w=0.75 l=0.5
X273 a_3441_n11595# a_3073_n10613# DVSS.t203 DVSS.t202 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X274 a_10618_2709# a_10180_3343# DVSS.t240 DVSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X275 VDD.t84 a_7064_n11635# a_6371_n10521# VDD.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X276 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t4 DVSS.t132 DVSS.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X277 B2.t1 a_10204_n8486.t9 B2.t0 VDD.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X278 a_1297_4914.t2 EF_AMUX2to1ISO_0.VO a_4503_4914.t0 VDD.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X279 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL SELA.t9 DVSS.t128 DVSS.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.214 ps=2.07 w=0.75 l=0.5
X280 VDD.t165 a_3173_n10525# a_3866_n11639# VDD.t164 sky130_fd_pr__pfet_g5v0d10v5 ad=0.111 pd=1.37 as=0.137 ps=1.49 w=0.42 l=1
X281 EF_R2RVCE_0.comparator_0.VBP.t3 EF_R2RVCE_0.comparator_0.VBP.t2 VDD.t29 VDD.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=1.45 ps=10.6 w=5 l=2
X282 EF_R2RVCE_0.comparator_0.VOUTANALOG.t7 a_4503_2982.t8 VDD.t198 VDD.t49 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X283 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t6 VDD.t139 VDD.t138 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X284 VDD.t127 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t5 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X285 VDD.t39 VDD.t36 VDD.t38 VDD.t37 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X286 VSS.t35 VSS.t34 a_1297_2982.t6 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X287 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_211_n4513# EF_AMUX2to1ISO_0.VO VDD.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X288 VDD.t191 EF_R2RVCE_0.comparator_0.VBP.t5 a_1297_4914.t11 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X289 a_10618_2709# a_10162_2241# VDD.t129 VDD.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0.214 pd=1.99 as=0.214 ps=1.99 w=0.42 l=1
X290 VDD.t114 a_1355_5983.t0 a_1355_5983.t1 VDD.t113 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X291 VSS.t33 VSS.t31 VSS.t32 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45 pd=10.6 as=0 ps=0 w=5 l=2
X292 VSS.t19 a_4503_4914.t4 a_4503_4914.t5 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X293 a_211_n4513# a_206_n3488.t9 VDD.t202 VDD.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X294 B1.t2 a_6809_n9511.t6 B1.t1 DVSS.t225 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X295 VDD.t145 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t5 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0.428 pd=3.57 as=0.21 ps=1.78 w=1.5 l=0.5
X296 EF_AMUX2to1ISO_1.VO a_6809_n4509# EF_AMUX2to1ISO_1.VO DVSS.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
D5 DVSS.t122 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X297 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10204_n3484.t9 EF_AMUX2to1ISO_1.VO DVSS.t37 sky130_fd_pr__nfet_g5v0d10v5 ad=0.29 pd=2.29 as=0.58 ps=4.58 w=2 l=0.5
X298 a_10039_n11591# a_9671_n10609# DVDD.t19 DVDD.t18 sky130_fd_pr__pfet_01v8_hvt ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X299 a_1297_2982.t8 EF_AMUX2to1ISO_1.VO a_1355_5983.t5 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X300 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t6 VDD.t171 VDD.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X301 DVDD.t17 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL a_9671_n10609# DVDD.t16 sky130_fd_pr__pfet_01v8_hvt ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X302 EF_AMUX2to1ISO_0.VO a_211_n4513# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN VDD.t136 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X303 A1.t1 a_206_n8490.t7 A1.t0 VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X304 a_3866_n11639# a_3441_n11595# DVSS.t44 DVSS.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X305 DVSS.t100 a_41_n11595# a_466_n11639# DVSS.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X306 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t6 VDD.t11 VDD.t10 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.428 ps=3.57 w=1.5 l=0.5
X307 a_5555_8917# a_10015_9447# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X308 VDD.t199 a_4503_2982.t9 EF_R2RVCE_0.comparator_0.VOUTANALOG.t8 VDD.t43 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X309 DVSS.t121 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6804_n3484.t2 DVSS.t120 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X310 a_206_n8490.t0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD.t87 VDD.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X311 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t15 a_6804_n8486.t9 B1.t4 DVSS.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X312 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t6 a_6809_n4509# EF_AMUX2to1ISO_1.VO VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X313 DVSS.t40 SELB.t8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL DVSS.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=0.214 pd=2.07 as=0.105 ps=1.03 w=0.75 l=0.5
X314 VSS.t30 VSS.t29 VSS.t30 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X315 VSS.t28 VSS.t27 VSS.t28 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X316 EF_AMUX2to1ISO_1.VO a_6804_n3484.t8 EF_AMUX2to1ISO_1.VO VDD.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X317 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL SELB.t9 DVDD.t5 DVDD.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X318 a_6809_n4509# a_6804_n3484.t9 VDD.t66 VDD.t65 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X319 VDD.t104 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10204_n3484.t0 VDD.t103 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X320 DVSS.t201 a_3073_n10613# a_3173_n10525# DVSS.t200 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X321 a_1755_1820.t1 a_1755_1820.t0 VDD.t116 VDD.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X322 a_10914_2086# a_10618_2709# VDD.t194 VDD.t132 sky130_fd_pr__pfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.244 ps=1.83 w=1.5 l=0.5
X323 a_1425_9823.t2 EF_R2RVCE_0.comparator_bias_0.down VDD.t151 VDD.t150 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=1.45 ps=10.6 w=5 l=2
X324 a_1355_5983.t4 EF_AMUX2to1ISO_1.VO a_1297_2982.t7 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X325 VSS.t23 a_1755_6080.t0 a_1755_6080.t1 VSS.t11 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X326 a_10039_n11591# a_9671_n10609# DVSS.t134 DVSS.t133 sky130_fd_pr__nfet_01v8 ad=0.248 pd=2.27 as=0.118 ps=1.12 w=0.84 l=0.15
X327 a_466_n11639# a_41_n11595# DVSS.t98 DVSS.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X328 VDD.t102 a_3606_n3488.t7 a_3611_n4513# VDD.t101 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X329 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3606_n3488.t8 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0 ps=0 w=1 l=0.5
X330 DVSS.t117 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL a_9671_n10609# DVSS.t116 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X331 DVSS.t42 a_3441_n11595# a_3866_n11639# DVSS.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X332 VDD.t35 VDD.t33 VDD.t35 VDD.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X333 VDD.t78 a_206_n8490.t8 a_211_n9515.t0 VDD.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X334 a_n227_n10525# a_n327_n10613# DVSS.t211 DVSS.t210 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X335 VDD.t163 a_3173_n10525# a_4380_n10861# VDD.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0.244 pd=1.83 as=0.398 ps=3.53 w=1.5 l=0.5
X336 a_10475_5424# a_10235_4600# DVSS.t155 DVSS.t154 sky130_fd_pr__nfet_g5v0d10v5 ad=0.199 pd=2.03 as=0.105 ps=1.03 w=0.75 l=0.5
X337 DVSS.t239 a_10180_3343# a_10136_2294# DVSS.t238 sky130_fd_pr__nfet_01v8 ad=0.118 pd=1.12 as=0.248 ps=2.27 w=0.84 l=0.15
X338 a_3606_n3488.t0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD.t93 VDD.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X339 EF_AMUX2to1ISO_1.VO a_10209_n4509# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD.t146 sky130_fd_pr__pfet_g5v0d10v5 ad=0.29 pd=2.58 as=0.145 ps=1.29 w=1 l=0.5
X340 a_3173_n10525# a_3073_n10613# DVSS.t199 DVSS.t198 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
X341 DVSS.t10 a_6271_n10609# a_6371_n10521# DVSS.t9 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X342 VSS.t26 VSS.t25 VSS.t26 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0 ps=0 w=5 l=2
X343 DVSS.t119 a_3606_n3488.t9 a_3611_n4513# DVSS.t118 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X344 DVSS.t92 a_206_n8490.t9 a_211_n9515.t2 DVSS.t91 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.58 ps=4.58 w=2 l=0.5
X345 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_8085_2982.t3 VDD.t76 VDD.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9 pd=20.6 as=1.45 ps=10.3 w=10 l=2
X346 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10209_n4509# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=4.2 ps=33.6 w=2 l=0.5
X347 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3606_n8490.t9 A2.t0 DVSS.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0.29 ps=2.29 w=2 l=0.5
X348 VDD.t169 a_1755_1820.t7 EF_R2RVCE_0.comparator_0.VOUTANALOG.t1 VDD.t3 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X349 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10209_n9511.t6 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN DVSS.t126 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X350 VDD.t149 EF_R2RVCE_0.comparator_bias_0.down a_1425_9823.t1 VDD.t148 sky130_fd_pr__pfet_g5v0d10v5 ad=1.45 pd=10.6 as=0.725 ps=5.29 w=5 l=2
X351 EF_R2RVCE_0.comparator_bias_0.down a_1425_9823.t9 EF_R2RVCE_0.comparator_0.VBN.t8 VDD.t185 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X352 VDD.t86 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_206_n3488.t0 VDD.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0.145 pd=1.29 as=0.29 ps=2.58 w=1 l=0.5
X353 DVSS.t259 a_n227_n10525# a_980_n10861# DVSS.t258 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X354 VDD.t176 a_10013_10507# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X355 a_5555_7857# a_10015_8387# DVSS sky130_fd_pr__res_high_po w=1.41 l=20.1
X356 a_1297_2982.t4 EF_AMUX2to1ISO_0.VO a_4503_2982.t0 VSS.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
D6 DVSS.t108 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X357 a_6371_n10521# a_6271_n10609# DVSS.t8 DVSS.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X358 a_10179_5308# a_10169_4802# DVSS.t1 DVSS.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0.105 pd=1.03 as=0.179 ps=1.26 w=0.75 l=0.5
X359 A1.t6 a_211_n9515.t6 A1.t5 DVSS.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0.58 pd=4.58 as=0 ps=0 w=2 l=0.5
X360 DVSS.t28 a_10039_n11591# a_10464_n11635# DVSS.t27 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.21 ps=1.78 w=1.5 l=0.5
X361 DVSS.t233 a_9771_n10521# a_10978_n10857# DVSS.t232 sky130_fd_pr__nfet_g5v0d10v5 ad=0.122 pd=1.08 as=0.199 ps=2.03 w=0.75 l=0.5
X362 a_1755_6080.t4 a_1355_5983.t9 VDD.t141 VDD.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0.725 pd=5.29 as=0.725 ps=5.29 w=5 l=2
X363 DVSS.t237 a_10180_3343# a_10618_2709# DVSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.398 pd=3.53 as=0.21 ps=1.78 w=1.5 l=0.5
X364 DVSS.t236 a_10180_3343# a_10618_2709# DVSS.t235 sky130_fd_pr__nfet_g5v0d10v5 ad=0.21 pd=1.78 as=0.398 ps=3.53 w=1.5 l=0.5
D7 DVSS.t75 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
R0 a_1297_4914.n93 a_1297_4914.n91 8.86963
R1 a_1297_4914.n90 a_1297_4914.n89 6.31679
R2 a_1297_4914.n0 a_1297_4914.n61 6.12797
R3 a_1297_4914.n7 a_1297_4914.n19 6.12763
R4 a_1297_4914.n36 a_1297_4914.n48 6.12763
R5 a_1297_4914.n21 a_1297_4914.n33 5.96676
R6 a_1297_4914.n62 a_1297_4914.n76 5.63002
R7 a_1297_4914.n80 a_1297_4914.n78 5.63
R8 a_1297_4914.n17 a_1297_4914.t3 5.5395
R9 a_1297_4914.n17 a_1297_4914.t2 5.5395
R10 a_1297_4914.n74 a_1297_4914.t1 5.5395
R11 a_1297_4914.n74 a_1297_4914.t7 5.5395
R12 a_1297_4914.n31 a_1297_4914.t4 5.5395
R13 a_1297_4914.n31 a_1297_4914.t6 5.5395
R14 a_1297_4914.n46 a_1297_4914.t5 5.5395
R15 a_1297_4914.n46 a_1297_4914.t9 5.5395
R16 a_1297_4914.n56 a_1297_4914.t11 5.5395
R17 a_1297_4914.n56 a_1297_4914.t10 5.5395
R18 a_1297_4914.n93 a_1297_4914.t8 5.5395
R19 a_1297_4914.t0 a_1297_4914.n93 5.5395
R20 a_1297_4914.n41 a_1297_4914.n44 4.5005
R21 a_1297_4914.n26 a_1297_4914.n29 4.5005
R22 a_1297_4914.n20 a_1297_4914.n25 4.5005
R23 a_1297_4914.n49 a_1297_4914.n53 4.5005
R24 a_1297_4914.n54 a_1297_4914.n60 4.5005
R25 a_1297_4914.n35 a_1297_4914.n40 4.5005
R26 a_1297_4914.n63 a_1297_4914.n68 4.5005
R27 a_1297_4914.n12 a_1297_4914.n15 4.5005
R28 a_1297_4914.n69 a_1297_4914.n72 4.5005
R29 a_1297_4914.n6 a_1297_4914.n11 4.5005
R30 a_1297_4914.n85 a_1297_4914.n87 4.5005
R31 a_1297_4914.n82 a_1297_4914.n84 4.5005
R32 a_1297_4914.n15 a_1297_4914.n13 3.76521
R33 a_1297_4914.n72 a_1297_4914.n70 3.76521
R34 a_1297_4914.n29 a_1297_4914.n27 3.76521
R35 a_1297_4914.n44 a_1297_4914.n42 3.76521
R36 a_1297_4914.n60 a_1297_4914.n58 3.76521
R37 a_1297_4914.n87 a_1297_4914.n86 3.76521
R38 a_1297_4914.n11 a_1297_4914.n9 3.38874
R39 a_1297_4914.n68 a_1297_4914.n66 3.38874
R40 a_1297_4914.n25 a_1297_4914.n23 3.38874
R41 a_1297_4914.n40 a_1297_4914.n38 3.38874
R42 a_1297_4914.n53 a_1297_4914.n51 3.38874
R43 a_1297_4914.n11 a_1297_4914.n8 3.01226
R44 a_1297_4914.n68 a_1297_4914.n65 3.01226
R45 a_1297_4914.n25 a_1297_4914.n22 3.01226
R46 a_1297_4914.n40 a_1297_4914.n37 3.01226
R47 a_1297_4914.n53 a_1297_4914.n50 3.01226
R48 a_1297_4914.n84 a_1297_4914.n83 3.01226
R49 a_1297_4914.n15 a_1297_4914.n14 2.63579
R50 a_1297_4914.n72 a_1297_4914.n71 2.63579
R51 a_1297_4914.n29 a_1297_4914.n28 2.63579
R52 a_1297_4914.n44 a_1297_4914.n43 2.63579
R53 a_1297_4914.n60 a_1297_4914.n59 2.63579
R54 a_1297_4914.n1 a_1297_4914.n0 2.2019
R55 a_1297_4914.n1 a_1297_4914.n36 1.48434
R56 a_1297_4914.n3 a_1297_4914.n21 1.48434
R57 a_1297_4914.n5 a_1297_4914.n7 1.48434
R58 a_1297_4914.n4 a_1297_4914.n64 1.48434
R59 a_1297_4914.n73 a_1297_4914.n75 1.4669
R60 a_1297_4914.n55 a_1297_4914.n57 1.4669
R61 a_1297_4914.n16 a_1297_4914.n18 1.46689
R62 a_1297_4914.n30 a_1297_4914.n32 1.46689
R63 a_1297_4914.n45 a_1297_4914.n47 1.46689
R64 a_1297_4914.n90 a_1297_4914.n88 1.46687
R65 a_1297_4914.n5 a_1297_4914.n4 0.718062
R66 a_1297_4914.n4 a_1297_4914.n3 0.700686
R67 a_1297_4914.n2 a_1297_4914.n1 0.699908
R68 a_1297_4914.n75 a_1297_4914.n74 0.400769
R69 a_1297_4914.n57 a_1297_4914.n56 0.400769
R70 a_1297_4914.n18 a_1297_4914.n17 0.400768
R71 a_1297_4914.n32 a_1297_4914.n31 0.400768
R72 a_1297_4914.n47 a_1297_4914.n46 0.400768
R73 a_1297_4914.n93 a_1297_4914.n90 0.40076
R74 a_1297_4914.n64 a_1297_4914.n62 0.337583
R75 a_1297_4914.n81 a_1297_4914.n80 0.337269
R76 a_1297_4914.n76 a_1297_4914.n77 0.161367
R77 a_1297_4914.n33 a_1297_4914.n34 0.161367
R78 a_1297_4914.n78 a_1297_4914.n79 0.161367
R79 a_1297_4914.n9 a_1297_4914.n10 0.150167
R80 a_1297_4914.n66 a_1297_4914.n67 0.150167
R81 a_1297_4914.n23 a_1297_4914.n24 0.150167
R82 a_1297_4914.n38 a_1297_4914.n39 0.150167
R83 a_1297_4914.n51 a_1297_4914.n52 0.150167
R84 a_1297_4914.n91 a_1297_4914.n92 0.14967
R85 a_1297_4914.n85 a_1297_4914.n82 0.142861
R86 a_1297_4914.n20 a_1297_4914.n26 0.142861
R87 a_1297_4914.n63 a_1297_4914.n69 0.142861
R88 a_1297_4914.n6 a_1297_4914.n12 0.142841
R89 a_1297_4914.n35 a_1297_4914.n41 0.142841
R90 a_1297_4914.n49 a_1297_4914.n54 0.142841
R91 a_1297_4914.n7 a_1297_4914.n6 0.078121
R92 a_1297_4914.n21 a_1297_4914.n20 0.078121
R93 a_1297_4914.n36 a_1297_4914.n35 0.078121
R94 a_1297_4914.n82 a_1297_4914.n81 0.078121
R95 a_1297_4914.n0 a_1297_4914.n49 0.0777794
R96 a_1297_4914.n64 a_1297_4914.n63 0.0777794
R97 a_1297_4914.n12 a_1297_4914.n16 0.0415156
R98 a_1297_4914.n26 a_1297_4914.n30 0.0415156
R99 a_1297_4914.n41 a_1297_4914.n45 0.0415156
R100 a_1297_4914.n54 a_1297_4914.n55 0.0415156
R101 a_1297_4914.n69 a_1297_4914.n73 0.0415156
R102 a_1297_4914.n88 a_1297_4914.n85 0.0415156
R103 a_1297_4914.n3 a_1297_4914.n2 0.0360311
R104 a_1297_4914.n81 a_1297_4914.n5 2.20191
R105 a_4503_4914.n56 a_4503_4914.t4 60.2505
R106 a_4503_4914.n33 a_4503_4914.t8 60.2505
R107 a_4503_4914.n10 a_4503_4914.t9 60.2505
R108 a_4503_4914.n70 a_4503_4914.t6 60.2505
R109 a_4503_4914.n7 a_4503_4914.n78 9.3005
R110 a_4503_4914.n80 a_4503_4914.n79 9.3005
R111 a_4503_4914.n7 a_4503_4914.n77 9.3005
R112 a_4503_4914.n77 a_4503_4914.n76 9.3005
R113 a_4503_4914.n44 a_4503_4914.n43 9.3005
R114 a_4503_4914.n1 a_4503_4914.n25 9.3005
R115 a_4503_4914.n20 a_4503_4914.n19 9.3005
R116 a_4503_4914.n0 a_4503_4914.n18 9.3005
R117 a_4503_4914.n0 a_4503_4914.n17 9.3005
R118 a_4503_4914.n17 a_4503_4914.n16 9.3005
R119 a_4503_4914.n2 a_4503_4914.n26 9.3005
R120 a_4503_4914.n2 a_4503_4914.n32 9.3005
R121 a_4503_4914.n32 a_4503_4914.n31 9.3005
R122 a_4503_4914.n3 a_4503_4914.n42 9.3005
R123 a_4503_4914.n3 a_4503_4914.n41 9.3005
R124 a_4503_4914.n41 a_4503_4914.n40 9.3005
R125 a_4503_4914.n4 a_4503_4914.n48 9.3005
R126 a_4503_4914.n5 a_4503_4914.n55 9.3005
R127 a_4503_4914.n55 a_4503_4914.n54 9.3005
R128 a_4503_4914.n5 a_4503_4914.n49 9.3005
R129 a_4503_4914.n6 a_4503_4914.n64 9.3005
R130 a_4503_4914.n64 a_4503_4914.n63 9.3005
R131 a_4503_4914.n67 a_4503_4914.n66 9.3005
R132 a_4503_4914.n6 a_4503_4914.n65 9.3005
R133 a_4503_4914.n34 a_4503_4914.n33 8.76429
R134 a_4503_4914.n57 a_4503_4914.n56 8.76429
R135 a_4503_4914.n15 a_4503_4914.n14 8.21641
R136 a_4503_4914.n30 a_4503_4914.n29 8.21641
R137 a_4503_4914.n39 a_4503_4914.n38 8.21641
R138 a_4503_4914.n75 a_4503_4914.n74 8.21641
R139 a_4503_4914.n53 a_4503_4914.n52 8.21641
R140 a_4503_4914.n62 a_4503_4914.n61 8.21641
R141 a_4503_4914.n11 a_4503_4914.n10 6.92242
R142 a_4503_4914.n71 a_4503_4914.n70 6.92012
R143 a_4503_4914.n13 a_4503_4914.n12 5.64756
R144 a_4503_4914.n28 a_4503_4914.n27 5.64756
R145 a_4503_4914.n37 a_4503_4914.n36 5.64756
R146 a_4503_4914.n73 a_4503_4914.n72 5.64756
R147 a_4503_4914.n51 a_4503_4914.n50 5.64756
R148 a_4503_4914.n60 a_4503_4914.n59 5.64756
R149 a_4503_4914.n104 a_4503_4914.t2 5.5395
R150 a_4503_4914.n104 a_4503_4914.t1 5.5395
R151 a_4503_4914.n130 a_4503_4914.t0 5.5395
R152 a_4503_4914.t3 a_4503_4914.n130 5.5395
R153 a_4503_4914.n84 a_4503_4914.n83 5.27461
R154 a_4503_4914.n22 a_4503_4914.n21 4.76425
R155 a_4503_4914.n24 a_4503_4914.n23 4.76425
R156 a_4503_4914.n46 a_4503_4914.n45 4.76425
R157 a_4503_4914.n81 a_4503_4914.n69 4.76425
R158 a_4503_4914.n47 a_4503_4914.n9 4.76425
R159 a_4503_4914.n68 a_4503_4914.n8 4.76425
R160 a_4503_4914.n35 a_4503_4914.n34 4.6505
R161 a_4503_4914.n58 a_4503_4914.n57 4.6505
R162 a_4503_4914.n114 a_4503_4914.n113 4.51815
R163 a_4503_4914.n121 a_4503_4914.n120 4.51815
R164 a_4503_4914.n85 a_4503_4914.n96 6.0005
R165 a_4503_4914.n86 a_4503_4914.n88 4.5005
R166 a_4503_4914.n102 a_4503_4914.n107 4.5005
R167 a_4503_4914.n103 a_4503_4914.n111 4.5005
R168 a_4503_4914.n100 a_4503_4914.n125 4.5005
R169 a_4503_4914.n98 a_4503_4914.n128 4.5005
R170 a_4503_4914.n111 a_4503_4914.n108 4.14168
R171 a_4503_4914.n125 a_4503_4914.n122 4.14168
R172 a_4503_4914.n7 a_4503_4914.n71 3.47756
R173 a_4503_4914.n0 a_4503_4914.n11 3.4767
R174 a_4503_4914.n96 a_4503_4914.n95 3.38238
R175 a_4503_4914.n117 a_4503_4914.t5 3.3065
R176 a_4503_4914.n117 a_4503_4914.t7 3.3065
R177 a_4503_4914.n90 a_4503_4914.n117 3.21134
R178 a_4503_4914.n112 a_4503_4914.n114 3.03311
R179 a_4503_4914.n99 a_4503_4914.n121 3.03311
R180 a_4503_4914.n130 a_4503_4914.n97 2.85325
R181 a_4503_4914.n106 a_4503_4914.n105 2.25932
R182 a_4503_4914.n127 a_4503_4914.n126 2.25932
R183 a_4503_4914.n111 a_4503_4914.n109 2.22452
R184 a_4503_4914.n125 a_4503_4914.n123 2.22452
R185 a_4503_4914.n118 a_4503_4914.n116 2.11721
R186 a_4503_4914.n96 a_4503_4914.n94 1.88285
R187 a_4503_4914.n130 a_4503_4914.n129 1.64452
R188 a_4503_4914.n89 a_4503_4914.n92 6.0005
R189 a_4503_4914.n119 a_4503_4914.n118 1.46063
R190 a_4503_4914.n92 a_4503_4914.n91 1.12991
R191 a_4503_4914.n16 a_4503_4914.n15 1.09595
R192 a_4503_4914.n31 a_4503_4914.n30 1.09595
R193 a_4503_4914.n40 a_4503_4914.n39 1.09595
R194 a_4503_4914.n76 a_4503_4914.n75 1.09595
R195 a_4503_4914.n54 a_4503_4914.n53 1.09595
R196 a_4503_4914.n63 a_4503_4914.n62 1.09595
R197 a_4503_4914.n17 a_4503_4914.n13 0.753441
R198 a_4503_4914.n32 a_4503_4914.n28 0.753441
R199 a_4503_4914.n41 a_4503_4914.n37 0.753441
R200 a_4503_4914.n77 a_4503_4914.n73 0.753441
R201 a_4503_4914.n55 a_4503_4914.n51 0.753441
R202 a_4503_4914.n64 a_4503_4914.n60 0.753441
R203 a_4503_4914.n94 a_4503_4914.n93 0.753441
R204 a_4503_4914.n107 a_4503_4914.n106 0.753441
R205 a_4503_4914.n128 a_4503_4914.n127 0.753441
R206 a_4503_4914.n116 a_4503_4914.n90 0.699656
R207 a_4503_4914.n118 a_4503_4914.n115 0.599941
R208 a_4503_4914.n115 a_4503_4914.n101 0.580288
R209 a_4503_4914.n102 a_4503_4914.n104 2.20064
R210 a_4503_4914.n24 a_4503_4914.n22 0.458354
R211 a_4503_4914.n47 a_4503_4914.n46 0.458354
R212 a_4503_4914.n88 a_4503_4914.n87 0.376971
R213 a_4503_4914.n82 a_4503_4914.n68 0.229427
R214 a_4503_4914.n82 a_4503_4914.n81 0.229427
R215 a_4503_4914.n84 a_4503_4914.n82 0.191391
R216 a_4503_4914.n35 a_4503_4914.n2 0.190717
R217 a_4503_4914.n3 a_4503_4914.n35 0.190717
R218 a_4503_4914.n58 a_4503_4914.n5 0.190717
R219 a_4503_4914.n6 a_4503_4914.n58 0.190717
R220 a_4503_4914.n22 a_4503_4914.n20 0.15935
R221 a_4503_4914.n1 a_4503_4914.n24 0.15935
R222 a_4503_4914.n46 a_4503_4914.n44 0.15935
R223 a_4503_4914.n4 a_4503_4914.n47 0.15935
R224 a_4503_4914.n68 a_4503_4914.n67 0.15935
R225 a_4503_4914.n81 a_4503_4914.n80 0.15935
R226 a_4503_4914.n89 a_4503_4914.n90 0.0960207
R227 a_4503_4914.n103 a_4503_4914.n102 0.0905117
R228 a_4503_4914.n98 a_4503_4914.n100 0.0900826
R229 a_4503_4914.n85 a_4503_4914.n89 0.0765135
R230 a_4503_4914.n86 a_4503_4914.n84 0.125375
R231 a_4503_4914.n99 a_4503_4914.n119 0.0595526
R232 a_4503_4914.n115 a_4503_4914.n112 0.0536977
R233 a_4503_4914.n100 a_4503_4914.n99 0.0454219
R234 a_4503_4914.n112 a_4503_4914.n103 0.0454219
R235 a_4503_4914.n86 a_4503_4914.n85 1.53935
R236 a_4503_4914.n80 a_4503_4914.n7 0.0466957
R237 a_4503_4914.n67 a_4503_4914.n6 0.0466957
R238 a_4503_4914.n5 a_4503_4914.n4 0.0466957
R239 a_4503_4914.n44 a_4503_4914.n3 0.0466957
R240 a_4503_4914.n2 a_4503_4914.n1 0.0466957
R241 a_4503_4914.n20 a_4503_4914.n0 0.0466957
R242 a_4503_4914.n109 a_4503_4914.n110 0.0303633
R243 a_4503_4914.n123 a_4503_4914.n124 0.0303633
R244 a_4503_4914.n129 a_4503_4914.n98 0.557389
R245 VDD.n10976 VDD.n9208 2851.48
R246 VDD.n10984 VDD.n9074 2851.48
R247 VDD.n10979 VDD.n9074 2851.48
R248 VDD.n9208 VDD.n8732 2823.94
R249 VDD.n6924 VDD.n6621 1758.86
R250 VDD.n12419 VDD.n6924 1758.86
R251 VDD.n10210 VDD.n6577 1758.86
R252 VDD.n10210 VDD.n6921 1758.86
R253 VDD.n12693 VDD.n12692 1299.66
R254 VDD.n9970 VDD.t206 840.188
R255 VDD.n9970 VDD.t142 840.188
R256 VDD.n12712 VDD.n12711 784.588
R257 VDD.n9194 VDD.n9193 783.936
R258 VDD.n8570 VDD.n8569 767.823
R259 VDD.n12709 VDD.n6602 737.648
R260 VDD.n8195 VDD.n8086 720.883
R261 VDD.n9191 VDD.n9076 644.766
R262 VDD.n6700 VDD.n6621 609.235
R263 VDD.n10055 VDD.n10054 585
R264 VDD.n10066 VDD.n10065 585
R265 VDD.n10075 VDD.n10074 585
R266 VDD.n10064 VDD.n10063 585
R267 VDD.n10073 VDD.n10025 585
R268 VDD.n10034 VDD.n10032 585
R269 VDD.n10045 VDD.n10039 585
R270 VDD.n10044 VDD.n10043 585
R271 VDD.n10041 VDD.n10038 585
R272 VDD.n10056 VDD.n10028 585
R273 VDD.n10614 VDD.n10613 585
R274 VDD.n10626 VDD.n10625 585
R275 VDD.n10635 VDD.n10634 585
R276 VDD.n10633 VDD.n10144 585
R277 VDD.n10624 VDD.n10586 585
R278 VDD.n10593 VDD.n10591 585
R279 VDD.n10604 VDD.n10598 585
R280 VDD.n10603 VDD.n10602 585
R281 VDD.n10600 VDD.n10597 585
R282 VDD.n10615 VDD.n10588 585
R283 VDD.n10521 VDD.n10520 585
R284 VDD.n10522 VDD.n10515 585
R285 VDD.n10563 VDD.n10501 585
R286 VDD.n10565 VDD.n10564 585
R287 VDD.n10537 VDD.n10534 585
R288 VDD.n10533 VDD.n10503 585
R289 VDD.n10544 VDD.n10543 585
R290 VDD.n10542 VDD.n10541 585
R291 VDD.n10551 VDD.n10550 585
R292 VDD.n10552 VDD.n10535 585
R293 VDD.n9592 VDD.n9584 585
R294 VDD.n9605 VDD.n9583 585
R295 VDD.n9574 VDD.n9573 585
R296 VDD.n9570 VDD.n9569 585
R297 VDD.n9565 VDD.n9564 585
R298 VDD.n9633 VDD.n9632 585
R299 VDD.n9604 VDD.n9603 585
R300 VDD.n9615 VDD.n9614 585
R301 VDD.n9634 VDD.n9561 585
R302 VDD.n9630 VDD.n9629 585
R303 VDD.n9622 VDD.n9621 585
R304 VDD.n9594 VDD.n9593 585
R305 VDD.n10763 VDD.n10701 585
R306 VDD.n10729 VDD.n10726 585
R307 VDD.n10739 VDD.n10738 585
R308 VDD.n10747 VDD.n10715 585
R309 VDD.n10720 VDD.n10719 585
R310 VDD.n10732 VDD.n10731 585
R311 VDD.n10737 VDD.n10725 585
R312 VDD.n10746 VDD.n10745 585
R313 VDD.n10721 VDD.n10714 585
R314 VDD.n10717 VDD.n10710 585
R315 VDD.n10706 VDD.n10702 585
R316 VDD.n10765 VDD.n10764 585
R317 VDD.n8933 VDD.n8928 585
R318 VDD.n8934 VDD.n8933 585
R319 VDD.n9049 VDD.n9048 585
R320 VDD.n9050 VDD.n9049 585
R321 VDD.n9033 VDD.n9032 585
R322 VDD.n9033 VDD.n8795 585
R323 VDD.n8910 VDD.n8909 585
R324 VDD.n8765 VDD.n8763 585
R325 VDD.n8915 VDD.n8914 585
R326 VDD.n8913 VDD.n8888 585
R327 VDD.n8904 VDD.n8903 585
R328 VDD.n8907 VDD.n8891 585
R329 VDD.n9311 VDD.n9310 585
R330 VDD.n9312 VDD.n9311 585
R331 VDD.n10924 VDD.n9328 585
R332 VDD.n9386 VDD.n9385 585
R333 VDD.n9388 VDD.n9361 585
R334 VDD.n9442 VDD.n9441 585
R335 VDD.n9378 VDD.n9362 585
R336 VDD.n9365 VDD.n9364 585
R337 VDD.n9368 VDD.n9367 585
R338 VDD.n9376 VDD.n9375 585
R339 VDD.n9431 VDD.n9396 585
R340 VDD.n9403 VDD.n9401 585
R341 VDD.n9433 VDD.n9432 585
R342 VDD.n9400 VDD.n9397 585
R343 VDD.n9440 VDD.n9439 585
R344 VDD.n10991 VDD.n8731 550.754
R345 VDD.n10963 VDD.n9218 550.754
R346 VDD.n9194 VDD.n9073 479.688
R347 VDD.n10984 VDD.n9073 479.688
R348 VDD.n10989 VDD.n10988 456.74
R349 VDD.n10961 VDD.n10960 456.74
R350 VDD.n6741 VDD.n6714 440.276
R351 VDD.n12679 VDD.n6715 440.276
R352 VDD.n6701 VDD.n6577 427.842
R353 VDD.n12424 VDD.n6906 426.517
R354 VDD.n12452 VDD.n6902 426.517
R355 VDD.n9905 VDD.t207 403.574
R356 VDD.n9904 VDD.t143 403.574
R357 VDD.n6261 VDD.n6258 373.449
R358 VDD.n6289 VDD.n6288 373.449
R359 VDD.n6366 VDD.n6365 373.449
R360 VDD.n6382 VDD.n5903 373.449
R361 VDD.n5407 VDD.n5404 373.449
R362 VDD.n5435 VDD.n5434 373.449
R363 VDD.n5512 VDD.n5511 373.449
R364 VDD.n5528 VDD.n5049 373.449
R365 VDD.n4621 VDD.n4618 373.449
R366 VDD.n4649 VDD.n4648 373.449
R367 VDD.n4726 VDD.n4725 373.449
R368 VDD.n4742 VDD.n4263 373.449
R369 VDD.n3767 VDD.n3764 373.449
R370 VDD.n3795 VDD.n3794 373.449
R371 VDD.n3872 VDD.n3871 373.449
R372 VDD.n3888 VDD.n3409 373.449
R373 VDD.n2981 VDD.n2978 373.449
R374 VDD.n3009 VDD.n3008 373.449
R375 VDD.n3086 VDD.n3085 373.449
R376 VDD.n3102 VDD.n2623 373.449
R377 VDD.n2126 VDD.n2123 373.449
R378 VDD.n2154 VDD.n2153 373.449
R379 VDD.n2231 VDD.n2230 373.449
R380 VDD.n2247 VDD.n1768 373.449
R381 VDD.n10975 VDD.n10974 357.288
R382 VDD.n10983 VDD.n10981 357.288
R383 VDD.n10981 VDD.n10980 357.288
R384 VDD.n10974 VDD.n8734 354.019
R385 VDD.n5959 VDD.n5919 351.829
R386 VDD.n5980 VDD.n5979 351.829
R387 VDD.n6545 VDD.n5793 351.829
R388 VDD.n6525 VDD.n5789 351.829
R389 VDD.n5105 VDD.n5065 351.829
R390 VDD.n5126 VDD.n5125 351.829
R391 VDD.n5691 VDD.n4939 351.829
R392 VDD.n5671 VDD.n4935 351.829
R393 VDD.n4319 VDD.n4279 351.829
R394 VDD.n4340 VDD.n4339 351.829
R395 VDD.n4905 VDD.n4153 351.829
R396 VDD.n4885 VDD.n4149 351.829
R397 VDD.n3465 VDD.n3425 351.829
R398 VDD.n3486 VDD.n3485 351.829
R399 VDD.n4051 VDD.n3299 351.829
R400 VDD.n4031 VDD.n3295 351.829
R401 VDD.n2679 VDD.n2639 351.829
R402 VDD.n2700 VDD.n2699 351.829
R403 VDD.n3265 VDD.n2513 351.829
R404 VDD.n3245 VDD.n2509 351.829
R405 VDD.n1824 VDD.n1784 351.829
R406 VDD.n1845 VDD.n1844 351.829
R407 VDD.n2410 VDD.n1658 351.829
R408 VDD.n2390 VDD.n1654 351.829
R409 VDD.n12694 VDD.n12693 340.084
R410 VDD.n9966 VDD.n9965 321.882
R411 VDD.n9961 VDD.n9909 321.882
R412 VDD.n9944 VDD.n9943 321.882
R413 VDD.n9939 VDD.n9917 321.882
R414 VDD.n9932 VDD.n9919 321.882
R415 VDD.n5761 VDD.n5743 321.882
R416 VDD.n5747 VDD.n5742 321.882
R417 VDD.n5724 VDD.n5716 321.882
R418 VDD.n5737 VDD.n5716 321.882
R419 VDD.n5737 VDD.n5714 321.882
R420 VDD.n5766 VDD.n5714 321.882
R421 VDD.n4121 VDD.n4103 321.882
R422 VDD.n4107 VDD.n4102 321.882
R423 VDD.n4084 VDD.n4076 321.882
R424 VDD.n4097 VDD.n4076 321.882
R425 VDD.n4097 VDD.n4074 321.882
R426 VDD.n4126 VDD.n4074 321.882
R427 VDD.n2481 VDD.n2462 321.882
R428 VDD.n2466 VDD.n2461 321.882
R429 VDD.n2443 VDD.n2435 321.882
R430 VDD.n2456 VDD.n2435 321.882
R431 VDD.n2456 VDD.n2433 321.882
R432 VDD.n2486 VDD.n2433 321.882
R433 VDD.n841 VDD.n822 321.882
R434 VDD.n826 VDD.n821 321.882
R435 VDD.n803 VDD.n795 321.882
R436 VDD.n816 VDD.n795 321.882
R437 VDD.n816 VDD.n793 321.882
R438 VDD.n846 VDD.n793 321.882
R439 VDD.n10428 VDD.n6921 300.546
R440 VDD.n9150 VDD.n9091 292.5
R441 VDD.n10110 VDD.n10099 291.75
R442 VDD.n10110 VDD.n10109 291.562
R443 VDD.n12127 VDD.n7354 271.43
R444 VDD.n11586 VDD.n11585 271.43
R445 VDD.n5765 VDD.n5764 266.731
R446 VDD.n4125 VDD.n4124 266.731
R447 VDD.n2485 VDD.n2484 266.731
R448 VDD.n845 VDD.n844 266.731
R449 VDD.n9178 VDD.n9173 247.893
R450 VDD.n9178 VDD.n8732 247.893
R451 VDD.n2471 VDD.t168 240.534
R452 VDD.n831 VDD.t131 240.534
R453 VDD.n6018 VDD.n5932 239.793
R454 VDD.n6333 VDD.n6018 239.793
R455 VDD.n6026 VDD.n5929 239.793
R456 VDD.n6026 VDD.n6023 239.793
R457 VDD.n6344 VDD.n5937 239.793
R458 VDD.n6300 VDD.n5781 239.793
R459 VDD.n6342 VDD.n5941 239.793
R460 VDD.n6294 VDD.n5785 239.793
R461 VDD.n5164 VDD.n5078 239.793
R462 VDD.n5479 VDD.n5164 239.793
R463 VDD.n5172 VDD.n5075 239.793
R464 VDD.n5172 VDD.n5169 239.793
R465 VDD.n5490 VDD.n5083 239.793
R466 VDD.n5446 VDD.n4927 239.793
R467 VDD.n5488 VDD.n5087 239.793
R468 VDD.n5440 VDD.n4931 239.793
R469 VDD.n4378 VDD.n4292 239.793
R470 VDD.n4693 VDD.n4378 239.793
R471 VDD.n4386 VDD.n4289 239.793
R472 VDD.n4386 VDD.n4383 239.793
R473 VDD.n4704 VDD.n4297 239.793
R474 VDD.n4660 VDD.n4141 239.793
R475 VDD.n4702 VDD.n4301 239.793
R476 VDD.n4654 VDD.n4145 239.793
R477 VDD.n3524 VDD.n3438 239.793
R478 VDD.n3839 VDD.n3524 239.793
R479 VDD.n3532 VDD.n3435 239.793
R480 VDD.n3532 VDD.n3529 239.793
R481 VDD.n3850 VDD.n3443 239.793
R482 VDD.n3806 VDD.n3287 239.793
R483 VDD.n3848 VDD.n3447 239.793
R484 VDD.n3800 VDD.n3291 239.793
R485 VDD.n2738 VDD.n2652 239.793
R486 VDD.n3053 VDD.n2738 239.793
R487 VDD.n2746 VDD.n2649 239.793
R488 VDD.n2746 VDD.n2743 239.793
R489 VDD.n3064 VDD.n2657 239.793
R490 VDD.n3020 VDD.n2501 239.793
R491 VDD.n3062 VDD.n2661 239.793
R492 VDD.n3014 VDD.n2505 239.793
R493 VDD.n1883 VDD.n1797 239.793
R494 VDD.n2198 VDD.n1883 239.793
R495 VDD.n1891 VDD.n1794 239.793
R496 VDD.n1891 VDD.n1888 239.793
R497 VDD.n2209 VDD.n1802 239.793
R498 VDD.n2165 VDD.n1646 239.793
R499 VDD.n2207 VDD.n1806 239.793
R500 VDD.n2159 VDD.n1650 239.793
R501 VDD.n4114 VDD.t84 239.755
R502 VDD.n5754 VDD.t22 239.697
R503 VDD.n9955 VDD.t129 237.577
R504 VDD.n9941 VDD.t208 233.279
R505 VDD.n8500 VDD.n7809 232.623
R506 VDD.n9061 VDD.n9060 231.905
R507 VDD.n10076 VDD.n10024 229.476
R508 VDD.n10636 VDD.n10143 229.476
R509 VDD.n10529 VDD.n10528 229.476
R510 VDD.n9423 VDD.n9422 228.99
R511 VDD.n12713 VDD.n12712 228
R512 VDD.n8574 VDD.n8573 228
R513 VDD.n8578 VDD.n8577 228
R514 VDD.n8582 VDD.n8581 228
R515 VDD.n8584 VDD.n7760 228
R516 VDD.n8588 VDD.n7753 228
R517 VDD.n8592 VDD.n7750 228
R518 VDD.n8597 VDD.n7750 228
R519 VDD.n8597 VDD.n7751 228
R520 VDD.n7751 VDD.n7730 228
R521 VDD.n11440 VDD.n7730 228
R522 VDD.n11440 VDD.n7731 228
R523 VDD.n11436 VDD.n7731 228
R524 VDD.n11436 VDD.n7734 228
R525 VDD.n8618 VDD.n7734 228
R526 VDD.n11421 VDD.n8618 228
R527 VDD.n11421 VDD.n8624 228
R528 VDD.n11417 VDD.n8624 228
R529 VDD.n11417 VDD.n8627 228
R530 VDD.n8649 VDD.n8627 228
R531 VDD.n11402 VDD.n8649 228
R532 VDD.n11402 VDD.n8655 228
R533 VDD.n11398 VDD.n8655 228
R534 VDD.n11398 VDD.n8658 228
R535 VDD.n8670 VDD.n8658 228
R536 VDD.n8695 VDD.n8670 228
R537 VDD.n8695 VDD.n8687 228
R538 VDD.n11377 VDD.n8687 228
R539 VDD.n11377 VDD.n8693 228
R540 VDD.n11373 VDD.n8693 228
R541 VDD.n11373 VDD.n8699 228
R542 VDD.n8722 VDD.n8699 228
R543 VDD.n11358 VDD.n8722 228
R544 VDD.n11358 VDD.n11029 228
R545 VDD.n11354 VDD.n11029 228
R546 VDD.n11354 VDD.n11032 228
R547 VDD.n11054 VDD.n11032 228
R548 VDD.n11339 VDD.n11054 228
R549 VDD.n11339 VDD.n11059 228
R550 VDD.n11335 VDD.n11059 228
R551 VDD.n11335 VDD.n11062 228
R552 VDD.n11324 VDD.n11062 228
R553 VDD.n11324 VDD.n11077 228
R554 VDD.n11320 VDD.n11077 228
R555 VDD.n11320 VDD.n11079 228
R556 VDD.n11107 VDD.n11079 228
R557 VDD.n11305 VDD.n11107 228
R558 VDD.n11305 VDD.n11113 228
R559 VDD.n11301 VDD.n11113 228
R560 VDD.n11301 VDD.n11116 228
R561 VDD.n11137 VDD.n11116 228
R562 VDD.n11286 VDD.n11137 228
R563 VDD.n11286 VDD.n11144 228
R564 VDD.n11282 VDD.n11144 228
R565 VDD.n11282 VDD.n11147 228
R566 VDD.n11169 VDD.n11147 228
R567 VDD.n11267 VDD.n11169 228
R568 VDD.n11267 VDD.n11175 228
R569 VDD.n11263 VDD.n11175 228
R570 VDD.n11263 VDD.n11178 228
R571 VDD.n11191 VDD.n11178 228
R572 VDD.n11236 VDD.n11191 228
R573 VDD.n11236 VDD.n11208 228
R574 VDD.n11242 VDD.n11208 228
R575 VDD.n11242 VDD.n11234 228
R576 VDD.n11234 VDD.n6597 228
R577 VDD.n12711 VDD.n6597 228
R578 VDD.n8204 VDD.n8086 228
R579 VDD.n8204 VDD.n8077 228
R580 VDD.n8215 VDD.n8077 228
R581 VDD.n8216 VDD.n8215 228
R582 VDD.n8216 VDD.n8071 228
R583 VDD.n8228 VDD.n8071 228
R584 VDD.n8228 VDD.n8064 228
R585 VDD.n8236 VDD.n8064 228
R586 VDD.n8236 VDD.n8058 228
R587 VDD.n8248 VDD.n8058 228
R588 VDD.n8248 VDD.n8049 228
R589 VDD.n8259 VDD.n8049 228
R590 VDD.n8260 VDD.n8259 228
R591 VDD.n8260 VDD.n8043 228
R592 VDD.n8272 VDD.n8043 228
R593 VDD.n8272 VDD.n8036 228
R594 VDD.n8280 VDD.n8036 228
R595 VDD.n8280 VDD.n8026 228
R596 VDD.n8290 VDD.n8026 228
R597 VDD.n8291 VDD.n8290 228
R598 VDD.n8291 VDD.n8020 228
R599 VDD.n8303 VDD.n8020 228
R600 VDD.n8303 VDD.n8013 228
R601 VDD.n8311 VDD.n8013 228
R602 VDD.n8311 VDD.n8007 228
R603 VDD.n8323 VDD.n8007 228
R604 VDD.n8323 VDD.n7998 228
R605 VDD.n8335 VDD.n7998 228
R606 VDD.n8336 VDD.n8335 228
R607 VDD.n8337 VDD.n8336 228
R608 VDD.n8489 VDD.n8337 228
R609 VDD.n8489 VDD.n8338 228
R610 VDD.n8482 VDD.n8338 228
R611 VDD.n8482 VDD.n8346 228
R612 VDD.n8474 VDD.n8346 228
R613 VDD.n8474 VDD.n8353 228
R614 VDD.n8467 VDD.n8353 228
R615 VDD.n8467 VDD.n8363 228
R616 VDD.n8460 VDD.n8363 228
R617 VDD.n8460 VDD.n8369 228
R618 VDD.n8453 VDD.n8369 228
R619 VDD.n8453 VDD.n8379 228
R620 VDD.n8445 VDD.n8379 228
R621 VDD.n8445 VDD.n8386 228
R622 VDD.n8438 VDD.n8386 228
R623 VDD.n8438 VDD.n8396 228
R624 VDD.n8430 VDD.n8396 228
R625 VDD.n8430 VDD.n8403 228
R626 VDD.n8423 VDD.n8403 228
R627 VDD.n8423 VDD.n7762 228
R628 VDD.n8569 VDD.n7762 228
R629 VDD.n8150 VDD.n7746 228
R630 VDD.n8599 VDD.n7746 228
R631 VDD.n8599 VDD.n7724 228
R632 VDD.n11443 VDD.n7724 228
R633 VDD.n11443 VDD.n11442 228
R634 VDD.n11442 VDD.n7725 228
R635 VDD.n11434 VDD.n7725 228
R636 VDD.n11434 VDD.n7737 228
R637 VDD.n11424 VDD.n7737 228
R638 VDD.n11424 VDD.n11423 228
R639 VDD.n11423 VDD.n8619 228
R640 VDD.n11415 VDD.n8619 228
R641 VDD.n11415 VDD.n8631 228
R642 VDD.n11405 VDD.n8631 228
R643 VDD.n11405 VDD.n11404 228
R644 VDD.n11404 VDD.n8650 228
R645 VDD.n11396 VDD.n8650 228
R646 VDD.n11396 VDD.n8661 228
R647 VDD.n11389 VDD.n8661 228
R648 VDD.n11389 VDD.n8671 228
R649 VDD.n11380 VDD.n8671 228
R650 VDD.n11380 VDD.n11379 228
R651 VDD.n11379 VDD.n8688 228
R652 VDD.n11371 VDD.n8688 228
R653 VDD.n11371 VDD.n8703 228
R654 VDD.n11361 VDD.n8703 228
R655 VDD.n11361 VDD.n11360 228
R656 VDD.n11360 VDD.n8723 228
R657 VDD.n11352 VDD.n8723 228
R658 VDD.n11352 VDD.n11036 228
R659 VDD.n11342 VDD.n11036 228
R660 VDD.n11342 VDD.n11341 228
R661 VDD.n11341 VDD.n11055 228
R662 VDD.n11333 VDD.n11055 228
R663 VDD.n11333 VDD.n11065 228
R664 VDD.n11326 VDD.n11065 228
R665 VDD.n11326 VDD.n11073 228
R666 VDD.n11318 VDD.n11073 228
R667 VDD.n11318 VDD.n11083 228
R668 VDD.n11308 VDD.n11083 228
R669 VDD.n11308 VDD.n11307 228
R670 VDD.n11307 VDD.n11108 228
R671 VDD.n11299 VDD.n11108 228
R672 VDD.n11299 VDD.n11120 228
R673 VDD.n11289 VDD.n11120 228
R674 VDD.n11289 VDD.n11288 228
R675 VDD.n11288 VDD.n11138 228
R676 VDD.n11280 VDD.n11138 228
R677 VDD.n11280 VDD.n11151 228
R678 VDD.n11270 VDD.n11151 228
R679 VDD.n11270 VDD.n11269 228
R680 VDD.n11269 VDD.n11170 228
R681 VDD.n11261 VDD.n11170 228
R682 VDD.n11261 VDD.n11182 228
R683 VDD.n11254 VDD.n11182 228
R684 VDD.n11254 VDD.n11192 228
R685 VDD.n11245 VDD.n11192 228
R686 VDD.n11245 VDD.n11244 228
R687 VDD.n11244 VDD.n11209 228
R688 VDD.n11209 VDD.n6601 228
R689 VDD.n12709 VDD.n6601 228
R690 VDD.n10427 VDD.n6576 220.383
R691 VDD.n6938 VDD.n6932 218.608
R692 VDD.n5937 VDD.n5936 218.173
R693 VDD.n6554 VDD.n5781 218.173
R694 VDD.n5985 VDD.n5941 218.173
R695 VDD.n6552 VDD.n5785 218.173
R696 VDD.n5083 VDD.n5082 218.173
R697 VDD.n5700 VDD.n4927 218.173
R698 VDD.n5131 VDD.n5087 218.173
R699 VDD.n5698 VDD.n4931 218.173
R700 VDD.n4297 VDD.n4296 218.173
R701 VDD.n4914 VDD.n4141 218.173
R702 VDD.n4345 VDD.n4301 218.173
R703 VDD.n4912 VDD.n4145 218.173
R704 VDD.n3443 VDD.n3442 218.173
R705 VDD.n4060 VDD.n3287 218.173
R706 VDD.n3491 VDD.n3447 218.173
R707 VDD.n4058 VDD.n3291 218.173
R708 VDD.n2657 VDD.n2656 218.173
R709 VDD.n3274 VDD.n2501 218.173
R710 VDD.n2705 VDD.n2661 218.173
R711 VDD.n3272 VDD.n2505 218.173
R712 VDD.n1802 VDD.n1801 218.173
R713 VDD.n2419 VDD.n1646 218.173
R714 VDD.n1850 VDD.n1806 218.173
R715 VDD.n2417 VDD.n1650 218.173
R716 VDD.n9963 VDD.t128 217.947
R717 VDD.n5763 VDD.t21 217.947
R718 VDD.n4123 VDD.t83 217.947
R719 VDD.n2483 VDD.t167 217.947
R720 VDD.n843 VDD.t130 217.947
R721 VDD.n12771 VDD.n6576 213.983
R722 VDD.n12326 VDD.n12325 205.079
R723 VDD.n12325 VDD.n7002 205.079
R724 VDD.n12316 VDD.n7002 205.079
R725 VDD.n12316 VDD.n12315 205.079
R726 VDD.n12315 VDD.n12314 205.079
R727 VDD.n12314 VDD.n7011 205.079
R728 VDD.n7021 VDD.n7011 205.079
R729 VDD.n12304 VDD.n7021 205.079
R730 VDD.n12304 VDD.n12303 205.079
R731 VDD.n12303 VDD.n12302 205.079
R732 VDD.n12302 VDD.n7022 205.079
R733 VDD.n12293 VDD.n7022 205.079
R734 VDD.n12293 VDD.n12292 205.079
R735 VDD.n12292 VDD.n12291 205.079
R736 VDD.n12291 VDD.n7031 205.079
R737 VDD.n12282 VDD.n7031 205.079
R738 VDD.n12282 VDD.n12281 205.079
R739 VDD.n12281 VDD.n12280 205.079
R740 VDD.n12280 VDD.n7040 205.079
R741 VDD.n12271 VDD.n7040 205.079
R742 VDD.n12271 VDD.n12270 205.079
R743 VDD.n12270 VDD.n12269 205.079
R744 VDD.n12269 VDD.n7049 205.079
R745 VDD.n7060 VDD.n7049 205.079
R746 VDD.n12260 VDD.n7060 205.079
R747 VDD.n12260 VDD.n12259 205.079
R748 VDD.n12259 VDD.n12258 205.079
R749 VDD.n12258 VDD.n7061 205.079
R750 VDD.n12249 VDD.n7061 205.079
R751 VDD.n12247 VDD.n7072 205.079
R752 VDD.n12238 VDD.n7072 205.079
R753 VDD.n12238 VDD.n12237 205.079
R754 VDD.n12237 VDD.n12236 205.079
R755 VDD.n12236 VDD.n7262 205.079
R756 VDD.n7273 VDD.n7262 205.079
R757 VDD.n12227 VDD.n7273 205.079
R758 VDD.n12227 VDD.n12226 205.079
R759 VDD.n12226 VDD.n12225 205.079
R760 VDD.n12225 VDD.n7274 205.079
R761 VDD.n12216 VDD.n7274 205.079
R762 VDD.n12216 VDD.n12215 205.079
R763 VDD.n12215 VDD.n12214 205.079
R764 VDD.n12214 VDD.n7283 205.079
R765 VDD.n12205 VDD.n7283 205.079
R766 VDD.n12205 VDD.n12204 205.079
R767 VDD.n12204 VDD.n12203 205.079
R768 VDD.n12203 VDD.n7292 205.079
R769 VDD.n12194 VDD.n7292 205.079
R770 VDD.n12194 VDD.n12193 205.079
R771 VDD.n12193 VDD.n12192 205.079
R772 VDD.n12192 VDD.n7301 205.079
R773 VDD.n12183 VDD.n7301 205.079
R774 VDD.n12183 VDD.n12182 205.079
R775 VDD.n12182 VDD.n12181 205.079
R776 VDD.n12181 VDD.n7310 205.079
R777 VDD.n12172 VDD.n7310 205.079
R778 VDD.n12172 VDD.n12171 205.079
R779 VDD.n12171 VDD.n12170 205.079
R780 VDD.n12170 VDD.n7317 205.079
R781 VDD.n12161 VDD.n7317 205.079
R782 VDD.n12161 VDD.n12160 205.079
R783 VDD.n12160 VDD.n12159 205.079
R784 VDD.n12159 VDD.n7326 205.079
R785 VDD.n12150 VDD.n7326 205.079
R786 VDD.n12150 VDD.n12149 205.079
R787 VDD.n12149 VDD.n12148 205.079
R788 VDD.n12148 VDD.n7335 205.079
R789 VDD.n12139 VDD.n7335 205.079
R790 VDD.n12139 VDD.n12138 205.079
R791 VDD.n12138 VDD.n12137 205.079
R792 VDD.n12137 VDD.n7344 205.079
R793 VDD.n7354 VDD.n7344 205.079
R794 VDD.n12127 VDD.n12126 205.079
R795 VDD.n12126 VDD.n12125 205.079
R796 VDD.n12125 VDD.n7355 205.079
R797 VDD.n12119 VDD.n7355 205.079
R798 VDD.n12119 VDD.n12118 205.079
R799 VDD.n12118 VDD.n12117 205.079
R800 VDD.n12117 VDD.n7359 205.079
R801 VDD.n12111 VDD.n7359 205.079
R802 VDD.n12111 VDD.n12110 205.079
R803 VDD.n12110 VDD.n12109 205.079
R804 VDD.n12109 VDD.n7363 205.079
R805 VDD.n12103 VDD.n7363 205.079
R806 VDD.n12103 VDD.n12102 205.079
R807 VDD.n12102 VDD.n12101 205.079
R808 VDD.n12101 VDD.n7367 205.079
R809 VDD.n12095 VDD.n7367 205.079
R810 VDD.n12095 VDD.n12094 205.079
R811 VDD.n11651 VDD.n11650 205.079
R812 VDD.n11652 VDD.n11651 205.079
R813 VDD.n11652 VDD.n7604 205.079
R814 VDD.n11663 VDD.n7604 205.079
R815 VDD.n11664 VDD.n11663 205.079
R816 VDD.n11665 VDD.n11664 205.079
R817 VDD.n11665 VDD.n7598 205.079
R818 VDD.n11675 VDD.n7598 205.079
R819 VDD.n11676 VDD.n11675 205.079
R820 VDD.n11677 VDD.n11676 205.079
R821 VDD.n11677 VDD.n7590 205.079
R822 VDD.n11687 VDD.n7590 205.079
R823 VDD.n11688 VDD.n11687 205.079
R824 VDD.n11689 VDD.n11688 205.079
R825 VDD.n11689 VDD.n7583 205.079
R826 VDD.n11700 VDD.n7583 205.079
R827 VDD.n11701 VDD.n11700 205.079
R828 VDD.n11702 VDD.n11701 205.079
R829 VDD.n11702 VDD.n7576 205.079
R830 VDD.n11713 VDD.n7576 205.079
R831 VDD.n11714 VDD.n11713 205.079
R832 VDD.n11715 VDD.n11714 205.079
R833 VDD.n11715 VDD.n7569 205.079
R834 VDD.n11726 VDD.n7569 205.079
R835 VDD.n11727 VDD.n11726 205.079
R836 VDD.n11728 VDD.n11727 205.079
R837 VDD.n11728 VDD.n7563 205.079
R838 VDD.n11738 VDD.n7563 205.079
R839 VDD.n11739 VDD.n11738 205.079
R840 VDD.n11740 VDD.n11739 205.079
R841 VDD.n11740 VDD.n7556 205.079
R842 VDD.n11751 VDD.n7556 205.079
R843 VDD.n11752 VDD.n11751 205.079
R844 VDD.n11753 VDD.n11752 205.079
R845 VDD.n11753 VDD.n7549 205.079
R846 VDD.n11764 VDD.n7549 205.079
R847 VDD.n11765 VDD.n11764 205.079
R848 VDD.n11766 VDD.n11765 205.079
R849 VDD.n11766 VDD.n7542 205.079
R850 VDD.n11777 VDD.n7542 205.079
R851 VDD.n11778 VDD.n11777 205.079
R852 VDD.n11779 VDD.n11778 205.079
R853 VDD.n11779 VDD.n7536 205.079
R854 VDD.n11789 VDD.n7536 205.079
R855 VDD.n11790 VDD.n11789 205.079
R856 VDD.n11791 VDD.n11790 205.079
R857 VDD.n11791 VDD.n7528 205.079
R858 VDD.n11801 VDD.n7528 205.079
R859 VDD.n11802 VDD.n11801 205.079
R860 VDD.n11803 VDD.n11802 205.079
R861 VDD.n11803 VDD.n7521 205.079
R862 VDD.n11814 VDD.n7521 205.079
R863 VDD.n11815 VDD.n11814 205.079
R864 VDD.n11816 VDD.n11815 205.079
R865 VDD.n11816 VDD.n7514 205.079
R866 VDD.n11827 VDD.n7514 205.079
R867 VDD.n11828 VDD.n11827 205.079
R868 VDD.n11829 VDD.n11828 205.079
R869 VDD.n11829 VDD.n7507 205.079
R870 VDD.n11840 VDD.n7507 205.079
R871 VDD.n11841 VDD.n11840 205.079
R872 VDD.n11842 VDD.n11841 205.079
R873 VDD.n11842 VDD.n7501 205.079
R874 VDD.n11852 VDD.n7501 205.079
R875 VDD.n11853 VDD.n11852 205.079
R876 VDD.n11854 VDD.n11853 205.079
R877 VDD.n11854 VDD.n7494 205.079
R878 VDD.n11865 VDD.n7494 205.079
R879 VDD.n11866 VDD.n11865 205.079
R880 VDD.n11867 VDD.n11866 205.079
R881 VDD.n11867 VDD.n7487 205.079
R882 VDD.n11878 VDD.n7487 205.079
R883 VDD.n11879 VDD.n11878 205.079
R884 VDD.n11880 VDD.n11879 205.079
R885 VDD.n11880 VDD.n7480 205.079
R886 VDD.n11891 VDD.n7480 205.079
R887 VDD.n11892 VDD.n11891 205.079
R888 VDD.n11893 VDD.n11892 205.079
R889 VDD.n11893 VDD.n7474 205.079
R890 VDD.n11903 VDD.n7474 205.079
R891 VDD.n11904 VDD.n11903 205.079
R892 VDD.n11905 VDD.n11904 205.079
R893 VDD.n11905 VDD.n7466 205.079
R894 VDD.n11915 VDD.n7466 205.079
R895 VDD.n11916 VDD.n11915 205.079
R896 VDD.n11917 VDD.n11916 205.079
R897 VDD.n11917 VDD.n7459 205.079
R898 VDD.n11928 VDD.n7459 205.079
R899 VDD.n11929 VDD.n11928 205.079
R900 VDD.n11930 VDD.n11929 205.079
R901 VDD.n11930 VDD.n7452 205.079
R902 VDD.n11941 VDD.n7452 205.079
R903 VDD.n11942 VDD.n11941 205.079
R904 VDD.n11943 VDD.n11942 205.079
R905 VDD.n11943 VDD.n7445 205.079
R906 VDD.n11954 VDD.n7445 205.079
R907 VDD.n11955 VDD.n11954 205.079
R908 VDD.n11956 VDD.n11955 205.079
R909 VDD.n11956 VDD.n7439 205.079
R910 VDD.n11966 VDD.n7439 205.079
R911 VDD.n11967 VDD.n11966 205.079
R912 VDD.n11968 VDD.n11967 205.079
R913 VDD.n11968 VDD.n7432 205.079
R914 VDD.n11979 VDD.n7432 205.079
R915 VDD.n11980 VDD.n11979 205.079
R916 VDD.n11981 VDD.n11980 205.079
R917 VDD.n11981 VDD.n7425 205.079
R918 VDD.n11992 VDD.n7425 205.079
R919 VDD.n11993 VDD.n11992 205.079
R920 VDD.n11994 VDD.n11993 205.079
R921 VDD.n11994 VDD.n7418 205.079
R922 VDD.n12005 VDD.n7418 205.079
R923 VDD.n12006 VDD.n12005 205.079
R924 VDD.n12007 VDD.n12006 205.079
R925 VDD.n12007 VDD.n7412 205.079
R926 VDD.n12017 VDD.n7412 205.079
R927 VDD.n12018 VDD.n12017 205.079
R928 VDD.n12019 VDD.n12018 205.079
R929 VDD.n12019 VDD.n7404 205.079
R930 VDD.n12029 VDD.n7404 205.079
R931 VDD.n12030 VDD.n12029 205.079
R932 VDD.n12031 VDD.n12030 205.079
R933 VDD.n12031 VDD.n7397 205.079
R934 VDD.n12042 VDD.n7397 205.079
R935 VDD.n12043 VDD.n12042 205.079
R936 VDD.n12044 VDD.n12043 205.079
R937 VDD.n12044 VDD.n7390 205.079
R938 VDD.n12055 VDD.n7390 205.079
R939 VDD.n12056 VDD.n12055 205.079
R940 VDD.n12057 VDD.n12056 205.079
R941 VDD.n12057 VDD.n7383 205.079
R942 VDD.n12068 VDD.n7383 205.079
R943 VDD.n12069 VDD.n12068 205.079
R944 VDD.n12070 VDD.n12069 205.079
R945 VDD.n12070 VDD.n7377 205.079
R946 VDD.n12083 VDD.n7377 205.079
R947 VDD.n12084 VDD.n12083 205.079
R948 VDD.n12085 VDD.n12084 205.079
R949 VDD.n12085 VDD.n7371 205.079
R950 VDD.n11450 VDD.n11449 205.079
R951 VDD.n11450 VDD.n7711 205.079
R952 VDD.n11461 VDD.n7711 205.079
R953 VDD.n11462 VDD.n11461 205.079
R954 VDD.n11463 VDD.n11462 205.079
R955 VDD.n11463 VDD.n7705 205.079
R956 VDD.n11473 VDD.n7705 205.079
R957 VDD.n11474 VDD.n11473 205.079
R958 VDD.n11475 VDD.n11474 205.079
R959 VDD.n11475 VDD.n7698 205.079
R960 VDD.n11485 VDD.n7698 205.079
R961 VDD.n11486 VDD.n11485 205.079
R962 VDD.n11487 VDD.n11486 205.079
R963 VDD.n11487 VDD.n7691 205.079
R964 VDD.n11498 VDD.n7691 205.079
R965 VDD.n11499 VDD.n11498 205.079
R966 VDD.n11500 VDD.n11499 205.079
R967 VDD.n11500 VDD.n7684 205.079
R968 VDD.n11511 VDD.n7684 205.079
R969 VDD.n11512 VDD.n11511 205.079
R970 VDD.n11513 VDD.n11512 205.079
R971 VDD.n11513 VDD.n7677 205.079
R972 VDD.n11524 VDD.n7677 205.079
R973 VDD.n11525 VDD.n11524 205.079
R974 VDD.n11526 VDD.n11525 205.079
R975 VDD.n11526 VDD.n7670 205.079
R976 VDD.n11534 VDD.n7670 205.079
R977 VDD.n11535 VDD.n11534 205.079
R978 VDD.n11536 VDD.n11535 205.079
R979 VDD.n11536 VDD.n7663 205.079
R980 VDD.n11547 VDD.n7663 205.079
R981 VDD.n11548 VDD.n11547 205.079
R982 VDD.n11549 VDD.n11548 205.079
R983 VDD.n11549 VDD.n7656 205.079
R984 VDD.n11560 VDD.n7656 205.079
R985 VDD.n11561 VDD.n11560 205.079
R986 VDD.n11562 VDD.n11561 205.079
R987 VDD.n11562 VDD.n7649 205.079
R988 VDD.n11573 VDD.n7649 205.079
R989 VDD.n11574 VDD.n11573 205.079
R990 VDD.n11575 VDD.n11574 205.079
R991 VDD.n11575 VDD.n7643 205.079
R992 VDD.n11585 VDD.n7643 205.079
R993 VDD.n11587 VDD.n11586 205.079
R994 VDD.n11587 VDD.n7636 205.079
R995 VDD.n11598 VDD.n7636 205.079
R996 VDD.n11599 VDD.n11598 205.079
R997 VDD.n11600 VDD.n11599 205.079
R998 VDD.n11600 VDD.n7629 205.079
R999 VDD.n11611 VDD.n7629 205.079
R1000 VDD.n11612 VDD.n11611 205.079
R1001 VDD.n11613 VDD.n11612 205.079
R1002 VDD.n11613 VDD.n7622 205.079
R1003 VDD.n11624 VDD.n7622 205.079
R1004 VDD.n11625 VDD.n11624 205.079
R1005 VDD.n11626 VDD.n11625 205.079
R1006 VDD.n11626 VDD.n7615 205.079
R1007 VDD.n11639 VDD.n7615 205.079
R1008 VDD.n11640 VDD.n11639 205.079
R1009 VDD.n11641 VDD.n11640 205.079
R1010 VDD.n6224 VDD.n6223 205.079
R1011 VDD.n6224 VDD.n6067 205.079
R1012 VDD.n6230 VDD.n6067 205.079
R1013 VDD.n6231 VDD.n6230 205.079
R1014 VDD.n6232 VDD.n6231 205.079
R1015 VDD.n6232 VDD.n6063 205.079
R1016 VDD.n6238 VDD.n6063 205.079
R1017 VDD.n6239 VDD.n6238 205.079
R1018 VDD.n6240 VDD.n6239 205.079
R1019 VDD.n6240 VDD.n6059 205.079
R1020 VDD.n6247 VDD.n6059 205.079
R1021 VDD.n6248 VDD.n6247 205.079
R1022 VDD.n6250 VDD.n6248 205.079
R1023 VDD.n6145 VDD.n6112 205.079
R1024 VDD.n6145 VDD.n6144 205.079
R1025 VDD.n6144 VDD.n6143 205.079
R1026 VDD.n6143 VDD.n6113 205.079
R1027 VDD.n6137 VDD.n6113 205.079
R1028 VDD.n6137 VDD.n6136 205.079
R1029 VDD.n6136 VDD.n6135 205.079
R1030 VDD.n6135 VDD.n6117 205.079
R1031 VDD.n6129 VDD.n6117 205.079
R1032 VDD.n6129 VDD.n6128 205.079
R1033 VDD.n6128 VDD.n6127 205.079
R1034 VDD.n6127 VDD.n6122 205.079
R1035 VDD.n6122 VDD.n6121 205.079
R1036 VDD.n6513 VDD.n5813 205.079
R1037 VDD.n6513 VDD.n6512 205.079
R1038 VDD.n6512 VDD.n6511 205.079
R1039 VDD.n6511 VDD.n5814 205.079
R1040 VDD.n6505 VDD.n5814 205.079
R1041 VDD.n6505 VDD.n6504 205.079
R1042 VDD.n6504 VDD.n6503 205.079
R1043 VDD.n6503 VDD.n5818 205.079
R1044 VDD.n6497 VDD.n5818 205.079
R1045 VDD.n6497 VDD.n6496 205.079
R1046 VDD.n6496 VDD.n6495 205.079
R1047 VDD.n6495 VDD.n5822 205.079
R1048 VDD.n6489 VDD.n5822 205.079
R1049 VDD.n6398 VDD.n5875 205.079
R1050 VDD.n6399 VDD.n6398 205.079
R1051 VDD.n6400 VDD.n6399 205.079
R1052 VDD.n6400 VDD.n5871 205.079
R1053 VDD.n6406 VDD.n5871 205.079
R1054 VDD.n6407 VDD.n6406 205.079
R1055 VDD.n6408 VDD.n6407 205.079
R1056 VDD.n6408 VDD.n5867 205.079
R1057 VDD.n6414 VDD.n5867 205.079
R1058 VDD.n6415 VDD.n6414 205.079
R1059 VDD.n6416 VDD.n6415 205.079
R1060 VDD.n6416 VDD.n5862 205.079
R1061 VDD.n6423 VDD.n5862 205.079
R1062 VDD.n5370 VDD.n5369 205.079
R1063 VDD.n5370 VDD.n5213 205.079
R1064 VDD.n5376 VDD.n5213 205.079
R1065 VDD.n5377 VDD.n5376 205.079
R1066 VDD.n5378 VDD.n5377 205.079
R1067 VDD.n5378 VDD.n5209 205.079
R1068 VDD.n5384 VDD.n5209 205.079
R1069 VDD.n5385 VDD.n5384 205.079
R1070 VDD.n5386 VDD.n5385 205.079
R1071 VDD.n5386 VDD.n5205 205.079
R1072 VDD.n5393 VDD.n5205 205.079
R1073 VDD.n5394 VDD.n5393 205.079
R1074 VDD.n5396 VDD.n5394 205.079
R1075 VDD.n5291 VDD.n5258 205.079
R1076 VDD.n5291 VDD.n5290 205.079
R1077 VDD.n5290 VDD.n5289 205.079
R1078 VDD.n5289 VDD.n5259 205.079
R1079 VDD.n5283 VDD.n5259 205.079
R1080 VDD.n5283 VDD.n5282 205.079
R1081 VDD.n5282 VDD.n5281 205.079
R1082 VDD.n5281 VDD.n5263 205.079
R1083 VDD.n5275 VDD.n5263 205.079
R1084 VDD.n5275 VDD.n5274 205.079
R1085 VDD.n5274 VDD.n5273 205.079
R1086 VDD.n5273 VDD.n5268 205.079
R1087 VDD.n5268 VDD.n5267 205.079
R1088 VDD.n5659 VDD.n4959 205.079
R1089 VDD.n5659 VDD.n5658 205.079
R1090 VDD.n5658 VDD.n5657 205.079
R1091 VDD.n5657 VDD.n4960 205.079
R1092 VDD.n5651 VDD.n4960 205.079
R1093 VDD.n5651 VDD.n5650 205.079
R1094 VDD.n5650 VDD.n5649 205.079
R1095 VDD.n5649 VDD.n4964 205.079
R1096 VDD.n5643 VDD.n4964 205.079
R1097 VDD.n5643 VDD.n5642 205.079
R1098 VDD.n5642 VDD.n5641 205.079
R1099 VDD.n5641 VDD.n4968 205.079
R1100 VDD.n5635 VDD.n4968 205.079
R1101 VDD.n5544 VDD.n5021 205.079
R1102 VDD.n5545 VDD.n5544 205.079
R1103 VDD.n5546 VDD.n5545 205.079
R1104 VDD.n5546 VDD.n5017 205.079
R1105 VDD.n5552 VDD.n5017 205.079
R1106 VDD.n5553 VDD.n5552 205.079
R1107 VDD.n5554 VDD.n5553 205.079
R1108 VDD.n5554 VDD.n5013 205.079
R1109 VDD.n5560 VDD.n5013 205.079
R1110 VDD.n5561 VDD.n5560 205.079
R1111 VDD.n5562 VDD.n5561 205.079
R1112 VDD.n5562 VDD.n5008 205.079
R1113 VDD.n5569 VDD.n5008 205.079
R1114 VDD.n4584 VDD.n4583 205.079
R1115 VDD.n4584 VDD.n4427 205.079
R1116 VDD.n4590 VDD.n4427 205.079
R1117 VDD.n4591 VDD.n4590 205.079
R1118 VDD.n4592 VDD.n4591 205.079
R1119 VDD.n4592 VDD.n4423 205.079
R1120 VDD.n4598 VDD.n4423 205.079
R1121 VDD.n4599 VDD.n4598 205.079
R1122 VDD.n4600 VDD.n4599 205.079
R1123 VDD.n4600 VDD.n4419 205.079
R1124 VDD.n4607 VDD.n4419 205.079
R1125 VDD.n4608 VDD.n4607 205.079
R1126 VDD.n4610 VDD.n4608 205.079
R1127 VDD.n4505 VDD.n4472 205.079
R1128 VDD.n4505 VDD.n4504 205.079
R1129 VDD.n4504 VDD.n4503 205.079
R1130 VDD.n4503 VDD.n4473 205.079
R1131 VDD.n4497 VDD.n4473 205.079
R1132 VDD.n4497 VDD.n4496 205.079
R1133 VDD.n4496 VDD.n4495 205.079
R1134 VDD.n4495 VDD.n4477 205.079
R1135 VDD.n4489 VDD.n4477 205.079
R1136 VDD.n4489 VDD.n4488 205.079
R1137 VDD.n4488 VDD.n4487 205.079
R1138 VDD.n4487 VDD.n4482 205.079
R1139 VDD.n4482 VDD.n4481 205.079
R1140 VDD.n4873 VDD.n4173 205.079
R1141 VDD.n4873 VDD.n4872 205.079
R1142 VDD.n4872 VDD.n4871 205.079
R1143 VDD.n4871 VDD.n4174 205.079
R1144 VDD.n4865 VDD.n4174 205.079
R1145 VDD.n4865 VDD.n4864 205.079
R1146 VDD.n4864 VDD.n4863 205.079
R1147 VDD.n4863 VDD.n4178 205.079
R1148 VDD.n4857 VDD.n4178 205.079
R1149 VDD.n4857 VDD.n4856 205.079
R1150 VDD.n4856 VDD.n4855 205.079
R1151 VDD.n4855 VDD.n4182 205.079
R1152 VDD.n4849 VDD.n4182 205.079
R1153 VDD.n4758 VDD.n4235 205.079
R1154 VDD.n4759 VDD.n4758 205.079
R1155 VDD.n4760 VDD.n4759 205.079
R1156 VDD.n4760 VDD.n4231 205.079
R1157 VDD.n4766 VDD.n4231 205.079
R1158 VDD.n4767 VDD.n4766 205.079
R1159 VDD.n4768 VDD.n4767 205.079
R1160 VDD.n4768 VDD.n4227 205.079
R1161 VDD.n4774 VDD.n4227 205.079
R1162 VDD.n4775 VDD.n4774 205.079
R1163 VDD.n4776 VDD.n4775 205.079
R1164 VDD.n4776 VDD.n4222 205.079
R1165 VDD.n4783 VDD.n4222 205.079
R1166 VDD.n3730 VDD.n3729 205.079
R1167 VDD.n3730 VDD.n3573 205.079
R1168 VDD.n3736 VDD.n3573 205.079
R1169 VDD.n3737 VDD.n3736 205.079
R1170 VDD.n3738 VDD.n3737 205.079
R1171 VDD.n3738 VDD.n3569 205.079
R1172 VDD.n3744 VDD.n3569 205.079
R1173 VDD.n3745 VDD.n3744 205.079
R1174 VDD.n3746 VDD.n3745 205.079
R1175 VDD.n3746 VDD.n3565 205.079
R1176 VDD.n3753 VDD.n3565 205.079
R1177 VDD.n3754 VDD.n3753 205.079
R1178 VDD.n3756 VDD.n3754 205.079
R1179 VDD.n3651 VDD.n3618 205.079
R1180 VDD.n3651 VDD.n3650 205.079
R1181 VDD.n3650 VDD.n3649 205.079
R1182 VDD.n3649 VDD.n3619 205.079
R1183 VDD.n3643 VDD.n3619 205.079
R1184 VDD.n3643 VDD.n3642 205.079
R1185 VDD.n3642 VDD.n3641 205.079
R1186 VDD.n3641 VDD.n3623 205.079
R1187 VDD.n3635 VDD.n3623 205.079
R1188 VDD.n3635 VDD.n3634 205.079
R1189 VDD.n3634 VDD.n3633 205.079
R1190 VDD.n3633 VDD.n3628 205.079
R1191 VDD.n3628 VDD.n3627 205.079
R1192 VDD.n4019 VDD.n3319 205.079
R1193 VDD.n4019 VDD.n4018 205.079
R1194 VDD.n4018 VDD.n4017 205.079
R1195 VDD.n4017 VDD.n3320 205.079
R1196 VDD.n4011 VDD.n3320 205.079
R1197 VDD.n4011 VDD.n4010 205.079
R1198 VDD.n4010 VDD.n4009 205.079
R1199 VDD.n4009 VDD.n3324 205.079
R1200 VDD.n4003 VDD.n3324 205.079
R1201 VDD.n4003 VDD.n4002 205.079
R1202 VDD.n4002 VDD.n4001 205.079
R1203 VDD.n4001 VDD.n3328 205.079
R1204 VDD.n3995 VDD.n3328 205.079
R1205 VDD.n3904 VDD.n3381 205.079
R1206 VDD.n3905 VDD.n3904 205.079
R1207 VDD.n3906 VDD.n3905 205.079
R1208 VDD.n3906 VDD.n3377 205.079
R1209 VDD.n3912 VDD.n3377 205.079
R1210 VDD.n3913 VDD.n3912 205.079
R1211 VDD.n3914 VDD.n3913 205.079
R1212 VDD.n3914 VDD.n3373 205.079
R1213 VDD.n3920 VDD.n3373 205.079
R1214 VDD.n3921 VDD.n3920 205.079
R1215 VDD.n3922 VDD.n3921 205.079
R1216 VDD.n3922 VDD.n3368 205.079
R1217 VDD.n3929 VDD.n3368 205.079
R1218 VDD.n2944 VDD.n2943 205.079
R1219 VDD.n2944 VDD.n2787 205.079
R1220 VDD.n2950 VDD.n2787 205.079
R1221 VDD.n2951 VDD.n2950 205.079
R1222 VDD.n2952 VDD.n2951 205.079
R1223 VDD.n2952 VDD.n2783 205.079
R1224 VDD.n2958 VDD.n2783 205.079
R1225 VDD.n2959 VDD.n2958 205.079
R1226 VDD.n2960 VDD.n2959 205.079
R1227 VDD.n2960 VDD.n2779 205.079
R1228 VDD.n2967 VDD.n2779 205.079
R1229 VDD.n2968 VDD.n2967 205.079
R1230 VDD.n2970 VDD.n2968 205.079
R1231 VDD.n2865 VDD.n2832 205.079
R1232 VDD.n2865 VDD.n2864 205.079
R1233 VDD.n2864 VDD.n2863 205.079
R1234 VDD.n2863 VDD.n2833 205.079
R1235 VDD.n2857 VDD.n2833 205.079
R1236 VDD.n2857 VDD.n2856 205.079
R1237 VDD.n2856 VDD.n2855 205.079
R1238 VDD.n2855 VDD.n2837 205.079
R1239 VDD.n2849 VDD.n2837 205.079
R1240 VDD.n2849 VDD.n2848 205.079
R1241 VDD.n2848 VDD.n2847 205.079
R1242 VDD.n2847 VDD.n2842 205.079
R1243 VDD.n2842 VDD.n2841 205.079
R1244 VDD.n3233 VDD.n2533 205.079
R1245 VDD.n3233 VDD.n3232 205.079
R1246 VDD.n3232 VDD.n3231 205.079
R1247 VDD.n3231 VDD.n2534 205.079
R1248 VDD.n3225 VDD.n2534 205.079
R1249 VDD.n3225 VDD.n3224 205.079
R1250 VDD.n3224 VDD.n3223 205.079
R1251 VDD.n3223 VDD.n2538 205.079
R1252 VDD.n3217 VDD.n2538 205.079
R1253 VDD.n3217 VDD.n3216 205.079
R1254 VDD.n3216 VDD.n3215 205.079
R1255 VDD.n3215 VDD.n2542 205.079
R1256 VDD.n3209 VDD.n2542 205.079
R1257 VDD.n3118 VDD.n2595 205.079
R1258 VDD.n3119 VDD.n3118 205.079
R1259 VDD.n3120 VDD.n3119 205.079
R1260 VDD.n3120 VDD.n2591 205.079
R1261 VDD.n3126 VDD.n2591 205.079
R1262 VDD.n3127 VDD.n3126 205.079
R1263 VDD.n3128 VDD.n3127 205.079
R1264 VDD.n3128 VDD.n2587 205.079
R1265 VDD.n3134 VDD.n2587 205.079
R1266 VDD.n3135 VDD.n3134 205.079
R1267 VDD.n3136 VDD.n3135 205.079
R1268 VDD.n3136 VDD.n2582 205.079
R1269 VDD.n3143 VDD.n2582 205.079
R1270 VDD.n2089 VDD.n2088 205.079
R1271 VDD.n2089 VDD.n1932 205.079
R1272 VDD.n2095 VDD.n1932 205.079
R1273 VDD.n2096 VDD.n2095 205.079
R1274 VDD.n2097 VDD.n2096 205.079
R1275 VDD.n2097 VDD.n1928 205.079
R1276 VDD.n2103 VDD.n1928 205.079
R1277 VDD.n2104 VDD.n2103 205.079
R1278 VDD.n2105 VDD.n2104 205.079
R1279 VDD.n2105 VDD.n1924 205.079
R1280 VDD.n2112 VDD.n1924 205.079
R1281 VDD.n2113 VDD.n2112 205.079
R1282 VDD.n2115 VDD.n2113 205.079
R1283 VDD.n2010 VDD.n1977 205.079
R1284 VDD.n2010 VDD.n2009 205.079
R1285 VDD.n2009 VDD.n2008 205.079
R1286 VDD.n2008 VDD.n1978 205.079
R1287 VDD.n2002 VDD.n1978 205.079
R1288 VDD.n2002 VDD.n2001 205.079
R1289 VDD.n2001 VDD.n2000 205.079
R1290 VDD.n2000 VDD.n1982 205.079
R1291 VDD.n1994 VDD.n1982 205.079
R1292 VDD.n1994 VDD.n1993 205.079
R1293 VDD.n1993 VDD.n1992 205.079
R1294 VDD.n1992 VDD.n1987 205.079
R1295 VDD.n1987 VDD.n1986 205.079
R1296 VDD.n2378 VDD.n1678 205.079
R1297 VDD.n2378 VDD.n2377 205.079
R1298 VDD.n2377 VDD.n2376 205.079
R1299 VDD.n2376 VDD.n1679 205.079
R1300 VDD.n2370 VDD.n1679 205.079
R1301 VDD.n2370 VDD.n2369 205.079
R1302 VDD.n2369 VDD.n2368 205.079
R1303 VDD.n2368 VDD.n1683 205.079
R1304 VDD.n2362 VDD.n1683 205.079
R1305 VDD.n2362 VDD.n2361 205.079
R1306 VDD.n2361 VDD.n2360 205.079
R1307 VDD.n2360 VDD.n1687 205.079
R1308 VDD.n2354 VDD.n1687 205.079
R1309 VDD.n2263 VDD.n1740 205.079
R1310 VDD.n2264 VDD.n2263 205.079
R1311 VDD.n2265 VDD.n2264 205.079
R1312 VDD.n2265 VDD.n1736 205.079
R1313 VDD.n2271 VDD.n1736 205.079
R1314 VDD.n2272 VDD.n2271 205.079
R1315 VDD.n2273 VDD.n2272 205.079
R1316 VDD.n2273 VDD.n1732 205.079
R1317 VDD.n2279 VDD.n1732 205.079
R1318 VDD.n2280 VDD.n2279 205.079
R1319 VDD.n2281 VDD.n2280 205.079
R1320 VDD.n2281 VDD.n1727 205.079
R1321 VDD.n2288 VDD.n1727 205.079
R1322 VDD.n6431 VDD.n5857 203.786
R1323 VDD.n6432 VDD.n6431 203.786
R1324 VDD.n6433 VDD.n6432 203.786
R1325 VDD.n6433 VDD.n5853 203.786
R1326 VDD.n6439 VDD.n5853 203.786
R1327 VDD.n6440 VDD.n6439 203.786
R1328 VDD.n6441 VDD.n6440 203.786
R1329 VDD.n6441 VDD.n5849 203.786
R1330 VDD.n6447 VDD.n5849 203.786
R1331 VDD.n6448 VDD.n6447 203.786
R1332 VDD.n6449 VDD.n6448 203.786
R1333 VDD.n6449 VDD.n5845 203.786
R1334 VDD.n6455 VDD.n5845 203.786
R1335 VDD.n6456 VDD.n6455 203.786
R1336 VDD.n6457 VDD.n6456 203.786
R1337 VDD.n6457 VDD.n5841 203.786
R1338 VDD.n6463 VDD.n5841 203.786
R1339 VDD.n6464 VDD.n6463 203.786
R1340 VDD.n6465 VDD.n6464 203.786
R1341 VDD.n6465 VDD.n5837 203.786
R1342 VDD.n6471 VDD.n5837 203.786
R1343 VDD.n6472 VDD.n6471 203.786
R1344 VDD.n6473 VDD.n6472 203.786
R1345 VDD.n6473 VDD.n5833 203.786
R1346 VDD.n6479 VDD.n5833 203.786
R1347 VDD.n6480 VDD.n6479 203.786
R1348 VDD.n6481 VDD.n6480 203.786
R1349 VDD.n6481 VDD.n5826 203.786
R1350 VDD.n5577 VDD.n5003 203.786
R1351 VDD.n5578 VDD.n5577 203.786
R1352 VDD.n5579 VDD.n5578 203.786
R1353 VDD.n5579 VDD.n4999 203.786
R1354 VDD.n5585 VDD.n4999 203.786
R1355 VDD.n5586 VDD.n5585 203.786
R1356 VDD.n5587 VDD.n5586 203.786
R1357 VDD.n5587 VDD.n4995 203.786
R1358 VDD.n5593 VDD.n4995 203.786
R1359 VDD.n5594 VDD.n5593 203.786
R1360 VDD.n5595 VDD.n5594 203.786
R1361 VDD.n5595 VDD.n4991 203.786
R1362 VDD.n5601 VDD.n4991 203.786
R1363 VDD.n5602 VDD.n5601 203.786
R1364 VDD.n5603 VDD.n5602 203.786
R1365 VDD.n5603 VDD.n4987 203.786
R1366 VDD.n5609 VDD.n4987 203.786
R1367 VDD.n5610 VDD.n5609 203.786
R1368 VDD.n5611 VDD.n5610 203.786
R1369 VDD.n5611 VDD.n4983 203.786
R1370 VDD.n5617 VDD.n4983 203.786
R1371 VDD.n5618 VDD.n5617 203.786
R1372 VDD.n5619 VDD.n5618 203.786
R1373 VDD.n5619 VDD.n4979 203.786
R1374 VDD.n5625 VDD.n4979 203.786
R1375 VDD.n5626 VDD.n5625 203.786
R1376 VDD.n5627 VDD.n5626 203.786
R1377 VDD.n5627 VDD.n4972 203.786
R1378 VDD.n4791 VDD.n4217 203.786
R1379 VDD.n4792 VDD.n4791 203.786
R1380 VDD.n4793 VDD.n4792 203.786
R1381 VDD.n4793 VDD.n4213 203.786
R1382 VDD.n4799 VDD.n4213 203.786
R1383 VDD.n4800 VDD.n4799 203.786
R1384 VDD.n4801 VDD.n4800 203.786
R1385 VDD.n4801 VDD.n4209 203.786
R1386 VDD.n4807 VDD.n4209 203.786
R1387 VDD.n4808 VDD.n4807 203.786
R1388 VDD.n4809 VDD.n4808 203.786
R1389 VDD.n4809 VDD.n4205 203.786
R1390 VDD.n4815 VDD.n4205 203.786
R1391 VDD.n4816 VDD.n4815 203.786
R1392 VDD.n4817 VDD.n4816 203.786
R1393 VDD.n4817 VDD.n4201 203.786
R1394 VDD.n4823 VDD.n4201 203.786
R1395 VDD.n4824 VDD.n4823 203.786
R1396 VDD.n4825 VDD.n4824 203.786
R1397 VDD.n4825 VDD.n4197 203.786
R1398 VDD.n4831 VDD.n4197 203.786
R1399 VDD.n4832 VDD.n4831 203.786
R1400 VDD.n4833 VDD.n4832 203.786
R1401 VDD.n4833 VDD.n4193 203.786
R1402 VDD.n4839 VDD.n4193 203.786
R1403 VDD.n4840 VDD.n4839 203.786
R1404 VDD.n4841 VDD.n4840 203.786
R1405 VDD.n4841 VDD.n4186 203.786
R1406 VDD.n3937 VDD.n3363 203.786
R1407 VDD.n3938 VDD.n3937 203.786
R1408 VDD.n3939 VDD.n3938 203.786
R1409 VDD.n3939 VDD.n3359 203.786
R1410 VDD.n3945 VDD.n3359 203.786
R1411 VDD.n3946 VDD.n3945 203.786
R1412 VDD.n3947 VDD.n3946 203.786
R1413 VDD.n3947 VDD.n3355 203.786
R1414 VDD.n3953 VDD.n3355 203.786
R1415 VDD.n3954 VDD.n3953 203.786
R1416 VDD.n3955 VDD.n3954 203.786
R1417 VDD.n3955 VDD.n3351 203.786
R1418 VDD.n3961 VDD.n3351 203.786
R1419 VDD.n3962 VDD.n3961 203.786
R1420 VDD.n3963 VDD.n3962 203.786
R1421 VDD.n3963 VDD.n3347 203.786
R1422 VDD.n3969 VDD.n3347 203.786
R1423 VDD.n3970 VDD.n3969 203.786
R1424 VDD.n3971 VDD.n3970 203.786
R1425 VDD.n3971 VDD.n3343 203.786
R1426 VDD.n3977 VDD.n3343 203.786
R1427 VDD.n3978 VDD.n3977 203.786
R1428 VDD.n3979 VDD.n3978 203.786
R1429 VDD.n3979 VDD.n3339 203.786
R1430 VDD.n3985 VDD.n3339 203.786
R1431 VDD.n3986 VDD.n3985 203.786
R1432 VDD.n3987 VDD.n3986 203.786
R1433 VDD.n3987 VDD.n3332 203.786
R1434 VDD.n3151 VDD.n2577 203.786
R1435 VDD.n3152 VDD.n3151 203.786
R1436 VDD.n3153 VDD.n3152 203.786
R1437 VDD.n3153 VDD.n2573 203.786
R1438 VDD.n3159 VDD.n2573 203.786
R1439 VDD.n3160 VDD.n3159 203.786
R1440 VDD.n3161 VDD.n3160 203.786
R1441 VDD.n3161 VDD.n2569 203.786
R1442 VDD.n3167 VDD.n2569 203.786
R1443 VDD.n3168 VDD.n3167 203.786
R1444 VDD.n3169 VDD.n3168 203.786
R1445 VDD.n3169 VDD.n2565 203.786
R1446 VDD.n3175 VDD.n2565 203.786
R1447 VDD.n3176 VDD.n3175 203.786
R1448 VDD.n3177 VDD.n3176 203.786
R1449 VDD.n3177 VDD.n2561 203.786
R1450 VDD.n3183 VDD.n2561 203.786
R1451 VDD.n3184 VDD.n3183 203.786
R1452 VDD.n3185 VDD.n3184 203.786
R1453 VDD.n3185 VDD.n2557 203.786
R1454 VDD.n3191 VDD.n2557 203.786
R1455 VDD.n3192 VDD.n3191 203.786
R1456 VDD.n3193 VDD.n3192 203.786
R1457 VDD.n3193 VDD.n2553 203.786
R1458 VDD.n3199 VDD.n2553 203.786
R1459 VDD.n3200 VDD.n3199 203.786
R1460 VDD.n3201 VDD.n3200 203.786
R1461 VDD.n3201 VDD.n2546 203.786
R1462 VDD.n2296 VDD.n1722 203.786
R1463 VDD.n2297 VDD.n2296 203.786
R1464 VDD.n2298 VDD.n2297 203.786
R1465 VDD.n2298 VDD.n1718 203.786
R1466 VDD.n2304 VDD.n1718 203.786
R1467 VDD.n2305 VDD.n2304 203.786
R1468 VDD.n2306 VDD.n2305 203.786
R1469 VDD.n2306 VDD.n1714 203.786
R1470 VDD.n2312 VDD.n1714 203.786
R1471 VDD.n2313 VDD.n2312 203.786
R1472 VDD.n2314 VDD.n2313 203.786
R1473 VDD.n2314 VDD.n1710 203.786
R1474 VDD.n2320 VDD.n1710 203.786
R1475 VDD.n2321 VDD.n2320 203.786
R1476 VDD.n2322 VDD.n2321 203.786
R1477 VDD.n2322 VDD.n1706 203.786
R1478 VDD.n2328 VDD.n1706 203.786
R1479 VDD.n2329 VDD.n2328 203.786
R1480 VDD.n2330 VDD.n2329 203.786
R1481 VDD.n2330 VDD.n1702 203.786
R1482 VDD.n2336 VDD.n1702 203.786
R1483 VDD.n2337 VDD.n2336 203.786
R1484 VDD.n2338 VDD.n2337 203.786
R1485 VDD.n2338 VDD.n1698 203.786
R1486 VDD.n2344 VDD.n1698 203.786
R1487 VDD.n2345 VDD.n2344 203.786
R1488 VDD.n2346 VDD.n2345 203.786
R1489 VDD.n2346 VDD.n1691 203.786
R1490 VDD.n11649 VDD.n7612 198.731
R1491 VDD.n12087 VDD.n7372 195.649
R1492 VDD.n11643 VDD.n7611 195.404
R1493 VDD.n12327 VDD.n12326 193.984
R1494 VDD.n12409 VDD.n6933 186.405
R1495 VDD.n9979 VDD.n9978 185
R1496 VDD.n9977 VDD.n9974 185
R1497 VDD.n9183 VDD.n9076 185
R1498 VDD.n9169 VDD.n9076 185
R1499 VDD.n9184 VDD.n9183 185
R1500 VDD.n9184 VDD.n9169 185
R1501 VDD.n9183 VDD.n9182 185
R1502 VDD.n10960 VDD.n10959 185
R1503 VDD.n10960 VDD.n9221 185
R1504 VDD.n10958 VDD.n9221 185
R1505 VDD.n10959 VDD.n10958 185
R1506 VDD.n10959 VDD.n9222 185
R1507 VDD.n9222 VDD.n9221 185
R1508 VDD.n9209 VDD.n7070 185
R1509 VDD.n9218 VDD.n7070 185
R1510 VDD.n9217 VDD.n7070 185
R1511 VDD.n11026 VDD.n8729 185
R1512 VDD.n8729 VDD.n8720 185
R1513 VDD.n11025 VDD.n8720 185
R1514 VDD.n8730 VDD.n8720 185
R1515 VDD.n10988 VDD.n8720 185
R1516 VDD.n11026 VDD.n8730 185
R1517 VDD.n8731 VDD.n8720 185
R1518 VDD.n8728 VDD.n8720 185
R1519 VDD.n10494 VDD.n10432 185
R1520 VDD.n10432 VDD.n10162 185
R1521 VDD.n10495 VDD.n10494 185
R1522 VDD.n10494 VDD.n10422 185
R1523 VDD.n10494 VDD.n10493 185
R1524 VDD.n10479 VDD.n10478 185
R1525 VDD.n10479 VDD.n10448 185
R1526 VDD.n10481 VDD.n10479 185
R1527 VDD.n10493 VDD.n10162 185
R1528 VDD.n10422 VDD.n10162 185
R1529 VDD.n10495 VDD.n10162 185
R1530 VDD.n6925 VDD.n6923 185
R1531 VDD.n12475 VDD.n12474 185
R1532 VDD.n12482 VDD.n12481 185
R1533 VDD.n12489 VDD.n6910 185
R1534 VDD.n12480 VDD.n12428 185
R1535 VDD.n12488 VDD.n12487 185
R1536 VDD.n12488 VDD.n12426 185
R1537 VDD.n6912 VDD.n6909 185
R1538 VDD.n12426 VDD.n6912 185
R1539 VDD.n12423 VDD.n12422 185
R1540 VDD.n12472 VDD.n12471 185
R1541 VDD.n12466 VDD.n12465 185
R1542 VDD.n12460 VDD.n12438 185
R1543 VDD.n12473 VDD.n12432 185
R1544 VDD.n12473 VDD.n12426 185
R1545 VDD.n12468 VDD.n12467 185
R1546 VDD.n12462 VDD.n12461 185
R1547 VDD.n12456 VDD.n12455 185
R1548 VDD.n12454 VDD.n12453 185
R1549 VDD.n12476 VDD.n12430 185
R1550 VDD.n6939 VDD.n6938 183.524
R1551 VDD.n12404 VDD.n6939 183.524
R1552 VDD.n12404 VDD.n12403 183.524
R1553 VDD.n12403 VDD.n12402 183.524
R1554 VDD.n12402 VDD.n6940 183.524
R1555 VDD.n12393 VDD.n6940 183.524
R1556 VDD.n12393 VDD.n12392 183.524
R1557 VDD.n12392 VDD.n12391 183.524
R1558 VDD.n12391 VDD.n6949 183.524
R1559 VDD.n12382 VDD.n6949 183.524
R1560 VDD.n12382 VDD.n12381 183.524
R1561 VDD.n12381 VDD.n12380 183.524
R1562 VDD.n12380 VDD.n6958 183.524
R1563 VDD.n12371 VDD.n12370 183.524
R1564 VDD.n12370 VDD.n12369 183.524
R1565 VDD.n12369 VDD.n6968 183.524
R1566 VDD.n12360 VDD.n6968 183.524
R1567 VDD.n12360 VDD.n12359 183.524
R1568 VDD.n12359 VDD.n12358 183.524
R1569 VDD.n12358 VDD.n6977 183.524
R1570 VDD.n12349 VDD.n6977 183.524
R1571 VDD.n12349 VDD.n12348 183.524
R1572 VDD.n12348 VDD.n12347 183.524
R1573 VDD.n12347 VDD.n6984 183.524
R1574 VDD.n12338 VDD.n6984 183.524
R1575 VDD.n12338 VDD.n12337 183.524
R1576 VDD.n12337 VDD.n12336 183.524
R1577 VDD.n12336 VDD.n6993 183.524
R1578 VDD.n12327 VDD.n6993 183.524
R1579 VDD.n10979 VDD.n9198 179.883
R1580 VDD.n5738 VDD.n5715 175.386
R1581 VDD.n5765 VDD.n5739 175.386
R1582 VDD.n4098 VDD.n4075 175.386
R1583 VDD.n4125 VDD.n4099 175.386
R1584 VDD.n2457 VDD.n2434 175.386
R1585 VDD.n2485 VDD.n2458 175.386
R1586 VDD.n817 VDD.n794 175.386
R1587 VDD.n845 VDD.n818 175.386
R1588 VDD.n10067 VDD.n10025 174.535
R1589 VDD.n10063 VDD.n10062 174.535
R1590 VDD.n10054 VDD.n10053 174.535
R1591 VDD.n10046 VDD.n10041 174.535
R1592 VDD.n10587 VDD.n10144 174.535
R1593 VDD.n10624 VDD.n10623 174.535
R1594 VDD.n10613 VDD.n10612 174.535
R1595 VDD.n10605 VDD.n10600 174.535
R1596 VDD.n10520 VDD.n10502 174.535
R1597 VDD.n10563 VDD.n10562 174.535
R1598 VDD.n10553 VDD.n10537 174.535
R1599 VDD.n10551 VDD.n10538 174.535
R1600 VDD.n9606 VDD.n9584 174.535
R1601 VDD.n9604 VDD.n9585 174.535
R1602 VDD.n9616 VDD.n9615 174.535
R1603 VDD.n9623 VDD.n9622 174.535
R1604 VDD.n9631 VDD.n9630 174.535
R1605 VDD.n10763 VDD.n10762 174.535
R1606 VDD.n10718 VDD.n10717 174.535
R1607 VDD.n10748 VDD.n10721 174.535
R1608 VDD.n10746 VDD.n10722 174.535
R1609 VDD.n10737 VDD.n10736 174.535
R1610 VDD.n8911 VDD.n8910 174.535
R1611 VDD.n8905 VDD.n8904 174.535
R1612 VDD.n9375 VDD.n9374 174.535
R1613 VDD.n9385 VDD.n9384 174.535
R1614 VDD.n9441 VDD.n9391 174.535
R1615 VDD.n9432 VDD.n9392 174.535
R1616 VDD.n9430 VDD.n9397 174.535
R1617 VDD.n5724 VDD.t144 171.452
R1618 VDD.n4084 VDD.t109 171.452
R1619 VDD.n2443 VDD.t23 171.452
R1620 VDD.n803 VDD.t126 171.452
R1621 VDD.n8538 VDD.n7783 171
R1622 VDD.n6249 VDD.n5813 168.889
R1623 VDD.n5879 VDD.n5875 168.889
R1624 VDD.n5395 VDD.n4959 168.889
R1625 VDD.n5025 VDD.n5021 168.889
R1626 VDD.n4609 VDD.n4173 168.889
R1627 VDD.n4239 VDD.n4235 168.889
R1628 VDD.n3755 VDD.n3319 168.889
R1629 VDD.n3385 VDD.n3381 168.889
R1630 VDD.n2969 VDD.n2533 168.889
R1631 VDD.n2599 VDD.n2595 168.889
R1632 VDD.n2114 VDD.n1678 168.889
R1633 VDD.n1744 VDD.n1740 168.889
R1634 VDD.n8121 VDD.n8112 167.919
R1635 VDD.n6967 VDD.n6958 167.331
R1636 VDD.n6425 VDD.n6424 164.827
R1637 VDD.n5571 VDD.n5570 164.827
R1638 VDD.n4785 VDD.n4784 164.827
R1639 VDD.n3931 VDD.n3930 164.827
R1640 VDD.n3145 VDD.n3144 164.827
R1641 VDD.n2290 VDD.n2289 164.827
R1642 VDD.n12093 VDD.n12092 162.857
R1643 VDD.n6489 VDD.n6488 162.857
R1644 VDD.n6424 VDD.n6423 162.857
R1645 VDD.n5635 VDD.n5634 162.857
R1646 VDD.n5570 VDD.n5569 162.857
R1647 VDD.n4849 VDD.n4848 162.857
R1648 VDD.n4784 VDD.n4783 162.857
R1649 VDD.n3995 VDD.n3994 162.857
R1650 VDD.n3930 VDD.n3929 162.857
R1651 VDD.n3209 VDD.n3208 162.857
R1652 VDD.n3144 VDD.n3143 162.857
R1653 VDD.n2354 VDD.n2353 162.857
R1654 VDD.n2289 VDD.n2288 162.857
R1655 VDD.n6488 VDD.n6487 161.831
R1656 VDD.n5634 VDD.n5633 161.831
R1657 VDD.n4848 VDD.n4847 161.831
R1658 VDD.n3994 VDD.n3993 161.831
R1659 VDD.n3208 VDD.n3207 161.831
R1660 VDD.n2353 VDD.n2352 161.831
R1661 VDD.n5727 VDD.t145 160.743
R1662 VDD.n4087 VDD.t110 160.743
R1663 VDD.n2446 VDD.t24 160.743
R1664 VDD.n806 VDD.t127 160.743
R1665 VDD.n9912 VDD.t209 160.742
R1666 VDD.n6380 VDD.n5879 160.256
R1667 VDD.n5526 VDD.n5025 160.256
R1668 VDD.n4740 VDD.n4239 160.256
R1669 VDD.n3886 VDD.n3385 160.256
R1670 VDD.n3100 VDD.n2599 160.256
R1671 VDD.n2245 VDD.n1744 160.256
R1672 VDD.n9928 VDD.t212 159.81
R1673 VDD.n9072 VDD.n8729 159.156
R1674 VDD.n6159 VDD.n6101 159.113
R1675 VDD.n6160 VDD.n6159 159.113
R1676 VDD.n6161 VDD.n6160 159.113
R1677 VDD.n6161 VDD.n6097 159.113
R1678 VDD.n6167 VDD.n6097 159.113
R1679 VDD.n6168 VDD.n6167 159.113
R1680 VDD.n6169 VDD.n6168 159.113
R1681 VDD.n6169 VDD.n6093 159.113
R1682 VDD.n6175 VDD.n6093 159.113
R1683 VDD.n6176 VDD.n6175 159.113
R1684 VDD.n6177 VDD.n6176 159.113
R1685 VDD.n6177 VDD.n6089 159.113
R1686 VDD.n6183 VDD.n6089 159.113
R1687 VDD.n6184 VDD.n6183 159.113
R1688 VDD.n6185 VDD.n6184 159.113
R1689 VDD.n6185 VDD.n6085 159.113
R1690 VDD.n6191 VDD.n6085 159.113
R1691 VDD.n6192 VDD.n6191 159.113
R1692 VDD.n6193 VDD.n6192 159.113
R1693 VDD.n6193 VDD.n6081 159.113
R1694 VDD.n6199 VDD.n6081 159.113
R1695 VDD.n6200 VDD.n6199 159.113
R1696 VDD.n6201 VDD.n6200 159.113
R1697 VDD.n6201 VDD.n6077 159.113
R1698 VDD.n6208 VDD.n6077 159.113
R1699 VDD.n6209 VDD.n6208 159.113
R1700 VDD.n6210 VDD.n6209 159.113
R1701 VDD.n6210 VDD.n6071 159.113
R1702 VDD.n5305 VDD.n5247 159.113
R1703 VDD.n5306 VDD.n5305 159.113
R1704 VDD.n5307 VDD.n5306 159.113
R1705 VDD.n5307 VDD.n5243 159.113
R1706 VDD.n5313 VDD.n5243 159.113
R1707 VDD.n5314 VDD.n5313 159.113
R1708 VDD.n5315 VDD.n5314 159.113
R1709 VDD.n5315 VDD.n5239 159.113
R1710 VDD.n5321 VDD.n5239 159.113
R1711 VDD.n5322 VDD.n5321 159.113
R1712 VDD.n5323 VDD.n5322 159.113
R1713 VDD.n5323 VDD.n5235 159.113
R1714 VDD.n5329 VDD.n5235 159.113
R1715 VDD.n5330 VDD.n5329 159.113
R1716 VDD.n5331 VDD.n5330 159.113
R1717 VDD.n5331 VDD.n5231 159.113
R1718 VDD.n5337 VDD.n5231 159.113
R1719 VDD.n5338 VDD.n5337 159.113
R1720 VDD.n5339 VDD.n5338 159.113
R1721 VDD.n5339 VDD.n5227 159.113
R1722 VDD.n5345 VDD.n5227 159.113
R1723 VDD.n5346 VDD.n5345 159.113
R1724 VDD.n5347 VDD.n5346 159.113
R1725 VDD.n5347 VDD.n5223 159.113
R1726 VDD.n5354 VDD.n5223 159.113
R1727 VDD.n5355 VDD.n5354 159.113
R1728 VDD.n5356 VDD.n5355 159.113
R1729 VDD.n5356 VDD.n5217 159.113
R1730 VDD.n4519 VDD.n4461 159.113
R1731 VDD.n4520 VDD.n4519 159.113
R1732 VDD.n4521 VDD.n4520 159.113
R1733 VDD.n4521 VDD.n4457 159.113
R1734 VDD.n4527 VDD.n4457 159.113
R1735 VDD.n4528 VDD.n4527 159.113
R1736 VDD.n4529 VDD.n4528 159.113
R1737 VDD.n4529 VDD.n4453 159.113
R1738 VDD.n4535 VDD.n4453 159.113
R1739 VDD.n4536 VDD.n4535 159.113
R1740 VDD.n4537 VDD.n4536 159.113
R1741 VDD.n4537 VDD.n4449 159.113
R1742 VDD.n4543 VDD.n4449 159.113
R1743 VDD.n4544 VDD.n4543 159.113
R1744 VDD.n4545 VDD.n4544 159.113
R1745 VDD.n4545 VDD.n4445 159.113
R1746 VDD.n4551 VDD.n4445 159.113
R1747 VDD.n4552 VDD.n4551 159.113
R1748 VDD.n4553 VDD.n4552 159.113
R1749 VDD.n4553 VDD.n4441 159.113
R1750 VDD.n4559 VDD.n4441 159.113
R1751 VDD.n4560 VDD.n4559 159.113
R1752 VDD.n4561 VDD.n4560 159.113
R1753 VDD.n4561 VDD.n4437 159.113
R1754 VDD.n4568 VDD.n4437 159.113
R1755 VDD.n4569 VDD.n4568 159.113
R1756 VDD.n4570 VDD.n4569 159.113
R1757 VDD.n4570 VDD.n4431 159.113
R1758 VDD.n3665 VDD.n3607 159.113
R1759 VDD.n3666 VDD.n3665 159.113
R1760 VDD.n3667 VDD.n3666 159.113
R1761 VDD.n3667 VDD.n3603 159.113
R1762 VDD.n3673 VDD.n3603 159.113
R1763 VDD.n3674 VDD.n3673 159.113
R1764 VDD.n3675 VDD.n3674 159.113
R1765 VDD.n3675 VDD.n3599 159.113
R1766 VDD.n3681 VDD.n3599 159.113
R1767 VDD.n3682 VDD.n3681 159.113
R1768 VDD.n3683 VDD.n3682 159.113
R1769 VDD.n3683 VDD.n3595 159.113
R1770 VDD.n3689 VDD.n3595 159.113
R1771 VDD.n3690 VDD.n3689 159.113
R1772 VDD.n3691 VDD.n3690 159.113
R1773 VDD.n3691 VDD.n3591 159.113
R1774 VDD.n3697 VDD.n3591 159.113
R1775 VDD.n3698 VDD.n3697 159.113
R1776 VDD.n3699 VDD.n3698 159.113
R1777 VDD.n3699 VDD.n3587 159.113
R1778 VDD.n3705 VDD.n3587 159.113
R1779 VDD.n3706 VDD.n3705 159.113
R1780 VDD.n3707 VDD.n3706 159.113
R1781 VDD.n3707 VDD.n3583 159.113
R1782 VDD.n3714 VDD.n3583 159.113
R1783 VDD.n3715 VDD.n3714 159.113
R1784 VDD.n3716 VDD.n3715 159.113
R1785 VDD.n3716 VDD.n3577 159.113
R1786 VDD.n2879 VDD.n2821 159.113
R1787 VDD.n2880 VDD.n2879 159.113
R1788 VDD.n2881 VDD.n2880 159.113
R1789 VDD.n2881 VDD.n2817 159.113
R1790 VDD.n2887 VDD.n2817 159.113
R1791 VDD.n2888 VDD.n2887 159.113
R1792 VDD.n2889 VDD.n2888 159.113
R1793 VDD.n2889 VDD.n2813 159.113
R1794 VDD.n2895 VDD.n2813 159.113
R1795 VDD.n2896 VDD.n2895 159.113
R1796 VDD.n2897 VDD.n2896 159.113
R1797 VDD.n2897 VDD.n2809 159.113
R1798 VDD.n2903 VDD.n2809 159.113
R1799 VDD.n2904 VDD.n2903 159.113
R1800 VDD.n2905 VDD.n2904 159.113
R1801 VDD.n2905 VDD.n2805 159.113
R1802 VDD.n2911 VDD.n2805 159.113
R1803 VDD.n2912 VDD.n2911 159.113
R1804 VDD.n2913 VDD.n2912 159.113
R1805 VDD.n2913 VDD.n2801 159.113
R1806 VDD.n2919 VDD.n2801 159.113
R1807 VDD.n2920 VDD.n2919 159.113
R1808 VDD.n2921 VDD.n2920 159.113
R1809 VDD.n2921 VDD.n2797 159.113
R1810 VDD.n2928 VDD.n2797 159.113
R1811 VDD.n2929 VDD.n2928 159.113
R1812 VDD.n2930 VDD.n2929 159.113
R1813 VDD.n2930 VDD.n2791 159.113
R1814 VDD.n2024 VDD.n1966 159.113
R1815 VDD.n2025 VDD.n2024 159.113
R1816 VDD.n2026 VDD.n2025 159.113
R1817 VDD.n2026 VDD.n1962 159.113
R1818 VDD.n2032 VDD.n1962 159.113
R1819 VDD.n2033 VDD.n2032 159.113
R1820 VDD.n2034 VDD.n2033 159.113
R1821 VDD.n2034 VDD.n1958 159.113
R1822 VDD.n2040 VDD.n1958 159.113
R1823 VDD.n2041 VDD.n2040 159.113
R1824 VDD.n2042 VDD.n2041 159.113
R1825 VDD.n2042 VDD.n1954 159.113
R1826 VDD.n2048 VDD.n1954 159.113
R1827 VDD.n2049 VDD.n2048 159.113
R1828 VDD.n2050 VDD.n2049 159.113
R1829 VDD.n2050 VDD.n1950 159.113
R1830 VDD.n2056 VDD.n1950 159.113
R1831 VDD.n2057 VDD.n2056 159.113
R1832 VDD.n2058 VDD.n2057 159.113
R1833 VDD.n2058 VDD.n1946 159.113
R1834 VDD.n2064 VDD.n1946 159.113
R1835 VDD.n2065 VDD.n2064 159.113
R1836 VDD.n2066 VDD.n2065 159.113
R1837 VDD.n2066 VDD.n1942 159.113
R1838 VDD.n2073 VDD.n1942 159.113
R1839 VDD.n2074 VDD.n2073 159.113
R1840 VDD.n2075 VDD.n2074 159.113
R1841 VDD.n2075 VDD.n1936 159.113
R1842 VDD.n5719 VDD.t11 158.225
R1843 VDD.n4079 VDD.t112 158.225
R1844 VDD.n2438 VDD.t139 158.225
R1845 VDD.n798 VDD.t171 158.225
R1846 VDD.n6249 VDD.n5807 154.488
R1847 VDD.n5395 VDD.n4953 154.488
R1848 VDD.n4609 VDD.n4167 154.488
R1849 VDD.n3755 VDD.n3313 154.488
R1850 VDD.n2969 VDD.n2527 154.488
R1851 VDD.n2114 VDD.n1672 154.488
R1852 VDD.n10481 VDD.n10480 153.975
R1853 VDD.n9650 VDD.n9647 152
R1854 VDD.n9649 VDD.n9648 152
R1855 VDD.n9667 VDD.n9661 152
R1856 VDD.n9666 VDD.n9665 152
R1857 VDD.n10793 VDD.n10790 152
R1858 VDD.n10792 VDD.n10791 152
R1859 VDD.n10810 VDD.n10804 152
R1860 VDD.n10809 VDD.n10808 152
R1861 VDD.n8869 VDD.n8866 152
R1862 VDD.n8868 VDD.n8867 152
R1863 VDD.n8967 VDD.n8966 152
R1864 VDD.n8962 VDD.n8860 152
R1865 VDD.n8961 VDD.n8960 152
R1866 VDD.n8965 VDD.n8964 152
R1867 VDD.n9005 VDD.n9004 152
R1868 VDD.n9006 VDD.n9000 152
R1869 VDD.n8987 VDD.n8986 152
R1870 VDD.n8984 VDD.n8983 152
R1871 VDD.n8985 VDD.n8832 152
R1872 VDD.n8988 VDD.n8833 152
R1873 VDD.n9279 VDD.n9278 152
R1874 VDD.n9281 VDD.n9280 152
R1875 VDD.n9409 VDD.n9408 152
R1876 VDD.n9411 VDD.n9410 152
R1877 VDD.t3 VDD.t4 151.181
R1878 VDD.t6 VDD.t3 151.181
R1879 VDD.t115 VDD.t160 151.181
R1880 VDD.t113 VDD.t115 151.181
R1881 VDD.t134 VDD.t113 151.181
R1882 VDD.t1 VDD.t134 151.181
R1883 VDD.t140 VDD.t1 151.181
R1884 VDD.t52 VDD.t140 151.181
R1885 VDD.t37 VDD.t52 151.181
R1886 VDD.n6154 VDD.n6102 141.731
R1887 VDD.n6213 VDD.n6212 141.731
R1888 VDD.n5300 VDD.n5248 141.731
R1889 VDD.n5359 VDD.n5358 141.731
R1890 VDD.n4514 VDD.n4462 141.731
R1891 VDD.n4573 VDD.n4572 141.731
R1892 VDD.n3660 VDD.n3608 141.731
R1893 VDD.n3719 VDD.n3718 141.731
R1894 VDD.n2874 VDD.n2822 141.731
R1895 VDD.n2933 VDD.n2932 141.731
R1896 VDD.n2019 VDD.n1967 141.731
R1897 VDD.n2078 VDD.n2077 141.731
R1898 VDD.n6426 VDD.n5858 140.19
R1899 VDD.n6486 VDD.n5829 140.19
R1900 VDD.n5572 VDD.n5004 140.19
R1901 VDD.n5632 VDD.n4975 140.19
R1902 VDD.n4786 VDD.n4218 140.19
R1903 VDD.n4846 VDD.n4189 140.19
R1904 VDD.n3932 VDD.n3364 140.19
R1905 VDD.n3992 VDD.n3335 140.19
R1906 VDD.n3146 VDD.n2578 140.19
R1907 VDD.n3206 VDD.n2549 140.19
R1908 VDD.n2291 VDD.n1723 140.19
R1909 VDD.n2351 VDD.n1694 140.19
R1910 VDD.n12128 VDD.n7352 138.649
R1911 VDD.n12091 VDD.n7370 138.649
R1912 VDD.n11584 VDD.n7642 138.649
R1913 VDD.n11644 VDD.n11642 138.649
R1914 VDD.n12692 VDD.n6701 137.311
R1915 VDD.n6723 VDD.n6714 133.655
R1916 VDD.n12673 VDD.n6723 133.655
R1917 VDD.n12673 VDD.n6724 133.655
R1918 VDD.n12669 VDD.n6724 133.655
R1919 VDD.n12669 VDD.n6746 133.655
R1920 VDD.n12661 VDD.n6746 133.655
R1921 VDD.n12661 VDD.n6755 133.655
R1922 VDD.n12657 VDD.n6755 133.655
R1923 VDD.n12657 VDD.n6757 133.655
R1924 VDD.n12649 VDD.n6757 133.655
R1925 VDD.n12649 VDD.n6766 133.655
R1926 VDD.n12645 VDD.n6766 133.655
R1927 VDD.n12645 VDD.n6768 133.655
R1928 VDD.n12637 VDD.n6768 133.655
R1929 VDD.n12637 VDD.n6778 133.655
R1930 VDD.n12633 VDD.n6778 133.655
R1931 VDD.n12633 VDD.n6780 133.655
R1932 VDD.n12625 VDD.n6780 133.655
R1933 VDD.n12625 VDD.n6790 133.655
R1934 VDD.n12621 VDD.n6790 133.655
R1935 VDD.n12621 VDD.n6792 133.655
R1936 VDD.n12613 VDD.n6792 133.655
R1937 VDD.n12613 VDD.n6800 133.655
R1938 VDD.n12609 VDD.n6800 133.655
R1939 VDD.n12609 VDD.n6802 133.655
R1940 VDD.n12601 VDD.n6802 133.655
R1941 VDD.n12601 VDD.n6812 133.655
R1942 VDD.n12597 VDD.n6812 133.655
R1943 VDD.n12597 VDD.n6814 133.655
R1944 VDD.n12589 VDD.n6814 133.655
R1945 VDD.n12589 VDD.n6821 133.655
R1946 VDD.n12585 VDD.n6821 133.655
R1947 VDD.n12585 VDD.n6823 133.655
R1948 VDD.n12577 VDD.n6823 133.655
R1949 VDD.n12577 VDD.n6832 133.655
R1950 VDD.n12573 VDD.n6832 133.655
R1951 VDD.n12573 VDD.n6834 133.655
R1952 VDD.n12565 VDD.n6834 133.655
R1953 VDD.n12565 VDD.n6844 133.655
R1954 VDD.n12561 VDD.n6844 133.655
R1955 VDD.n12561 VDD.n6846 133.655
R1956 VDD.n12553 VDD.n6846 133.655
R1957 VDD.n12553 VDD.n6854 133.655
R1958 VDD.n12549 VDD.n6854 133.655
R1959 VDD.n12549 VDD.n6856 133.655
R1960 VDD.n12541 VDD.n6856 133.655
R1961 VDD.n12541 VDD.n6866 133.655
R1962 VDD.n12537 VDD.n6866 133.655
R1963 VDD.n12537 VDD.n6868 133.655
R1964 VDD.n12529 VDD.n6868 133.655
R1965 VDD.n12529 VDD.n6876 133.655
R1966 VDD.n12525 VDD.n6876 133.655
R1967 VDD.n12525 VDD.n6878 133.655
R1968 VDD.n12517 VDD.n6878 133.655
R1969 VDD.n12517 VDD.n6888 133.655
R1970 VDD.n12513 VDD.n6888 133.655
R1971 VDD.n12513 VDD.n6890 133.655
R1972 VDD.n12505 VDD.n6890 133.655
R1973 VDD.n12505 VDD.n6900 133.655
R1974 VDD.n12501 VDD.n6900 133.655
R1975 VDD.n12501 VDD.n6902 133.655
R1976 VDD.n6732 VDD.n6729 133.655
R1977 VDD.n6735 VDD.n6734 133.655
R1978 VDD.n6739 VDD.n6738 133.655
R1979 VDD.n12679 VDD.n6716 133.655
R1980 VDD.n12675 VDD.n6716 133.655
R1981 VDD.n12675 VDD.n6719 133.655
R1982 VDD.n12667 VDD.n6719 133.655
R1983 VDD.n12667 VDD.n6750 133.655
R1984 VDD.n12663 VDD.n6750 133.655
R1985 VDD.n12663 VDD.n6752 133.655
R1986 VDD.n12655 VDD.n6752 133.655
R1987 VDD.n12655 VDD.n6760 133.655
R1988 VDD.n12651 VDD.n6760 133.655
R1989 VDD.n12651 VDD.n6762 133.655
R1990 VDD.n12643 VDD.n6762 133.655
R1991 VDD.n12643 VDD.n6772 133.655
R1992 VDD.n12639 VDD.n6772 133.655
R1993 VDD.n12639 VDD.n6774 133.655
R1994 VDD.n12631 VDD.n6774 133.655
R1995 VDD.n12631 VDD.n6784 133.655
R1996 VDD.n12627 VDD.n6784 133.655
R1997 VDD.n12627 VDD.n6786 133.655
R1998 VDD.n12619 VDD.n6786 133.655
R1999 VDD.n12619 VDD.n6794 133.655
R2000 VDD.n12615 VDD.n6794 133.655
R2001 VDD.n12615 VDD.n6796 133.655
R2002 VDD.n12607 VDD.n6796 133.655
R2003 VDD.n12607 VDD.n6806 133.655
R2004 VDD.n12603 VDD.n6806 133.655
R2005 VDD.n12603 VDD.n6808 133.655
R2006 VDD.n12595 VDD.n6808 133.655
R2007 VDD.n12595 VDD.n6817 133.655
R2008 VDD.n12591 VDD.n6817 133.655
R2009 VDD.n12591 VDD.n6819 133.655
R2010 VDD.n12583 VDD.n6819 133.655
R2011 VDD.n12583 VDD.n6826 133.655
R2012 VDD.n12579 VDD.n6826 133.655
R2013 VDD.n12579 VDD.n6828 133.655
R2014 VDD.n12571 VDD.n6828 133.655
R2015 VDD.n12571 VDD.n6838 133.655
R2016 VDD.n12567 VDD.n6838 133.655
R2017 VDD.n12567 VDD.n6840 133.655
R2018 VDD.n12559 VDD.n6840 133.655
R2019 VDD.n12559 VDD.n6850 133.655
R2020 VDD.n12555 VDD.n6850 133.655
R2021 VDD.n12555 VDD.n6852 133.655
R2022 VDD.n12547 VDD.n6852 133.655
R2023 VDD.n12547 VDD.n6860 133.655
R2024 VDD.n12543 VDD.n6860 133.655
R2025 VDD.n12543 VDD.n6862 133.655
R2026 VDD.n12535 VDD.n6862 133.655
R2027 VDD.n12535 VDD.n6871 133.655
R2028 VDD.n12531 VDD.n6871 133.655
R2029 VDD.n12531 VDD.n6873 133.655
R2030 VDD.n12523 VDD.n6873 133.655
R2031 VDD.n12523 VDD.n6882 133.655
R2032 VDD.n12519 VDD.n6882 133.655
R2033 VDD.n12519 VDD.n6884 133.655
R2034 VDD.n12511 VDD.n6884 133.655
R2035 VDD.n12511 VDD.n6894 133.655
R2036 VDD.n12507 VDD.n6894 133.655
R2037 VDD.n12507 VDD.n6896 133.655
R2038 VDD.n12499 VDD.n6896 133.655
R2039 VDD.n12499 VDD.n6906 133.655
R2040 VDD.n5990 VDD.n5937 133.655
R2041 VDD.n6001 VDD.n5941 133.655
R2042 VDD.n6039 VDD.n6026 133.655
R2043 VDD.n6037 VDD.n6036 133.655
R2044 VDD.n6033 VDD.n6032 133.655
R2045 VDD.n6030 VDD.n6018 133.655
R2046 VDD.n6288 VDD.n6046 133.655
R2047 VDD.n6365 VDD.n5915 133.655
R2048 VDD.n6357 VDD.n5915 133.655
R2049 VDD.n6357 VDD.n5922 133.655
R2050 VDD.n6349 VDD.n5922 133.655
R2051 VDD.n6349 VDD.n5932 133.655
R2052 VDD.n6333 VDD.n6332 133.655
R2053 VDD.n6332 VDD.n6019 133.655
R2054 VDD.n6324 VDD.n6019 133.655
R2055 VDD.n6324 VDD.n6290 133.655
R2056 VDD.n6290 VDD.n6289 133.655
R2057 VDD.n6378 VDD.n5904 133.655
R2058 VDD.n6370 VDD.n5910 133.655
R2059 VDD.n5925 VDD.n5903 133.655
R2060 VDD.n6355 VDD.n5925 133.655
R2061 VDD.n6355 VDD.n5926 133.655
R2062 VDD.n6351 VDD.n5926 133.655
R2063 VDD.n6351 VDD.n5929 133.655
R2064 VDD.n6330 VDD.n6023 133.655
R2065 VDD.n6330 VDD.n6024 133.655
R2066 VDD.n6326 VDD.n6024 133.655
R2067 VDD.n6326 VDD.n6044 133.655
R2068 VDD.n6258 VDD.n6044 133.655
R2069 VDD.n5965 VDD.n5964 133.655
R2070 VDD.n5971 VDD.n5970 133.655
R2071 VDD.n6362 VDD.n5919 133.655
R2072 VDD.n6362 VDD.n5920 133.655
R2073 VDD.n5936 VDD.n5920 133.655
R2074 VDD.n6344 VDD.n5938 133.655
R2075 VDD.n6336 VDD.n5938 133.655
R2076 VDD.n6336 VDD.n6008 133.655
R2077 VDD.n6299 VDD.n6008 133.655
R2078 VDD.n6300 VDD.n6299 133.655
R2079 VDD.n6554 VDD.n5782 133.655
R2080 VDD.n6546 VDD.n6545 133.655
R2081 VDD.n6536 VDD.n6535 133.655
R2082 VDD.n6527 VDD.n5806 133.655
R2083 VDD.n5980 VDD.n5918 133.655
R2084 VDD.n5984 VDD.n5918 133.655
R2085 VDD.n5985 VDD.n5984 133.655
R2086 VDD.n6342 VDD.n5942 133.655
R2087 VDD.n6338 VDD.n5942 133.655
R2088 VDD.n6338 VDD.n6005 133.655
R2089 VDD.n6297 VDD.n6005 133.655
R2090 VDD.n6297 VDD.n6294 133.655
R2091 VDD.n6552 VDD.n5786 133.655
R2092 VDD.n6548 VDD.n5786 133.655
R2093 VDD.n6548 VDD.n5789 133.655
R2094 VDD.n6319 VDD.n5781 133.655
R2095 VDD.n6308 VDD.n5785 133.655
R2096 VDD.n5136 VDD.n5083 133.655
R2097 VDD.n5147 VDD.n5087 133.655
R2098 VDD.n5185 VDD.n5172 133.655
R2099 VDD.n5183 VDD.n5182 133.655
R2100 VDD.n5179 VDD.n5178 133.655
R2101 VDD.n5176 VDD.n5164 133.655
R2102 VDD.n5434 VDD.n5192 133.655
R2103 VDD.n5511 VDD.n5061 133.655
R2104 VDD.n5503 VDD.n5061 133.655
R2105 VDD.n5503 VDD.n5068 133.655
R2106 VDD.n5495 VDD.n5068 133.655
R2107 VDD.n5495 VDD.n5078 133.655
R2108 VDD.n5479 VDD.n5478 133.655
R2109 VDD.n5478 VDD.n5165 133.655
R2110 VDD.n5470 VDD.n5165 133.655
R2111 VDD.n5470 VDD.n5436 133.655
R2112 VDD.n5436 VDD.n5435 133.655
R2113 VDD.n5524 VDD.n5050 133.655
R2114 VDD.n5516 VDD.n5056 133.655
R2115 VDD.n5071 VDD.n5049 133.655
R2116 VDD.n5501 VDD.n5071 133.655
R2117 VDD.n5501 VDD.n5072 133.655
R2118 VDD.n5497 VDD.n5072 133.655
R2119 VDD.n5497 VDD.n5075 133.655
R2120 VDD.n5476 VDD.n5169 133.655
R2121 VDD.n5476 VDD.n5170 133.655
R2122 VDD.n5472 VDD.n5170 133.655
R2123 VDD.n5472 VDD.n5190 133.655
R2124 VDD.n5404 VDD.n5190 133.655
R2125 VDD.n5111 VDD.n5110 133.655
R2126 VDD.n5117 VDD.n5116 133.655
R2127 VDD.n5508 VDD.n5065 133.655
R2128 VDD.n5508 VDD.n5066 133.655
R2129 VDD.n5082 VDD.n5066 133.655
R2130 VDD.n5490 VDD.n5084 133.655
R2131 VDD.n5482 VDD.n5084 133.655
R2132 VDD.n5482 VDD.n5154 133.655
R2133 VDD.n5445 VDD.n5154 133.655
R2134 VDD.n5446 VDD.n5445 133.655
R2135 VDD.n5700 VDD.n4928 133.655
R2136 VDD.n5692 VDD.n5691 133.655
R2137 VDD.n5682 VDD.n5681 133.655
R2138 VDD.n5673 VDD.n4952 133.655
R2139 VDD.n5126 VDD.n5064 133.655
R2140 VDD.n5130 VDD.n5064 133.655
R2141 VDD.n5131 VDD.n5130 133.655
R2142 VDD.n5488 VDD.n5088 133.655
R2143 VDD.n5484 VDD.n5088 133.655
R2144 VDD.n5484 VDD.n5151 133.655
R2145 VDD.n5443 VDD.n5151 133.655
R2146 VDD.n5443 VDD.n5440 133.655
R2147 VDD.n5698 VDD.n4932 133.655
R2148 VDD.n5694 VDD.n4932 133.655
R2149 VDD.n5694 VDD.n4935 133.655
R2150 VDD.n5465 VDD.n4927 133.655
R2151 VDD.n5454 VDD.n4931 133.655
R2152 VDD.n4350 VDD.n4297 133.655
R2153 VDD.n4361 VDD.n4301 133.655
R2154 VDD.n4399 VDD.n4386 133.655
R2155 VDD.n4397 VDD.n4396 133.655
R2156 VDD.n4393 VDD.n4392 133.655
R2157 VDD.n4390 VDD.n4378 133.655
R2158 VDD.n4648 VDD.n4406 133.655
R2159 VDD.n4725 VDD.n4275 133.655
R2160 VDD.n4717 VDD.n4275 133.655
R2161 VDD.n4717 VDD.n4282 133.655
R2162 VDD.n4709 VDD.n4282 133.655
R2163 VDD.n4709 VDD.n4292 133.655
R2164 VDD.n4693 VDD.n4692 133.655
R2165 VDD.n4692 VDD.n4379 133.655
R2166 VDD.n4684 VDD.n4379 133.655
R2167 VDD.n4684 VDD.n4650 133.655
R2168 VDD.n4650 VDD.n4649 133.655
R2169 VDD.n4738 VDD.n4264 133.655
R2170 VDD.n4730 VDD.n4270 133.655
R2171 VDD.n4285 VDD.n4263 133.655
R2172 VDD.n4715 VDD.n4285 133.655
R2173 VDD.n4715 VDD.n4286 133.655
R2174 VDD.n4711 VDD.n4286 133.655
R2175 VDD.n4711 VDD.n4289 133.655
R2176 VDD.n4690 VDD.n4383 133.655
R2177 VDD.n4690 VDD.n4384 133.655
R2178 VDD.n4686 VDD.n4384 133.655
R2179 VDD.n4686 VDD.n4404 133.655
R2180 VDD.n4618 VDD.n4404 133.655
R2181 VDD.n4325 VDD.n4324 133.655
R2182 VDD.n4331 VDD.n4330 133.655
R2183 VDD.n4722 VDD.n4279 133.655
R2184 VDD.n4722 VDD.n4280 133.655
R2185 VDD.n4296 VDD.n4280 133.655
R2186 VDD.n4704 VDD.n4298 133.655
R2187 VDD.n4696 VDD.n4298 133.655
R2188 VDD.n4696 VDD.n4368 133.655
R2189 VDD.n4659 VDD.n4368 133.655
R2190 VDD.n4660 VDD.n4659 133.655
R2191 VDD.n4914 VDD.n4142 133.655
R2192 VDD.n4906 VDD.n4905 133.655
R2193 VDD.n4896 VDD.n4895 133.655
R2194 VDD.n4887 VDD.n4166 133.655
R2195 VDD.n4340 VDD.n4278 133.655
R2196 VDD.n4344 VDD.n4278 133.655
R2197 VDD.n4345 VDD.n4344 133.655
R2198 VDD.n4702 VDD.n4302 133.655
R2199 VDD.n4698 VDD.n4302 133.655
R2200 VDD.n4698 VDD.n4365 133.655
R2201 VDD.n4657 VDD.n4365 133.655
R2202 VDD.n4657 VDD.n4654 133.655
R2203 VDD.n4912 VDD.n4146 133.655
R2204 VDD.n4908 VDD.n4146 133.655
R2205 VDD.n4908 VDD.n4149 133.655
R2206 VDD.n4679 VDD.n4141 133.655
R2207 VDD.n4668 VDD.n4145 133.655
R2208 VDD.n3496 VDD.n3443 133.655
R2209 VDD.n3507 VDD.n3447 133.655
R2210 VDD.n3545 VDD.n3532 133.655
R2211 VDD.n3543 VDD.n3542 133.655
R2212 VDD.n3539 VDD.n3538 133.655
R2213 VDD.n3536 VDD.n3524 133.655
R2214 VDD.n3794 VDD.n3552 133.655
R2215 VDD.n3871 VDD.n3421 133.655
R2216 VDD.n3863 VDD.n3421 133.655
R2217 VDD.n3863 VDD.n3428 133.655
R2218 VDD.n3855 VDD.n3428 133.655
R2219 VDD.n3855 VDD.n3438 133.655
R2220 VDD.n3839 VDD.n3838 133.655
R2221 VDD.n3838 VDD.n3525 133.655
R2222 VDD.n3830 VDD.n3525 133.655
R2223 VDD.n3830 VDD.n3796 133.655
R2224 VDD.n3796 VDD.n3795 133.655
R2225 VDD.n3884 VDD.n3410 133.655
R2226 VDD.n3876 VDD.n3416 133.655
R2227 VDD.n3431 VDD.n3409 133.655
R2228 VDD.n3861 VDD.n3431 133.655
R2229 VDD.n3861 VDD.n3432 133.655
R2230 VDD.n3857 VDD.n3432 133.655
R2231 VDD.n3857 VDD.n3435 133.655
R2232 VDD.n3836 VDD.n3529 133.655
R2233 VDD.n3836 VDD.n3530 133.655
R2234 VDD.n3832 VDD.n3530 133.655
R2235 VDD.n3832 VDD.n3550 133.655
R2236 VDD.n3764 VDD.n3550 133.655
R2237 VDD.n3471 VDD.n3470 133.655
R2238 VDD.n3477 VDD.n3476 133.655
R2239 VDD.n3868 VDD.n3425 133.655
R2240 VDD.n3868 VDD.n3426 133.655
R2241 VDD.n3442 VDD.n3426 133.655
R2242 VDD.n3850 VDD.n3444 133.655
R2243 VDD.n3842 VDD.n3444 133.655
R2244 VDD.n3842 VDD.n3514 133.655
R2245 VDD.n3805 VDD.n3514 133.655
R2246 VDD.n3806 VDD.n3805 133.655
R2247 VDD.n4060 VDD.n3288 133.655
R2248 VDD.n4052 VDD.n4051 133.655
R2249 VDD.n4042 VDD.n4041 133.655
R2250 VDD.n4033 VDD.n3312 133.655
R2251 VDD.n3486 VDD.n3424 133.655
R2252 VDD.n3490 VDD.n3424 133.655
R2253 VDD.n3491 VDD.n3490 133.655
R2254 VDD.n3848 VDD.n3448 133.655
R2255 VDD.n3844 VDD.n3448 133.655
R2256 VDD.n3844 VDD.n3511 133.655
R2257 VDD.n3803 VDD.n3511 133.655
R2258 VDD.n3803 VDD.n3800 133.655
R2259 VDD.n4058 VDD.n3292 133.655
R2260 VDD.n4054 VDD.n3292 133.655
R2261 VDD.n4054 VDD.n3295 133.655
R2262 VDD.n3825 VDD.n3287 133.655
R2263 VDD.n3814 VDD.n3291 133.655
R2264 VDD.n2710 VDD.n2657 133.655
R2265 VDD.n2721 VDD.n2661 133.655
R2266 VDD.n2759 VDD.n2746 133.655
R2267 VDD.n2757 VDD.n2756 133.655
R2268 VDD.n2753 VDD.n2752 133.655
R2269 VDD.n2750 VDD.n2738 133.655
R2270 VDD.n3008 VDD.n2766 133.655
R2271 VDD.n3085 VDD.n2635 133.655
R2272 VDD.n3077 VDD.n2635 133.655
R2273 VDD.n3077 VDD.n2642 133.655
R2274 VDD.n3069 VDD.n2642 133.655
R2275 VDD.n3069 VDD.n2652 133.655
R2276 VDD.n3053 VDD.n3052 133.655
R2277 VDD.n3052 VDD.n2739 133.655
R2278 VDD.n3044 VDD.n2739 133.655
R2279 VDD.n3044 VDD.n3010 133.655
R2280 VDD.n3010 VDD.n3009 133.655
R2281 VDD.n3098 VDD.n2624 133.655
R2282 VDD.n3090 VDD.n2630 133.655
R2283 VDD.n2645 VDD.n2623 133.655
R2284 VDD.n3075 VDD.n2645 133.655
R2285 VDD.n3075 VDD.n2646 133.655
R2286 VDD.n3071 VDD.n2646 133.655
R2287 VDD.n3071 VDD.n2649 133.655
R2288 VDD.n3050 VDD.n2743 133.655
R2289 VDD.n3050 VDD.n2744 133.655
R2290 VDD.n3046 VDD.n2744 133.655
R2291 VDD.n3046 VDD.n2764 133.655
R2292 VDD.n2978 VDD.n2764 133.655
R2293 VDD.n2685 VDD.n2684 133.655
R2294 VDD.n2691 VDD.n2690 133.655
R2295 VDD.n3082 VDD.n2639 133.655
R2296 VDD.n3082 VDD.n2640 133.655
R2297 VDD.n2656 VDD.n2640 133.655
R2298 VDD.n3064 VDD.n2658 133.655
R2299 VDD.n3056 VDD.n2658 133.655
R2300 VDD.n3056 VDD.n2728 133.655
R2301 VDD.n3019 VDD.n2728 133.655
R2302 VDD.n3020 VDD.n3019 133.655
R2303 VDD.n3274 VDD.n2502 133.655
R2304 VDD.n3266 VDD.n3265 133.655
R2305 VDD.n3256 VDD.n3255 133.655
R2306 VDD.n3247 VDD.n2526 133.655
R2307 VDD.n2700 VDD.n2638 133.655
R2308 VDD.n2704 VDD.n2638 133.655
R2309 VDD.n2705 VDD.n2704 133.655
R2310 VDD.n3062 VDD.n2662 133.655
R2311 VDD.n3058 VDD.n2662 133.655
R2312 VDD.n3058 VDD.n2725 133.655
R2313 VDD.n3017 VDD.n2725 133.655
R2314 VDD.n3017 VDD.n3014 133.655
R2315 VDD.n3272 VDD.n2506 133.655
R2316 VDD.n3268 VDD.n2506 133.655
R2317 VDD.n3268 VDD.n2509 133.655
R2318 VDD.n3039 VDD.n2501 133.655
R2319 VDD.n3028 VDD.n2505 133.655
R2320 VDD.n1855 VDD.n1802 133.655
R2321 VDD.n1866 VDD.n1806 133.655
R2322 VDD.n1904 VDD.n1891 133.655
R2323 VDD.n1902 VDD.n1901 133.655
R2324 VDD.n1898 VDD.n1897 133.655
R2325 VDD.n1895 VDD.n1883 133.655
R2326 VDD.n2153 VDD.n1911 133.655
R2327 VDD.n2230 VDD.n1780 133.655
R2328 VDD.n2222 VDD.n1780 133.655
R2329 VDD.n2222 VDD.n1787 133.655
R2330 VDD.n2214 VDD.n1787 133.655
R2331 VDD.n2214 VDD.n1797 133.655
R2332 VDD.n2198 VDD.n2197 133.655
R2333 VDD.n2197 VDD.n1884 133.655
R2334 VDD.n2189 VDD.n1884 133.655
R2335 VDD.n2189 VDD.n2155 133.655
R2336 VDD.n2155 VDD.n2154 133.655
R2337 VDD.n2243 VDD.n1769 133.655
R2338 VDD.n2235 VDD.n1775 133.655
R2339 VDD.n1790 VDD.n1768 133.655
R2340 VDD.n2220 VDD.n1790 133.655
R2341 VDD.n2220 VDD.n1791 133.655
R2342 VDD.n2216 VDD.n1791 133.655
R2343 VDD.n2216 VDD.n1794 133.655
R2344 VDD.n2195 VDD.n1888 133.655
R2345 VDD.n2195 VDD.n1889 133.655
R2346 VDD.n2191 VDD.n1889 133.655
R2347 VDD.n2191 VDD.n1909 133.655
R2348 VDD.n2123 VDD.n1909 133.655
R2349 VDD.n1830 VDD.n1829 133.655
R2350 VDD.n1836 VDD.n1835 133.655
R2351 VDD.n2227 VDD.n1784 133.655
R2352 VDD.n2227 VDD.n1785 133.655
R2353 VDD.n1801 VDD.n1785 133.655
R2354 VDD.n2209 VDD.n1803 133.655
R2355 VDD.n2201 VDD.n1803 133.655
R2356 VDD.n2201 VDD.n1873 133.655
R2357 VDD.n2164 VDD.n1873 133.655
R2358 VDD.n2165 VDD.n2164 133.655
R2359 VDD.n2419 VDD.n1647 133.655
R2360 VDD.n2411 VDD.n2410 133.655
R2361 VDD.n2401 VDD.n2400 133.655
R2362 VDD.n2392 VDD.n1671 133.655
R2363 VDD.n1845 VDD.n1783 133.655
R2364 VDD.n1849 VDD.n1783 133.655
R2365 VDD.n1850 VDD.n1849 133.655
R2366 VDD.n2207 VDD.n1807 133.655
R2367 VDD.n2203 VDD.n1807 133.655
R2368 VDD.n2203 VDD.n1870 133.655
R2369 VDD.n2162 VDD.n1870 133.655
R2370 VDD.n2162 VDD.n2159 133.655
R2371 VDD.n2417 VDD.n1651 133.655
R2372 VDD.n2413 VDD.n1651 133.655
R2373 VDD.n2413 VDD.n1654 133.655
R2374 VDD.n2184 VDD.n1646 133.655
R2375 VDD.n2173 VDD.n1650 133.655
R2376 VDD.n1259 VDD.n1255 133.655
R2377 VDD.n1514 VDD.n1513 133.655
R2378 VDD.n860 VDD.n859 133.655
R2379 VDD.n1242 VDD.n1241 133.655
R2380 VDD.n1213 VDD.n1210 133.655
R2381 VDD.n1129 VDD.n1128 133.655
R2382 VDD.n31 VDD.n27 133.655
R2383 VDD.n286 VDD.n285 133.655
R2384 VDD.n414 VDD.n413 133.655
R2385 VDD.n14 VDD.n13 133.655
R2386 VDD.n767 VDD.n764 133.655
R2387 VDD.n683 VDD.n682 133.655
R2388 VDD.n6152 VDD.n6106 128.696
R2389 VDD.n5298 VDD.n5252 128.696
R2390 VDD.n4512 VDD.n4466 128.696
R2391 VDD.n3658 VDD.n3612 128.696
R2392 VDD.n2872 VDD.n2826 128.696
R2393 VDD.n2017 VDD.n1971 128.696
R2394 VDD.n9221 VDD.t37 126.425
R2395 VDD.n6222 VDD.n6221 126.356
R2396 VDD.n5368 VDD.n5367 126.356
R2397 VDD.n4582 VDD.n4581 126.356
R2398 VDD.n3728 VDD.n3727 126.356
R2399 VDD.n2942 VDD.n2941 126.356
R2400 VDD.n2087 VDD.n2086 126.356
R2401 VDD.n12249 VDD.n12248 123.651
R2402 VDD.n9963 VDD.t195 117.838
R2403 VDD.t187 VDD.n5763 117.838
R2404 VDD.t73 VDD.n4123 117.838
R2405 VDD.t164 VDD.n2483 117.838
R2406 VDD.t204 VDD.n843 117.838
R2407 VDD.n11650 VDD.n7611 117.62
R2408 VDD.n10042 VDD.t149 116.841
R2409 VDD.n10601 VDD.t151 116.841
R2410 VDD.n9369 VDD.t47 116.841
R2411 VDD.t29 VDD.n10540 116.841
R2412 VDD.t35 VDD.n9635 116.841
R2413 VDD.n10733 VDD.t39 116.841
R2414 VDD.t41 VDD.n8887 116.841
R2415 VDD.t195 VDD.t132 112.624
R2416 VDD.n12405 VDD.n6936 104.757
R2417 VDD.n12405 VDD.n6937 104.757
R2418 VDD.n12401 VDD.n6937 104.757
R2419 VDD.n12401 VDD.n6941 104.757
R2420 VDD.n12394 VDD.n6941 104.757
R2421 VDD.n12394 VDD.n6948 104.757
R2422 VDD.n12390 VDD.n6948 104.757
R2423 VDD.n12390 VDD.n6950 104.757
R2424 VDD.n12383 VDD.n6950 104.757
R2425 VDD.n12383 VDD.n6957 104.757
R2426 VDD.n12379 VDD.n6957 104.757
R2427 VDD.n12379 VDD.n6959 104.757
R2428 VDD.n12372 VDD.n6959 104.757
R2429 VDD.n12372 VDD.n6966 104.757
R2430 VDD.n12368 VDD.n6966 104.757
R2431 VDD.n12368 VDD.n6969 104.757
R2432 VDD.n12361 VDD.n6969 104.757
R2433 VDD.n12361 VDD.n6976 104.757
R2434 VDD.n12357 VDD.n6976 104.757
R2435 VDD.n12357 VDD.n6978 104.757
R2436 VDD.n12350 VDD.n6978 104.757
R2437 VDD.n12350 VDD.n6983 104.757
R2438 VDD.n12346 VDD.n6983 104.757
R2439 VDD.n12346 VDD.n6985 104.757
R2440 VDD.n12339 VDD.n6985 104.757
R2441 VDD.n12339 VDD.n6992 104.757
R2442 VDD.n12335 VDD.n6992 104.757
R2443 VDD.n12335 VDD.n6994 104.757
R2444 VDD.n12328 VDD.n6994 104.757
R2445 VDD.n12328 VDD.n7001 104.757
R2446 VDD.n12324 VDD.n7001 104.757
R2447 VDD.n12324 VDD.n7003 104.757
R2448 VDD.n12317 VDD.n7003 104.757
R2449 VDD.n12317 VDD.n7010 104.757
R2450 VDD.n12313 VDD.n7010 104.757
R2451 VDD.n12313 VDD.n7012 104.757
R2452 VDD.n7019 VDD.n7012 104.757
R2453 VDD.n12305 VDD.n7019 104.757
R2454 VDD.n12305 VDD.n7020 104.757
R2455 VDD.n12301 VDD.n7020 104.757
R2456 VDD.n12301 VDD.n7023 104.757
R2457 VDD.n12294 VDD.n7023 104.757
R2458 VDD.n12294 VDD.n7030 104.757
R2459 VDD.n12290 VDD.n7030 104.757
R2460 VDD.n12290 VDD.n7032 104.757
R2461 VDD.n12283 VDD.n7032 104.757
R2462 VDD.n12283 VDD.n7039 104.757
R2463 VDD.n12279 VDD.n7039 104.757
R2464 VDD.n12279 VDD.n7041 104.757
R2465 VDD.n12272 VDD.n7041 104.757
R2466 VDD.n12272 VDD.n7048 104.757
R2467 VDD.n12268 VDD.n7048 104.757
R2468 VDD.n12268 VDD.n7050 104.757
R2469 VDD.n7058 VDD.n7050 104.757
R2470 VDD.n12261 VDD.n7058 104.757
R2471 VDD.n12261 VDD.n7059 104.757
R2472 VDD.n12257 VDD.n7059 104.757
R2473 VDD.n12257 VDD.n7062 104.757
R2474 VDD.n12250 VDD.n7062 104.757
R2475 VDD.n12250 VDD.n7069 104.757
R2476 VDD.n7134 VDD.n7132 104.757
R2477 VDD.n7141 VDD.n7123 104.757
R2478 VDD.n7144 VDD.n7143 104.757
R2479 VDD.n7153 VDD.n7151 104.757
R2480 VDD.n7161 VDD.n7115 104.757
R2481 VDD.n7165 VDD.n7163 104.757
R2482 VDD.n7172 VDD.n7111 104.757
R2483 VDD.n7175 VDD.n7174 104.757
R2484 VDD.n7184 VDD.n7182 104.757
R2485 VDD.n7191 VDD.n7103 104.757
R2486 VDD.n7194 VDD.n7193 104.757
R2487 VDD.n7203 VDD.n7201 104.757
R2488 VDD.n7210 VDD.n7095 104.757
R2489 VDD.n7214 VDD.n7213 104.757
R2490 VDD.n7222 VDD.n7091 104.757
R2491 VDD.n7225 VDD.n7224 104.757
R2492 VDD.n7234 VDD.n7232 104.757
R2493 VDD.n7241 VDD.n7083 104.757
R2494 VDD.n7244 VDD.n7243 104.757
R2495 VDD.n7253 VDD.n7251 104.757
R2496 VDD.n12246 VDD.n7073 104.757
R2497 VDD.n12246 VDD.n7074 104.757
R2498 VDD.n12239 VDD.n7074 104.757
R2499 VDD.n12239 VDD.n7261 104.757
R2500 VDD.n12235 VDD.n7261 104.757
R2501 VDD.n12235 VDD.n7263 104.757
R2502 VDD.n7271 VDD.n7263 104.757
R2503 VDD.n12228 VDD.n7271 104.757
R2504 VDD.n12228 VDD.n7272 104.757
R2505 VDD.n12224 VDD.n7272 104.757
R2506 VDD.n12224 VDD.n7275 104.757
R2507 VDD.n12217 VDD.n7275 104.757
R2508 VDD.n12217 VDD.n7282 104.757
R2509 VDD.n12213 VDD.n7282 104.757
R2510 VDD.n12213 VDD.n7284 104.757
R2511 VDD.n12206 VDD.n7284 104.757
R2512 VDD.n12206 VDD.n7291 104.757
R2513 VDD.n12202 VDD.n7291 104.757
R2514 VDD.n12202 VDD.n7293 104.757
R2515 VDD.n12195 VDD.n7293 104.757
R2516 VDD.n12195 VDD.n7300 104.757
R2517 VDD.n12191 VDD.n7300 104.757
R2518 VDD.n12191 VDD.n7302 104.757
R2519 VDD.n12184 VDD.n7302 104.757
R2520 VDD.n12184 VDD.n7309 104.757
R2521 VDD.n12180 VDD.n7309 104.757
R2522 VDD.n12180 VDD.n7311 104.757
R2523 VDD.n12173 VDD.n7311 104.757
R2524 VDD.n12173 VDD.n7316 104.757
R2525 VDD.n12169 VDD.n7316 104.757
R2526 VDD.n12169 VDD.n7318 104.757
R2527 VDD.n12162 VDD.n7318 104.757
R2528 VDD.n12162 VDD.n7325 104.757
R2529 VDD.n12158 VDD.n7325 104.757
R2530 VDD.n12158 VDD.n7327 104.757
R2531 VDD.n12151 VDD.n7327 104.757
R2532 VDD.n12151 VDD.n7334 104.757
R2533 VDD.n12147 VDD.n7334 104.757
R2534 VDD.n12147 VDD.n7336 104.757
R2535 VDD.n12140 VDD.n7336 104.757
R2536 VDD.n12140 VDD.n7343 104.757
R2537 VDD.n12136 VDD.n7343 104.757
R2538 VDD.n12136 VDD.n7345 104.757
R2539 VDD.n7352 VDD.n7345 104.757
R2540 VDD.n12128 VDD.n7353 104.757
R2541 VDD.n12124 VDD.n7353 104.757
R2542 VDD.n12124 VDD.n7356 104.757
R2543 VDD.n12120 VDD.n7356 104.757
R2544 VDD.n12120 VDD.n7358 104.757
R2545 VDD.n12116 VDD.n7358 104.757
R2546 VDD.n12116 VDD.n7360 104.757
R2547 VDD.n12112 VDD.n7360 104.757
R2548 VDD.n12112 VDD.n7362 104.757
R2549 VDD.n12108 VDD.n7362 104.757
R2550 VDD.n12108 VDD.n7364 104.757
R2551 VDD.n12104 VDD.n7364 104.757
R2552 VDD.n12104 VDD.n7366 104.757
R2553 VDD.n12100 VDD.n7366 104.757
R2554 VDD.n12100 VDD.n7368 104.757
R2555 VDD.n12096 VDD.n7368 104.757
R2556 VDD.n12096 VDD.n7370 104.757
R2557 VDD.n11653 VDD.n7610 104.757
R2558 VDD.n11653 VDD.n7605 104.757
R2559 VDD.n11662 VDD.n7605 104.757
R2560 VDD.n11662 VDD.n7603 104.757
R2561 VDD.n11666 VDD.n7603 104.757
R2562 VDD.n11666 VDD.n7599 104.757
R2563 VDD.n11674 VDD.n7599 104.757
R2564 VDD.n11674 VDD.n7597 104.757
R2565 VDD.n11678 VDD.n7597 104.757
R2566 VDD.n11678 VDD.n7591 104.757
R2567 VDD.n11686 VDD.n7591 104.757
R2568 VDD.n11686 VDD.n7589 104.757
R2569 VDD.n11690 VDD.n7589 104.757
R2570 VDD.n11690 VDD.n7584 104.757
R2571 VDD.n11699 VDD.n7584 104.757
R2572 VDD.n11699 VDD.n7582 104.757
R2573 VDD.n11703 VDD.n7582 104.757
R2574 VDD.n11703 VDD.n7577 104.757
R2575 VDD.n11712 VDD.n7577 104.757
R2576 VDD.n11712 VDD.n7575 104.757
R2577 VDD.n11716 VDD.n7575 104.757
R2578 VDD.n11716 VDD.n7570 104.757
R2579 VDD.n11725 VDD.n7570 104.757
R2580 VDD.n11725 VDD.n7568 104.757
R2581 VDD.n11729 VDD.n7568 104.757
R2582 VDD.n11729 VDD.n7564 104.757
R2583 VDD.n11737 VDD.n7564 104.757
R2584 VDD.n11737 VDD.n7562 104.757
R2585 VDD.n11741 VDD.n7562 104.757
R2586 VDD.n11741 VDD.n7557 104.757
R2587 VDD.n11750 VDD.n7557 104.757
R2588 VDD.n11750 VDD.n7555 104.757
R2589 VDD.n11754 VDD.n7555 104.757
R2590 VDD.n11754 VDD.n7550 104.757
R2591 VDD.n11763 VDD.n7550 104.757
R2592 VDD.n11763 VDD.n7548 104.757
R2593 VDD.n11767 VDD.n7548 104.757
R2594 VDD.n11767 VDD.n7543 104.757
R2595 VDD.n11776 VDD.n7543 104.757
R2596 VDD.n11776 VDD.n7541 104.757
R2597 VDD.n11780 VDD.n7541 104.757
R2598 VDD.n11780 VDD.n7537 104.757
R2599 VDD.n11788 VDD.n7537 104.757
R2600 VDD.n11788 VDD.n7535 104.757
R2601 VDD.n11792 VDD.n7535 104.757
R2602 VDD.n11792 VDD.n7529 104.757
R2603 VDD.n11800 VDD.n7529 104.757
R2604 VDD.n11800 VDD.n7527 104.757
R2605 VDD.n11804 VDD.n7527 104.757
R2606 VDD.n11804 VDD.n7522 104.757
R2607 VDD.n11813 VDD.n7522 104.757
R2608 VDD.n11813 VDD.n7520 104.757
R2609 VDD.n11817 VDD.n7520 104.757
R2610 VDD.n11817 VDD.n7515 104.757
R2611 VDD.n11826 VDD.n7515 104.757
R2612 VDD.n11826 VDD.n7513 104.757
R2613 VDD.n11830 VDD.n7513 104.757
R2614 VDD.n11830 VDD.n7508 104.757
R2615 VDD.n11839 VDD.n7508 104.757
R2616 VDD.n11839 VDD.n7506 104.757
R2617 VDD.n11843 VDD.n7506 104.757
R2618 VDD.n11843 VDD.n7502 104.757
R2619 VDD.n11851 VDD.n7502 104.757
R2620 VDD.n11851 VDD.n7500 104.757
R2621 VDD.n11855 VDD.n7500 104.757
R2622 VDD.n11855 VDD.n7495 104.757
R2623 VDD.n11864 VDD.n7495 104.757
R2624 VDD.n11864 VDD.n7493 104.757
R2625 VDD.n11868 VDD.n7493 104.757
R2626 VDD.n11868 VDD.n7488 104.757
R2627 VDD.n11877 VDD.n7488 104.757
R2628 VDD.n11877 VDD.n7486 104.757
R2629 VDD.n11881 VDD.n7486 104.757
R2630 VDD.n11881 VDD.n7481 104.757
R2631 VDD.n11890 VDD.n7481 104.757
R2632 VDD.n11890 VDD.n7479 104.757
R2633 VDD.n11894 VDD.n7479 104.757
R2634 VDD.n11894 VDD.n7475 104.757
R2635 VDD.n11902 VDD.n7475 104.757
R2636 VDD.n11902 VDD.n7473 104.757
R2637 VDD.n11906 VDD.n7473 104.757
R2638 VDD.n11906 VDD.n7467 104.757
R2639 VDD.n11914 VDD.n7467 104.757
R2640 VDD.n11914 VDD.n7465 104.757
R2641 VDD.n11918 VDD.n7465 104.757
R2642 VDD.n11918 VDD.n7460 104.757
R2643 VDD.n11927 VDD.n7460 104.757
R2644 VDD.n11927 VDD.n7458 104.757
R2645 VDD.n11931 VDD.n7458 104.757
R2646 VDD.n11931 VDD.n7453 104.757
R2647 VDD.n11940 VDD.n7453 104.757
R2648 VDD.n11940 VDD.n7451 104.757
R2649 VDD.n11944 VDD.n7451 104.757
R2650 VDD.n11944 VDD.n7446 104.757
R2651 VDD.n11953 VDD.n7446 104.757
R2652 VDD.n11953 VDD.n7444 104.757
R2653 VDD.n11957 VDD.n7444 104.757
R2654 VDD.n11957 VDD.n7440 104.757
R2655 VDD.n11965 VDD.n7440 104.757
R2656 VDD.n11965 VDD.n7438 104.757
R2657 VDD.n11969 VDD.n7438 104.757
R2658 VDD.n11969 VDD.n7433 104.757
R2659 VDD.n11978 VDD.n7433 104.757
R2660 VDD.n11978 VDD.n7431 104.757
R2661 VDD.n11982 VDD.n7431 104.757
R2662 VDD.n11982 VDD.n7426 104.757
R2663 VDD.n11991 VDD.n7426 104.757
R2664 VDD.n11991 VDD.n7424 104.757
R2665 VDD.n11995 VDD.n7424 104.757
R2666 VDD.n11995 VDD.n7419 104.757
R2667 VDD.n12004 VDD.n7419 104.757
R2668 VDD.n12004 VDD.n7417 104.757
R2669 VDD.n12008 VDD.n7417 104.757
R2670 VDD.n12008 VDD.n7413 104.757
R2671 VDD.n12016 VDD.n7413 104.757
R2672 VDD.n12016 VDD.n7411 104.757
R2673 VDD.n12020 VDD.n7411 104.757
R2674 VDD.n12020 VDD.n7405 104.757
R2675 VDD.n12028 VDD.n7405 104.757
R2676 VDD.n12028 VDD.n7403 104.757
R2677 VDD.n12032 VDD.n7403 104.757
R2678 VDD.n12032 VDD.n7398 104.757
R2679 VDD.n12041 VDD.n7398 104.757
R2680 VDD.n12041 VDD.n7396 104.757
R2681 VDD.n12045 VDD.n7396 104.757
R2682 VDD.n12045 VDD.n7391 104.757
R2683 VDD.n12054 VDD.n7391 104.757
R2684 VDD.n12054 VDD.n7389 104.757
R2685 VDD.n12058 VDD.n7389 104.757
R2686 VDD.n12058 VDD.n7384 104.757
R2687 VDD.n12067 VDD.n7384 104.757
R2688 VDD.n12067 VDD.n7382 104.757
R2689 VDD.n12071 VDD.n7382 104.757
R2690 VDD.n12071 VDD.n7378 104.757
R2691 VDD.n12082 VDD.n7378 104.757
R2692 VDD.n12082 VDD.n7375 104.757
R2693 VDD.n12086 VDD.n7375 104.757
R2694 VDD.n12087 VDD.n12086 104.757
R2695 VDD.n7835 VDD.n7831 104.757
R2696 VDD.n7947 VDD.n7835 104.757
R2697 VDD.n7945 VDD.n7836 104.757
R2698 VDD.n7938 VDD.n7937 104.757
R2699 VDD.n7935 VDD.n7842 104.757
R2700 VDD.n7901 VDD.n7866 104.757
R2701 VDD.n7899 VDD.n7868 104.757
R2702 VDD.n7892 VDD.n7891 104.757
R2703 VDD.n7889 VDD.n7874 104.757
R2704 VDD.n7882 VDD.n7717 104.757
R2705 VDD.n11451 VDD.n7717 104.757
R2706 VDD.n11451 VDD.n7712 104.757
R2707 VDD.n11460 VDD.n7712 104.757
R2708 VDD.n11460 VDD.n7710 104.757
R2709 VDD.n11464 VDD.n7710 104.757
R2710 VDD.n11464 VDD.n7706 104.757
R2711 VDD.n11472 VDD.n7706 104.757
R2712 VDD.n11472 VDD.n7704 104.757
R2713 VDD.n11476 VDD.n7704 104.757
R2714 VDD.n11476 VDD.n7699 104.757
R2715 VDD.n11484 VDD.n7699 104.757
R2716 VDD.n11484 VDD.n7697 104.757
R2717 VDD.n11488 VDD.n7697 104.757
R2718 VDD.n11488 VDD.n7692 104.757
R2719 VDD.n11497 VDD.n7692 104.757
R2720 VDD.n11497 VDD.n7690 104.757
R2721 VDD.n11501 VDD.n7690 104.757
R2722 VDD.n11501 VDD.n7685 104.757
R2723 VDD.n11510 VDD.n7685 104.757
R2724 VDD.n11510 VDD.n7683 104.757
R2725 VDD.n11514 VDD.n7683 104.757
R2726 VDD.n11514 VDD.n7678 104.757
R2727 VDD.n11523 VDD.n7678 104.757
R2728 VDD.n11523 VDD.n7676 104.757
R2729 VDD.n11527 VDD.n7676 104.757
R2730 VDD.n11527 VDD.n7671 104.757
R2731 VDD.n11533 VDD.n7671 104.757
R2732 VDD.n11533 VDD.n7669 104.757
R2733 VDD.n11537 VDD.n7669 104.757
R2734 VDD.n11537 VDD.n7664 104.757
R2735 VDD.n11546 VDD.n7664 104.757
R2736 VDD.n11546 VDD.n7662 104.757
R2737 VDD.n11550 VDD.n7662 104.757
R2738 VDD.n11550 VDD.n7657 104.757
R2739 VDD.n11559 VDD.n7657 104.757
R2740 VDD.n11559 VDD.n7655 104.757
R2741 VDD.n11563 VDD.n7655 104.757
R2742 VDD.n11563 VDD.n7650 104.757
R2743 VDD.n11572 VDD.n7650 104.757
R2744 VDD.n11572 VDD.n7648 104.757
R2745 VDD.n11576 VDD.n7648 104.757
R2746 VDD.n11576 VDD.n7644 104.757
R2747 VDD.n11584 VDD.n7644 104.757
R2748 VDD.n11588 VDD.n7642 104.757
R2749 VDD.n11588 VDD.n7637 104.757
R2750 VDD.n11597 VDD.n7637 104.757
R2751 VDD.n11597 VDD.n7635 104.757
R2752 VDD.n11601 VDD.n7635 104.757
R2753 VDD.n11601 VDD.n7630 104.757
R2754 VDD.n11610 VDD.n7630 104.757
R2755 VDD.n11610 VDD.n7628 104.757
R2756 VDD.n11614 VDD.n7628 104.757
R2757 VDD.n11614 VDD.n7623 104.757
R2758 VDD.n11623 VDD.n7623 104.757
R2759 VDD.n11623 VDD.n7621 104.757
R2760 VDD.n11627 VDD.n7621 104.757
R2761 VDD.n11627 VDD.n7616 104.757
R2762 VDD.n11638 VDD.n7616 104.757
R2763 VDD.n11638 VDD.n7614 104.757
R2764 VDD.n11642 VDD.n7614 104.757
R2765 VDD.n8536 VDD.n8535 104.757
R2766 VDD.n8528 VDD.n7792 104.757
R2767 VDD.n8526 VDD.n7793 104.757
R2768 VDD.n8519 VDD.n8518 104.757
R2769 VDD.n8516 VDD.n7798 104.757
R2770 VDD.n8509 VDD.n8508 104.757
R2771 VDD.n8501 VDD.n7808 104.757
R2772 VDD.n8501 VDD.n8500 104.757
R2773 VDD.n8121 VDD.n8088 104.757
R2774 VDD.n8199 VDD.n8088 104.757
R2775 VDD.n8200 VDD.n8199 104.757
R2776 VDD.n8200 VDD.n8082 104.757
R2777 VDD.n8212 VDD.n8082 104.757
R2778 VDD.n8212 VDD.n8075 104.757
R2779 VDD.n8220 VDD.n8075 104.757
R2780 VDD.n8220 VDD.n8066 104.757
R2781 VDD.n8231 VDD.n8066 104.757
R2782 VDD.n8232 VDD.n8231 104.757
R2783 VDD.n8232 VDD.n8060 104.757
R2784 VDD.n8244 VDD.n8060 104.757
R2785 VDD.n8244 VDD.n8054 104.757
R2786 VDD.n8256 VDD.n8054 104.757
R2787 VDD.n8256 VDD.n8047 104.757
R2788 VDD.n8264 VDD.n8047 104.757
R2789 VDD.n8264 VDD.n8038 104.757
R2790 VDD.n8275 VDD.n8038 104.757
R2791 VDD.n8276 VDD.n8275 104.757
R2792 VDD.n8276 VDD.n8031 104.757
R2793 VDD.n8287 VDD.n8031 104.757
R2794 VDD.n8287 VDD.n8024 104.757
R2795 VDD.n8295 VDD.n8024 104.757
R2796 VDD.n8295 VDD.n8015 104.757
R2797 VDD.n8306 VDD.n8015 104.757
R2798 VDD.n8307 VDD.n8306 104.757
R2799 VDD.n8307 VDD.n8009 104.757
R2800 VDD.n8319 VDD.n8009 104.757
R2801 VDD.n8319 VDD.n8003 104.757
R2802 VDD.n8331 VDD.n8003 104.757
R2803 VDD.n8331 VDD.n7990 104.757
R2804 VDD.n8496 VDD.n7990 104.757
R2805 VDD.n8496 VDD.n7991 104.757
R2806 VDD.n8486 VDD.n7991 104.757
R2807 VDD.n8486 VDD.n8485 104.757
R2808 VDD.n8485 VDD.n8341 104.757
R2809 VDD.n8357 VDD.n8341 104.757
R2810 VDD.n8471 VDD.n8357 104.757
R2811 VDD.n8471 VDD.n8470 104.757
R2812 VDD.n8470 VDD.n8358 104.757
R2813 VDD.n8373 VDD.n8358 104.757
R2814 VDD.n8457 VDD.n8373 104.757
R2815 VDD.n8457 VDD.n8456 104.757
R2816 VDD.n8456 VDD.n8374 104.757
R2817 VDD.n8390 VDD.n8374 104.757
R2818 VDD.n8442 VDD.n8390 104.757
R2819 VDD.n8442 VDD.n8441 104.757
R2820 VDD.n8441 VDD.n8391 104.757
R2821 VDD.n8407 VDD.n8391 104.757
R2822 VDD.n8427 VDD.n8407 104.757
R2823 VDD.n8427 VDD.n8426 104.757
R2824 VDD.n8426 VDD.n8408 104.757
R2825 VDD.n8408 VDD.n7765 104.757
R2826 VDD.n8566 VDD.n7765 104.757
R2827 VDD.n8566 VDD.n7766 104.757
R2828 VDD.n8559 VDD.n7766 104.757
R2829 VDD.n8559 VDD.n8558 104.757
R2830 VDD.n8558 VDD.n7771 104.757
R2831 VDD.n8554 VDD.n7771 104.757
R2832 VDD.n8554 VDD.n7774 104.757
R2833 VDD.n8547 VDD.n7774 104.757
R2834 VDD.n8547 VDD.n7781 104.757
R2835 VDD.n8543 VDD.n7781 104.757
R2836 VDD.n8116 VDD.n8115 104.757
R2837 VDD.n8188 VDD.n8111 104.757
R2838 VDD.n8186 VDD.n8126 104.757
R2839 VDD.n8177 VDD.n8176 104.757
R2840 VDD.n8167 VDD.n8143 104.757
R2841 VDD.n8165 VDD.n8144 104.757
R2842 VDD.n8155 VDD.n8153 104.757
R2843 VDD.n8155 VDD.n8154 104.757
R2844 VDD.n8154 VDD.n7720 104.757
R2845 VDD.n11446 VDD.n7720 104.757
R2846 VDD.n11446 VDD.n7721 104.757
R2847 VDD.n8612 VDD.n7721 104.757
R2848 VDD.n8613 VDD.n8612 104.757
R2849 VDD.n8614 VDD.n8613 104.757
R2850 VDD.n11427 VDD.n8614 104.757
R2851 VDD.n11427 VDD.n8615 104.757
R2852 VDD.n8643 VDD.n8615 104.757
R2853 VDD.n8644 VDD.n8643 104.757
R2854 VDD.n8645 VDD.n8644 104.757
R2855 VDD.n11408 VDD.n8645 104.757
R2856 VDD.n11408 VDD.n8646 104.757
R2857 VDD.n8675 VDD.n8646 104.757
R2858 VDD.n8675 VDD.n8664 104.757
R2859 VDD.n11393 VDD.n8664 104.757
R2860 VDD.n11393 VDD.n11392 104.757
R2861 VDD.n11392 VDD.n8665 104.757
R2862 VDD.n11383 VDD.n8665 104.757
R2863 VDD.n11383 VDD.n8684 104.757
R2864 VDD.n8715 VDD.n8684 104.757
R2865 VDD.n8716 VDD.n8715 104.757
R2866 VDD.n8717 VDD.n8716 104.757
R2867 VDD.n11364 VDD.n8717 104.757
R2868 VDD.n11364 VDD.n8718 104.757
R2869 VDD.n11048 VDD.n8718 104.757
R2870 VDD.n11049 VDD.n11048 104.757
R2871 VDD.n11050 VDD.n11049 104.757
R2872 VDD.n11345 VDD.n11050 104.757
R2873 VDD.n11345 VDD.n11051 104.757
R2874 VDD.n11097 VDD.n11051 104.757
R2875 VDD.n11098 VDD.n11097 104.757
R2876 VDD.n11099 VDD.n11098 104.757
R2877 VDD.n11100 VDD.n11099 104.757
R2878 VDD.n11101 VDD.n11100 104.757
R2879 VDD.n11102 VDD.n11101 104.757
R2880 VDD.n11103 VDD.n11102 104.757
R2881 VDD.n11311 VDD.n11103 104.757
R2882 VDD.n11311 VDD.n11104 104.757
R2883 VDD.n11132 VDD.n11104 104.757
R2884 VDD.n11133 VDD.n11132 104.757
R2885 VDD.n11134 VDD.n11133 104.757
R2886 VDD.n11292 VDD.n11134 104.757
R2887 VDD.n11292 VDD.n11135 104.757
R2888 VDD.n11163 VDD.n11135 104.757
R2889 VDD.n11164 VDD.n11163 104.757
R2890 VDD.n11165 VDD.n11164 104.757
R2891 VDD.n11273 VDD.n11165 104.757
R2892 VDD.n11273 VDD.n11166 104.757
R2893 VDD.n11196 VDD.n11166 104.757
R2894 VDD.n11196 VDD.n11185 104.757
R2895 VDD.n11258 VDD.n11185 104.757
R2896 VDD.n11258 VDD.n11257 104.757
R2897 VDD.n11257 VDD.n11186 104.757
R2898 VDD.n11248 VDD.n11186 104.757
R2899 VDD.n11248 VDD.n11205 104.757
R2900 VDD.n11215 VDD.n11205 104.757
R2901 VDD.n11231 VDD.n11215 104.757
R2902 VDD.n11231 VDD.n11221 104.757
R2903 VDD.n11221 VDD.n11220 104.757
R2904 VDD.n11220 VDD.n11219 104.757
R2905 VDD.n11216 VDD.n6620 104.757
R2906 VDD.n12696 VDD.n12695 104.757
R2907 VDD.n12695 VDD.n6614 104.757
R2908 VDD.n12689 VDD.n6614 104.757
R2909 VDD.n12689 VDD.n6703 104.757
R2910 VDD.n12682 VDD.n6703 104.757
R2911 VDD.n12682 VDD.n6711 104.757
R2912 VDD.n10257 VDD.n6711 104.757
R2913 VDD.n10258 VDD.n10257 104.757
R2914 VDD.n10258 VDD.n10249 104.757
R2915 VDD.n10265 VDD.n10249 104.757
R2916 VDD.n10266 VDD.n10265 104.757
R2917 VDD.n10266 VDD.n10245 104.757
R2918 VDD.n10273 VDD.n10245 104.757
R2919 VDD.n10274 VDD.n10273 104.757
R2920 VDD.n10274 VDD.n10239 104.757
R2921 VDD.n10282 VDD.n10239 104.757
R2922 VDD.n10283 VDD.n10282 104.757
R2923 VDD.n10284 VDD.n10283 104.757
R2924 VDD.n10284 VDD.n10235 104.757
R2925 VDD.n10291 VDD.n10235 104.757
R2926 VDD.n10292 VDD.n10291 104.757
R2927 VDD.n10292 VDD.n10231 104.757
R2928 VDD.n10299 VDD.n10231 104.757
R2929 VDD.n10300 VDD.n10299 104.757
R2930 VDD.n10300 VDD.n10227 104.757
R2931 VDD.n10307 VDD.n10227 104.757
R2932 VDD.n10308 VDD.n10307 104.757
R2933 VDD.n10308 VDD.n10221 104.757
R2934 VDD.n10315 VDD.n10221 104.757
R2935 VDD.n10316 VDD.n10315 104.757
R2936 VDD.n10316 VDD.n10217 104.757
R2937 VDD.n10323 VDD.n10217 104.757
R2938 VDD.n10324 VDD.n10323 104.757
R2939 VDD.n10324 VDD.n10213 104.757
R2940 VDD.n10333 VDD.n10213 104.757
R2941 VDD.n10336 VDD.n10333 104.757
R2942 VDD.n10337 VDD.n10336 104.757
R2943 VDD.n10337 VDD.n10206 104.757
R2944 VDD.n10344 VDD.n10206 104.757
R2945 VDD.n10345 VDD.n10344 104.757
R2946 VDD.n10345 VDD.n10202 104.757
R2947 VDD.n10352 VDD.n10202 104.757
R2948 VDD.n10353 VDD.n10352 104.757
R2949 VDD.n10353 VDD.n10198 104.757
R2950 VDD.n10360 VDD.n10198 104.757
R2951 VDD.n10361 VDD.n10360 104.757
R2952 VDD.n10361 VDD.n10194 104.757
R2953 VDD.n10368 VDD.n10194 104.757
R2954 VDD.n10369 VDD.n10368 104.757
R2955 VDD.n10369 VDD.n10188 104.757
R2956 VDD.n10376 VDD.n10188 104.757
R2957 VDD.n10378 VDD.n10376 104.757
R2958 VDD.n10378 VDD.n10377 104.757
R2959 VDD.n10377 VDD.n10184 104.757
R2960 VDD.n10386 VDD.n10184 104.757
R2961 VDD.n10387 VDD.n10386 104.757
R2962 VDD.n10387 VDD.n10178 104.757
R2963 VDD.n10394 VDD.n10178 104.757
R2964 VDD.n10395 VDD.n10394 104.757
R2965 VDD.n10395 VDD.n10174 104.757
R2966 VDD.n10402 VDD.n10174 104.757
R2967 VDD.n10403 VDD.n10402 104.757
R2968 VDD.n10403 VDD.n10170 104.757
R2969 VDD.n10410 VDD.n10170 104.757
R2970 VDD.n10411 VDD.n10410 104.757
R2971 VDD.n10411 VDD.n10165 104.757
R2972 VDD.n10419 VDD.n10165 104.757
R2973 VDD.n10419 VDD.n10166 104.757
R2974 VDD.n10166 VDD.n6931 104.757
R2975 VDD.n12412 VDD.n6931 104.757
R2976 VDD.n12410 VDD.n12409 104.757
R2977 VDD.n6158 VDD.n6100 104.757
R2978 VDD.n6162 VDD.n6100 104.757
R2979 VDD.n6162 VDD.n6098 104.757
R2980 VDD.n6166 VDD.n6098 104.757
R2981 VDD.n6166 VDD.n6096 104.757
R2982 VDD.n6170 VDD.n6096 104.757
R2983 VDD.n6170 VDD.n6094 104.757
R2984 VDD.n6174 VDD.n6094 104.757
R2985 VDD.n6174 VDD.n6092 104.757
R2986 VDD.n6178 VDD.n6092 104.757
R2987 VDD.n6178 VDD.n6090 104.757
R2988 VDD.n6182 VDD.n6090 104.757
R2989 VDD.n6182 VDD.n6088 104.757
R2990 VDD.n6186 VDD.n6088 104.757
R2991 VDD.n6186 VDD.n6086 104.757
R2992 VDD.n6190 VDD.n6086 104.757
R2993 VDD.n6190 VDD.n6084 104.757
R2994 VDD.n6194 VDD.n6084 104.757
R2995 VDD.n6194 VDD.n6082 104.757
R2996 VDD.n6198 VDD.n6082 104.757
R2997 VDD.n6198 VDD.n6080 104.757
R2998 VDD.n6202 VDD.n6080 104.757
R2999 VDD.n6202 VDD.n6078 104.757
R3000 VDD.n6207 VDD.n6078 104.757
R3001 VDD.n6207 VDD.n6075 104.757
R3002 VDD.n6211 VDD.n6075 104.757
R3003 VDD.n6212 VDD.n6211 104.757
R3004 VDD.n6150 VDD.n6108 104.757
R3005 VDD.n6146 VDD.n6108 104.757
R3006 VDD.n6146 VDD.n6111 104.757
R3007 VDD.n6142 VDD.n6111 104.757
R3008 VDD.n6142 VDD.n6114 104.757
R3009 VDD.n6138 VDD.n6114 104.757
R3010 VDD.n6138 VDD.n6116 104.757
R3011 VDD.n6134 VDD.n6116 104.757
R3012 VDD.n6134 VDD.n6118 104.757
R3013 VDD.n6130 VDD.n6118 104.757
R3014 VDD.n6130 VDD.n6120 104.757
R3015 VDD.n6126 VDD.n6120 104.757
R3016 VDD.n6126 VDD.n6123 104.757
R3017 VDD.n6123 VDD.n5898 104.757
R3018 VDD.n6389 VDD.n5898 104.757
R3019 VDD.n6368 VDD.n5890 104.757
R3020 VDD.n5949 VDD.n5890 104.757
R3021 VDD.n5953 VDD.n5952 104.757
R3022 VDD.n6393 VDD.n5876 104.757
R3023 VDD.n6397 VDD.n5876 104.757
R3024 VDD.n6397 VDD.n5874 104.757
R3025 VDD.n6401 VDD.n5874 104.757
R3026 VDD.n6401 VDD.n5872 104.757
R3027 VDD.n6405 VDD.n5872 104.757
R3028 VDD.n6405 VDD.n5870 104.757
R3029 VDD.n6409 VDD.n5870 104.757
R3030 VDD.n6409 VDD.n5868 104.757
R3031 VDD.n6413 VDD.n5868 104.757
R3032 VDD.n6413 VDD.n5866 104.757
R3033 VDD.n6417 VDD.n5866 104.757
R3034 VDD.n6417 VDD.n5863 104.757
R3035 VDD.n6422 VDD.n5863 104.757
R3036 VDD.n6422 VDD.n5864 104.757
R3037 VDD.n6426 VDD.n5860 104.757
R3038 VDD.n6430 VDD.n5858 104.757
R3039 VDD.n6430 VDD.n5856 104.757
R3040 VDD.n6434 VDD.n5856 104.757
R3041 VDD.n6434 VDD.n5854 104.757
R3042 VDD.n6438 VDD.n5854 104.757
R3043 VDD.n6438 VDD.n5852 104.757
R3044 VDD.n6442 VDD.n5852 104.757
R3045 VDD.n6442 VDD.n5850 104.757
R3046 VDD.n6446 VDD.n5850 104.757
R3047 VDD.n6446 VDD.n5848 104.757
R3048 VDD.n6450 VDD.n5848 104.757
R3049 VDD.n6450 VDD.n5846 104.757
R3050 VDD.n6454 VDD.n5846 104.757
R3051 VDD.n6454 VDD.n5844 104.757
R3052 VDD.n6458 VDD.n5844 104.757
R3053 VDD.n6458 VDD.n5842 104.757
R3054 VDD.n6462 VDD.n5842 104.757
R3055 VDD.n6462 VDD.n5840 104.757
R3056 VDD.n6466 VDD.n5840 104.757
R3057 VDD.n6466 VDD.n5838 104.757
R3058 VDD.n6470 VDD.n5838 104.757
R3059 VDD.n6470 VDD.n5836 104.757
R3060 VDD.n6474 VDD.n5836 104.757
R3061 VDD.n6474 VDD.n5834 104.757
R3062 VDD.n6478 VDD.n5834 104.757
R3063 VDD.n6478 VDD.n5832 104.757
R3064 VDD.n6482 VDD.n5832 104.757
R3065 VDD.n6482 VDD.n5829 104.757
R3066 VDD.n6215 VDD.n6073 104.757
R3067 VDD.n6219 VDD.n6070 104.757
R3068 VDD.n6225 VDD.n6070 104.757
R3069 VDD.n6225 VDD.n6068 104.757
R3070 VDD.n6229 VDD.n6068 104.757
R3071 VDD.n6229 VDD.n6066 104.757
R3072 VDD.n6233 VDD.n6066 104.757
R3073 VDD.n6233 VDD.n6064 104.757
R3074 VDD.n6237 VDD.n6064 104.757
R3075 VDD.n6237 VDD.n6062 104.757
R3076 VDD.n6241 VDD.n6062 104.757
R3077 VDD.n6241 VDD.n6060 104.757
R3078 VDD.n6246 VDD.n6060 104.757
R3079 VDD.n6246 VDD.n6057 104.757
R3080 VDD.n6251 VDD.n6057 104.757
R3081 VDD.n6252 VDD.n6251 104.757
R3082 VDD.n6264 VDD.n6053 104.757
R3083 VDD.n6267 VDD.n6266 104.757
R3084 VDD.n6278 VDD.n6277 104.757
R3085 VDD.n6285 VDD.n6284 104.757
R3086 VDD.n6540 VDD.n6539 104.757
R3087 VDD.n6532 VDD.n5803 104.757
R3088 VDD.n6530 VDD.n5804 104.757
R3089 VDD.n6522 VDD.n6521 104.757
R3090 VDD.n6519 VDD.n5810 104.757
R3091 VDD.n6514 VDD.n5810 104.757
R3092 VDD.n6514 VDD.n5812 104.757
R3093 VDD.n6510 VDD.n5812 104.757
R3094 VDD.n6510 VDD.n5815 104.757
R3095 VDD.n6506 VDD.n5815 104.757
R3096 VDD.n6506 VDD.n5817 104.757
R3097 VDD.n6502 VDD.n5817 104.757
R3098 VDD.n6502 VDD.n5819 104.757
R3099 VDD.n6498 VDD.n5819 104.757
R3100 VDD.n6498 VDD.n5821 104.757
R3101 VDD.n6494 VDD.n5821 104.757
R3102 VDD.n6494 VDD.n5823 104.757
R3103 VDD.n6490 VDD.n5823 104.757
R3104 VDD.n6490 VDD.n5825 104.757
R3105 VDD.n6486 VDD.n5828 104.757
R3106 VDD.n5304 VDD.n5246 104.757
R3107 VDD.n5308 VDD.n5246 104.757
R3108 VDD.n5308 VDD.n5244 104.757
R3109 VDD.n5312 VDD.n5244 104.757
R3110 VDD.n5312 VDD.n5242 104.757
R3111 VDD.n5316 VDD.n5242 104.757
R3112 VDD.n5316 VDD.n5240 104.757
R3113 VDD.n5320 VDD.n5240 104.757
R3114 VDD.n5320 VDD.n5238 104.757
R3115 VDD.n5324 VDD.n5238 104.757
R3116 VDD.n5324 VDD.n5236 104.757
R3117 VDD.n5328 VDD.n5236 104.757
R3118 VDD.n5328 VDD.n5234 104.757
R3119 VDD.n5332 VDD.n5234 104.757
R3120 VDD.n5332 VDD.n5232 104.757
R3121 VDD.n5336 VDD.n5232 104.757
R3122 VDD.n5336 VDD.n5230 104.757
R3123 VDD.n5340 VDD.n5230 104.757
R3124 VDD.n5340 VDD.n5228 104.757
R3125 VDD.n5344 VDD.n5228 104.757
R3126 VDD.n5344 VDD.n5226 104.757
R3127 VDD.n5348 VDD.n5226 104.757
R3128 VDD.n5348 VDD.n5224 104.757
R3129 VDD.n5353 VDD.n5224 104.757
R3130 VDD.n5353 VDD.n5221 104.757
R3131 VDD.n5357 VDD.n5221 104.757
R3132 VDD.n5358 VDD.n5357 104.757
R3133 VDD.n5296 VDD.n5254 104.757
R3134 VDD.n5292 VDD.n5254 104.757
R3135 VDD.n5292 VDD.n5257 104.757
R3136 VDD.n5288 VDD.n5257 104.757
R3137 VDD.n5288 VDD.n5260 104.757
R3138 VDD.n5284 VDD.n5260 104.757
R3139 VDD.n5284 VDD.n5262 104.757
R3140 VDD.n5280 VDD.n5262 104.757
R3141 VDD.n5280 VDD.n5264 104.757
R3142 VDD.n5276 VDD.n5264 104.757
R3143 VDD.n5276 VDD.n5266 104.757
R3144 VDD.n5272 VDD.n5266 104.757
R3145 VDD.n5272 VDD.n5269 104.757
R3146 VDD.n5269 VDD.n5044 104.757
R3147 VDD.n5535 VDD.n5044 104.757
R3148 VDD.n5514 VDD.n5036 104.757
R3149 VDD.n5095 VDD.n5036 104.757
R3150 VDD.n5099 VDD.n5098 104.757
R3151 VDD.n5539 VDD.n5022 104.757
R3152 VDD.n5543 VDD.n5022 104.757
R3153 VDD.n5543 VDD.n5020 104.757
R3154 VDD.n5547 VDD.n5020 104.757
R3155 VDD.n5547 VDD.n5018 104.757
R3156 VDD.n5551 VDD.n5018 104.757
R3157 VDD.n5551 VDD.n5016 104.757
R3158 VDD.n5555 VDD.n5016 104.757
R3159 VDD.n5555 VDD.n5014 104.757
R3160 VDD.n5559 VDD.n5014 104.757
R3161 VDD.n5559 VDD.n5012 104.757
R3162 VDD.n5563 VDD.n5012 104.757
R3163 VDD.n5563 VDD.n5009 104.757
R3164 VDD.n5568 VDD.n5009 104.757
R3165 VDD.n5568 VDD.n5010 104.757
R3166 VDD.n5572 VDD.n5006 104.757
R3167 VDD.n5576 VDD.n5004 104.757
R3168 VDD.n5576 VDD.n5002 104.757
R3169 VDD.n5580 VDD.n5002 104.757
R3170 VDD.n5580 VDD.n5000 104.757
R3171 VDD.n5584 VDD.n5000 104.757
R3172 VDD.n5584 VDD.n4998 104.757
R3173 VDD.n5588 VDD.n4998 104.757
R3174 VDD.n5588 VDD.n4996 104.757
R3175 VDD.n5592 VDD.n4996 104.757
R3176 VDD.n5592 VDD.n4994 104.757
R3177 VDD.n5596 VDD.n4994 104.757
R3178 VDD.n5596 VDD.n4992 104.757
R3179 VDD.n5600 VDD.n4992 104.757
R3180 VDD.n5600 VDD.n4990 104.757
R3181 VDD.n5604 VDD.n4990 104.757
R3182 VDD.n5604 VDD.n4988 104.757
R3183 VDD.n5608 VDD.n4988 104.757
R3184 VDD.n5608 VDD.n4986 104.757
R3185 VDD.n5612 VDD.n4986 104.757
R3186 VDD.n5612 VDD.n4984 104.757
R3187 VDD.n5616 VDD.n4984 104.757
R3188 VDD.n5616 VDD.n4982 104.757
R3189 VDD.n5620 VDD.n4982 104.757
R3190 VDD.n5620 VDD.n4980 104.757
R3191 VDD.n5624 VDD.n4980 104.757
R3192 VDD.n5624 VDD.n4978 104.757
R3193 VDD.n5628 VDD.n4978 104.757
R3194 VDD.n5628 VDD.n4975 104.757
R3195 VDD.n5361 VDD.n5219 104.757
R3196 VDD.n5365 VDD.n5216 104.757
R3197 VDD.n5371 VDD.n5216 104.757
R3198 VDD.n5371 VDD.n5214 104.757
R3199 VDD.n5375 VDD.n5214 104.757
R3200 VDD.n5375 VDD.n5212 104.757
R3201 VDD.n5379 VDD.n5212 104.757
R3202 VDD.n5379 VDD.n5210 104.757
R3203 VDD.n5383 VDD.n5210 104.757
R3204 VDD.n5383 VDD.n5208 104.757
R3205 VDD.n5387 VDD.n5208 104.757
R3206 VDD.n5387 VDD.n5206 104.757
R3207 VDD.n5392 VDD.n5206 104.757
R3208 VDD.n5392 VDD.n5203 104.757
R3209 VDD.n5397 VDD.n5203 104.757
R3210 VDD.n5398 VDD.n5397 104.757
R3211 VDD.n5410 VDD.n5199 104.757
R3212 VDD.n5413 VDD.n5412 104.757
R3213 VDD.n5424 VDD.n5423 104.757
R3214 VDD.n5431 VDD.n5430 104.757
R3215 VDD.n5686 VDD.n5685 104.757
R3216 VDD.n5678 VDD.n4949 104.757
R3217 VDD.n5676 VDD.n4950 104.757
R3218 VDD.n5668 VDD.n5667 104.757
R3219 VDD.n5665 VDD.n4956 104.757
R3220 VDD.n5660 VDD.n4956 104.757
R3221 VDD.n5660 VDD.n4958 104.757
R3222 VDD.n5656 VDD.n4958 104.757
R3223 VDD.n5656 VDD.n4961 104.757
R3224 VDD.n5652 VDD.n4961 104.757
R3225 VDD.n5652 VDD.n4963 104.757
R3226 VDD.n5648 VDD.n4963 104.757
R3227 VDD.n5648 VDD.n4965 104.757
R3228 VDD.n5644 VDD.n4965 104.757
R3229 VDD.n5644 VDD.n4967 104.757
R3230 VDD.n5640 VDD.n4967 104.757
R3231 VDD.n5640 VDD.n4969 104.757
R3232 VDD.n5636 VDD.n4969 104.757
R3233 VDD.n5636 VDD.n4971 104.757
R3234 VDD.n5632 VDD.n4974 104.757
R3235 VDD.n4518 VDD.n4460 104.757
R3236 VDD.n4522 VDD.n4460 104.757
R3237 VDD.n4522 VDD.n4458 104.757
R3238 VDD.n4526 VDD.n4458 104.757
R3239 VDD.n4526 VDD.n4456 104.757
R3240 VDD.n4530 VDD.n4456 104.757
R3241 VDD.n4530 VDD.n4454 104.757
R3242 VDD.n4534 VDD.n4454 104.757
R3243 VDD.n4534 VDD.n4452 104.757
R3244 VDD.n4538 VDD.n4452 104.757
R3245 VDD.n4538 VDD.n4450 104.757
R3246 VDD.n4542 VDD.n4450 104.757
R3247 VDD.n4542 VDD.n4448 104.757
R3248 VDD.n4546 VDD.n4448 104.757
R3249 VDD.n4546 VDD.n4446 104.757
R3250 VDD.n4550 VDD.n4446 104.757
R3251 VDD.n4550 VDD.n4444 104.757
R3252 VDD.n4554 VDD.n4444 104.757
R3253 VDD.n4554 VDD.n4442 104.757
R3254 VDD.n4558 VDD.n4442 104.757
R3255 VDD.n4558 VDD.n4440 104.757
R3256 VDD.n4562 VDD.n4440 104.757
R3257 VDD.n4562 VDD.n4438 104.757
R3258 VDD.n4567 VDD.n4438 104.757
R3259 VDD.n4567 VDD.n4435 104.757
R3260 VDD.n4571 VDD.n4435 104.757
R3261 VDD.n4572 VDD.n4571 104.757
R3262 VDD.n4510 VDD.n4468 104.757
R3263 VDD.n4506 VDD.n4468 104.757
R3264 VDD.n4506 VDD.n4471 104.757
R3265 VDD.n4502 VDD.n4471 104.757
R3266 VDD.n4502 VDD.n4474 104.757
R3267 VDD.n4498 VDD.n4474 104.757
R3268 VDD.n4498 VDD.n4476 104.757
R3269 VDD.n4494 VDD.n4476 104.757
R3270 VDD.n4494 VDD.n4478 104.757
R3271 VDD.n4490 VDD.n4478 104.757
R3272 VDD.n4490 VDD.n4480 104.757
R3273 VDD.n4486 VDD.n4480 104.757
R3274 VDD.n4486 VDD.n4483 104.757
R3275 VDD.n4483 VDD.n4258 104.757
R3276 VDD.n4749 VDD.n4258 104.757
R3277 VDD.n4728 VDD.n4250 104.757
R3278 VDD.n4309 VDD.n4250 104.757
R3279 VDD.n4313 VDD.n4312 104.757
R3280 VDD.n4753 VDD.n4236 104.757
R3281 VDD.n4757 VDD.n4236 104.757
R3282 VDD.n4757 VDD.n4234 104.757
R3283 VDD.n4761 VDD.n4234 104.757
R3284 VDD.n4761 VDD.n4232 104.757
R3285 VDD.n4765 VDD.n4232 104.757
R3286 VDD.n4765 VDD.n4230 104.757
R3287 VDD.n4769 VDD.n4230 104.757
R3288 VDD.n4769 VDD.n4228 104.757
R3289 VDD.n4773 VDD.n4228 104.757
R3290 VDD.n4773 VDD.n4226 104.757
R3291 VDD.n4777 VDD.n4226 104.757
R3292 VDD.n4777 VDD.n4223 104.757
R3293 VDD.n4782 VDD.n4223 104.757
R3294 VDD.n4782 VDD.n4224 104.757
R3295 VDD.n4786 VDD.n4220 104.757
R3296 VDD.n4790 VDD.n4218 104.757
R3297 VDD.n4790 VDD.n4216 104.757
R3298 VDD.n4794 VDD.n4216 104.757
R3299 VDD.n4794 VDD.n4214 104.757
R3300 VDD.n4798 VDD.n4214 104.757
R3301 VDD.n4798 VDD.n4212 104.757
R3302 VDD.n4802 VDD.n4212 104.757
R3303 VDD.n4802 VDD.n4210 104.757
R3304 VDD.n4806 VDD.n4210 104.757
R3305 VDD.n4806 VDD.n4208 104.757
R3306 VDD.n4810 VDD.n4208 104.757
R3307 VDD.n4810 VDD.n4206 104.757
R3308 VDD.n4814 VDD.n4206 104.757
R3309 VDD.n4814 VDD.n4204 104.757
R3310 VDD.n4818 VDD.n4204 104.757
R3311 VDD.n4818 VDD.n4202 104.757
R3312 VDD.n4822 VDD.n4202 104.757
R3313 VDD.n4822 VDD.n4200 104.757
R3314 VDD.n4826 VDD.n4200 104.757
R3315 VDD.n4826 VDD.n4198 104.757
R3316 VDD.n4830 VDD.n4198 104.757
R3317 VDD.n4830 VDD.n4196 104.757
R3318 VDD.n4834 VDD.n4196 104.757
R3319 VDD.n4834 VDD.n4194 104.757
R3320 VDD.n4838 VDD.n4194 104.757
R3321 VDD.n4838 VDD.n4192 104.757
R3322 VDD.n4842 VDD.n4192 104.757
R3323 VDD.n4842 VDD.n4189 104.757
R3324 VDD.n4575 VDD.n4433 104.757
R3325 VDD.n4579 VDD.n4430 104.757
R3326 VDD.n4585 VDD.n4430 104.757
R3327 VDD.n4585 VDD.n4428 104.757
R3328 VDD.n4589 VDD.n4428 104.757
R3329 VDD.n4589 VDD.n4426 104.757
R3330 VDD.n4593 VDD.n4426 104.757
R3331 VDD.n4593 VDD.n4424 104.757
R3332 VDD.n4597 VDD.n4424 104.757
R3333 VDD.n4597 VDD.n4422 104.757
R3334 VDD.n4601 VDD.n4422 104.757
R3335 VDD.n4601 VDD.n4420 104.757
R3336 VDD.n4606 VDD.n4420 104.757
R3337 VDD.n4606 VDD.n4417 104.757
R3338 VDD.n4611 VDD.n4417 104.757
R3339 VDD.n4612 VDD.n4611 104.757
R3340 VDD.n4624 VDD.n4413 104.757
R3341 VDD.n4627 VDD.n4626 104.757
R3342 VDD.n4638 VDD.n4637 104.757
R3343 VDD.n4645 VDD.n4644 104.757
R3344 VDD.n4900 VDD.n4899 104.757
R3345 VDD.n4892 VDD.n4163 104.757
R3346 VDD.n4890 VDD.n4164 104.757
R3347 VDD.n4882 VDD.n4881 104.757
R3348 VDD.n4879 VDD.n4170 104.757
R3349 VDD.n4874 VDD.n4170 104.757
R3350 VDD.n4874 VDD.n4172 104.757
R3351 VDD.n4870 VDD.n4172 104.757
R3352 VDD.n4870 VDD.n4175 104.757
R3353 VDD.n4866 VDD.n4175 104.757
R3354 VDD.n4866 VDD.n4177 104.757
R3355 VDD.n4862 VDD.n4177 104.757
R3356 VDD.n4862 VDD.n4179 104.757
R3357 VDD.n4858 VDD.n4179 104.757
R3358 VDD.n4858 VDD.n4181 104.757
R3359 VDD.n4854 VDD.n4181 104.757
R3360 VDD.n4854 VDD.n4183 104.757
R3361 VDD.n4850 VDD.n4183 104.757
R3362 VDD.n4850 VDD.n4185 104.757
R3363 VDD.n4846 VDD.n4188 104.757
R3364 VDD.n3664 VDD.n3606 104.757
R3365 VDD.n3668 VDD.n3606 104.757
R3366 VDD.n3668 VDD.n3604 104.757
R3367 VDD.n3672 VDD.n3604 104.757
R3368 VDD.n3672 VDD.n3602 104.757
R3369 VDD.n3676 VDD.n3602 104.757
R3370 VDD.n3676 VDD.n3600 104.757
R3371 VDD.n3680 VDD.n3600 104.757
R3372 VDD.n3680 VDD.n3598 104.757
R3373 VDD.n3684 VDD.n3598 104.757
R3374 VDD.n3684 VDD.n3596 104.757
R3375 VDD.n3688 VDD.n3596 104.757
R3376 VDD.n3688 VDD.n3594 104.757
R3377 VDD.n3692 VDD.n3594 104.757
R3378 VDD.n3692 VDD.n3592 104.757
R3379 VDD.n3696 VDD.n3592 104.757
R3380 VDD.n3696 VDD.n3590 104.757
R3381 VDD.n3700 VDD.n3590 104.757
R3382 VDD.n3700 VDD.n3588 104.757
R3383 VDD.n3704 VDD.n3588 104.757
R3384 VDD.n3704 VDD.n3586 104.757
R3385 VDD.n3708 VDD.n3586 104.757
R3386 VDD.n3708 VDD.n3584 104.757
R3387 VDD.n3713 VDD.n3584 104.757
R3388 VDD.n3713 VDD.n3581 104.757
R3389 VDD.n3717 VDD.n3581 104.757
R3390 VDD.n3718 VDD.n3717 104.757
R3391 VDD.n3656 VDD.n3614 104.757
R3392 VDD.n3652 VDD.n3614 104.757
R3393 VDD.n3652 VDD.n3617 104.757
R3394 VDD.n3648 VDD.n3617 104.757
R3395 VDD.n3648 VDD.n3620 104.757
R3396 VDD.n3644 VDD.n3620 104.757
R3397 VDD.n3644 VDD.n3622 104.757
R3398 VDD.n3640 VDD.n3622 104.757
R3399 VDD.n3640 VDD.n3624 104.757
R3400 VDD.n3636 VDD.n3624 104.757
R3401 VDD.n3636 VDD.n3626 104.757
R3402 VDD.n3632 VDD.n3626 104.757
R3403 VDD.n3632 VDD.n3629 104.757
R3404 VDD.n3629 VDD.n3404 104.757
R3405 VDD.n3895 VDD.n3404 104.757
R3406 VDD.n3874 VDD.n3396 104.757
R3407 VDD.n3455 VDD.n3396 104.757
R3408 VDD.n3459 VDD.n3458 104.757
R3409 VDD.n3899 VDD.n3382 104.757
R3410 VDD.n3903 VDD.n3382 104.757
R3411 VDD.n3903 VDD.n3380 104.757
R3412 VDD.n3907 VDD.n3380 104.757
R3413 VDD.n3907 VDD.n3378 104.757
R3414 VDD.n3911 VDD.n3378 104.757
R3415 VDD.n3911 VDD.n3376 104.757
R3416 VDD.n3915 VDD.n3376 104.757
R3417 VDD.n3915 VDD.n3374 104.757
R3418 VDD.n3919 VDD.n3374 104.757
R3419 VDD.n3919 VDD.n3372 104.757
R3420 VDD.n3923 VDD.n3372 104.757
R3421 VDD.n3923 VDD.n3369 104.757
R3422 VDD.n3928 VDD.n3369 104.757
R3423 VDD.n3928 VDD.n3370 104.757
R3424 VDD.n3932 VDD.n3366 104.757
R3425 VDD.n3936 VDD.n3364 104.757
R3426 VDD.n3936 VDD.n3362 104.757
R3427 VDD.n3940 VDD.n3362 104.757
R3428 VDD.n3940 VDD.n3360 104.757
R3429 VDD.n3944 VDD.n3360 104.757
R3430 VDD.n3944 VDD.n3358 104.757
R3431 VDD.n3948 VDD.n3358 104.757
R3432 VDD.n3948 VDD.n3356 104.757
R3433 VDD.n3952 VDD.n3356 104.757
R3434 VDD.n3952 VDD.n3354 104.757
R3435 VDD.n3956 VDD.n3354 104.757
R3436 VDD.n3956 VDD.n3352 104.757
R3437 VDD.n3960 VDD.n3352 104.757
R3438 VDD.n3960 VDD.n3350 104.757
R3439 VDD.n3964 VDD.n3350 104.757
R3440 VDD.n3964 VDD.n3348 104.757
R3441 VDD.n3968 VDD.n3348 104.757
R3442 VDD.n3968 VDD.n3346 104.757
R3443 VDD.n3972 VDD.n3346 104.757
R3444 VDD.n3972 VDD.n3344 104.757
R3445 VDD.n3976 VDD.n3344 104.757
R3446 VDD.n3976 VDD.n3342 104.757
R3447 VDD.n3980 VDD.n3342 104.757
R3448 VDD.n3980 VDD.n3340 104.757
R3449 VDD.n3984 VDD.n3340 104.757
R3450 VDD.n3984 VDD.n3338 104.757
R3451 VDD.n3988 VDD.n3338 104.757
R3452 VDD.n3988 VDD.n3335 104.757
R3453 VDD.n3721 VDD.n3579 104.757
R3454 VDD.n3725 VDD.n3576 104.757
R3455 VDD.n3731 VDD.n3576 104.757
R3456 VDD.n3731 VDD.n3574 104.757
R3457 VDD.n3735 VDD.n3574 104.757
R3458 VDD.n3735 VDD.n3572 104.757
R3459 VDD.n3739 VDD.n3572 104.757
R3460 VDD.n3739 VDD.n3570 104.757
R3461 VDD.n3743 VDD.n3570 104.757
R3462 VDD.n3743 VDD.n3568 104.757
R3463 VDD.n3747 VDD.n3568 104.757
R3464 VDD.n3747 VDD.n3566 104.757
R3465 VDD.n3752 VDD.n3566 104.757
R3466 VDD.n3752 VDD.n3563 104.757
R3467 VDD.n3757 VDD.n3563 104.757
R3468 VDD.n3758 VDD.n3757 104.757
R3469 VDD.n3770 VDD.n3559 104.757
R3470 VDD.n3773 VDD.n3772 104.757
R3471 VDD.n3784 VDD.n3783 104.757
R3472 VDD.n3791 VDD.n3790 104.757
R3473 VDD.n4046 VDD.n4045 104.757
R3474 VDD.n4038 VDD.n3309 104.757
R3475 VDD.n4036 VDD.n3310 104.757
R3476 VDD.n4028 VDD.n4027 104.757
R3477 VDD.n4025 VDD.n3316 104.757
R3478 VDD.n4020 VDD.n3316 104.757
R3479 VDD.n4020 VDD.n3318 104.757
R3480 VDD.n4016 VDD.n3318 104.757
R3481 VDD.n4016 VDD.n3321 104.757
R3482 VDD.n4012 VDD.n3321 104.757
R3483 VDD.n4012 VDD.n3323 104.757
R3484 VDD.n4008 VDD.n3323 104.757
R3485 VDD.n4008 VDD.n3325 104.757
R3486 VDD.n4004 VDD.n3325 104.757
R3487 VDD.n4004 VDD.n3327 104.757
R3488 VDD.n4000 VDD.n3327 104.757
R3489 VDD.n4000 VDD.n3329 104.757
R3490 VDD.n3996 VDD.n3329 104.757
R3491 VDD.n3996 VDD.n3331 104.757
R3492 VDD.n3992 VDD.n3334 104.757
R3493 VDD.n2878 VDD.n2820 104.757
R3494 VDD.n2882 VDD.n2820 104.757
R3495 VDD.n2882 VDD.n2818 104.757
R3496 VDD.n2886 VDD.n2818 104.757
R3497 VDD.n2886 VDD.n2816 104.757
R3498 VDD.n2890 VDD.n2816 104.757
R3499 VDD.n2890 VDD.n2814 104.757
R3500 VDD.n2894 VDD.n2814 104.757
R3501 VDD.n2894 VDD.n2812 104.757
R3502 VDD.n2898 VDD.n2812 104.757
R3503 VDD.n2898 VDD.n2810 104.757
R3504 VDD.n2902 VDD.n2810 104.757
R3505 VDD.n2902 VDD.n2808 104.757
R3506 VDD.n2906 VDD.n2808 104.757
R3507 VDD.n2906 VDD.n2806 104.757
R3508 VDD.n2910 VDD.n2806 104.757
R3509 VDD.n2910 VDD.n2804 104.757
R3510 VDD.n2914 VDD.n2804 104.757
R3511 VDD.n2914 VDD.n2802 104.757
R3512 VDD.n2918 VDD.n2802 104.757
R3513 VDD.n2918 VDD.n2800 104.757
R3514 VDD.n2922 VDD.n2800 104.757
R3515 VDD.n2922 VDD.n2798 104.757
R3516 VDD.n2927 VDD.n2798 104.757
R3517 VDD.n2927 VDD.n2795 104.757
R3518 VDD.n2931 VDD.n2795 104.757
R3519 VDD.n2932 VDD.n2931 104.757
R3520 VDD.n2870 VDD.n2828 104.757
R3521 VDD.n2866 VDD.n2828 104.757
R3522 VDD.n2866 VDD.n2831 104.757
R3523 VDD.n2862 VDD.n2831 104.757
R3524 VDD.n2862 VDD.n2834 104.757
R3525 VDD.n2858 VDD.n2834 104.757
R3526 VDD.n2858 VDD.n2836 104.757
R3527 VDD.n2854 VDD.n2836 104.757
R3528 VDD.n2854 VDD.n2838 104.757
R3529 VDD.n2850 VDD.n2838 104.757
R3530 VDD.n2850 VDD.n2840 104.757
R3531 VDD.n2846 VDD.n2840 104.757
R3532 VDD.n2846 VDD.n2843 104.757
R3533 VDD.n2843 VDD.n2618 104.757
R3534 VDD.n3109 VDD.n2618 104.757
R3535 VDD.n3088 VDD.n2610 104.757
R3536 VDD.n2669 VDD.n2610 104.757
R3537 VDD.n2673 VDD.n2672 104.757
R3538 VDD.n3113 VDD.n2596 104.757
R3539 VDD.n3117 VDD.n2596 104.757
R3540 VDD.n3117 VDD.n2594 104.757
R3541 VDD.n3121 VDD.n2594 104.757
R3542 VDD.n3121 VDD.n2592 104.757
R3543 VDD.n3125 VDD.n2592 104.757
R3544 VDD.n3125 VDD.n2590 104.757
R3545 VDD.n3129 VDD.n2590 104.757
R3546 VDD.n3129 VDD.n2588 104.757
R3547 VDD.n3133 VDD.n2588 104.757
R3548 VDD.n3133 VDD.n2586 104.757
R3549 VDD.n3137 VDD.n2586 104.757
R3550 VDD.n3137 VDD.n2583 104.757
R3551 VDD.n3142 VDD.n2583 104.757
R3552 VDD.n3142 VDD.n2584 104.757
R3553 VDD.n3146 VDD.n2580 104.757
R3554 VDD.n3150 VDD.n2578 104.757
R3555 VDD.n3150 VDD.n2576 104.757
R3556 VDD.n3154 VDD.n2576 104.757
R3557 VDD.n3154 VDD.n2574 104.757
R3558 VDD.n3158 VDD.n2574 104.757
R3559 VDD.n3158 VDD.n2572 104.757
R3560 VDD.n3162 VDD.n2572 104.757
R3561 VDD.n3162 VDD.n2570 104.757
R3562 VDD.n3166 VDD.n2570 104.757
R3563 VDD.n3166 VDD.n2568 104.757
R3564 VDD.n3170 VDD.n2568 104.757
R3565 VDD.n3170 VDD.n2566 104.757
R3566 VDD.n3174 VDD.n2566 104.757
R3567 VDD.n3174 VDD.n2564 104.757
R3568 VDD.n3178 VDD.n2564 104.757
R3569 VDD.n3178 VDD.n2562 104.757
R3570 VDD.n3182 VDD.n2562 104.757
R3571 VDD.n3182 VDD.n2560 104.757
R3572 VDD.n3186 VDD.n2560 104.757
R3573 VDD.n3186 VDD.n2558 104.757
R3574 VDD.n3190 VDD.n2558 104.757
R3575 VDD.n3190 VDD.n2556 104.757
R3576 VDD.n3194 VDD.n2556 104.757
R3577 VDD.n3194 VDD.n2554 104.757
R3578 VDD.n3198 VDD.n2554 104.757
R3579 VDD.n3198 VDD.n2552 104.757
R3580 VDD.n3202 VDD.n2552 104.757
R3581 VDD.n3202 VDD.n2549 104.757
R3582 VDD.n2935 VDD.n2793 104.757
R3583 VDD.n2939 VDD.n2790 104.757
R3584 VDD.n2945 VDD.n2790 104.757
R3585 VDD.n2945 VDD.n2788 104.757
R3586 VDD.n2949 VDD.n2788 104.757
R3587 VDD.n2949 VDD.n2786 104.757
R3588 VDD.n2953 VDD.n2786 104.757
R3589 VDD.n2953 VDD.n2784 104.757
R3590 VDD.n2957 VDD.n2784 104.757
R3591 VDD.n2957 VDD.n2782 104.757
R3592 VDD.n2961 VDD.n2782 104.757
R3593 VDD.n2961 VDD.n2780 104.757
R3594 VDD.n2966 VDD.n2780 104.757
R3595 VDD.n2966 VDD.n2777 104.757
R3596 VDD.n2971 VDD.n2777 104.757
R3597 VDD.n2972 VDD.n2971 104.757
R3598 VDD.n2984 VDD.n2773 104.757
R3599 VDD.n2987 VDD.n2986 104.757
R3600 VDD.n2998 VDD.n2997 104.757
R3601 VDD.n3005 VDD.n3004 104.757
R3602 VDD.n3260 VDD.n3259 104.757
R3603 VDD.n3252 VDD.n2523 104.757
R3604 VDD.n3250 VDD.n2524 104.757
R3605 VDD.n3242 VDD.n3241 104.757
R3606 VDD.n3239 VDD.n2530 104.757
R3607 VDD.n3234 VDD.n2530 104.757
R3608 VDD.n3234 VDD.n2532 104.757
R3609 VDD.n3230 VDD.n2532 104.757
R3610 VDD.n3230 VDD.n2535 104.757
R3611 VDD.n3226 VDD.n2535 104.757
R3612 VDD.n3226 VDD.n2537 104.757
R3613 VDD.n3222 VDD.n2537 104.757
R3614 VDD.n3222 VDD.n2539 104.757
R3615 VDD.n3218 VDD.n2539 104.757
R3616 VDD.n3218 VDD.n2541 104.757
R3617 VDD.n3214 VDD.n2541 104.757
R3618 VDD.n3214 VDD.n2543 104.757
R3619 VDD.n3210 VDD.n2543 104.757
R3620 VDD.n3210 VDD.n2545 104.757
R3621 VDD.n3206 VDD.n2548 104.757
R3622 VDD.n2023 VDD.n1965 104.757
R3623 VDD.n2027 VDD.n1965 104.757
R3624 VDD.n2027 VDD.n1963 104.757
R3625 VDD.n2031 VDD.n1963 104.757
R3626 VDD.n2031 VDD.n1961 104.757
R3627 VDD.n2035 VDD.n1961 104.757
R3628 VDD.n2035 VDD.n1959 104.757
R3629 VDD.n2039 VDD.n1959 104.757
R3630 VDD.n2039 VDD.n1957 104.757
R3631 VDD.n2043 VDD.n1957 104.757
R3632 VDD.n2043 VDD.n1955 104.757
R3633 VDD.n2047 VDD.n1955 104.757
R3634 VDD.n2047 VDD.n1953 104.757
R3635 VDD.n2051 VDD.n1953 104.757
R3636 VDD.n2051 VDD.n1951 104.757
R3637 VDD.n2055 VDD.n1951 104.757
R3638 VDD.n2055 VDD.n1949 104.757
R3639 VDD.n2059 VDD.n1949 104.757
R3640 VDD.n2059 VDD.n1947 104.757
R3641 VDD.n2063 VDD.n1947 104.757
R3642 VDD.n2063 VDD.n1945 104.757
R3643 VDD.n2067 VDD.n1945 104.757
R3644 VDD.n2067 VDD.n1943 104.757
R3645 VDD.n2072 VDD.n1943 104.757
R3646 VDD.n2072 VDD.n1940 104.757
R3647 VDD.n2076 VDD.n1940 104.757
R3648 VDD.n2077 VDD.n2076 104.757
R3649 VDD.n2015 VDD.n1973 104.757
R3650 VDD.n2011 VDD.n1973 104.757
R3651 VDD.n2011 VDD.n1976 104.757
R3652 VDD.n2007 VDD.n1976 104.757
R3653 VDD.n2007 VDD.n1979 104.757
R3654 VDD.n2003 VDD.n1979 104.757
R3655 VDD.n2003 VDD.n1981 104.757
R3656 VDD.n1999 VDD.n1981 104.757
R3657 VDD.n1999 VDD.n1983 104.757
R3658 VDD.n1995 VDD.n1983 104.757
R3659 VDD.n1995 VDD.n1985 104.757
R3660 VDD.n1991 VDD.n1985 104.757
R3661 VDD.n1991 VDD.n1988 104.757
R3662 VDD.n1988 VDD.n1763 104.757
R3663 VDD.n2254 VDD.n1763 104.757
R3664 VDD.n2233 VDD.n1755 104.757
R3665 VDD.n1814 VDD.n1755 104.757
R3666 VDD.n1818 VDD.n1817 104.757
R3667 VDD.n2258 VDD.n1741 104.757
R3668 VDD.n2262 VDD.n1741 104.757
R3669 VDD.n2262 VDD.n1739 104.757
R3670 VDD.n2266 VDD.n1739 104.757
R3671 VDD.n2266 VDD.n1737 104.757
R3672 VDD.n2270 VDD.n1737 104.757
R3673 VDD.n2270 VDD.n1735 104.757
R3674 VDD.n2274 VDD.n1735 104.757
R3675 VDD.n2274 VDD.n1733 104.757
R3676 VDD.n2278 VDD.n1733 104.757
R3677 VDD.n2278 VDD.n1731 104.757
R3678 VDD.n2282 VDD.n1731 104.757
R3679 VDD.n2282 VDD.n1728 104.757
R3680 VDD.n2287 VDD.n1728 104.757
R3681 VDD.n2287 VDD.n1729 104.757
R3682 VDD.n2291 VDD.n1725 104.757
R3683 VDD.n2295 VDD.n1723 104.757
R3684 VDD.n2295 VDD.n1721 104.757
R3685 VDD.n2299 VDD.n1721 104.757
R3686 VDD.n2299 VDD.n1719 104.757
R3687 VDD.n2303 VDD.n1719 104.757
R3688 VDD.n2303 VDD.n1717 104.757
R3689 VDD.n2307 VDD.n1717 104.757
R3690 VDD.n2307 VDD.n1715 104.757
R3691 VDD.n2311 VDD.n1715 104.757
R3692 VDD.n2311 VDD.n1713 104.757
R3693 VDD.n2315 VDD.n1713 104.757
R3694 VDD.n2315 VDD.n1711 104.757
R3695 VDD.n2319 VDD.n1711 104.757
R3696 VDD.n2319 VDD.n1709 104.757
R3697 VDD.n2323 VDD.n1709 104.757
R3698 VDD.n2323 VDD.n1707 104.757
R3699 VDD.n2327 VDD.n1707 104.757
R3700 VDD.n2327 VDD.n1705 104.757
R3701 VDD.n2331 VDD.n1705 104.757
R3702 VDD.n2331 VDD.n1703 104.757
R3703 VDD.n2335 VDD.n1703 104.757
R3704 VDD.n2335 VDD.n1701 104.757
R3705 VDD.n2339 VDD.n1701 104.757
R3706 VDD.n2339 VDD.n1699 104.757
R3707 VDD.n2343 VDD.n1699 104.757
R3708 VDD.n2343 VDD.n1697 104.757
R3709 VDD.n2347 VDD.n1697 104.757
R3710 VDD.n2347 VDD.n1694 104.757
R3711 VDD.n2080 VDD.n1938 104.757
R3712 VDD.n2084 VDD.n1935 104.757
R3713 VDD.n2090 VDD.n1935 104.757
R3714 VDD.n2090 VDD.n1933 104.757
R3715 VDD.n2094 VDD.n1933 104.757
R3716 VDD.n2094 VDD.n1931 104.757
R3717 VDD.n2098 VDD.n1931 104.757
R3718 VDD.n2098 VDD.n1929 104.757
R3719 VDD.n2102 VDD.n1929 104.757
R3720 VDD.n2102 VDD.n1927 104.757
R3721 VDD.n2106 VDD.n1927 104.757
R3722 VDD.n2106 VDD.n1925 104.757
R3723 VDD.n2111 VDD.n1925 104.757
R3724 VDD.n2111 VDD.n1922 104.757
R3725 VDD.n2116 VDD.n1922 104.757
R3726 VDD.n2117 VDD.n2116 104.757
R3727 VDD.n2129 VDD.n1918 104.757
R3728 VDD.n2132 VDD.n2131 104.757
R3729 VDD.n2143 VDD.n2142 104.757
R3730 VDD.n2150 VDD.n2149 104.757
R3731 VDD.n2405 VDD.n2404 104.757
R3732 VDD.n2397 VDD.n1668 104.757
R3733 VDD.n2395 VDD.n1669 104.757
R3734 VDD.n2387 VDD.n2386 104.757
R3735 VDD.n2384 VDD.n1675 104.757
R3736 VDD.n2379 VDD.n1675 104.757
R3737 VDD.n2379 VDD.n1677 104.757
R3738 VDD.n2375 VDD.n1677 104.757
R3739 VDD.n2375 VDD.n1680 104.757
R3740 VDD.n2371 VDD.n1680 104.757
R3741 VDD.n2371 VDD.n1682 104.757
R3742 VDD.n2367 VDD.n1682 104.757
R3743 VDD.n2367 VDD.n1684 104.757
R3744 VDD.n2363 VDD.n1684 104.757
R3745 VDD.n2363 VDD.n1686 104.757
R3746 VDD.n2359 VDD.n1686 104.757
R3747 VDD.n2359 VDD.n1688 104.757
R3748 VDD.n2355 VDD.n1688 104.757
R3749 VDD.n2355 VDD.n1690 104.757
R3750 VDD.n2351 VDD.n1693 104.757
R3751 VDD.n12491 VDD.n6912 104.172
R3752 VDD.n12488 VDD.n12427 104.172
R3753 VDD.n12469 VDD.n12468 104.172
R3754 VDD.n12458 VDD.n12456 104.172
R3755 VDD.n9195 VDD.n9075 98.9686
R3756 VDD.n6212 VDD.n6074 96.8641
R3757 VDD.n5358 VDD.n5220 96.8641
R3758 VDD.n4572 VDD.n4434 96.8641
R3759 VDD.n3718 VDD.n3580 96.8641
R3760 VDD.n2932 VDD.n2794 96.8641
R3761 VDD.n2077 VDD.n1939 96.8641
R3762 VDD.n924 VDD.n881 96.8641
R3763 VDD.n478 VDD.n435 96.8641
R3764 VDD.t10 VDD.n5738 96.8274
R3765 VDD.t111 VDD.n4098 96.8274
R3766 VDD.t138 VDD.n2457 96.8274
R3767 VDD.t170 VDD.n817 96.8274
R3768 VDD.n6223 VDD.n6222 96.5084
R3769 VDD.n6112 VDD.n6106 96.5084
R3770 VDD.n5369 VDD.n5368 96.5084
R3771 VDD.n5258 VDD.n5252 96.5084
R3772 VDD.n4583 VDD.n4582 96.5084
R3773 VDD.n4472 VDD.n4466 96.5084
R3774 VDD.n3729 VDD.n3728 96.5084
R3775 VDD.n3618 VDD.n3612 96.5084
R3776 VDD.n2943 VDD.n2942 96.5084
R3777 VDD.n2832 VDD.n2826 96.5084
R3778 VDD.n2088 VDD.n2087 96.5084
R3779 VDD.n1977 VDD.n1971 96.5084
R3780 VDD.n9950 VDD.t196 92.7485
R3781 VDD.n8118 VDD.n8116 92.5005
R3782 VDD.n8115 VDD.n8104 92.5005
R3783 VDD.n8111 VDD.n8105 92.5005
R3784 VDD.n8189 VDD.n8188 92.5005
R3785 VDD.n8186 VDD.n8185 92.5005
R3786 VDD.n8128 VDD.n8126 92.5005
R3787 VDD.n8178 VDD.n8177 92.5005
R3788 VDD.n8176 VDD.n8175 92.5005
R3789 VDD.n8143 VDD.n8137 92.5005
R3790 VDD.n8168 VDD.n8167 92.5005
R3791 VDD.n8165 VDD.n8164 92.5005
R3792 VDD.n8146 VDD.n8144 92.5005
R3793 VDD.n8153 VDD.n8149 92.5005
R3794 VDD.n8156 VDD.n8155 92.5005
R3795 VDD.n8155 VDD.n8125 92.5005
R3796 VDD.n8157 VDD.n8150 92.5005
R3797 VDD.n8148 VDD.n8147 92.5005
R3798 VDD.n8163 VDD.n8162 92.5005
R3799 VDD.n8142 VDD.n8141 92.5005
R3800 VDD.n8140 VDD.n8139 92.5005
R3801 VDD.n8174 VDD.n8173 92.5005
R3802 VDD.n8133 VDD.n8132 92.5005
R3803 VDD.n8131 VDD.n8130 92.5005
R3804 VDD.n8184 VDD.n8183 92.5005
R3805 VDD.n8110 VDD.n8109 92.5005
R3806 VDD.n8108 VDD.n8103 92.5005
R3807 VDD.n8195 VDD.n8194 92.5005
R3808 VDD.n8154 VDD.n7745 92.5005
R3809 VDD.n8154 VDD.n7747 92.5005
R3810 VDD.n8602 VDD.n7720 92.5005
R3811 VDD.n7748 VDD.n7720 92.5005
R3812 VDD.n11446 VDD.n11445 92.5005
R3813 VDD.n11447 VDD.n11446 92.5005
R3814 VDD.n7726 VDD.n7721 92.5005
R3815 VDD.n7728 VDD.n7721 92.5005
R3816 VDD.n8612 VDD.n8611 92.5005
R3817 VDD.n8612 VDD.n7729 92.5005
R3818 VDD.n8613 VDD.n7738 92.5005
R3819 VDD.n8613 VDD.n7735 92.5005
R3820 VDD.n8614 VDD.n7739 92.5005
R3821 VDD.n9168 VDD.n8614 92.5005
R3822 VDD.n11428 VDD.n11427 92.5005
R3823 VDD.n11427 VDD.n11426 92.5005
R3824 VDD.n8621 VDD.n8615 92.5005
R3825 VDD.n8617 VDD.n8615 92.5005
R3826 VDD.n8643 VDD.n8642 92.5005
R3827 VDD.n8643 VDD.n8623 92.5005
R3828 VDD.n8644 VDD.n8632 92.5005
R3829 VDD.n8644 VDD.n8629 92.5005
R3830 VDD.n8645 VDD.n8633 92.5005
R3831 VDD.n8645 VDD.n8630 92.5005
R3832 VDD.n11409 VDD.n11408 92.5005
R3833 VDD.n11408 VDD.n11407 92.5005
R3834 VDD.n8652 VDD.n8646 92.5005
R3835 VDD.n8648 VDD.n8646 92.5005
R3836 VDD.n8676 VDD.n8675 92.5005
R3837 VDD.n8675 VDD.n8654 92.5005
R3838 VDD.n8664 VDD.n8662 92.5005
R3839 VDD.n8664 VDD.n8659 92.5005
R3840 VDD.n11394 VDD.n11393 92.5005
R3841 VDD.n11393 VDD.n8660 92.5005
R3842 VDD.n11392 VDD.n8667 92.5005
R3843 VDD.n11392 VDD.n11391 92.5005
R3844 VDD.n8672 VDD.n8665 92.5005
R3845 VDD.n8669 VDD.n8665 92.5005
R3846 VDD.n11384 VDD.n11383 92.5005
R3847 VDD.n11383 VDD.n11382 92.5005
R3848 VDD.n8690 VDD.n8684 92.5005
R3849 VDD.n8686 VDD.n8684 92.5005
R3850 VDD.n8715 VDD.n8714 92.5005
R3851 VDD.n8715 VDD.n8692 92.5005
R3852 VDD.n8716 VDD.n8704 92.5005
R3853 VDD.n8716 VDD.n8701 92.5005
R3854 VDD.n8717 VDD.n8705 92.5005
R3855 VDD.n8717 VDD.n8702 92.5005
R3856 VDD.n11365 VDD.n11364 92.5005
R3857 VDD.n11364 VDD.n11363 92.5005
R3858 VDD.n8725 VDD.n8718 92.5005
R3859 VDD.n11027 VDD.n8718 92.5005
R3860 VDD.n11048 VDD.n11047 92.5005
R3861 VDD.n11048 VDD.n11028 92.5005
R3862 VDD.n11049 VDD.n11037 92.5005
R3863 VDD.n11049 VDD.n11034 92.5005
R3864 VDD.n11050 VDD.n11038 92.5005
R3865 VDD.n11050 VDD.n11035 92.5005
R3866 VDD.n11346 VDD.n11345 92.5005
R3867 VDD.n11345 VDD.n11344 92.5005
R3868 VDD.n11057 VDD.n11051 92.5005
R3869 VDD.n11053 VDD.n11051 92.5005
R3870 VDD.n11097 VDD.n11094 92.5005
R3871 VDD.n11097 VDD.n11096 92.5005
R3872 VDD.n11098 VDD.n11066 92.5005
R3873 VDD.n11098 VDD.n11063 92.5005
R3874 VDD.n11099 VDD.n11067 92.5005
R3875 VDD.n11099 VDD.n11064 92.5005
R3876 VDD.n11100 VDD.n11071 92.5005
R3877 VDD.n11100 VDD.n11075 92.5005
R3878 VDD.n11101 VDD.n11072 92.5005
R3879 VDD.n11101 VDD.n11076 92.5005
R3880 VDD.n11102 VDD.n11085 92.5005
R3881 VDD.n11102 VDD.n11081 92.5005
R3882 VDD.n11103 VDD.n11086 92.5005
R3883 VDD.n11103 VDD.n11082 92.5005
R3884 VDD.n11312 VDD.n11311 92.5005
R3885 VDD.n11311 VDD.n11310 92.5005
R3886 VDD.n11110 VDD.n11104 92.5005
R3887 VDD.n11106 VDD.n11104 92.5005
R3888 VDD.n11132 VDD.n11131 92.5005
R3889 VDD.n11132 VDD.n11112 92.5005
R3890 VDD.n11133 VDD.n11121 92.5005
R3891 VDD.n11133 VDD.n11118 92.5005
R3892 VDD.n11134 VDD.n11122 92.5005
R3893 VDD.n11134 VDD.n11119 92.5005
R3894 VDD.n11293 VDD.n11292 92.5005
R3895 VDD.n11292 VDD.n11291 92.5005
R3896 VDD.n11140 VDD.n11135 92.5005
R3897 VDD.n11142 VDD.n11135 92.5005
R3898 VDD.n11163 VDD.n11162 92.5005
R3899 VDD.n11163 VDD.n11143 92.5005
R3900 VDD.n11164 VDD.n11152 92.5005
R3901 VDD.n11164 VDD.n11149 92.5005
R3902 VDD.n11165 VDD.n11153 92.5005
R3903 VDD.n11165 VDD.n11150 92.5005
R3904 VDD.n11274 VDD.n11273 92.5005
R3905 VDD.n11273 VDD.n11272 92.5005
R3906 VDD.n11172 VDD.n11166 92.5005
R3907 VDD.n11168 VDD.n11166 92.5005
R3908 VDD.n11197 VDD.n11196 92.5005
R3909 VDD.n11196 VDD.n11174 92.5005
R3910 VDD.n11185 VDD.n11183 92.5005
R3911 VDD.n11185 VDD.n11180 92.5005
R3912 VDD.n11259 VDD.n11258 92.5005
R3913 VDD.n11258 VDD.n11181 92.5005
R3914 VDD.n11257 VDD.n11188 92.5005
R3915 VDD.n11257 VDD.n11256 92.5005
R3916 VDD.n11193 VDD.n11186 92.5005
R3917 VDD.n11190 VDD.n11186 92.5005
R3918 VDD.n11249 VDD.n11248 92.5005
R3919 VDD.n11248 VDD.n11247 92.5005
R3920 VDD.n11211 VDD.n11205 92.5005
R3921 VDD.n11207 VDD.n11205 92.5005
R3922 VDD.n11223 VDD.n11215 92.5005
R3923 VDD.n11215 VDD.n11213 92.5005
R3924 VDD.n11231 VDD.n11230 92.5005
R3925 VDD.n11232 VDD.n11231 92.5005
R3926 VDD.n11221 VDD.n6603 92.5005
R3927 VDD.n11221 VDD.n6599 92.5005
R3928 VDD.n11220 VDD.n6604 92.5005
R3929 VDD.n11220 VDD.n6600 92.5005
R3930 VDD.n12709 VDD.n12708 92.5005
R3931 VDD.n12710 VDD.n12709 92.5005
R3932 VDD.n11229 VDD.n6601 92.5005
R3933 VDD.n11214 VDD.n6601 92.5005
R3934 VDD.n11222 VDD.n11209 92.5005
R3935 VDD.n11233 VDD.n11209 92.5005
R3936 VDD.n11244 VDD.n11212 92.5005
R3937 VDD.n11244 VDD.n11243 92.5005
R3938 VDD.n11245 VDD.n11204 92.5005
R3939 VDD.n11246 VDD.n11245 92.5005
R3940 VDD.n11203 VDD.n11192 92.5005
R3941 VDD.n11206 VDD.n11192 92.5005
R3942 VDD.n11254 VDD.n11253 92.5005
R3943 VDD.n11255 VDD.n11254 92.5005
R3944 VDD.n11187 VDD.n11182 92.5005
R3945 VDD.n11189 VDD.n11182 92.5005
R3946 VDD.n11261 VDD.n11260 92.5005
R3947 VDD.n11262 VDD.n11261 92.5005
R3948 VDD.n11198 VDD.n11170 92.5005
R3949 VDD.n11179 VDD.n11170 92.5005
R3950 VDD.n11269 VDD.n11173 92.5005
R3951 VDD.n11269 VDD.n11268 92.5005
R3952 VDD.n11270 VDD.n11157 92.5005
R3953 VDD.n11271 VDD.n11270 92.5005
R3954 VDD.n11156 VDD.n11151 92.5005
R3955 VDD.n11167 VDD.n11151 92.5005
R3956 VDD.n11280 VDD.n11279 92.5005
R3957 VDD.n11281 VDD.n11280 92.5005
R3958 VDD.n11161 VDD.n11138 92.5005
R3959 VDD.n11148 VDD.n11138 92.5005
R3960 VDD.n11288 VDD.n11141 92.5005
R3961 VDD.n11288 VDD.n11287 92.5005
R3962 VDD.n11289 VDD.n11126 92.5005
R3963 VDD.n11290 VDD.n11289 92.5005
R3964 VDD.n11125 VDD.n11120 92.5005
R3965 VDD.n11136 VDD.n11120 92.5005
R3966 VDD.n11299 VDD.n11298 92.5005
R3967 VDD.n11300 VDD.n11299 92.5005
R3968 VDD.n11130 VDD.n11108 92.5005
R3969 VDD.n11117 VDD.n11108 92.5005
R3970 VDD.n11307 VDD.n11111 92.5005
R3971 VDD.n11307 VDD.n11306 92.5005
R3972 VDD.n11308 VDD.n11089 92.5005
R3973 VDD.n11309 VDD.n11308 92.5005
R3974 VDD.n11088 VDD.n11083 92.5005
R3975 VDD.n11105 VDD.n11083 92.5005
R3976 VDD.n11318 VDD.n11317 92.5005
R3977 VDD.n11319 VDD.n11318 92.5005
R3978 VDD.n11084 VDD.n11073 92.5005
R3979 VDD.n11080 VDD.n11073 92.5005
R3980 VDD.n11327 VDD.n11326 92.5005
R3981 VDD.n11326 VDD.n11325 92.5005
R3982 VDD.n11070 VDD.n11065 92.5005
R3983 VDD.n11074 VDD.n11065 92.5005
R3984 VDD.n11333 VDD.n11332 92.5005
R3985 VDD.n11334 VDD.n11333 92.5005
R3986 VDD.n11093 VDD.n11055 92.5005
R3987 VDD.n11095 VDD.n11055 92.5005
R3988 VDD.n11341 VDD.n11058 92.5005
R3989 VDD.n11341 VDD.n11340 92.5005
R3990 VDD.n11342 VDD.n11042 92.5005
R3991 VDD.n11343 VDD.n11342 92.5005
R3992 VDD.n11041 VDD.n11036 92.5005
R3993 VDD.n11052 VDD.n11036 92.5005
R3994 VDD.n11352 VDD.n11351 92.5005
R3995 VDD.n11353 VDD.n11352 92.5005
R3996 VDD.n11046 VDD.n8723 92.5005
R3997 VDD.n11033 VDD.n8723 92.5005
R3998 VDD.n11360 VDD.n8726 92.5005
R3999 VDD.n11360 VDD.n11359 92.5005
R4000 VDD.n11361 VDD.n8709 92.5005
R4001 VDD.n11362 VDD.n11361 92.5005
R4002 VDD.n8708 VDD.n8703 92.5005
R4003 VDD.n8719 VDD.n8703 92.5005
R4004 VDD.n11371 VDD.n11370 92.5005
R4005 VDD.n11372 VDD.n11371 92.5005
R4006 VDD.n8713 VDD.n8688 92.5005
R4007 VDD.n8700 VDD.n8688 92.5005
R4008 VDD.n11379 VDD.n8691 92.5005
R4009 VDD.n11379 VDD.n11378 92.5005
R4010 VDD.n11380 VDD.n8683 92.5005
R4011 VDD.n11381 VDD.n11380 92.5005
R4012 VDD.n8682 VDD.n8671 92.5005
R4013 VDD.n8685 VDD.n8671 92.5005
R4014 VDD.n11389 VDD.n11388 92.5005
R4015 VDD.n11390 VDD.n11389 92.5005
R4016 VDD.n8666 VDD.n8661 92.5005
R4017 VDD.n8668 VDD.n8661 92.5005
R4018 VDD.n11396 VDD.n11395 92.5005
R4019 VDD.n11397 VDD.n11396 92.5005
R4020 VDD.n8677 VDD.n8650 92.5005
R4021 VDD.n9176 VDD.n8650 92.5005
R4022 VDD.n11404 VDD.n8653 92.5005
R4023 VDD.n11404 VDD.n11403 92.5005
R4024 VDD.n11405 VDD.n8637 92.5005
R4025 VDD.n11406 VDD.n11405 92.5005
R4026 VDD.n8636 VDD.n8631 92.5005
R4027 VDD.n8647 VDD.n8631 92.5005
R4028 VDD.n11415 VDD.n11414 92.5005
R4029 VDD.n11416 VDD.n11415 92.5005
R4030 VDD.n8641 VDD.n8619 92.5005
R4031 VDD.n8628 VDD.n8619 92.5005
R4032 VDD.n11423 VDD.n8622 92.5005
R4033 VDD.n11423 VDD.n11422 92.5005
R4034 VDD.n11424 VDD.n7743 92.5005
R4035 VDD.n11425 VDD.n11424 92.5005
R4036 VDD.n7742 VDD.n7737 92.5005
R4037 VDD.n8616 VDD.n7737 92.5005
R4038 VDD.n11434 VDD.n11433 92.5005
R4039 VDD.n11435 VDD.n11434 92.5005
R4040 VDD.n8610 VDD.n7725 92.5005
R4041 VDD.n9172 VDD.n7725 92.5005
R4042 VDD.n11442 VDD.n7727 92.5005
R4043 VDD.n11442 VDD.n11441 92.5005
R4044 VDD.n11444 VDD.n11443 92.5005
R4045 VDD.n11443 VDD.n7719 92.5005
R4046 VDD.n8601 VDD.n7724 92.5005
R4047 VDD.n7724 VDD.n7718 92.5005
R4048 VDD.n8600 VDD.n8599 92.5005
R4049 VDD.n8599 VDD.n8598 92.5005
R4050 VDD.n8151 VDD.n7746 92.5005
R4051 VDD.n8499 VDD.n7746 92.5005
R4052 VDD.n12413 VDD.n12412 92.5005
R4053 VDD.n12410 VDD.n6930 92.5005
R4054 VDD.n12409 VDD.n12408 92.5005
R4055 VDD.n12409 VDD.n6932 92.5005
R4056 VDD.n6938 VDD.n6933 92.5005
R4057 VDD.n6939 VDD.n6936 92.5005
R4058 VDD.n12406 VDD.n12405 92.5005
R4059 VDD.n12405 VDD.n12404 92.5005
R4060 VDD.n6942 VDD.n6937 92.5005
R4061 VDD.n12403 VDD.n6937 92.5005
R4062 VDD.n12401 VDD.n12400 92.5005
R4063 VDD.n12402 VDD.n12401 92.5005
R4064 VDD.n6944 VDD.n6941 92.5005
R4065 VDD.n6941 VDD.n6940 92.5005
R4066 VDD.n12395 VDD.n12394 92.5005
R4067 VDD.n12394 VDD.n12393 92.5005
R4068 VDD.n6951 VDD.n6948 92.5005
R4069 VDD.n12392 VDD.n6948 92.5005
R4070 VDD.n12390 VDD.n12389 92.5005
R4071 VDD.n12391 VDD.n12390 92.5005
R4072 VDD.n6953 VDD.n6950 92.5005
R4073 VDD.n6950 VDD.n6949 92.5005
R4074 VDD.n12384 VDD.n12383 92.5005
R4075 VDD.n12383 VDD.n12382 92.5005
R4076 VDD.n6960 VDD.n6957 92.5005
R4077 VDD.n12381 VDD.n6957 92.5005
R4078 VDD.n12379 VDD.n12378 92.5005
R4079 VDD.n12380 VDD.n12379 92.5005
R4080 VDD.n6962 VDD.n6959 92.5005
R4081 VDD.n6959 VDD.n6958 92.5005
R4082 VDD.n12373 VDD.n12372 92.5005
R4083 VDD.n12372 VDD.n12371 92.5005
R4084 VDD.n6970 VDD.n6966 92.5005
R4085 VDD.n12370 VDD.n6966 92.5005
R4086 VDD.n12368 VDD.n12367 92.5005
R4087 VDD.n12369 VDD.n12368 92.5005
R4088 VDD.n6972 VDD.n6969 92.5005
R4089 VDD.n6969 VDD.n6968 92.5005
R4090 VDD.n12362 VDD.n12361 92.5005
R4091 VDD.n12361 VDD.n12360 92.5005
R4092 VDD.n6976 VDD.n6975 92.5005
R4093 VDD.n12359 VDD.n6976 92.5005
R4094 VDD.n12357 VDD.n12356 92.5005
R4095 VDD.n12358 VDD.n12357 92.5005
R4096 VDD.n6980 VDD.n6978 92.5005
R4097 VDD.n6978 VDD.n6977 92.5005
R4098 VDD.n12351 VDD.n12350 92.5005
R4099 VDD.n12350 VDD.n12349 92.5005
R4100 VDD.n6986 VDD.n6983 92.5005
R4101 VDD.n12348 VDD.n6983 92.5005
R4102 VDD.n12346 VDD.n12345 92.5005
R4103 VDD.n12347 VDD.n12346 92.5005
R4104 VDD.n6988 VDD.n6985 92.5005
R4105 VDD.n6985 VDD.n6984 92.5005
R4106 VDD.n12340 VDD.n12339 92.5005
R4107 VDD.n12339 VDD.n12338 92.5005
R4108 VDD.n6995 VDD.n6992 92.5005
R4109 VDD.n12337 VDD.n6992 92.5005
R4110 VDD.n12335 VDD.n12334 92.5005
R4111 VDD.n12336 VDD.n12335 92.5005
R4112 VDD.n6997 VDD.n6994 92.5005
R4113 VDD.n6994 VDD.n6993 92.5005
R4114 VDD.n12329 VDD.n12328 92.5005
R4115 VDD.n12328 VDD.n12327 92.5005
R4116 VDD.n7004 VDD.n7001 92.5005
R4117 VDD.n12326 VDD.n7001 92.5005
R4118 VDD.n12324 VDD.n12323 92.5005
R4119 VDD.n12325 VDD.n12324 92.5005
R4120 VDD.n7006 VDD.n7003 92.5005
R4121 VDD.n7003 VDD.n7002 92.5005
R4122 VDD.n12318 VDD.n12317 92.5005
R4123 VDD.n12317 VDD.n12316 92.5005
R4124 VDD.n7013 VDD.n7010 92.5005
R4125 VDD.n12315 VDD.n7010 92.5005
R4126 VDD.n12313 VDD.n12312 92.5005
R4127 VDD.n12314 VDD.n12313 92.5005
R4128 VDD.n12311 VDD.n7012 92.5005
R4129 VDD.n7012 VDD.n7011 92.5005
R4130 VDD.n7019 VDD.n7015 92.5005
R4131 VDD.n7021 VDD.n7019 92.5005
R4132 VDD.n12306 VDD.n12305 92.5005
R4133 VDD.n12305 VDD.n12304 92.5005
R4134 VDD.n7024 VDD.n7020 92.5005
R4135 VDD.n12303 VDD.n7020 92.5005
R4136 VDD.n12301 VDD.n12300 92.5005
R4137 VDD.n12302 VDD.n12301 92.5005
R4138 VDD.n7026 VDD.n7023 92.5005
R4139 VDD.n7023 VDD.n7022 92.5005
R4140 VDD.n12295 VDD.n12294 92.5005
R4141 VDD.n12294 VDD.n12293 92.5005
R4142 VDD.n7033 VDD.n7030 92.5005
R4143 VDD.n12292 VDD.n7030 92.5005
R4144 VDD.n12290 VDD.n12289 92.5005
R4145 VDD.n12291 VDD.n12290 92.5005
R4146 VDD.n7035 VDD.n7032 92.5005
R4147 VDD.n7032 VDD.n7031 92.5005
R4148 VDD.n12284 VDD.n12283 92.5005
R4149 VDD.n12283 VDD.n12282 92.5005
R4150 VDD.n7042 VDD.n7039 92.5005
R4151 VDD.n12281 VDD.n7039 92.5005
R4152 VDD.n12279 VDD.n12278 92.5005
R4153 VDD.n12280 VDD.n12279 92.5005
R4154 VDD.n7044 VDD.n7041 92.5005
R4155 VDD.n7041 VDD.n7040 92.5005
R4156 VDD.n12273 VDD.n12272 92.5005
R4157 VDD.n12272 VDD.n12271 92.5005
R4158 VDD.n7051 VDD.n7048 92.5005
R4159 VDD.n12270 VDD.n7048 92.5005
R4160 VDD.n12268 VDD.n12267 92.5005
R4161 VDD.n12269 VDD.n12268 92.5005
R4162 VDD.n7053 VDD.n7050 92.5005
R4163 VDD.n7050 VDD.n7049 92.5005
R4164 VDD.n7058 VDD.n7056 92.5005
R4165 VDD.n7060 VDD.n7058 92.5005
R4166 VDD.n12262 VDD.n12261 92.5005
R4167 VDD.n12261 VDD.n12260 92.5005
R4168 VDD.n7063 VDD.n7059 92.5005
R4169 VDD.n12259 VDD.n7059 92.5005
R4170 VDD.n12257 VDD.n12256 92.5005
R4171 VDD.n12258 VDD.n12257 92.5005
R4172 VDD.n7065 VDD.n7062 92.5005
R4173 VDD.n7062 VDD.n7061 92.5005
R4174 VDD.n12251 VDD.n12250 92.5005
R4175 VDD.n12250 VDD.n12249 92.5005
R4176 VDD.n7128 VDD.n7069 92.5005
R4177 VDD.n7132 VDD.n7131 92.5005
R4178 VDD.n7135 VDD.n7134 92.5005
R4179 VDD.n7124 VDD.n7123 92.5005
R4180 VDD.n7141 VDD.n7140 92.5005
R4181 VDD.n7145 VDD.n7144 92.5005
R4182 VDD.n7143 VDD.n7120 92.5005
R4183 VDD.n7151 VDD.n7150 92.5005
R4184 VDD.n7154 VDD.n7153 92.5005
R4185 VDD.n7116 VDD.n7115 92.5005
R4186 VDD.n7161 VDD.n7160 92.5005
R4187 VDD.n7163 VDD.n7114 92.5005
R4188 VDD.n7166 VDD.n7165 92.5005
R4189 VDD.n7112 VDD.n7111 92.5005
R4190 VDD.n7172 VDD.n7171 92.5005
R4191 VDD.n7176 VDD.n7175 92.5005
R4192 VDD.n7174 VDD.n7108 92.5005
R4193 VDD.n7182 VDD.n7181 92.5005
R4194 VDD.n7185 VDD.n7184 92.5005
R4195 VDD.n7104 VDD.n7103 92.5005
R4196 VDD.n7191 VDD.n7190 92.5005
R4197 VDD.n7195 VDD.n7194 92.5005
R4198 VDD.n7193 VDD.n7100 92.5005
R4199 VDD.n7201 VDD.n7200 92.5005
R4200 VDD.n7204 VDD.n7203 92.5005
R4201 VDD.n7096 VDD.n7095 92.5005
R4202 VDD.n7210 VDD.n7209 92.5005
R4203 VDD.n7215 VDD.n7214 92.5005
R4204 VDD.n7213 VDD.n7092 92.5005
R4205 VDD.n7220 VDD.n7091 92.5005
R4206 VDD.n7222 VDD.n7221 92.5005
R4207 VDD.n7226 VDD.n7225 92.5005
R4208 VDD.n7224 VDD.n7088 92.5005
R4209 VDD.n7232 VDD.n7231 92.5005
R4210 VDD.n7235 VDD.n7234 92.5005
R4211 VDD.n7084 VDD.n7083 92.5005
R4212 VDD.n7241 VDD.n7240 92.5005
R4213 VDD.n7245 VDD.n7244 92.5005
R4214 VDD.n7243 VDD.n7080 92.5005
R4215 VDD.n7251 VDD.n7250 92.5005
R4216 VDD.n7254 VDD.n7253 92.5005
R4217 VDD.n7255 VDD.n7073 92.5005
R4218 VDD.n12246 VDD.n12245 92.5005
R4219 VDD.n12247 VDD.n12246 92.5005
R4220 VDD.n7076 VDD.n7074 92.5005
R4221 VDD.n7074 VDD.n7072 92.5005
R4222 VDD.n12240 VDD.n12239 92.5005
R4223 VDD.n12239 VDD.n12238 92.5005
R4224 VDD.n7264 VDD.n7261 92.5005
R4225 VDD.n12237 VDD.n7261 92.5005
R4226 VDD.n12235 VDD.n12234 92.5005
R4227 VDD.n12236 VDD.n12235 92.5005
R4228 VDD.n7266 VDD.n7263 92.5005
R4229 VDD.n7263 VDD.n7262 92.5005
R4230 VDD.n7271 VDD.n7269 92.5005
R4231 VDD.n7273 VDD.n7271 92.5005
R4232 VDD.n12229 VDD.n12228 92.5005
R4233 VDD.n12228 VDD.n12227 92.5005
R4234 VDD.n7276 VDD.n7272 92.5005
R4235 VDD.n12226 VDD.n7272 92.5005
R4236 VDD.n12224 VDD.n12223 92.5005
R4237 VDD.n12225 VDD.n12224 92.5005
R4238 VDD.n7278 VDD.n7275 92.5005
R4239 VDD.n7275 VDD.n7274 92.5005
R4240 VDD.n12218 VDD.n12217 92.5005
R4241 VDD.n12217 VDD.n12216 92.5005
R4242 VDD.n7285 VDD.n7282 92.5005
R4243 VDD.n12215 VDD.n7282 92.5005
R4244 VDD.n12213 VDD.n12212 92.5005
R4245 VDD.n12214 VDD.n12213 92.5005
R4246 VDD.n7287 VDD.n7284 92.5005
R4247 VDD.n7284 VDD.n7283 92.5005
R4248 VDD.n12207 VDD.n12206 92.5005
R4249 VDD.n12206 VDD.n12205 92.5005
R4250 VDD.n7294 VDD.n7291 92.5005
R4251 VDD.n12204 VDD.n7291 92.5005
R4252 VDD.n12202 VDD.n12201 92.5005
R4253 VDD.n12203 VDD.n12202 92.5005
R4254 VDD.n7296 VDD.n7293 92.5005
R4255 VDD.n7293 VDD.n7292 92.5005
R4256 VDD.n12196 VDD.n12195 92.5005
R4257 VDD.n12195 VDD.n12194 92.5005
R4258 VDD.n7303 VDD.n7300 92.5005
R4259 VDD.n12193 VDD.n7300 92.5005
R4260 VDD.n12191 VDD.n12190 92.5005
R4261 VDD.n12192 VDD.n12191 92.5005
R4262 VDD.n7305 VDD.n7302 92.5005
R4263 VDD.n7302 VDD.n7301 92.5005
R4264 VDD.n12185 VDD.n12184 92.5005
R4265 VDD.n12184 VDD.n12183 92.5005
R4266 VDD.n7309 VDD.n7308 92.5005
R4267 VDD.n12182 VDD.n7309 92.5005
R4268 VDD.n12180 VDD.n12179 92.5005
R4269 VDD.n12181 VDD.n12180 92.5005
R4270 VDD.n7313 VDD.n7311 92.5005
R4271 VDD.n7311 VDD.n7310 92.5005
R4272 VDD.n12174 VDD.n12173 92.5005
R4273 VDD.n12173 VDD.n12172 92.5005
R4274 VDD.n7319 VDD.n7316 92.5005
R4275 VDD.n12171 VDD.n7316 92.5005
R4276 VDD.n12169 VDD.n12168 92.5005
R4277 VDD.n12170 VDD.n12169 92.5005
R4278 VDD.n7321 VDD.n7318 92.5005
R4279 VDD.n7318 VDD.n7317 92.5005
R4280 VDD.n12163 VDD.n12162 92.5005
R4281 VDD.n12162 VDD.n12161 92.5005
R4282 VDD.n7328 VDD.n7325 92.5005
R4283 VDD.n12160 VDD.n7325 92.5005
R4284 VDD.n12158 VDD.n12157 92.5005
R4285 VDD.n12159 VDD.n12158 92.5005
R4286 VDD.n7330 VDD.n7327 92.5005
R4287 VDD.n7327 VDD.n7326 92.5005
R4288 VDD.n12152 VDD.n12151 92.5005
R4289 VDD.n12151 VDD.n12150 92.5005
R4290 VDD.n7337 VDD.n7334 92.5005
R4291 VDD.n12149 VDD.n7334 92.5005
R4292 VDD.n12147 VDD.n12146 92.5005
R4293 VDD.n12148 VDD.n12147 92.5005
R4294 VDD.n7339 VDD.n7336 92.5005
R4295 VDD.n7336 VDD.n7335 92.5005
R4296 VDD.n12141 VDD.n12140 92.5005
R4297 VDD.n12140 VDD.n12139 92.5005
R4298 VDD.n7346 VDD.n7343 92.5005
R4299 VDD.n12138 VDD.n7343 92.5005
R4300 VDD.n12136 VDD.n12135 92.5005
R4301 VDD.n12137 VDD.n12136 92.5005
R4302 VDD.n12134 VDD.n7345 92.5005
R4303 VDD.n7345 VDD.n7344 92.5005
R4304 VDD.n7352 VDD.n7348 92.5005
R4305 VDD.n7354 VDD.n7352 92.5005
R4306 VDD.n12129 VDD.n12128 92.5005
R4307 VDD.n12128 VDD.n12127 92.5005
R4308 VDD.n7353 VDD.n7351 92.5005
R4309 VDD.n12126 VDD.n7353 92.5005
R4310 VDD.n12124 VDD.n12123 92.5005
R4311 VDD.n12125 VDD.n12124 92.5005
R4312 VDD.n12122 VDD.n7356 92.5005
R4313 VDD.n7356 VDD.n7355 92.5005
R4314 VDD.n12121 VDD.n12120 92.5005
R4315 VDD.n12120 VDD.n12119 92.5005
R4316 VDD.n7358 VDD.n7357 92.5005
R4317 VDD.n12118 VDD.n7358 92.5005
R4318 VDD.n12116 VDD.n12115 92.5005
R4319 VDD.n12117 VDD.n12116 92.5005
R4320 VDD.n12114 VDD.n7360 92.5005
R4321 VDD.n7360 VDD.n7359 92.5005
R4322 VDD.n12113 VDD.n12112 92.5005
R4323 VDD.n12112 VDD.n12111 92.5005
R4324 VDD.n7362 VDD.n7361 92.5005
R4325 VDD.n12110 VDD.n7362 92.5005
R4326 VDD.n12108 VDD.n12107 92.5005
R4327 VDD.n12109 VDD.n12108 92.5005
R4328 VDD.n12106 VDD.n7364 92.5005
R4329 VDD.n7364 VDD.n7363 92.5005
R4330 VDD.n12105 VDD.n12104 92.5005
R4331 VDD.n12104 VDD.n12103 92.5005
R4332 VDD.n7366 VDD.n7365 92.5005
R4333 VDD.n12102 VDD.n7366 92.5005
R4334 VDD.n12100 VDD.n12099 92.5005
R4335 VDD.n12101 VDD.n12100 92.5005
R4336 VDD.n12098 VDD.n7368 92.5005
R4337 VDD.n7368 VDD.n7367 92.5005
R4338 VDD.n12097 VDD.n12096 92.5005
R4339 VDD.n12096 VDD.n12095 92.5005
R4340 VDD.n7370 VDD.n7369 92.5005
R4341 VDD.n12094 VDD.n7370 92.5005
R4342 VDD.n12092 VDD.n7372 92.5005
R4343 VDD.n12092 VDD.n12091 92.5005
R4344 VDD.n12088 VDD.n12087 92.5005
R4345 VDD.n12087 VDD.n7371 92.5005
R4346 VDD.n12086 VDD.n7376 92.5005
R4347 VDD.n12086 VDD.n12085 92.5005
R4348 VDD.n12080 VDD.n7375 92.5005
R4349 VDD.n12084 VDD.n7375 92.5005
R4350 VDD.n12082 VDD.n12081 92.5005
R4351 VDD.n12083 VDD.n12082 92.5005
R4352 VDD.n12073 VDD.n7378 92.5005
R4353 VDD.n7378 VDD.n7377 92.5005
R4354 VDD.n12072 VDD.n12071 92.5005
R4355 VDD.n12071 VDD.n12070 92.5005
R4356 VDD.n7386 VDD.n7382 92.5005
R4357 VDD.n12069 VDD.n7382 92.5005
R4358 VDD.n12067 VDD.n12066 92.5005
R4359 VDD.n12068 VDD.n12067 92.5005
R4360 VDD.n12060 VDD.n7384 92.5005
R4361 VDD.n7384 VDD.n7383 92.5005
R4362 VDD.n12059 VDD.n12058 92.5005
R4363 VDD.n12058 VDD.n12057 92.5005
R4364 VDD.n7393 VDD.n7389 92.5005
R4365 VDD.n12056 VDD.n7389 92.5005
R4366 VDD.n12054 VDD.n12053 92.5005
R4367 VDD.n12055 VDD.n12054 92.5005
R4368 VDD.n12047 VDD.n7391 92.5005
R4369 VDD.n7391 VDD.n7390 92.5005
R4370 VDD.n12046 VDD.n12045 92.5005
R4371 VDD.n12045 VDD.n12044 92.5005
R4372 VDD.n7400 VDD.n7396 92.5005
R4373 VDD.n12043 VDD.n7396 92.5005
R4374 VDD.n12041 VDD.n12040 92.5005
R4375 VDD.n12042 VDD.n12041 92.5005
R4376 VDD.n12034 VDD.n7398 92.5005
R4377 VDD.n7398 VDD.n7397 92.5005
R4378 VDD.n12033 VDD.n12032 92.5005
R4379 VDD.n12032 VDD.n12031 92.5005
R4380 VDD.n7407 VDD.n7403 92.5005
R4381 VDD.n12030 VDD.n7403 92.5005
R4382 VDD.n12028 VDD.n12027 92.5005
R4383 VDD.n12029 VDD.n12028 92.5005
R4384 VDD.n7410 VDD.n7405 92.5005
R4385 VDD.n7405 VDD.n7404 92.5005
R4386 VDD.n12021 VDD.n12020 92.5005
R4387 VDD.n12020 VDD.n12019 92.5005
R4388 VDD.n7411 VDD.n7409 92.5005
R4389 VDD.n12018 VDD.n7411 92.5005
R4390 VDD.n12016 VDD.n12015 92.5005
R4391 VDD.n12017 VDD.n12016 92.5005
R4392 VDD.n7414 VDD.n7413 92.5005
R4393 VDD.n7413 VDD.n7412 92.5005
R4394 VDD.n12009 VDD.n12008 92.5005
R4395 VDD.n12008 VDD.n12007 92.5005
R4396 VDD.n7421 VDD.n7417 92.5005
R4397 VDD.n12006 VDD.n7417 92.5005
R4398 VDD.n12004 VDD.n12003 92.5005
R4399 VDD.n12005 VDD.n12004 92.5005
R4400 VDD.n11997 VDD.n7419 92.5005
R4401 VDD.n7419 VDD.n7418 92.5005
R4402 VDD.n11996 VDD.n11995 92.5005
R4403 VDD.n11995 VDD.n11994 92.5005
R4404 VDD.n7428 VDD.n7424 92.5005
R4405 VDD.n11993 VDD.n7424 92.5005
R4406 VDD.n11991 VDD.n11990 92.5005
R4407 VDD.n11992 VDD.n11991 92.5005
R4408 VDD.n11984 VDD.n7426 92.5005
R4409 VDD.n7426 VDD.n7425 92.5005
R4410 VDD.n11983 VDD.n11982 92.5005
R4411 VDD.n11982 VDD.n11981 92.5005
R4412 VDD.n7435 VDD.n7431 92.5005
R4413 VDD.n11980 VDD.n7431 92.5005
R4414 VDD.n11978 VDD.n11977 92.5005
R4415 VDD.n11979 VDD.n11978 92.5005
R4416 VDD.n11971 VDD.n7433 92.5005
R4417 VDD.n7433 VDD.n7432 92.5005
R4418 VDD.n11970 VDD.n11969 92.5005
R4419 VDD.n11969 VDD.n11968 92.5005
R4420 VDD.n11963 VDD.n7438 92.5005
R4421 VDD.n11967 VDD.n7438 92.5005
R4422 VDD.n11965 VDD.n11964 92.5005
R4423 VDD.n11966 VDD.n11965 92.5005
R4424 VDD.n7441 VDD.n7440 92.5005
R4425 VDD.n7440 VDD.n7439 92.5005
R4426 VDD.n11958 VDD.n11957 92.5005
R4427 VDD.n11957 VDD.n11956 92.5005
R4428 VDD.n7448 VDD.n7444 92.5005
R4429 VDD.n11955 VDD.n7444 92.5005
R4430 VDD.n11953 VDD.n11952 92.5005
R4431 VDD.n11954 VDD.n11953 92.5005
R4432 VDD.n11946 VDD.n7446 92.5005
R4433 VDD.n7446 VDD.n7445 92.5005
R4434 VDD.n11945 VDD.n11944 92.5005
R4435 VDD.n11944 VDD.n11943 92.5005
R4436 VDD.n7455 VDD.n7451 92.5005
R4437 VDD.n11942 VDD.n7451 92.5005
R4438 VDD.n11940 VDD.n11939 92.5005
R4439 VDD.n11941 VDD.n11940 92.5005
R4440 VDD.n11933 VDD.n7453 92.5005
R4441 VDD.n7453 VDD.n7452 92.5005
R4442 VDD.n11932 VDD.n11931 92.5005
R4443 VDD.n11931 VDD.n11930 92.5005
R4444 VDD.n7462 VDD.n7458 92.5005
R4445 VDD.n11929 VDD.n7458 92.5005
R4446 VDD.n11927 VDD.n11926 92.5005
R4447 VDD.n11928 VDD.n11927 92.5005
R4448 VDD.n11920 VDD.n7460 92.5005
R4449 VDD.n7460 VDD.n7459 92.5005
R4450 VDD.n11919 VDD.n11918 92.5005
R4451 VDD.n11918 VDD.n11917 92.5005
R4452 VDD.n7469 VDD.n7465 92.5005
R4453 VDD.n11916 VDD.n7465 92.5005
R4454 VDD.n11914 VDD.n11913 92.5005
R4455 VDD.n11915 VDD.n11914 92.5005
R4456 VDD.n7472 VDD.n7467 92.5005
R4457 VDD.n7467 VDD.n7466 92.5005
R4458 VDD.n11907 VDD.n11906 92.5005
R4459 VDD.n11906 VDD.n11905 92.5005
R4460 VDD.n7473 VDD.n7471 92.5005
R4461 VDD.n11904 VDD.n7473 92.5005
R4462 VDD.n11902 VDD.n11901 92.5005
R4463 VDD.n11903 VDD.n11902 92.5005
R4464 VDD.n7476 VDD.n7475 92.5005
R4465 VDD.n7475 VDD.n7474 92.5005
R4466 VDD.n11895 VDD.n11894 92.5005
R4467 VDD.n11894 VDD.n11893 92.5005
R4468 VDD.n7483 VDD.n7479 92.5005
R4469 VDD.n11892 VDD.n7479 92.5005
R4470 VDD.n11890 VDD.n11889 92.5005
R4471 VDD.n11891 VDD.n11890 92.5005
R4472 VDD.n11883 VDD.n7481 92.5005
R4473 VDD.n7481 VDD.n7480 92.5005
R4474 VDD.n11882 VDD.n11881 92.5005
R4475 VDD.n11881 VDD.n11880 92.5005
R4476 VDD.n7490 VDD.n7486 92.5005
R4477 VDD.n11879 VDD.n7486 92.5005
R4478 VDD.n11877 VDD.n11876 92.5005
R4479 VDD.n11878 VDD.n11877 92.5005
R4480 VDD.n11870 VDD.n7488 92.5005
R4481 VDD.n7488 VDD.n7487 92.5005
R4482 VDD.n11869 VDD.n11868 92.5005
R4483 VDD.n11868 VDD.n11867 92.5005
R4484 VDD.n7497 VDD.n7493 92.5005
R4485 VDD.n11866 VDD.n7493 92.5005
R4486 VDD.n11864 VDD.n11863 92.5005
R4487 VDD.n11865 VDD.n11864 92.5005
R4488 VDD.n11857 VDD.n7495 92.5005
R4489 VDD.n7495 VDD.n7494 92.5005
R4490 VDD.n11856 VDD.n11855 92.5005
R4491 VDD.n11855 VDD.n11854 92.5005
R4492 VDD.n11849 VDD.n7500 92.5005
R4493 VDD.n11853 VDD.n7500 92.5005
R4494 VDD.n11851 VDD.n11850 92.5005
R4495 VDD.n11852 VDD.n11851 92.5005
R4496 VDD.n7503 VDD.n7502 92.5005
R4497 VDD.n7502 VDD.n7501 92.5005
R4498 VDD.n11844 VDD.n11843 92.5005
R4499 VDD.n11843 VDD.n11842 92.5005
R4500 VDD.n7510 VDD.n7506 92.5005
R4501 VDD.n11841 VDD.n7506 92.5005
R4502 VDD.n11839 VDD.n11838 92.5005
R4503 VDD.n11840 VDD.n11839 92.5005
R4504 VDD.n11832 VDD.n7508 92.5005
R4505 VDD.n7508 VDD.n7507 92.5005
R4506 VDD.n11831 VDD.n11830 92.5005
R4507 VDD.n11830 VDD.n11829 92.5005
R4508 VDD.n7517 VDD.n7513 92.5005
R4509 VDD.n11828 VDD.n7513 92.5005
R4510 VDD.n11826 VDD.n11825 92.5005
R4511 VDD.n11827 VDD.n11826 92.5005
R4512 VDD.n11819 VDD.n7515 92.5005
R4513 VDD.n7515 VDD.n7514 92.5005
R4514 VDD.n11818 VDD.n11817 92.5005
R4515 VDD.n11817 VDD.n11816 92.5005
R4516 VDD.n7524 VDD.n7520 92.5005
R4517 VDD.n11815 VDD.n7520 92.5005
R4518 VDD.n11813 VDD.n11812 92.5005
R4519 VDD.n11814 VDD.n11813 92.5005
R4520 VDD.n11806 VDD.n7522 92.5005
R4521 VDD.n7522 VDD.n7521 92.5005
R4522 VDD.n11805 VDD.n11804 92.5005
R4523 VDD.n11804 VDD.n11803 92.5005
R4524 VDD.n7531 VDD.n7527 92.5005
R4525 VDD.n11802 VDD.n7527 92.5005
R4526 VDD.n11800 VDD.n11799 92.5005
R4527 VDD.n11801 VDD.n11800 92.5005
R4528 VDD.n7534 VDD.n7529 92.5005
R4529 VDD.n7529 VDD.n7528 92.5005
R4530 VDD.n11793 VDD.n11792 92.5005
R4531 VDD.n11792 VDD.n11791 92.5005
R4532 VDD.n7535 VDD.n7533 92.5005
R4533 VDD.n11790 VDD.n7535 92.5005
R4534 VDD.n11788 VDD.n11787 92.5005
R4535 VDD.n11789 VDD.n11788 92.5005
R4536 VDD.n7538 VDD.n7537 92.5005
R4537 VDD.n7537 VDD.n7536 92.5005
R4538 VDD.n11781 VDD.n11780 92.5005
R4539 VDD.n11780 VDD.n11779 92.5005
R4540 VDD.n7545 VDD.n7541 92.5005
R4541 VDD.n11778 VDD.n7541 92.5005
R4542 VDD.n11776 VDD.n11775 92.5005
R4543 VDD.n11777 VDD.n11776 92.5005
R4544 VDD.n11769 VDD.n7543 92.5005
R4545 VDD.n7543 VDD.n7542 92.5005
R4546 VDD.n11768 VDD.n11767 92.5005
R4547 VDD.n11767 VDD.n11766 92.5005
R4548 VDD.n7552 VDD.n7548 92.5005
R4549 VDD.n11765 VDD.n7548 92.5005
R4550 VDD.n11763 VDD.n11762 92.5005
R4551 VDD.n11764 VDD.n11763 92.5005
R4552 VDD.n11756 VDD.n7550 92.5005
R4553 VDD.n7550 VDD.n7549 92.5005
R4554 VDD.n11755 VDD.n11754 92.5005
R4555 VDD.n11754 VDD.n11753 92.5005
R4556 VDD.n7559 VDD.n7555 92.5005
R4557 VDD.n11752 VDD.n7555 92.5005
R4558 VDD.n11750 VDD.n11749 92.5005
R4559 VDD.n11751 VDD.n11750 92.5005
R4560 VDD.n11743 VDD.n7557 92.5005
R4561 VDD.n7557 VDD.n7556 92.5005
R4562 VDD.n11742 VDD.n11741 92.5005
R4563 VDD.n11741 VDD.n11740 92.5005
R4564 VDD.n11735 VDD.n7562 92.5005
R4565 VDD.n11739 VDD.n7562 92.5005
R4566 VDD.n11737 VDD.n11736 92.5005
R4567 VDD.n11738 VDD.n11737 92.5005
R4568 VDD.n7565 VDD.n7564 92.5005
R4569 VDD.n7564 VDD.n7563 92.5005
R4570 VDD.n11730 VDD.n11729 92.5005
R4571 VDD.n11729 VDD.n11728 92.5005
R4572 VDD.n7572 VDD.n7568 92.5005
R4573 VDD.n11727 VDD.n7568 92.5005
R4574 VDD.n11725 VDD.n11724 92.5005
R4575 VDD.n11726 VDD.n11725 92.5005
R4576 VDD.n11718 VDD.n7570 92.5005
R4577 VDD.n7570 VDD.n7569 92.5005
R4578 VDD.n11717 VDD.n11716 92.5005
R4579 VDD.n11716 VDD.n11715 92.5005
R4580 VDD.n7579 VDD.n7575 92.5005
R4581 VDD.n11714 VDD.n7575 92.5005
R4582 VDD.n11712 VDD.n11711 92.5005
R4583 VDD.n11713 VDD.n11712 92.5005
R4584 VDD.n11705 VDD.n7577 92.5005
R4585 VDD.n7577 VDD.n7576 92.5005
R4586 VDD.n11704 VDD.n11703 92.5005
R4587 VDD.n11703 VDD.n11702 92.5005
R4588 VDD.n7586 VDD.n7582 92.5005
R4589 VDD.n11701 VDD.n7582 92.5005
R4590 VDD.n11699 VDD.n11698 92.5005
R4591 VDD.n11700 VDD.n11699 92.5005
R4592 VDD.n11692 VDD.n7584 92.5005
R4593 VDD.n7584 VDD.n7583 92.5005
R4594 VDD.n11691 VDD.n11690 92.5005
R4595 VDD.n11690 VDD.n11689 92.5005
R4596 VDD.n7593 VDD.n7589 92.5005
R4597 VDD.n11688 VDD.n7589 92.5005
R4598 VDD.n11686 VDD.n11685 92.5005
R4599 VDD.n11687 VDD.n11686 92.5005
R4600 VDD.n7596 VDD.n7591 92.5005
R4601 VDD.n7591 VDD.n7590 92.5005
R4602 VDD.n11679 VDD.n11678 92.5005
R4603 VDD.n11678 VDD.n11677 92.5005
R4604 VDD.n7597 VDD.n7595 92.5005
R4605 VDD.n11676 VDD.n7597 92.5005
R4606 VDD.n11674 VDD.n11673 92.5005
R4607 VDD.n11675 VDD.n11674 92.5005
R4608 VDD.n7600 VDD.n7599 92.5005
R4609 VDD.n7599 VDD.n7598 92.5005
R4610 VDD.n11667 VDD.n11666 92.5005
R4611 VDD.n11666 VDD.n11665 92.5005
R4612 VDD.n7607 VDD.n7603 92.5005
R4613 VDD.n11664 VDD.n7603 92.5005
R4614 VDD.n11662 VDD.n11661 92.5005
R4615 VDD.n11663 VDD.n11662 92.5005
R4616 VDD.n11655 VDD.n7605 92.5005
R4617 VDD.n7605 VDD.n7604 92.5005
R4618 VDD.n11654 VDD.n11653 92.5005
R4619 VDD.n11653 VDD.n11652 92.5005
R4620 VDD.n11642 VDD.n7613 92.5005
R4621 VDD.n11642 VDD.n11641 92.5005
R4622 VDD.n7618 VDD.n7614 92.5005
R4623 VDD.n11640 VDD.n7614 92.5005
R4624 VDD.n11638 VDD.n11637 92.5005
R4625 VDD.n11639 VDD.n11638 92.5005
R4626 VDD.n11629 VDD.n7616 92.5005
R4627 VDD.n7616 VDD.n7615 92.5005
R4628 VDD.n11628 VDD.n11627 92.5005
R4629 VDD.n11627 VDD.n11626 92.5005
R4630 VDD.n7625 VDD.n7621 92.5005
R4631 VDD.n11625 VDD.n7621 92.5005
R4632 VDD.n11623 VDD.n11622 92.5005
R4633 VDD.n11624 VDD.n11623 92.5005
R4634 VDD.n11616 VDD.n7623 92.5005
R4635 VDD.n7623 VDD.n7622 92.5005
R4636 VDD.n7642 VDD.n7641 92.5005
R4637 VDD.n11586 VDD.n7642 92.5005
R4638 VDD.n11584 VDD.n11583 92.5005
R4639 VDD.n11585 VDD.n11584 92.5005
R4640 VDD.n7645 VDD.n7644 92.5005
R4641 VDD.n7644 VDD.n7643 92.5005
R4642 VDD.n11577 VDD.n11576 92.5005
R4643 VDD.n11576 VDD.n11575 92.5005
R4644 VDD.n7652 VDD.n7648 92.5005
R4645 VDD.n11574 VDD.n7648 92.5005
R4646 VDD.n11572 VDD.n11571 92.5005
R4647 VDD.n11573 VDD.n11572 92.5005
R4648 VDD.n11565 VDD.n7650 92.5005
R4649 VDD.n7650 VDD.n7649 92.5005
R4650 VDD.n11564 VDD.n11563 92.5005
R4651 VDD.n11563 VDD.n11562 92.5005
R4652 VDD.n7659 VDD.n7655 92.5005
R4653 VDD.n11561 VDD.n7655 92.5005
R4654 VDD.n11533 VDD.n11532 92.5005
R4655 VDD.n11534 VDD.n11533 92.5005
R4656 VDD.n7672 VDD.n7671 92.5005
R4657 VDD.n7671 VDD.n7670 92.5005
R4658 VDD.n11528 VDD.n11527 92.5005
R4659 VDD.n11527 VDD.n11526 92.5005
R4660 VDD.n7680 VDD.n7676 92.5005
R4661 VDD.n11525 VDD.n7676 92.5005
R4662 VDD.n11523 VDD.n11522 92.5005
R4663 VDD.n11524 VDD.n11523 92.5005
R4664 VDD.n11516 VDD.n7678 92.5005
R4665 VDD.n7678 VDD.n7677 92.5005
R4666 VDD.n11515 VDD.n11514 92.5005
R4667 VDD.n11514 VDD.n11513 92.5005
R4668 VDD.n7687 VDD.n7683 92.5005
R4669 VDD.n11512 VDD.n7683 92.5005
R4670 VDD.n11510 VDD.n11509 92.5005
R4671 VDD.n11511 VDD.n11510 92.5005
R4672 VDD.n11503 VDD.n7685 92.5005
R4673 VDD.n7685 VDD.n7684 92.5005
R4674 VDD.n11478 VDD.n11476 92.5005
R4675 VDD.n11476 VDD.n11475 92.5005
R4676 VDD.n7704 VDD.n7703 92.5005
R4677 VDD.n11474 VDD.n7704 92.5005
R4678 VDD.n11472 VDD.n11471 92.5005
R4679 VDD.n11473 VDD.n11472 92.5005
R4680 VDD.n7707 VDD.n7706 92.5005
R4681 VDD.n7706 VDD.n7705 92.5005
R4682 VDD.n11465 VDD.n11464 92.5005
R4683 VDD.n11464 VDD.n11463 92.5005
R4684 VDD.n7714 VDD.n7710 92.5005
R4685 VDD.n11462 VDD.n7710 92.5005
R4686 VDD.n11460 VDD.n11459 92.5005
R4687 VDD.n11461 VDD.n11460 92.5005
R4688 VDD.n11453 VDD.n7712 92.5005
R4689 VDD.n7712 VDD.n7711 92.5005
R4690 VDD.n11452 VDD.n11451 92.5005
R4691 VDD.n11451 VDD.n11450 92.5005
R4692 VDD.n7879 VDD.n7717 92.5005
R4693 VDD.n11449 VDD.n7717 92.5005
R4694 VDD.n7903 VDD.n7866 92.5005
R4695 VDD.n7864 VDD.n7862 92.5005
R4696 VDD.n7908 VDD.n7907 92.5005
R4697 VDD.n7911 VDD.n7910 92.5005
R4698 VDD.n7859 VDD.n7856 92.5005
R4699 VDD.n7917 VDD.n7916 92.5005
R4700 VDD.n7920 VDD.n7919 92.5005
R4701 VDD.n7853 VDD.n7850 92.5005
R4702 VDD.n7926 VDD.n7925 92.5005
R4703 VDD.n7929 VDD.n7928 92.5005
R4704 VDD.n7952 VDD.n7831 92.5005
R4705 VDD.n7954 VDD.n7953 92.5005
R4706 VDD.n7957 VDD.n7956 92.5005
R4707 VDD.n7828 VDD.n7825 92.5005
R4708 VDD.n7963 VDD.n7962 92.5005
R4709 VDD.n7966 VDD.n7965 92.5005
R4710 VDD.n7822 VDD.n7819 92.5005
R4711 VDD.n7972 VDD.n7971 92.5005
R4712 VDD.n7975 VDD.n7974 92.5005
R4713 VDD.n7816 VDD.n7812 92.5005
R4714 VDD.n7980 VDD.n7809 92.5005
R4715 VDD.n7835 VDD.n7832 92.5005
R4716 VDD.n7835 VDD.n7749 92.5005
R4717 VDD.n7948 VDD.n7947 92.5005
R4718 VDD.n7945 VDD.n7944 92.5005
R4719 VDD.n7837 VDD.n7836 92.5005
R4720 VDD.n7939 VDD.n7938 92.5005
R4721 VDD.n7937 VDD.n7841 92.5005
R4722 VDD.n7935 VDD.n7934 92.5005
R4723 VDD.n7844 VDD.n7842 92.5005
R4724 VDD.n7902 VDD.n7901 92.5005
R4725 VDD.n7899 VDD.n7898 92.5005
R4726 VDD.n7869 VDD.n7868 92.5005
R4727 VDD.n7893 VDD.n7892 92.5005
R4728 VDD.n7891 VDD.n7873 92.5005
R4729 VDD.n7889 VDD.n7888 92.5005
R4730 VDD.n7876 VDD.n7874 92.5005
R4731 VDD.n7883 VDD.n7882 92.5005
R4732 VDD.n11477 VDD.n7699 92.5005
R4733 VDD.n7699 VDD.n7698 92.5005
R4734 VDD.n11484 VDD.n11483 92.5005
R4735 VDD.n11485 VDD.n11484 92.5005
R4736 VDD.n7701 VDD.n7697 92.5005
R4737 VDD.n11486 VDD.n7697 92.5005
R4738 VDD.n11489 VDD.n11488 92.5005
R4739 VDD.n11488 VDD.n11487 92.5005
R4740 VDD.n11490 VDD.n7692 92.5005
R4741 VDD.n7692 VDD.n7691 92.5005
R4742 VDD.n11497 VDD.n11496 92.5005
R4743 VDD.n11498 VDD.n11497 92.5005
R4744 VDD.n7694 VDD.n7690 92.5005
R4745 VDD.n11499 VDD.n7690 92.5005
R4746 VDD.n11502 VDD.n11501 92.5005
R4747 VDD.n11501 VDD.n11500 92.5005
R4748 VDD.n7673 VDD.n7669 92.5005
R4749 VDD.n11535 VDD.n7669 92.5005
R4750 VDD.n11538 VDD.n11537 92.5005
R4751 VDD.n11537 VDD.n11536 92.5005
R4752 VDD.n11539 VDD.n7664 92.5005
R4753 VDD.n7664 VDD.n7663 92.5005
R4754 VDD.n11546 VDD.n11545 92.5005
R4755 VDD.n11547 VDD.n11546 92.5005
R4756 VDD.n7666 VDD.n7662 92.5005
R4757 VDD.n11548 VDD.n7662 92.5005
R4758 VDD.n11551 VDD.n11550 92.5005
R4759 VDD.n11550 VDD.n11549 92.5005
R4760 VDD.n11552 VDD.n7657 92.5005
R4761 VDD.n7657 VDD.n7656 92.5005
R4762 VDD.n11559 VDD.n11558 92.5005
R4763 VDD.n11560 VDD.n11559 92.5005
R4764 VDD.n11589 VDD.n11588 92.5005
R4765 VDD.n11588 VDD.n11587 92.5005
R4766 VDD.n11590 VDD.n7637 92.5005
R4767 VDD.n7637 VDD.n7636 92.5005
R4768 VDD.n11597 VDD.n11596 92.5005
R4769 VDD.n11598 VDD.n11597 92.5005
R4770 VDD.n7639 VDD.n7635 92.5005
R4771 VDD.n11599 VDD.n7635 92.5005
R4772 VDD.n11602 VDD.n11601 92.5005
R4773 VDD.n11601 VDD.n11600 92.5005
R4774 VDD.n11603 VDD.n7630 92.5005
R4775 VDD.n7630 VDD.n7629 92.5005
R4776 VDD.n11610 VDD.n11609 92.5005
R4777 VDD.n11611 VDD.n11610 92.5005
R4778 VDD.n7632 VDD.n7628 92.5005
R4779 VDD.n11612 VDD.n7628 92.5005
R4780 VDD.n11615 VDD.n11614 92.5005
R4781 VDD.n11614 VDD.n11613 92.5005
R4782 VDD.n11645 VDD.n11644 92.5005
R4783 VDD.n11651 VDD.n7610 92.5005
R4784 VDD.n11650 VDD.n11649 92.5005
R4785 VDD.n11647 VDD.n7612 92.5005
R4786 VDD.n7783 VDD.n7782 92.5005
R4787 VDD.n8544 VDD.n8543 92.5005
R4788 VDD.n8539 VDD.n8538 92.5005
R4789 VDD.n8536 VDD.n7784 92.5005
R4790 VDD.n8535 VDD.n8534 92.5005
R4791 VDD.n7792 VDD.n7788 92.5005
R4792 VDD.n8529 VDD.n8528 92.5005
R4793 VDD.n8526 VDD.n8525 92.5005
R4794 VDD.n7794 VDD.n7793 92.5005
R4795 VDD.n8520 VDD.n8519 92.5005
R4796 VDD.n8518 VDD.n7796 92.5005
R4797 VDD.n8516 VDD.n8515 92.5005
R4798 VDD.n7800 VDD.n7798 92.5005
R4799 VDD.n8510 VDD.n8509 92.5005
R4800 VDD.n8508 VDD.n8507 92.5005
R4801 VDD.n7808 VDD.n7805 92.5005
R4802 VDD.n8502 VDD.n8501 92.5005
R4803 VDD.n8501 VDD.n7785 92.5005
R4804 VDD.n8500 VDD.n7987 92.5005
R4805 VDD.n8500 VDD.n8499 92.5005
R4806 VDD.n8540 VDD.n7781 92.5005
R4807 VDD.n8545 VDD.n7781 92.5005
R4808 VDD.n7775 VDD.n7771 92.5005
R4809 VDD.n8556 VDD.n7771 92.5005
R4810 VDD.n8558 VDD.n7772 92.5005
R4811 VDD.n8558 VDD.n8557 92.5005
R4812 VDD.n8554 VDD.n8553 92.5005
R4813 VDD.n8555 VDD.n8554 92.5005
R4814 VDD.n7776 VDD.n7774 92.5005
R4815 VDD.n7774 VDD.n7773 92.5005
R4816 VDD.n8548 VDD.n8547 92.5005
R4817 VDD.n8547 VDD.n8546 92.5005
R4818 VDD.n8560 VDD.n8559 92.5005
R4819 VDD.n8559 VDD.n7755 92.5005
R4820 VDD.n8566 VDD.n8565 92.5005
R4821 VDD.n8567 VDD.n8566 92.5005
R4822 VDD.n8421 VDD.n8408 92.5005
R4823 VDD.n8413 VDD.n8408 92.5005
R4824 VDD.n8427 VDD.n8402 92.5005
R4825 VDD.n8428 VDD.n8427 92.5005
R4826 VDD.n8442 VDD.n8385 92.5005
R4827 VDD.n8443 VDD.n8442 92.5005
R4828 VDD.n8451 VDD.n8374 92.5005
R4829 VDD.n8378 VDD.n8374 92.5005
R4830 VDD.n8457 VDD.n8368 92.5005
R4831 VDD.n8458 VDD.n8457 92.5005
R4832 VDD.n8364 VDD.n8358 92.5005
R4833 VDD.n8362 VDD.n8358 92.5005
R4834 VDD.n8471 VDD.n8352 92.5005
R4835 VDD.n8472 VDD.n8471 92.5005
R4836 VDD.n8480 VDD.n8341 92.5005
R4837 VDD.n8345 VDD.n8341 92.5005
R4838 VDD.n8486 VDD.n7997 92.5005
R4839 VDD.n8487 VDD.n8486 92.5005
R4840 VDD.n8496 VDD.n8495 92.5005
R4841 VDD.n8497 VDD.n8496 92.5005
R4842 VDD.n8319 VDD.n8318 92.5005
R4843 VDD.n8320 VDD.n8319 92.5005
R4844 VDD.n8307 VDD.n8012 92.5005
R4845 VDD.n8308 VDD.n8307 92.5005
R4846 VDD.n8021 VDD.n8015 92.5005
R4847 VDD.n8019 VDD.n8015 92.5005
R4848 VDD.n8027 VDD.n8024 92.5005
R4849 VDD.n8025 VDD.n8024 92.5005
R4850 VDD.n8035 VDD.n8031 92.5005
R4851 VDD.n8278 VDD.n8031 92.5005
R4852 VDD.n8275 VDD.n8041 92.5005
R4853 VDD.n8275 VDD.n8274 92.5005
R4854 VDD.n8265 VDD.n8264 92.5005
R4855 VDD.n8264 VDD.n8263 92.5005
R4856 VDD.n8256 VDD.n8255 92.5005
R4857 VDD.n8257 VDD.n8256 92.5005
R4858 VDD.n8232 VDD.n8063 92.5005
R4859 VDD.n8233 VDD.n8232 92.5005
R4860 VDD.n8072 VDD.n8066 92.5005
R4861 VDD.n8070 VDD.n8066 92.5005
R4862 VDD.n8079 VDD.n8075 92.5005
R4863 VDD.n8076 VDD.n8075 92.5005
R4864 VDD.n8206 VDD.n8082 92.5005
R4865 VDD.n8202 VDD.n8082 92.5005
R4866 VDD.n8199 VDD.n8091 92.5005
R4867 VDD.n8199 VDD.n8198 92.5005
R4868 VDD.n8119 VDD.n8088 92.5005
R4869 VDD.n8092 VDD.n8088 92.5005
R4870 VDD.n8125 VDD.n8112 92.5005
R4871 VDD.n8122 VDD.n8121 92.5005
R4872 VDD.n8121 VDD.n8114 92.5005
R4873 VDD.n8200 VDD.n8085 92.5005
R4874 VDD.n8201 VDD.n8200 92.5005
R4875 VDD.n8090 VDD.n8086 92.5005
R4876 VDD.n8087 VDD.n8086 92.5005
R4877 VDD.n8205 VDD.n8204 92.5005
R4878 VDD.n8204 VDD.n8203 92.5005
R4879 VDD.n8212 VDD.n8211 92.5005
R4880 VDD.n8213 VDD.n8212 92.5005
R4881 VDD.n8083 VDD.n8077 92.5005
R4882 VDD.n8081 VDD.n8077 92.5005
R4883 VDD.n8215 VDD.n8080 92.5005
R4884 VDD.n8215 VDD.n8214 92.5005
R4885 VDD.n8221 VDD.n8220 92.5005
R4886 VDD.n8220 VDD.n8219 92.5005
R4887 VDD.n8216 VDD.n8074 92.5005
R4888 VDD.n8217 VDD.n8216 92.5005
R4889 VDD.n8222 VDD.n8071 92.5005
R4890 VDD.n8218 VDD.n8071 92.5005
R4891 VDD.n8231 VDD.n8069 92.5005
R4892 VDD.n8231 VDD.n8230 92.5005
R4893 VDD.n8228 VDD.n8227 92.5005
R4894 VDD.n8229 VDD.n8228 92.5005
R4895 VDD.n8067 VDD.n8064 92.5005
R4896 VDD.n8065 VDD.n8064 92.5005
R4897 VDD.n8061 VDD.n8060 92.5005
R4898 VDD.n8234 VDD.n8060 92.5005
R4899 VDD.n8237 VDD.n8236 92.5005
R4900 VDD.n8236 VDD.n8235 92.5005
R4901 VDD.n8242 VDD.n8058 92.5005
R4902 VDD.n8059 VDD.n8058 92.5005
R4903 VDD.n8244 VDD.n8243 92.5005
R4904 VDD.n8245 VDD.n8244 92.5005
R4905 VDD.n8250 VDD.n8054 92.5005
R4906 VDD.n8246 VDD.n8054 92.5005
R4907 VDD.n8249 VDD.n8248 92.5005
R4908 VDD.n8248 VDD.n8247 92.5005
R4909 VDD.n8055 VDD.n8049 92.5005
R4910 VDD.n8053 VDD.n8049 92.5005
R4911 VDD.n8051 VDD.n8047 92.5005
R4912 VDD.n8048 VDD.n8047 92.5005
R4913 VDD.n8259 VDD.n8052 92.5005
R4914 VDD.n8259 VDD.n8258 92.5005
R4915 VDD.n8260 VDD.n8046 92.5005
R4916 VDD.n8261 VDD.n8260 92.5005
R4917 VDD.n8044 VDD.n8038 92.5005
R4918 VDD.n8042 VDD.n8038 92.5005
R4919 VDD.n8266 VDD.n8043 92.5005
R4920 VDD.n8262 VDD.n8043 92.5005
R4921 VDD.n8272 VDD.n8271 92.5005
R4922 VDD.n8273 VDD.n8272 92.5005
R4923 VDD.n8276 VDD.n8034 92.5005
R4924 VDD.n8277 VDD.n8276 92.5005
R4925 VDD.n8039 VDD.n8036 92.5005
R4926 VDD.n8037 VDD.n8036 92.5005
R4927 VDD.n8281 VDD.n8280 92.5005
R4928 VDD.n8280 VDD.n8279 92.5005
R4929 VDD.n8287 VDD.n8286 92.5005
R4930 VDD.n8288 VDD.n8287 92.5005
R4931 VDD.n8032 VDD.n8026 92.5005
R4932 VDD.n8030 VDD.n8026 92.5005
R4933 VDD.n8290 VDD.n8029 92.5005
R4934 VDD.n8290 VDD.n8289 92.5005
R4935 VDD.n8296 VDD.n8295 92.5005
R4936 VDD.n8295 VDD.n8294 92.5005
R4937 VDD.n8291 VDD.n8023 92.5005
R4938 VDD.n8292 VDD.n8291 92.5005
R4939 VDD.n8297 VDD.n8020 92.5005
R4940 VDD.n8293 VDD.n8020 92.5005
R4941 VDD.n8306 VDD.n8018 92.5005
R4942 VDD.n8306 VDD.n8305 92.5005
R4943 VDD.n8303 VDD.n8302 92.5005
R4944 VDD.n8304 VDD.n8303 92.5005
R4945 VDD.n8016 VDD.n8013 92.5005
R4946 VDD.n8014 VDD.n8013 92.5005
R4947 VDD.n8010 VDD.n8009 92.5005
R4948 VDD.n8309 VDD.n8009 92.5005
R4949 VDD.n8312 VDD.n8311 92.5005
R4950 VDD.n8311 VDD.n8310 92.5005
R4951 VDD.n8317 VDD.n8007 92.5005
R4952 VDD.n8008 VDD.n8007 92.5005
R4953 VDD.n8325 VDD.n8003 92.5005
R4954 VDD.n8321 VDD.n8003 92.5005
R4955 VDD.n8324 VDD.n8323 92.5005
R4956 VDD.n8323 VDD.n8322 92.5005
R4957 VDD.n8004 VDD.n7998 92.5005
R4958 VDD.n8002 VDD.n7998 92.5005
R4959 VDD.n8331 VDD.n8330 92.5005
R4960 VDD.n8332 VDD.n8331 92.5005
R4961 VDD.n8000 VDD.n7990 92.5005
R4962 VDD.n8333 VDD.n7990 92.5005
R4963 VDD.n8335 VDD.n8001 92.5005
R4964 VDD.n8335 VDD.n8334 92.5005
R4965 VDD.n8336 VDD.n7992 92.5005
R4966 VDD.n8336 VDD.n7988 92.5005
R4967 VDD.n7996 VDD.n7991 92.5005
R4968 VDD.n8339 VDD.n7991 92.5005
R4969 VDD.n8337 VDD.n7993 92.5005
R4970 VDD.n8337 VDD.n7989 92.5005
R4971 VDD.n8490 VDD.n8489 92.5005
R4972 VDD.n8489 VDD.n8488 92.5005
R4973 VDD.n8485 VDD.n8344 92.5005
R4974 VDD.n8485 VDD.n8484 92.5005
R4975 VDD.n8343 VDD.n8338 92.5005
R4976 VDD.n8340 VDD.n8338 92.5005
R4977 VDD.n8482 VDD.n8481 92.5005
R4978 VDD.n8483 VDD.n8482 92.5005
R4979 VDD.n8357 VDD.n8351 92.5005
R4980 VDD.n8357 VDD.n8355 92.5005
R4981 VDD.n8348 VDD.n8346 92.5005
R4982 VDD.n8354 VDD.n8346 92.5005
R4983 VDD.n8475 VDD.n8474 92.5005
R4984 VDD.n8474 VDD.n8473 92.5005
R4985 VDD.n8470 VDD.n8361 92.5005
R4986 VDD.n8470 VDD.n8469 92.5005
R4987 VDD.n8359 VDD.n8353 92.5005
R4988 VDD.n8356 VDD.n8353 92.5005
R4989 VDD.n8467 VDD.n8466 92.5005
R4990 VDD.n8468 VDD.n8467 92.5005
R4991 VDD.n8373 VDD.n8367 92.5005
R4992 VDD.n8373 VDD.n8371 92.5005
R4993 VDD.n8366 VDD.n8363 92.5005
R4994 VDD.n8370 VDD.n8363 92.5005
R4995 VDD.n8461 VDD.n8460 92.5005
R4996 VDD.n8460 VDD.n8459 92.5005
R4997 VDD.n8456 VDD.n8377 92.5005
R4998 VDD.n8456 VDD.n8455 92.5005
R4999 VDD.n8376 VDD.n8369 92.5005
R5000 VDD.n8372 VDD.n8369 92.5005
R5001 VDD.n8453 VDD.n8452 92.5005
R5002 VDD.n8454 VDD.n8453 92.5005
R5003 VDD.n8390 VDD.n8384 92.5005
R5004 VDD.n8390 VDD.n8388 92.5005
R5005 VDD.n8381 VDD.n8379 92.5005
R5006 VDD.n8387 VDD.n8379 92.5005
R5007 VDD.n8446 VDD.n8445 92.5005
R5008 VDD.n8445 VDD.n8444 92.5005
R5009 VDD.n8441 VDD.n8394 92.5005
R5010 VDD.n8441 VDD.n8440 92.5005
R5011 VDD.n8393 VDD.n8386 92.5005
R5012 VDD.n8389 VDD.n8386 92.5005
R5013 VDD.n8438 VDD.n8437 92.5005
R5014 VDD.n8439 VDD.n8438 92.5005
R5015 VDD.n8436 VDD.n8391 92.5005
R5016 VDD.n8395 VDD.n8391 92.5005
R5017 VDD.n8407 VDD.n8401 92.5005
R5018 VDD.n8407 VDD.n8405 92.5005
R5019 VDD.n8398 VDD.n8396 92.5005
R5020 VDD.n8404 VDD.n8396 92.5005
R5021 VDD.n8431 VDD.n8430 92.5005
R5022 VDD.n8430 VDD.n8429 92.5005
R5023 VDD.n8426 VDD.n8411 92.5005
R5024 VDD.n8426 VDD.n8425 92.5005
R5025 VDD.n8410 VDD.n8403 92.5005
R5026 VDD.n8406 VDD.n8403 92.5005
R5027 VDD.n8423 VDD.n8422 92.5005
R5028 VDD.n8424 VDD.n8423 92.5005
R5029 VDD.n8416 VDD.n7765 92.5005
R5030 VDD.n7765 VDD.n7764 92.5005
R5031 VDD.n8417 VDD.n7762 92.5005
R5032 VDD.n8412 VDD.n7762 92.5005
R5033 VDD.n8569 VDD.n7763 92.5005
R5034 VDD.n8569 VDD.n8568 92.5005
R5035 VDD.n7767 VDD.n7766 92.5005
R5036 VDD.n7766 VDD.n7754 92.5005
R5037 VDD.n8571 VDD.n8570 92.5005
R5038 VDD.n8573 VDD.n8572 92.5005
R5039 VDD.n8575 VDD.n8574 92.5005
R5040 VDD.n8577 VDD.n8576 92.5005
R5041 VDD.n8579 VDD.n8578 92.5005
R5042 VDD.n8581 VDD.n8580 92.5005
R5043 VDD.n8583 VDD.n8582 92.5005
R5044 VDD.n8585 VDD.n8584 92.5005
R5045 VDD.n8586 VDD.n7760 92.5005
R5046 VDD.n8588 VDD.n8587 92.5005
R5047 VDD.n7753 VDD.n7752 92.5005
R5048 VDD.n8593 VDD.n8592 92.5005
R5049 VDD.n8594 VDD.n7750 92.5005
R5050 VDD.n8499 VDD.n7750 92.5005
R5051 VDD.n8597 VDD.n8596 92.5005
R5052 VDD.n8598 VDD.n8597 92.5005
R5053 VDD.n8595 VDD.n7751 92.5005
R5054 VDD.n7751 VDD.n7718 92.5005
R5055 VDD.n7732 VDD.n7730 92.5005
R5056 VDD.n7730 VDD.n7719 92.5005
R5057 VDD.n11440 VDD.n11439 92.5005
R5058 VDD.n11441 VDD.n11440 92.5005
R5059 VDD.n11438 VDD.n7731 92.5005
R5060 VDD.n9172 VDD.n7731 92.5005
R5061 VDD.n11437 VDD.n11436 92.5005
R5062 VDD.n11436 VDD.n11435 92.5005
R5063 VDD.n7734 VDD.n7733 92.5005
R5064 VDD.n8616 VDD.n7734 92.5005
R5065 VDD.n8625 VDD.n8618 92.5005
R5066 VDD.n11425 VDD.n8618 92.5005
R5067 VDD.n11421 VDD.n11420 92.5005
R5068 VDD.n11422 VDD.n11421 92.5005
R5069 VDD.n11419 VDD.n8624 92.5005
R5070 VDD.n8628 VDD.n8624 92.5005
R5071 VDD.n11418 VDD.n11417 92.5005
R5072 VDD.n11417 VDD.n11416 92.5005
R5073 VDD.n8627 VDD.n8626 92.5005
R5074 VDD.n8647 VDD.n8627 92.5005
R5075 VDD.n8656 VDD.n8649 92.5005
R5076 VDD.n11406 VDD.n8649 92.5005
R5077 VDD.n11402 VDD.n11401 92.5005
R5078 VDD.n11403 VDD.n11402 92.5005
R5079 VDD.n11400 VDD.n8655 92.5005
R5080 VDD.n9176 VDD.n8655 92.5005
R5081 VDD.n11399 VDD.n11398 92.5005
R5082 VDD.n11398 VDD.n11397 92.5005
R5083 VDD.n8658 VDD.n8657 92.5005
R5084 VDD.n8668 VDD.n8658 92.5005
R5085 VDD.n8694 VDD.n8670 92.5005
R5086 VDD.n11390 VDD.n8670 92.5005
R5087 VDD.n8696 VDD.n8695 92.5005
R5088 VDD.n8695 VDD.n8685 92.5005
R5089 VDD.n8697 VDD.n8687 92.5005
R5090 VDD.n11381 VDD.n8687 92.5005
R5091 VDD.n11377 VDD.n11376 92.5005
R5092 VDD.n11378 VDD.n11377 92.5005
R5093 VDD.n11375 VDD.n8693 92.5005
R5094 VDD.n8700 VDD.n8693 92.5005
R5095 VDD.n11374 VDD.n11373 92.5005
R5096 VDD.n11373 VDD.n11372 92.5005
R5097 VDD.n8699 VDD.n8698 92.5005
R5098 VDD.n8719 VDD.n8699 92.5005
R5099 VDD.n11030 VDD.n8722 92.5005
R5100 VDD.n11362 VDD.n8722 92.5005
R5101 VDD.n11358 VDD.n11357 92.5005
R5102 VDD.n11359 VDD.n11358 92.5005
R5103 VDD.n11356 VDD.n11029 92.5005
R5104 VDD.n11033 VDD.n11029 92.5005
R5105 VDD.n11355 VDD.n11354 92.5005
R5106 VDD.n11354 VDD.n11353 92.5005
R5107 VDD.n11032 VDD.n11031 92.5005
R5108 VDD.n11052 VDD.n11032 92.5005
R5109 VDD.n11060 VDD.n11054 92.5005
R5110 VDD.n11343 VDD.n11054 92.5005
R5111 VDD.n11339 VDD.n11338 92.5005
R5112 VDD.n11340 VDD.n11339 92.5005
R5113 VDD.n11337 VDD.n11059 92.5005
R5114 VDD.n11095 VDD.n11059 92.5005
R5115 VDD.n11336 VDD.n11335 92.5005
R5116 VDD.n11335 VDD.n11334 92.5005
R5117 VDD.n11062 VDD.n11061 92.5005
R5118 VDD.n11074 VDD.n11062 92.5005
R5119 VDD.n11324 VDD.n11323 92.5005
R5120 VDD.n11325 VDD.n11324 92.5005
R5121 VDD.n11322 VDD.n11077 92.5005
R5122 VDD.n11080 VDD.n11077 92.5005
R5123 VDD.n11321 VDD.n11320 92.5005
R5124 VDD.n11320 VDD.n11319 92.5005
R5125 VDD.n11079 VDD.n11078 92.5005
R5126 VDD.n11105 VDD.n11079 92.5005
R5127 VDD.n11114 VDD.n11107 92.5005
R5128 VDD.n11309 VDD.n11107 92.5005
R5129 VDD.n11305 VDD.n11304 92.5005
R5130 VDD.n11306 VDD.n11305 92.5005
R5131 VDD.n11303 VDD.n11113 92.5005
R5132 VDD.n11117 VDD.n11113 92.5005
R5133 VDD.n11302 VDD.n11301 92.5005
R5134 VDD.n11301 VDD.n11300 92.5005
R5135 VDD.n11116 VDD.n11115 92.5005
R5136 VDD.n11136 VDD.n11116 92.5005
R5137 VDD.n11145 VDD.n11137 92.5005
R5138 VDD.n11290 VDD.n11137 92.5005
R5139 VDD.n11286 VDD.n11285 92.5005
R5140 VDD.n11287 VDD.n11286 92.5005
R5141 VDD.n11284 VDD.n11144 92.5005
R5142 VDD.n11148 VDD.n11144 92.5005
R5143 VDD.n11283 VDD.n11282 92.5005
R5144 VDD.n11282 VDD.n11281 92.5005
R5145 VDD.n11147 VDD.n11146 92.5005
R5146 VDD.n11167 VDD.n11147 92.5005
R5147 VDD.n11176 VDD.n11169 92.5005
R5148 VDD.n11271 VDD.n11169 92.5005
R5149 VDD.n11267 VDD.n11266 92.5005
R5150 VDD.n11268 VDD.n11267 92.5005
R5151 VDD.n11265 VDD.n11175 92.5005
R5152 VDD.n11179 VDD.n11175 92.5005
R5153 VDD.n11264 VDD.n11263 92.5005
R5154 VDD.n11263 VDD.n11262 92.5005
R5155 VDD.n11178 VDD.n11177 92.5005
R5156 VDD.n11189 VDD.n11178 92.5005
R5157 VDD.n11235 VDD.n11191 92.5005
R5158 VDD.n11255 VDD.n11191 92.5005
R5159 VDD.n11237 VDD.n11236 92.5005
R5160 VDD.n11236 VDD.n11206 92.5005
R5161 VDD.n11238 VDD.n11208 92.5005
R5162 VDD.n11246 VDD.n11208 92.5005
R5163 VDD.n11242 VDD.n11241 92.5005
R5164 VDD.n11243 VDD.n11242 92.5005
R5165 VDD.n11240 VDD.n11234 92.5005
R5166 VDD.n11234 VDD.n11233 92.5005
R5167 VDD.n11239 VDD.n6597 92.5005
R5168 VDD.n11214 VDD.n6597 92.5005
R5169 VDD.n12711 VDD.n6598 92.5005
R5170 VDD.n12711 VDD.n12710 92.5005
R5171 VDD.n12714 VDD.n12713 92.5005
R5172 VDD.n12716 VDD.n12715 92.5005
R5173 VDD.n12718 VDD.n6594 92.5005
R5174 VDD.n12721 VDD.n12720 92.5005
R5175 VDD.n12723 VDD.n12722 92.5005
R5176 VDD.n12725 VDD.n6592 92.5005
R5177 VDD.n12728 VDD.n12727 92.5005
R5178 VDD.n12730 VDD.n12729 92.5005
R5179 VDD.n12732 VDD.n6590 92.5005
R5180 VDD.n12735 VDD.n12734 92.5005
R5181 VDD.n12737 VDD.n12736 92.5005
R5182 VDD.n12739 VDD.n6588 92.5005
R5183 VDD.n12742 VDD.n12741 92.5005
R5184 VDD.n12744 VDD.n12743 92.5005
R5185 VDD.n12746 VDD.n6586 92.5005
R5186 VDD.n12749 VDD.n12748 92.5005
R5187 VDD.n12751 VDD.n12750 92.5005
R5188 VDD.n12753 VDD.n6584 92.5005
R5189 VDD.n12756 VDD.n12755 92.5005
R5190 VDD.n12758 VDD.n12757 92.5005
R5191 VDD.n12760 VDD.n6582 92.5005
R5192 VDD.n12763 VDD.n12762 92.5005
R5193 VDD.n12765 VDD.n12764 92.5005
R5194 VDD.n12767 VDD.n6578 92.5005
R5195 VDD.n12712 VDD.n6596 92.5005
R5196 VDD.n12712 VDD.n6580 92.5005
R5197 VDD.n11219 VDD.n11218 92.5005
R5198 VDD.n11216 VDD.n6622 92.5005
R5199 VDD.n12770 VDD.n12769 92.5005
R5200 VDD.n6669 VDD.n6575 92.5005
R5201 VDD.n6672 VDD.n6671 92.5005
R5202 VDD.n6674 VDD.n6668 92.5005
R5203 VDD.n6677 VDD.n6676 92.5005
R5204 VDD.n6679 VDD.n6678 92.5005
R5205 VDD.n6681 VDD.n6666 92.5005
R5206 VDD.n6684 VDD.n6683 92.5005
R5207 VDD.n6686 VDD.n6685 92.5005
R5208 VDD.n6688 VDD.n6664 92.5005
R5209 VDD.n6691 VDD.n6690 92.5005
R5210 VDD.n6693 VDD.n6692 92.5005
R5211 VDD.n6695 VDD.n6624 92.5005
R5212 VDD.n6698 VDD.n6697 92.5005
R5213 VDD.n6661 VDD.n6623 92.5005
R5214 VDD.n6659 VDD.n6658 92.5005
R5215 VDD.n6657 VDD.n6656 92.5005
R5216 VDD.n6654 VDD.n6626 92.5005
R5217 VDD.n6652 VDD.n6651 92.5005
R5218 VDD.n6650 VDD.n6649 92.5005
R5219 VDD.n6647 VDD.n6628 92.5005
R5220 VDD.n6645 VDD.n6644 92.5005
R5221 VDD.n6643 VDD.n6642 92.5005
R5222 VDD.n6640 VDD.n6630 92.5005
R5223 VDD.n6638 VDD.n6637 92.5005
R5224 VDD.n6636 VDD.n6635 92.5005
R5225 VDD.n6633 VDD.n6602 92.5005
R5226 VDD.n12694 VDD.n6620 92.5005
R5227 VDD.n12697 VDD.n12696 92.5005
R5228 VDD.n12695 VDD.n6612 92.5005
R5229 VDD.n12695 VDD.n12694 92.5005
R5230 VDD.n6705 VDD.n6614 92.5005
R5231 VDD.n12691 VDD.n6614 92.5005
R5232 VDD.n12689 VDD.n12688 92.5005
R5233 VDD.n12690 VDD.n12689 92.5005
R5234 VDD.n6707 VDD.n6703 92.5005
R5235 VDD.n6712 VDD.n6703 92.5005
R5236 VDD.n12683 VDD.n12682 92.5005
R5237 VDD.n12682 VDD.n12681 92.5005
R5238 VDD.n10253 VDD.n6711 92.5005
R5239 VDD.n6713 VDD.n6711 92.5005
R5240 VDD.n10257 VDD.n10256 92.5005
R5241 VDD.n10257 VDD.n6720 92.5005
R5242 VDD.n10259 VDD.n10258 92.5005
R5243 VDD.n10258 VDD.n6721 92.5005
R5244 VDD.n10250 VDD.n10249 92.5005
R5245 VDD.n10249 VDD.n6748 92.5005
R5246 VDD.n10265 VDD.n10264 92.5005
R5247 VDD.n10265 VDD.n6749 92.5005
R5248 VDD.n10267 VDD.n10266 92.5005
R5249 VDD.n10266 VDD.n6754 92.5005
R5250 VDD.n10246 VDD.n10245 92.5005
R5251 VDD.n10245 VDD.n10244 92.5005
R5252 VDD.n10273 VDD.n10272 92.5005
R5253 VDD.n10273 VDD.n6758 92.5005
R5254 VDD.n10275 VDD.n10274 92.5005
R5255 VDD.n10274 VDD.n6759 92.5005
R5256 VDD.n10240 VDD.n10239 92.5005
R5257 VDD.n10239 VDD.n6764 92.5005
R5258 VDD.n10282 VDD.n10281 92.5005
R5259 VDD.n10282 VDD.n6765 92.5005
R5260 VDD.n10283 VDD.n10238 92.5005
R5261 VDD.n10283 VDD.n6770 92.5005
R5262 VDD.n10285 VDD.n10284 92.5005
R5263 VDD.n10284 VDD.n6771 92.5005
R5264 VDD.n10236 VDD.n10235 92.5005
R5265 VDD.n10235 VDD.n6776 92.5005
R5266 VDD.n10291 VDD.n10290 92.5005
R5267 VDD.n10291 VDD.n6777 92.5005
R5268 VDD.n10293 VDD.n10292 92.5005
R5269 VDD.n10292 VDD.n6782 92.5005
R5270 VDD.n10232 VDD.n10231 92.5005
R5271 VDD.n10231 VDD.n6783 92.5005
R5272 VDD.n10299 VDD.n10298 92.5005
R5273 VDD.n10299 VDD.n6788 92.5005
R5274 VDD.n10301 VDD.n10300 92.5005
R5275 VDD.n10300 VDD.n6789 92.5005
R5276 VDD.n10228 VDD.n10227 92.5005
R5277 VDD.n10227 VDD.n10226 92.5005
R5278 VDD.n10307 VDD.n10306 92.5005
R5279 VDD.n10307 VDD.n6793 92.5005
R5280 VDD.n10309 VDD.n10308 92.5005
R5281 VDD.n10308 VDD.n6798 92.5005
R5282 VDD.n10222 VDD.n10221 92.5005
R5283 VDD.n10221 VDD.n6799 92.5005
R5284 VDD.n10315 VDD.n10314 92.5005
R5285 VDD.n10315 VDD.n6804 92.5005
R5286 VDD.n10317 VDD.n10316 92.5005
R5287 VDD.n10316 VDD.n6805 92.5005
R5288 VDD.n10218 VDD.n10217 92.5005
R5289 VDD.n10217 VDD.n6810 92.5005
R5290 VDD.n10323 VDD.n10322 92.5005
R5291 VDD.n10323 VDD.n6811 92.5005
R5292 VDD.n10325 VDD.n10324 92.5005
R5293 VDD.n10324 VDD.n6816 92.5005
R5294 VDD.n10214 VDD.n10213 92.5005
R5295 VDD.n10213 VDD.n10212 92.5005
R5296 VDD.n10333 VDD.n10332 92.5005
R5297 VDD.n10333 VDD.n6820 92.5005
R5298 VDD.n10336 VDD.n10209 92.5005
R5299 VDD.n10336 VDD.n10335 92.5005
R5300 VDD.n10338 VDD.n10337 92.5005
R5301 VDD.n10337 VDD.n6824 92.5005
R5302 VDD.n10207 VDD.n10206 92.5005
R5303 VDD.n10206 VDD.n6825 92.5005
R5304 VDD.n10344 VDD.n10343 92.5005
R5305 VDD.n10344 VDD.n6830 92.5005
R5306 VDD.n10346 VDD.n10345 92.5005
R5307 VDD.n10345 VDD.n6831 92.5005
R5308 VDD.n10203 VDD.n10202 92.5005
R5309 VDD.n10202 VDD.n6836 92.5005
R5310 VDD.n10352 VDD.n10351 92.5005
R5311 VDD.n10352 VDD.n6837 92.5005
R5312 VDD.n10354 VDD.n10353 92.5005
R5313 VDD.n10353 VDD.n6842 92.5005
R5314 VDD.n10199 VDD.n10198 92.5005
R5315 VDD.n10198 VDD.n6843 92.5005
R5316 VDD.n10360 VDD.n10359 92.5005
R5317 VDD.n10360 VDD.n6848 92.5005
R5318 VDD.n10362 VDD.n10361 92.5005
R5319 VDD.n10361 VDD.n6849 92.5005
R5320 VDD.n10195 VDD.n10194 92.5005
R5321 VDD.n10194 VDD.n10193 92.5005
R5322 VDD.n10368 VDD.n10367 92.5005
R5323 VDD.n10368 VDD.n6853 92.5005
R5324 VDD.n10370 VDD.n10369 92.5005
R5325 VDD.n10369 VDD.n6858 92.5005
R5326 VDD.n10189 VDD.n10188 92.5005
R5327 VDD.n10188 VDD.n6859 92.5005
R5328 VDD.n10376 VDD.n10375 92.5005
R5329 VDD.n10376 VDD.n6864 92.5005
R5330 VDD.n10379 VDD.n10378 92.5005
R5331 VDD.n10378 VDD.n6865 92.5005
R5332 VDD.n10377 VDD.n10185 92.5005
R5333 VDD.n10377 VDD.n6870 92.5005
R5334 VDD.n10384 VDD.n10184 92.5005
R5335 VDD.n10184 VDD.n10183 92.5005
R5336 VDD.n10386 VDD.n10385 92.5005
R5337 VDD.n10386 VDD.n6874 92.5005
R5338 VDD.n10388 VDD.n10387 92.5005
R5339 VDD.n10387 VDD.n6875 92.5005
R5340 VDD.n10179 VDD.n10178 92.5005
R5341 VDD.n10178 VDD.n6880 92.5005
R5342 VDD.n10394 VDD.n10393 92.5005
R5343 VDD.n10394 VDD.n6881 92.5005
R5344 VDD.n10396 VDD.n10395 92.5005
R5345 VDD.n10395 VDD.n6886 92.5005
R5346 VDD.n10175 VDD.n10174 92.5005
R5347 VDD.n10174 VDD.n6887 92.5005
R5348 VDD.n10402 VDD.n10401 92.5005
R5349 VDD.n10402 VDD.n6892 92.5005
R5350 VDD.n10404 VDD.n10403 92.5005
R5351 VDD.n10403 VDD.n6893 92.5005
R5352 VDD.n10171 VDD.n10170 92.5005
R5353 VDD.n10170 VDD.n6898 92.5005
R5354 VDD.n10410 VDD.n10409 92.5005
R5355 VDD.n10410 VDD.n6899 92.5005
R5356 VDD.n10412 VDD.n10411 92.5005
R5357 VDD.n10411 VDD.n6904 92.5005
R5358 VDD.n10167 VDD.n10165 92.5005
R5359 VDD.n10165 VDD.n6905 92.5005
R5360 VDD.n10419 VDD.n10418 92.5005
R5361 VDD.n10420 VDD.n10419 92.5005
R5362 VDD.n10166 VDD.n6926 92.5005
R5363 VDD.n10166 VDD.n6913 92.5005
R5364 VDD.n6931 VDD.n6927 92.5005
R5365 VDD.n10479 VDD.n6931 92.5005
R5366 VDD.n12679 VDD.n12678 92.5005
R5367 VDD.n12680 VDD.n12679 92.5005
R5368 VDD.n12677 VDD.n6716 92.5005
R5369 VDD.n6722 VDD.n6716 92.5005
R5370 VDD.n12676 VDD.n12675 92.5005
R5371 VDD.n12675 VDD.n12674 92.5005
R5372 VDD.n6719 VDD.n6718 92.5005
R5373 VDD.n6747 VDD.n6719 92.5005
R5374 VDD.n12667 VDD.n12666 92.5005
R5375 VDD.n12668 VDD.n12667 92.5005
R5376 VDD.n12665 VDD.n6750 92.5005
R5377 VDD.n6753 VDD.n6750 92.5005
R5378 VDD.n12664 VDD.n12663 92.5005
R5379 VDD.n12663 VDD.n12662 92.5005
R5380 VDD.n6752 VDD.n6751 92.5005
R5381 VDD.n10243 VDD.n6752 92.5005
R5382 VDD.n12655 VDD.n12654 92.5005
R5383 VDD.n12656 VDD.n12655 92.5005
R5384 VDD.n12653 VDD.n6760 92.5005
R5385 VDD.n6763 VDD.n6760 92.5005
R5386 VDD.n12652 VDD.n12651 92.5005
R5387 VDD.n12651 VDD.n12650 92.5005
R5388 VDD.n6762 VDD.n6761 92.5005
R5389 VDD.n6769 VDD.n6762 92.5005
R5390 VDD.n12643 VDD.n12642 92.5005
R5391 VDD.n12644 VDD.n12643 92.5005
R5392 VDD.n12641 VDD.n6772 92.5005
R5393 VDD.n6775 VDD.n6772 92.5005
R5394 VDD.n12640 VDD.n12639 92.5005
R5395 VDD.n12639 VDD.n12638 92.5005
R5396 VDD.n6774 VDD.n6773 92.5005
R5397 VDD.n6781 VDD.n6774 92.5005
R5398 VDD.n12631 VDD.n12630 92.5005
R5399 VDD.n12632 VDD.n12631 92.5005
R5400 VDD.n12629 VDD.n6784 92.5005
R5401 VDD.n6787 VDD.n6784 92.5005
R5402 VDD.n12628 VDD.n12627 92.5005
R5403 VDD.n12627 VDD.n12626 92.5005
R5404 VDD.n6786 VDD.n6785 92.5005
R5405 VDD.n10225 VDD.n6786 92.5005
R5406 VDD.n12619 VDD.n12618 92.5005
R5407 VDD.n12620 VDD.n12619 92.5005
R5408 VDD.n12617 VDD.n6794 92.5005
R5409 VDD.n6797 VDD.n6794 92.5005
R5410 VDD.n12616 VDD.n12615 92.5005
R5411 VDD.n12615 VDD.n12614 92.5005
R5412 VDD.n6796 VDD.n6795 92.5005
R5413 VDD.n6803 VDD.n6796 92.5005
R5414 VDD.n12607 VDD.n12606 92.5005
R5415 VDD.n12608 VDD.n12607 92.5005
R5416 VDD.n12605 VDD.n6806 92.5005
R5417 VDD.n6809 VDD.n6806 92.5005
R5418 VDD.n12604 VDD.n12603 92.5005
R5419 VDD.n12603 VDD.n12602 92.5005
R5420 VDD.n6808 VDD.n6807 92.5005
R5421 VDD.n6815 VDD.n6808 92.5005
R5422 VDD.n12595 VDD.n12594 92.5005
R5423 VDD.n12596 VDD.n12595 92.5005
R5424 VDD.n12593 VDD.n6817 92.5005
R5425 VDD.n10211 VDD.n6817 92.5005
R5426 VDD.n12592 VDD.n12591 92.5005
R5427 VDD.n12591 VDD.n12590 92.5005
R5428 VDD.n6819 VDD.n6818 92.5005
R5429 VDD.n10334 VDD.n6819 92.5005
R5430 VDD.n12583 VDD.n12582 92.5005
R5431 VDD.n12584 VDD.n12583 92.5005
R5432 VDD.n12581 VDD.n6826 92.5005
R5433 VDD.n6829 VDD.n6826 92.5005
R5434 VDD.n12580 VDD.n12579 92.5005
R5435 VDD.n12579 VDD.n12578 92.5005
R5436 VDD.n6828 VDD.n6827 92.5005
R5437 VDD.n6835 VDD.n6828 92.5005
R5438 VDD.n12571 VDD.n12570 92.5005
R5439 VDD.n12572 VDD.n12571 92.5005
R5440 VDD.n12569 VDD.n6838 92.5005
R5441 VDD.n6841 VDD.n6838 92.5005
R5442 VDD.n12568 VDD.n12567 92.5005
R5443 VDD.n12567 VDD.n12566 92.5005
R5444 VDD.n6840 VDD.n6839 92.5005
R5445 VDD.n6847 VDD.n6840 92.5005
R5446 VDD.n12559 VDD.n12558 92.5005
R5447 VDD.n12560 VDD.n12559 92.5005
R5448 VDD.n12557 VDD.n6850 92.5005
R5449 VDD.n10192 VDD.n6850 92.5005
R5450 VDD.n12556 VDD.n12555 92.5005
R5451 VDD.n12555 VDD.n12554 92.5005
R5452 VDD.n6852 VDD.n6851 92.5005
R5453 VDD.n6857 VDD.n6852 92.5005
R5454 VDD.n12547 VDD.n12546 92.5005
R5455 VDD.n12548 VDD.n12547 92.5005
R5456 VDD.n12545 VDD.n6860 92.5005
R5457 VDD.n6863 VDD.n6860 92.5005
R5458 VDD.n12544 VDD.n12543 92.5005
R5459 VDD.n12543 VDD.n12542 92.5005
R5460 VDD.n6862 VDD.n6861 92.5005
R5461 VDD.n6869 VDD.n6862 92.5005
R5462 VDD.n12535 VDD.n12534 92.5005
R5463 VDD.n12536 VDD.n12535 92.5005
R5464 VDD.n12533 VDD.n6871 92.5005
R5465 VDD.n10182 VDD.n6871 92.5005
R5466 VDD.n12532 VDD.n12531 92.5005
R5467 VDD.n12531 VDD.n12530 92.5005
R5468 VDD.n6873 VDD.n6872 92.5005
R5469 VDD.n6879 VDD.n6873 92.5005
R5470 VDD.n12523 VDD.n12522 92.5005
R5471 VDD.n12524 VDD.n12523 92.5005
R5472 VDD.n12521 VDD.n6882 92.5005
R5473 VDD.n6885 VDD.n6882 92.5005
R5474 VDD.n12520 VDD.n12519 92.5005
R5475 VDD.n12519 VDD.n12518 92.5005
R5476 VDD.n6884 VDD.n6883 92.5005
R5477 VDD.n6891 VDD.n6884 92.5005
R5478 VDD.n12511 VDD.n12510 92.5005
R5479 VDD.n12512 VDD.n12511 92.5005
R5480 VDD.n12509 VDD.n6894 92.5005
R5481 VDD.n6897 VDD.n6894 92.5005
R5482 VDD.n12508 VDD.n12507 92.5005
R5483 VDD.n12507 VDD.n12506 92.5005
R5484 VDD.n6896 VDD.n6895 92.5005
R5485 VDD.n6903 VDD.n6896 92.5005
R5486 VDD.n12499 VDD.n12498 92.5005
R5487 VDD.n12500 VDD.n12499 92.5005
R5488 VDD.n12497 VDD.n6906 92.5005
R5489 VDD.n10164 VDD.n6906 92.5005
R5490 VDD.n6730 VDD.n6729 92.5005
R5491 VDD.n6732 VDD.n6731 92.5005
R5492 VDD.n6734 VDD.n6727 92.5005
R5493 VDD.n6736 VDD.n6735 92.5005
R5494 VDD.n6738 VDD.n6737 92.5005
R5495 VDD.n6739 VDD.n6725 92.5005
R5496 VDD.n6742 VDD.n6741 92.5005
R5497 VDD.n6717 VDD.n6715 92.5005
R5498 VDD.n6902 VDD.n6901 92.5005
R5499 VDD.n10164 VDD.n6902 92.5005
R5500 VDD.n12502 VDD.n12501 92.5005
R5501 VDD.n12501 VDD.n12500 92.5005
R5502 VDD.n12503 VDD.n6900 92.5005
R5503 VDD.n6903 VDD.n6900 92.5005
R5504 VDD.n12505 VDD.n12504 92.5005
R5505 VDD.n12506 VDD.n12505 92.5005
R5506 VDD.n6890 VDD.n6889 92.5005
R5507 VDD.n6897 VDD.n6890 92.5005
R5508 VDD.n12514 VDD.n12513 92.5005
R5509 VDD.n12513 VDD.n12512 92.5005
R5510 VDD.n12515 VDD.n6888 92.5005
R5511 VDD.n6891 VDD.n6888 92.5005
R5512 VDD.n12517 VDD.n12516 92.5005
R5513 VDD.n12518 VDD.n12517 92.5005
R5514 VDD.n6878 VDD.n6877 92.5005
R5515 VDD.n6885 VDD.n6878 92.5005
R5516 VDD.n12526 VDD.n12525 92.5005
R5517 VDD.n12525 VDD.n12524 92.5005
R5518 VDD.n12527 VDD.n6876 92.5005
R5519 VDD.n6879 VDD.n6876 92.5005
R5520 VDD.n12529 VDD.n12528 92.5005
R5521 VDD.n12530 VDD.n12529 92.5005
R5522 VDD.n6868 VDD.n6867 92.5005
R5523 VDD.n10182 VDD.n6868 92.5005
R5524 VDD.n12538 VDD.n12537 92.5005
R5525 VDD.n12537 VDD.n12536 92.5005
R5526 VDD.n12539 VDD.n6866 92.5005
R5527 VDD.n6869 VDD.n6866 92.5005
R5528 VDD.n12541 VDD.n12540 92.5005
R5529 VDD.n12542 VDD.n12541 92.5005
R5530 VDD.n6856 VDD.n6855 92.5005
R5531 VDD.n6863 VDD.n6856 92.5005
R5532 VDD.n12550 VDD.n12549 92.5005
R5533 VDD.n12549 VDD.n12548 92.5005
R5534 VDD.n12551 VDD.n6854 92.5005
R5535 VDD.n6857 VDD.n6854 92.5005
R5536 VDD.n12553 VDD.n12552 92.5005
R5537 VDD.n12554 VDD.n12553 92.5005
R5538 VDD.n6846 VDD.n6845 92.5005
R5539 VDD.n10192 VDD.n6846 92.5005
R5540 VDD.n12562 VDD.n12561 92.5005
R5541 VDD.n12561 VDD.n12560 92.5005
R5542 VDD.n12563 VDD.n6844 92.5005
R5543 VDD.n6847 VDD.n6844 92.5005
R5544 VDD.n12565 VDD.n12564 92.5005
R5545 VDD.n12566 VDD.n12565 92.5005
R5546 VDD.n6834 VDD.n6833 92.5005
R5547 VDD.n6841 VDD.n6834 92.5005
R5548 VDD.n12574 VDD.n12573 92.5005
R5549 VDD.n12573 VDD.n12572 92.5005
R5550 VDD.n12575 VDD.n6832 92.5005
R5551 VDD.n6835 VDD.n6832 92.5005
R5552 VDD.n12577 VDD.n12576 92.5005
R5553 VDD.n12578 VDD.n12577 92.5005
R5554 VDD.n6823 VDD.n6822 92.5005
R5555 VDD.n6829 VDD.n6823 92.5005
R5556 VDD.n12586 VDD.n12585 92.5005
R5557 VDD.n12585 VDD.n12584 92.5005
R5558 VDD.n12587 VDD.n6821 92.5005
R5559 VDD.n10334 VDD.n6821 92.5005
R5560 VDD.n12589 VDD.n12588 92.5005
R5561 VDD.n12590 VDD.n12589 92.5005
R5562 VDD.n6814 VDD.n6813 92.5005
R5563 VDD.n10211 VDD.n6814 92.5005
R5564 VDD.n12598 VDD.n12597 92.5005
R5565 VDD.n12597 VDD.n12596 92.5005
R5566 VDD.n12599 VDD.n6812 92.5005
R5567 VDD.n6815 VDD.n6812 92.5005
R5568 VDD.n12601 VDD.n12600 92.5005
R5569 VDD.n12602 VDD.n12601 92.5005
R5570 VDD.n6802 VDD.n6801 92.5005
R5571 VDD.n6809 VDD.n6802 92.5005
R5572 VDD.n12610 VDD.n12609 92.5005
R5573 VDD.n12609 VDD.n12608 92.5005
R5574 VDD.n12611 VDD.n6800 92.5005
R5575 VDD.n6803 VDD.n6800 92.5005
R5576 VDD.n12613 VDD.n12612 92.5005
R5577 VDD.n12614 VDD.n12613 92.5005
R5578 VDD.n6792 VDD.n6791 92.5005
R5579 VDD.n6797 VDD.n6792 92.5005
R5580 VDD.n12622 VDD.n12621 92.5005
R5581 VDD.n12621 VDD.n12620 92.5005
R5582 VDD.n12623 VDD.n6790 92.5005
R5583 VDD.n10225 VDD.n6790 92.5005
R5584 VDD.n12625 VDD.n12624 92.5005
R5585 VDD.n12626 VDD.n12625 92.5005
R5586 VDD.n6780 VDD.n6779 92.5005
R5587 VDD.n6787 VDD.n6780 92.5005
R5588 VDD.n12634 VDD.n12633 92.5005
R5589 VDD.n12633 VDD.n12632 92.5005
R5590 VDD.n12635 VDD.n6778 92.5005
R5591 VDD.n6781 VDD.n6778 92.5005
R5592 VDD.n12637 VDD.n12636 92.5005
R5593 VDD.n12638 VDD.n12637 92.5005
R5594 VDD.n6768 VDD.n6767 92.5005
R5595 VDD.n6775 VDD.n6768 92.5005
R5596 VDD.n12646 VDD.n12645 92.5005
R5597 VDD.n12645 VDD.n12644 92.5005
R5598 VDD.n12647 VDD.n6766 92.5005
R5599 VDD.n6769 VDD.n6766 92.5005
R5600 VDD.n12649 VDD.n12648 92.5005
R5601 VDD.n12650 VDD.n12649 92.5005
R5602 VDD.n6757 VDD.n6756 92.5005
R5603 VDD.n6763 VDD.n6757 92.5005
R5604 VDD.n12658 VDD.n12657 92.5005
R5605 VDD.n12657 VDD.n12656 92.5005
R5606 VDD.n12659 VDD.n6755 92.5005
R5607 VDD.n10243 VDD.n6755 92.5005
R5608 VDD.n12661 VDD.n12660 92.5005
R5609 VDD.n12662 VDD.n12661 92.5005
R5610 VDD.n6746 VDD.n6745 92.5005
R5611 VDD.n6753 VDD.n6746 92.5005
R5612 VDD.n12670 VDD.n12669 92.5005
R5613 VDD.n12669 VDD.n12668 92.5005
R5614 VDD.n12671 VDD.n6724 92.5005
R5615 VDD.n6747 VDD.n6724 92.5005
R5616 VDD.n12673 VDD.n12672 92.5005
R5617 VDD.n12674 VDD.n12673 92.5005
R5618 VDD.n6744 VDD.n6723 92.5005
R5619 VDD.n6723 VDD.n6722 92.5005
R5620 VDD.n12680 VDD.n6714 92.5005
R5621 VDD.n6743 VDD.n6714 92.5005
R5622 VDD.n5903 VDD.n5900 92.5005
R5623 VDD.n6364 VDD.n5903 92.5005
R5624 VDD.n6258 VDD.n6257 92.5005
R5625 VDD.n6258 VDD.n5783 92.5005
R5626 VDD.n6044 VDD.n6043 92.5005
R5627 VDD.n6304 VDD.n6044 92.5005
R5628 VDD.n6327 VDD.n6326 92.5005
R5629 VDD.n6326 VDD.n6325 92.5005
R5630 VDD.n6328 VDD.n6024 92.5005
R5631 VDD.n6293 VDD.n6024 92.5005
R5632 VDD.n6330 VDD.n6329 92.5005
R5633 VDD.n6331 VDD.n6330 92.5005
R5634 VDD.n6042 VDD.n6023 92.5005
R5635 VDD.n6023 VDD.n6007 92.5005
R5636 VDD.n6037 VDD.n6025 92.5005
R5637 VDD.n6036 VDD.n6035 92.5005
R5638 VDD.n6034 VDD.n6033 92.5005
R5639 VDD.n6032 VDD.n6028 92.5005
R5640 VDD.n6030 VDD.n6029 92.5005
R5641 VDD.n6040 VDD.n6039 92.5005
R5642 VDD.n5929 VDD.n5928 92.5005
R5643 VDD.n5939 VDD.n5929 92.5005
R5644 VDD.n6352 VDD.n6351 92.5005
R5645 VDD.n6351 VDD.n6350 92.5005
R5646 VDD.n6353 VDD.n5926 92.5005
R5647 VDD.n5930 VDD.n5926 92.5005
R5648 VDD.n6355 VDD.n6354 92.5005
R5649 VDD.n6356 VDD.n6355 92.5005
R5650 VDD.n5927 VDD.n5925 92.5005
R5651 VDD.n5925 VDD.n5917 92.5005
R5652 VDD.n6395 VDD.n5876 92.5005
R5653 VDD.n5876 VDD.n5875 92.5005
R5654 VDD.n6418 VDD.n6417 92.5005
R5655 VDD.n6417 VDD.n6416 92.5005
R5656 VDD.n5866 VDD.n5865 92.5005
R5657 VDD.n6415 VDD.n5866 92.5005
R5658 VDD.n6413 VDD.n6412 92.5005
R5659 VDD.n6414 VDD.n6413 92.5005
R5660 VDD.n6411 VDD.n5868 92.5005
R5661 VDD.n5868 VDD.n5867 92.5005
R5662 VDD.n6410 VDD.n6409 92.5005
R5663 VDD.n6409 VDD.n6408 92.5005
R5664 VDD.n5870 VDD.n5869 92.5005
R5665 VDD.n6407 VDD.n5870 92.5005
R5666 VDD.n6405 VDD.n6404 92.5005
R5667 VDD.n6406 VDD.n6405 92.5005
R5668 VDD.n6403 VDD.n5872 92.5005
R5669 VDD.n5872 VDD.n5871 92.5005
R5670 VDD.n6402 VDD.n6401 92.5005
R5671 VDD.n6401 VDD.n6400 92.5005
R5672 VDD.n5874 VDD.n5873 92.5005
R5673 VDD.n6399 VDD.n5874 92.5005
R5674 VDD.n6397 VDD.n6396 92.5005
R5675 VDD.n6398 VDD.n6397 92.5005
R5676 VDD.n6419 VDD.n5863 92.5005
R5677 VDD.n5863 VDD.n5862 92.5005
R5678 VDD.n6422 VDD.n6421 92.5005
R5679 VDD.n6423 VDD.n6422 92.5005
R5680 VDD.n6420 VDD.n5864 92.5005
R5681 VDD.n5860 VDD.n5859 92.5005
R5682 VDD.n6427 VDD.n6426 92.5005
R5683 VDD.n6426 VDD.n6425 92.5005
R5684 VDD.n6430 VDD.n6429 92.5005
R5685 VDD.n6431 VDD.n6430 92.5005
R5686 VDD.n5856 VDD.n5855 92.5005
R5687 VDD.n6432 VDD.n5856 92.5005
R5688 VDD.n6435 VDD.n6434 92.5005
R5689 VDD.n6434 VDD.n6433 92.5005
R5690 VDD.n6436 VDD.n5854 92.5005
R5691 VDD.n5854 VDD.n5853 92.5005
R5692 VDD.n6438 VDD.n6437 92.5005
R5693 VDD.n6439 VDD.n6438 92.5005
R5694 VDD.n5852 VDD.n5851 92.5005
R5695 VDD.n6440 VDD.n5852 92.5005
R5696 VDD.n6443 VDD.n6442 92.5005
R5697 VDD.n6442 VDD.n6441 92.5005
R5698 VDD.n6444 VDD.n5850 92.5005
R5699 VDD.n5850 VDD.n5849 92.5005
R5700 VDD.n6446 VDD.n6445 92.5005
R5701 VDD.n6447 VDD.n6446 92.5005
R5702 VDD.n5848 VDD.n5847 92.5005
R5703 VDD.n6448 VDD.n5848 92.5005
R5704 VDD.n6451 VDD.n6450 92.5005
R5705 VDD.n6450 VDD.n6449 92.5005
R5706 VDD.n6452 VDD.n5846 92.5005
R5707 VDD.n5846 VDD.n5845 92.5005
R5708 VDD.n6454 VDD.n6453 92.5005
R5709 VDD.n6455 VDD.n6454 92.5005
R5710 VDD.n5844 VDD.n5843 92.5005
R5711 VDD.n6456 VDD.n5844 92.5005
R5712 VDD.n6459 VDD.n6458 92.5005
R5713 VDD.n6458 VDD.n6457 92.5005
R5714 VDD.n6460 VDD.n5842 92.5005
R5715 VDD.n5842 VDD.n5841 92.5005
R5716 VDD.n6462 VDD.n6461 92.5005
R5717 VDD.n6463 VDD.n6462 92.5005
R5718 VDD.n5840 VDD.n5839 92.5005
R5719 VDD.n6464 VDD.n5840 92.5005
R5720 VDD.n6467 VDD.n6466 92.5005
R5721 VDD.n6466 VDD.n6465 92.5005
R5722 VDD.n6468 VDD.n5838 92.5005
R5723 VDD.n5838 VDD.n5837 92.5005
R5724 VDD.n6470 VDD.n6469 92.5005
R5725 VDD.n6471 VDD.n6470 92.5005
R5726 VDD.n5836 VDD.n5835 92.5005
R5727 VDD.n6472 VDD.n5836 92.5005
R5728 VDD.n6475 VDD.n6474 92.5005
R5729 VDD.n6474 VDD.n6473 92.5005
R5730 VDD.n6476 VDD.n5834 92.5005
R5731 VDD.n5834 VDD.n5833 92.5005
R5732 VDD.n6478 VDD.n6477 92.5005
R5733 VDD.n6479 VDD.n6478 92.5005
R5734 VDD.n5832 VDD.n5831 92.5005
R5735 VDD.n6480 VDD.n5832 92.5005
R5736 VDD.n6483 VDD.n6482 92.5005
R5737 VDD.n6482 VDD.n6481 92.5005
R5738 VDD.n6484 VDD.n5829 92.5005
R5739 VDD.n5829 VDD.n5826 92.5005
R5740 VDD.n6428 VDD.n5858 92.5005
R5741 VDD.n5858 VDD.n5857 92.5005
R5742 VDD.n5821 VDD.n5820 92.5005
R5743 VDD.n6496 VDD.n5821 92.5005
R5744 VDD.n6499 VDD.n6498 92.5005
R5745 VDD.n6498 VDD.n6497 92.5005
R5746 VDD.n6500 VDD.n5819 92.5005
R5747 VDD.n5819 VDD.n5818 92.5005
R5748 VDD.n6502 VDD.n6501 92.5005
R5749 VDD.n6503 VDD.n6502 92.5005
R5750 VDD.n5817 VDD.n5816 92.5005
R5751 VDD.n6504 VDD.n5817 92.5005
R5752 VDD.n6507 VDD.n6506 92.5005
R5753 VDD.n6506 VDD.n6505 92.5005
R5754 VDD.n6508 VDD.n5815 92.5005
R5755 VDD.n5815 VDD.n5814 92.5005
R5756 VDD.n6510 VDD.n6509 92.5005
R5757 VDD.n6511 VDD.n6510 92.5005
R5758 VDD.n5812 VDD.n5811 92.5005
R5759 VDD.n6512 VDD.n5812 92.5005
R5760 VDD.n6515 VDD.n6514 92.5005
R5761 VDD.n6514 VDD.n6513 92.5005
R5762 VDD.n6516 VDD.n5810 92.5005
R5763 VDD.n5813 VDD.n5810 92.5005
R5764 VDD.n6492 VDD.n5823 92.5005
R5765 VDD.n5823 VDD.n5822 92.5005
R5766 VDD.n6491 VDD.n6490 92.5005
R5767 VDD.n6490 VDD.n6489 92.5005
R5768 VDD.n5825 VDD.n5824 92.5005
R5769 VDD.n5830 VDD.n5828 92.5005
R5770 VDD.n6486 VDD.n6485 92.5005
R5771 VDD.n6487 VDD.n6486 92.5005
R5772 VDD.n6494 VDD.n6493 92.5005
R5773 VDD.n6495 VDD.n6494 92.5005
R5774 VDD.n6519 VDD.n6518 92.5005
R5775 VDD.n6540 VDD.n5794 92.5005
R5776 VDD.n6539 VDD.n6538 92.5005
R5777 VDD.n5803 VDD.n5799 92.5005
R5778 VDD.n6533 VDD.n6532 92.5005
R5779 VDD.n6530 VDD.n6529 92.5005
R5780 VDD.n5805 VDD.n5804 92.5005
R5781 VDD.n6523 VDD.n6522 92.5005
R5782 VDD.n6521 VDD.n5808 92.5005
R5783 VDD.n6543 VDD.n6542 92.5005
R5784 VDD.n6280 VDD.n5779 92.5005
R5785 VDD.n6282 VDD.n5778 92.5005
R5786 VDD.n6054 VDD.n6053 92.5005
R5787 VDD.n6264 VDD.n6263 92.5005
R5788 VDD.n6268 VDD.n6267 92.5005
R5789 VDD.n6266 VDD.n6050 92.5005
R5790 VDD.n6277 VDD.n6276 92.5005
R5791 VDD.n6278 VDD.n6047 92.5005
R5792 VDD.n6275 VDD.n6046 92.5005
R5793 VDD.n6274 VDD.n6273 92.5005
R5794 VDD.n6270 VDD.n6269 92.5005
R5795 VDD.n6259 VDD.n6052 92.5005
R5796 VDD.n6262 VDD.n6261 92.5005
R5797 VDD.n6252 VDD.n6055 92.5005
R5798 VDD.n6255 VDD.n6254 92.5005
R5799 VDD.n6288 VDD.n6287 92.5005
R5800 VDD.n6288 VDD.n5784 92.5005
R5801 VDD.n6286 VDD.n6285 92.5005
R5802 VDD.n6284 VDD.n6048 92.5005
R5803 VDD.n6212 VDD.n6071 92.5005
R5804 VDD.n6214 VDD.n6213 92.5005
R5805 VDD.n6216 VDD.n6215 92.5005
R5806 VDD.n6217 VDD.n6073 92.5005
R5807 VDD.n6219 VDD.n6218 92.5005
R5808 VDD.n6070 VDD.n6069 92.5005
R5809 VDD.n6223 VDD.n6070 92.5005
R5810 VDD.n6226 VDD.n6225 92.5005
R5811 VDD.n6225 VDD.n6224 92.5005
R5812 VDD.n6227 VDD.n6068 92.5005
R5813 VDD.n6068 VDD.n6067 92.5005
R5814 VDD.n6229 VDD.n6228 92.5005
R5815 VDD.n6230 VDD.n6229 92.5005
R5816 VDD.n6066 VDD.n6065 92.5005
R5817 VDD.n6231 VDD.n6066 92.5005
R5818 VDD.n6234 VDD.n6233 92.5005
R5819 VDD.n6233 VDD.n6232 92.5005
R5820 VDD.n6235 VDD.n6064 92.5005
R5821 VDD.n6064 VDD.n6063 92.5005
R5822 VDD.n6237 VDD.n6236 92.5005
R5823 VDD.n6238 VDD.n6237 92.5005
R5824 VDD.n6062 VDD.n6061 92.5005
R5825 VDD.n6239 VDD.n6062 92.5005
R5826 VDD.n6242 VDD.n6241 92.5005
R5827 VDD.n6241 VDD.n6240 92.5005
R5828 VDD.n6243 VDD.n6060 92.5005
R5829 VDD.n6060 VDD.n6059 92.5005
R5830 VDD.n6246 VDD.n6245 92.5005
R5831 VDD.n6247 VDD.n6246 92.5005
R5832 VDD.n6244 VDD.n6057 92.5005
R5833 VDD.n6248 VDD.n6057 92.5005
R5834 VDD.n6251 VDD.n6058 92.5005
R5835 VDD.n6251 VDD.n6250 92.5005
R5836 VDD.n6100 VDD.n6099 92.5005
R5837 VDD.n6160 VDD.n6100 92.5005
R5838 VDD.n6163 VDD.n6162 92.5005
R5839 VDD.n6162 VDD.n6161 92.5005
R5840 VDD.n6164 VDD.n6098 92.5005
R5841 VDD.n6098 VDD.n6097 92.5005
R5842 VDD.n6166 VDD.n6165 92.5005
R5843 VDD.n6167 VDD.n6166 92.5005
R5844 VDD.n6096 VDD.n6095 92.5005
R5845 VDD.n6168 VDD.n6096 92.5005
R5846 VDD.n6171 VDD.n6170 92.5005
R5847 VDD.n6170 VDD.n6169 92.5005
R5848 VDD.n6172 VDD.n6094 92.5005
R5849 VDD.n6094 VDD.n6093 92.5005
R5850 VDD.n6174 VDD.n6173 92.5005
R5851 VDD.n6175 VDD.n6174 92.5005
R5852 VDD.n6092 VDD.n6091 92.5005
R5853 VDD.n6176 VDD.n6092 92.5005
R5854 VDD.n6179 VDD.n6178 92.5005
R5855 VDD.n6178 VDD.n6177 92.5005
R5856 VDD.n6180 VDD.n6090 92.5005
R5857 VDD.n6090 VDD.n6089 92.5005
R5858 VDD.n6182 VDD.n6181 92.5005
R5859 VDD.n6183 VDD.n6182 92.5005
R5860 VDD.n6088 VDD.n6087 92.5005
R5861 VDD.n6184 VDD.n6088 92.5005
R5862 VDD.n6187 VDD.n6186 92.5005
R5863 VDD.n6186 VDD.n6185 92.5005
R5864 VDD.n6188 VDD.n6086 92.5005
R5865 VDD.n6086 VDD.n6085 92.5005
R5866 VDD.n6190 VDD.n6189 92.5005
R5867 VDD.n6191 VDD.n6190 92.5005
R5868 VDD.n6084 VDD.n6083 92.5005
R5869 VDD.n6192 VDD.n6084 92.5005
R5870 VDD.n6195 VDD.n6194 92.5005
R5871 VDD.n6194 VDD.n6193 92.5005
R5872 VDD.n6196 VDD.n6082 92.5005
R5873 VDD.n6082 VDD.n6081 92.5005
R5874 VDD.n6198 VDD.n6197 92.5005
R5875 VDD.n6199 VDD.n6198 92.5005
R5876 VDD.n6080 VDD.n6079 92.5005
R5877 VDD.n6200 VDD.n6080 92.5005
R5878 VDD.n6203 VDD.n6202 92.5005
R5879 VDD.n6202 VDD.n6201 92.5005
R5880 VDD.n6204 VDD.n6078 92.5005
R5881 VDD.n6078 VDD.n6077 92.5005
R5882 VDD.n6207 VDD.n6206 92.5005
R5883 VDD.n6208 VDD.n6207 92.5005
R5884 VDD.n6205 VDD.n6075 92.5005
R5885 VDD.n6209 VDD.n6075 92.5005
R5886 VDD.n6211 VDD.n6076 92.5005
R5887 VDD.n6211 VDD.n6210 92.5005
R5888 VDD.n6155 VDD.n6154 92.5005
R5889 VDD.n6102 VDD.n6101 92.5005
R5890 VDD.n6159 VDD.n6158 92.5005
R5891 VDD.n5899 VDD.n5898 92.5005
R5892 VDD.n6121 VDD.n5898 92.5005
R5893 VDD.n6124 VDD.n6123 92.5005
R5894 VDD.n6123 VDD.n6122 92.5005
R5895 VDD.n6126 VDD.n6125 92.5005
R5896 VDD.n6127 VDD.n6126 92.5005
R5897 VDD.n6120 VDD.n6119 92.5005
R5898 VDD.n6128 VDD.n6120 92.5005
R5899 VDD.n6131 VDD.n6130 92.5005
R5900 VDD.n6130 VDD.n6129 92.5005
R5901 VDD.n6132 VDD.n6118 92.5005
R5902 VDD.n6118 VDD.n6117 92.5005
R5903 VDD.n6134 VDD.n6133 92.5005
R5904 VDD.n6135 VDD.n6134 92.5005
R5905 VDD.n6116 VDD.n6115 92.5005
R5906 VDD.n6136 VDD.n6116 92.5005
R5907 VDD.n6139 VDD.n6138 92.5005
R5908 VDD.n6138 VDD.n6137 92.5005
R5909 VDD.n6140 VDD.n6114 92.5005
R5910 VDD.n6114 VDD.n6113 92.5005
R5911 VDD.n6142 VDD.n6141 92.5005
R5912 VDD.n6143 VDD.n6142 92.5005
R5913 VDD.n6111 VDD.n6110 92.5005
R5914 VDD.n6144 VDD.n6111 92.5005
R5915 VDD.n6147 VDD.n6146 92.5005
R5916 VDD.n6146 VDD.n6145 92.5005
R5917 VDD.n6148 VDD.n6108 92.5005
R5918 VDD.n6112 VDD.n6108 92.5005
R5919 VDD.n6150 VDD.n6149 92.5005
R5920 VDD.n6109 VDD.n6107 92.5005
R5921 VDD.n6104 VDD.n6103 92.5005
R5922 VDD.n6394 VDD.n6393 92.5005
R5923 VDD.n5975 VDD.n5878 92.5005
R5924 VDD.n5977 VDD.n5976 92.5005
R5925 VDD.n5974 VDD.n5973 92.5005
R5926 VDD.n5944 VDD.n5943 92.5005
R5927 VDD.n5968 VDD.n5967 92.5005
R5928 VDD.n5946 VDD.n5945 92.5005
R5929 VDD.n5962 VDD.n5961 92.5005
R5930 VDD.n5958 VDD.n5957 92.5005
R5931 VDD.n5956 VDD.n5955 92.5005
R5932 VDD.n6369 VDD.n6368 92.5005
R5933 VDD.n6373 VDD.n6372 92.5005
R5934 VDD.n6376 VDD.n6375 92.5005
R5935 VDD.n5913 VDD.n5912 92.5005
R5936 VDD.n5902 VDD.n5901 92.5005
R5937 VDD.n6385 VDD.n6384 92.5005
R5938 VDD.n6386 VDD.n5897 92.5005
R5939 VDD.n6389 VDD.n6388 92.5005
R5940 VDD.n6383 VDD.n6382 92.5005
R5941 VDD.n5911 VDD.n5904 92.5005
R5942 VDD.n6378 VDD.n6377 92.5005
R5943 VDD.n6374 VDD.n5910 92.5005
R5944 VDD.n6371 VDD.n6370 92.5005
R5945 VDD.n5914 VDD.n5890 92.5005
R5946 VDD.n6391 VDD.n5890 92.5005
R5947 VDD.n6367 VDD.n6366 92.5005
R5948 VDD.n5950 VDD.n5949 92.5005
R5949 VDD.n5952 VDD.n5951 92.5005
R5950 VDD.n5954 VDD.n5953 92.5005
R5951 VDD.n5960 VDD.n5959 92.5005
R5952 VDD.n5979 VDD.n5978 92.5005
R5953 VDD.n5972 VDD.n5971 92.5005
R5954 VDD.n5970 VDD.n5969 92.5005
R5955 VDD.n5966 VDD.n5965 92.5005
R5956 VDD.n5964 VDD.n5963 92.5005
R5957 VDD.n5790 VDD.n5782 92.5005
R5958 VDD.n6547 VDD.n6546 92.5005
R5959 VDD.n6545 VDD.n6544 92.5005
R5960 VDD.n6545 VDD.n5791 92.5005
R5961 VDD.n6537 VDD.n6536 92.5005
R5962 VDD.n6535 VDD.n6534 92.5005
R5963 VDD.n5806 VDD.n5802 92.5005
R5964 VDD.n6528 VDD.n6527 92.5005
R5965 VDD.n6525 VDD.n6524 92.5005
R5966 VDD.n5798 VDD.n5793 92.5005
R5967 VDD.n6309 VDD.n6308 92.5005
R5968 VDD.n6311 VDD.n6310 92.5005
R5969 VDD.n6313 VDD.n6312 92.5005
R5970 VDD.n6315 VDD.n6314 92.5005
R5971 VDD.n6303 VDD.n6302 92.5005
R5972 VDD.n6320 VDD.n6319 92.5005
R5973 VDD.n5789 VDD.n5788 92.5005
R5974 VDD.n5791 VDD.n5789 92.5005
R5975 VDD.n6549 VDD.n6548 92.5005
R5976 VDD.n6548 VDD.n6547 92.5005
R5977 VDD.n6550 VDD.n5786 92.5005
R5978 VDD.n5790 VDD.n5786 92.5005
R5979 VDD.n6552 VDD.n6551 92.5005
R5980 VDD.n6553 VDD.n6552 92.5005
R5981 VDD.n6295 VDD.n6294 92.5005
R5982 VDD.n6294 VDD.n6045 92.5005
R5983 VDD.n6297 VDD.n6296 92.5005
R5984 VDD.n6298 VDD.n6297 92.5005
R5985 VDD.n6005 VDD.n6004 92.5005
R5986 VDD.n6022 VDD.n6005 92.5005
R5987 VDD.n6339 VDD.n6338 92.5005
R5988 VDD.n6338 VDD.n6337 92.5005
R5989 VDD.n6340 VDD.n5942 92.5005
R5990 VDD.n6006 VDD.n5942 92.5005
R5991 VDD.n6342 VDD.n6341 92.5005
R5992 VDD.n6343 VDD.n6342 92.5005
R5993 VDD.n5986 VDD.n5985 92.5005
R5994 VDD.n5985 VDD.n5924 92.5005
R5995 VDD.n5984 VDD.n5983 92.5005
R5996 VDD.n5984 VDD.n5923 92.5005
R5997 VDD.n5982 VDD.n5918 92.5005
R5998 VDD.n6363 VDD.n5918 92.5005
R5999 VDD.n5981 VDD.n5980 92.5005
R6000 VDD.n5980 VDD.n5905 92.5005
R6001 VDD.n6002 VDD.n6001 92.5005
R6002 VDD.n5999 VDD.n5987 92.5005
R6003 VDD.n5997 VDD.n5996 92.5005
R6004 VDD.n5995 VDD.n5994 92.5005
R6005 VDD.n5992 VDD.n5989 92.5005
R6006 VDD.n5990 VDD.n5934 92.5005
R6007 VDD.n5947 VDD.n5919 92.5005
R6008 VDD.n5919 VDD.n5905 92.5005
R6009 VDD.n6362 VDD.n6361 92.5005
R6010 VDD.n6363 VDD.n6362 92.5005
R6011 VDD.n6359 VDD.n5920 92.5005
R6012 VDD.n5923 VDD.n5920 92.5005
R6013 VDD.n5936 VDD.n5921 92.5005
R6014 VDD.n5936 VDD.n5924 92.5005
R6015 VDD.n6345 VDD.n6344 92.5005
R6016 VDD.n6344 VDD.n6343 92.5005
R6017 VDD.n6009 VDD.n5938 92.5005
R6018 VDD.n6006 VDD.n5938 92.5005
R6019 VDD.n6336 VDD.n6335 92.5005
R6020 VDD.n6337 VDD.n6336 92.5005
R6021 VDD.n6020 VDD.n6008 92.5005
R6022 VDD.n6022 VDD.n6008 92.5005
R6023 VDD.n6299 VDD.n6292 92.5005
R6024 VDD.n6299 VDD.n6298 92.5005
R6025 VDD.n6301 VDD.n6300 92.5005
R6026 VDD.n6300 VDD.n6045 92.5005
R6027 VDD.n6555 VDD.n6554 92.5005
R6028 VDD.n6554 VDD.n6553 92.5005
R6029 VDD.n6360 VDD.n5915 92.5005
R6030 VDD.n5917 VDD.n5915 92.5005
R6031 VDD.n6358 VDD.n6357 92.5005
R6032 VDD.n6357 VDD.n6356 92.5005
R6033 VDD.n5933 VDD.n5922 92.5005
R6034 VDD.n5930 VDD.n5922 92.5005
R6035 VDD.n6349 VDD.n6348 92.5005
R6036 VDD.n6350 VDD.n6349 92.5005
R6037 VDD.n6346 VDD.n5932 92.5005
R6038 VDD.n5939 VDD.n5932 92.5005
R6039 VDD.n6334 VDD.n6333 92.5005
R6040 VDD.n6333 VDD.n6007 92.5005
R6041 VDD.n6332 VDD.n6021 92.5005
R6042 VDD.n6332 VDD.n6331 92.5005
R6043 VDD.n6291 VDD.n6019 92.5005
R6044 VDD.n6293 VDD.n6019 92.5005
R6045 VDD.n6324 VDD.n6323 92.5005
R6046 VDD.n6325 VDD.n6324 92.5005
R6047 VDD.n6322 VDD.n6290 92.5005
R6048 VDD.n6304 VDD.n6290 92.5005
R6049 VDD.n6289 VDD.n5780 92.5005
R6050 VDD.n6289 VDD.n5783 92.5005
R6051 VDD.n6365 VDD.n5916 92.5005
R6052 VDD.n6365 VDD.n6364 92.5005
R6053 VDD.n5049 VDD.n5046 92.5005
R6054 VDD.n5510 VDD.n5049 92.5005
R6055 VDD.n5404 VDD.n5403 92.5005
R6056 VDD.n5404 VDD.n4929 92.5005
R6057 VDD.n5190 VDD.n5189 92.5005
R6058 VDD.n5450 VDD.n5190 92.5005
R6059 VDD.n5473 VDD.n5472 92.5005
R6060 VDD.n5472 VDD.n5471 92.5005
R6061 VDD.n5474 VDD.n5170 92.5005
R6062 VDD.n5439 VDD.n5170 92.5005
R6063 VDD.n5476 VDD.n5475 92.5005
R6064 VDD.n5477 VDD.n5476 92.5005
R6065 VDD.n5188 VDD.n5169 92.5005
R6066 VDD.n5169 VDD.n5153 92.5005
R6067 VDD.n5183 VDD.n5171 92.5005
R6068 VDD.n5182 VDD.n5181 92.5005
R6069 VDD.n5180 VDD.n5179 92.5005
R6070 VDD.n5178 VDD.n5174 92.5005
R6071 VDD.n5176 VDD.n5175 92.5005
R6072 VDD.n5186 VDD.n5185 92.5005
R6073 VDD.n5075 VDD.n5074 92.5005
R6074 VDD.n5085 VDD.n5075 92.5005
R6075 VDD.n5498 VDD.n5497 92.5005
R6076 VDD.n5497 VDD.n5496 92.5005
R6077 VDD.n5499 VDD.n5072 92.5005
R6078 VDD.n5076 VDD.n5072 92.5005
R6079 VDD.n5501 VDD.n5500 92.5005
R6080 VDD.n5502 VDD.n5501 92.5005
R6081 VDD.n5073 VDD.n5071 92.5005
R6082 VDD.n5071 VDD.n5063 92.5005
R6083 VDD.n5541 VDD.n5022 92.5005
R6084 VDD.n5022 VDD.n5021 92.5005
R6085 VDD.n5564 VDD.n5563 92.5005
R6086 VDD.n5563 VDD.n5562 92.5005
R6087 VDD.n5012 VDD.n5011 92.5005
R6088 VDD.n5561 VDD.n5012 92.5005
R6089 VDD.n5559 VDD.n5558 92.5005
R6090 VDD.n5560 VDD.n5559 92.5005
R6091 VDD.n5557 VDD.n5014 92.5005
R6092 VDD.n5014 VDD.n5013 92.5005
R6093 VDD.n5556 VDD.n5555 92.5005
R6094 VDD.n5555 VDD.n5554 92.5005
R6095 VDD.n5016 VDD.n5015 92.5005
R6096 VDD.n5553 VDD.n5016 92.5005
R6097 VDD.n5551 VDD.n5550 92.5005
R6098 VDD.n5552 VDD.n5551 92.5005
R6099 VDD.n5549 VDD.n5018 92.5005
R6100 VDD.n5018 VDD.n5017 92.5005
R6101 VDD.n5548 VDD.n5547 92.5005
R6102 VDD.n5547 VDD.n5546 92.5005
R6103 VDD.n5020 VDD.n5019 92.5005
R6104 VDD.n5545 VDD.n5020 92.5005
R6105 VDD.n5543 VDD.n5542 92.5005
R6106 VDD.n5544 VDD.n5543 92.5005
R6107 VDD.n5565 VDD.n5009 92.5005
R6108 VDD.n5009 VDD.n5008 92.5005
R6109 VDD.n5568 VDD.n5567 92.5005
R6110 VDD.n5569 VDD.n5568 92.5005
R6111 VDD.n5566 VDD.n5010 92.5005
R6112 VDD.n5006 VDD.n5005 92.5005
R6113 VDD.n5573 VDD.n5572 92.5005
R6114 VDD.n5572 VDD.n5571 92.5005
R6115 VDD.n5576 VDD.n5575 92.5005
R6116 VDD.n5577 VDD.n5576 92.5005
R6117 VDD.n5002 VDD.n5001 92.5005
R6118 VDD.n5578 VDD.n5002 92.5005
R6119 VDD.n5581 VDD.n5580 92.5005
R6120 VDD.n5580 VDD.n5579 92.5005
R6121 VDD.n5582 VDD.n5000 92.5005
R6122 VDD.n5000 VDD.n4999 92.5005
R6123 VDD.n5584 VDD.n5583 92.5005
R6124 VDD.n5585 VDD.n5584 92.5005
R6125 VDD.n4998 VDD.n4997 92.5005
R6126 VDD.n5586 VDD.n4998 92.5005
R6127 VDD.n5589 VDD.n5588 92.5005
R6128 VDD.n5588 VDD.n5587 92.5005
R6129 VDD.n5590 VDD.n4996 92.5005
R6130 VDD.n4996 VDD.n4995 92.5005
R6131 VDD.n5592 VDD.n5591 92.5005
R6132 VDD.n5593 VDD.n5592 92.5005
R6133 VDD.n4994 VDD.n4993 92.5005
R6134 VDD.n5594 VDD.n4994 92.5005
R6135 VDD.n5597 VDD.n5596 92.5005
R6136 VDD.n5596 VDD.n5595 92.5005
R6137 VDD.n5598 VDD.n4992 92.5005
R6138 VDD.n4992 VDD.n4991 92.5005
R6139 VDD.n5600 VDD.n5599 92.5005
R6140 VDD.n5601 VDD.n5600 92.5005
R6141 VDD.n4990 VDD.n4989 92.5005
R6142 VDD.n5602 VDD.n4990 92.5005
R6143 VDD.n5605 VDD.n5604 92.5005
R6144 VDD.n5604 VDD.n5603 92.5005
R6145 VDD.n5606 VDD.n4988 92.5005
R6146 VDD.n4988 VDD.n4987 92.5005
R6147 VDD.n5608 VDD.n5607 92.5005
R6148 VDD.n5609 VDD.n5608 92.5005
R6149 VDD.n4986 VDD.n4985 92.5005
R6150 VDD.n5610 VDD.n4986 92.5005
R6151 VDD.n5613 VDD.n5612 92.5005
R6152 VDD.n5612 VDD.n5611 92.5005
R6153 VDD.n5614 VDD.n4984 92.5005
R6154 VDD.n4984 VDD.n4983 92.5005
R6155 VDD.n5616 VDD.n5615 92.5005
R6156 VDD.n5617 VDD.n5616 92.5005
R6157 VDD.n4982 VDD.n4981 92.5005
R6158 VDD.n5618 VDD.n4982 92.5005
R6159 VDD.n5621 VDD.n5620 92.5005
R6160 VDD.n5620 VDD.n5619 92.5005
R6161 VDD.n5622 VDD.n4980 92.5005
R6162 VDD.n4980 VDD.n4979 92.5005
R6163 VDD.n5624 VDD.n5623 92.5005
R6164 VDD.n5625 VDD.n5624 92.5005
R6165 VDD.n4978 VDD.n4977 92.5005
R6166 VDD.n5626 VDD.n4978 92.5005
R6167 VDD.n5629 VDD.n5628 92.5005
R6168 VDD.n5628 VDD.n5627 92.5005
R6169 VDD.n5630 VDD.n4975 92.5005
R6170 VDD.n4975 VDD.n4972 92.5005
R6171 VDD.n5574 VDD.n5004 92.5005
R6172 VDD.n5004 VDD.n5003 92.5005
R6173 VDD.n4967 VDD.n4966 92.5005
R6174 VDD.n5642 VDD.n4967 92.5005
R6175 VDD.n5645 VDD.n5644 92.5005
R6176 VDD.n5644 VDD.n5643 92.5005
R6177 VDD.n5646 VDD.n4965 92.5005
R6178 VDD.n4965 VDD.n4964 92.5005
R6179 VDD.n5648 VDD.n5647 92.5005
R6180 VDD.n5649 VDD.n5648 92.5005
R6181 VDD.n4963 VDD.n4962 92.5005
R6182 VDD.n5650 VDD.n4963 92.5005
R6183 VDD.n5653 VDD.n5652 92.5005
R6184 VDD.n5652 VDD.n5651 92.5005
R6185 VDD.n5654 VDD.n4961 92.5005
R6186 VDD.n4961 VDD.n4960 92.5005
R6187 VDD.n5656 VDD.n5655 92.5005
R6188 VDD.n5657 VDD.n5656 92.5005
R6189 VDD.n4958 VDD.n4957 92.5005
R6190 VDD.n5658 VDD.n4958 92.5005
R6191 VDD.n5661 VDD.n5660 92.5005
R6192 VDD.n5660 VDD.n5659 92.5005
R6193 VDD.n5662 VDD.n4956 92.5005
R6194 VDD.n4959 VDD.n4956 92.5005
R6195 VDD.n5638 VDD.n4969 92.5005
R6196 VDD.n4969 VDD.n4968 92.5005
R6197 VDD.n5637 VDD.n5636 92.5005
R6198 VDD.n5636 VDD.n5635 92.5005
R6199 VDD.n4971 VDD.n4970 92.5005
R6200 VDD.n4976 VDD.n4974 92.5005
R6201 VDD.n5632 VDD.n5631 92.5005
R6202 VDD.n5633 VDD.n5632 92.5005
R6203 VDD.n5640 VDD.n5639 92.5005
R6204 VDD.n5641 VDD.n5640 92.5005
R6205 VDD.n5665 VDD.n5664 92.5005
R6206 VDD.n5686 VDD.n4940 92.5005
R6207 VDD.n5685 VDD.n5684 92.5005
R6208 VDD.n4949 VDD.n4945 92.5005
R6209 VDD.n5679 VDD.n5678 92.5005
R6210 VDD.n5676 VDD.n5675 92.5005
R6211 VDD.n4951 VDD.n4950 92.5005
R6212 VDD.n5669 VDD.n5668 92.5005
R6213 VDD.n5667 VDD.n4954 92.5005
R6214 VDD.n5689 VDD.n5688 92.5005
R6215 VDD.n5426 VDD.n4925 92.5005
R6216 VDD.n5428 VDD.n4924 92.5005
R6217 VDD.n5200 VDD.n5199 92.5005
R6218 VDD.n5410 VDD.n5409 92.5005
R6219 VDD.n5414 VDD.n5413 92.5005
R6220 VDD.n5412 VDD.n5196 92.5005
R6221 VDD.n5423 VDD.n5422 92.5005
R6222 VDD.n5424 VDD.n5193 92.5005
R6223 VDD.n5421 VDD.n5192 92.5005
R6224 VDD.n5420 VDD.n5419 92.5005
R6225 VDD.n5416 VDD.n5415 92.5005
R6226 VDD.n5405 VDD.n5198 92.5005
R6227 VDD.n5408 VDD.n5407 92.5005
R6228 VDD.n5398 VDD.n5201 92.5005
R6229 VDD.n5401 VDD.n5400 92.5005
R6230 VDD.n5434 VDD.n5433 92.5005
R6231 VDD.n5434 VDD.n4930 92.5005
R6232 VDD.n5432 VDD.n5431 92.5005
R6233 VDD.n5430 VDD.n5194 92.5005
R6234 VDD.n5358 VDD.n5217 92.5005
R6235 VDD.n5360 VDD.n5359 92.5005
R6236 VDD.n5362 VDD.n5361 92.5005
R6237 VDD.n5363 VDD.n5219 92.5005
R6238 VDD.n5365 VDD.n5364 92.5005
R6239 VDD.n5216 VDD.n5215 92.5005
R6240 VDD.n5369 VDD.n5216 92.5005
R6241 VDD.n5372 VDD.n5371 92.5005
R6242 VDD.n5371 VDD.n5370 92.5005
R6243 VDD.n5373 VDD.n5214 92.5005
R6244 VDD.n5214 VDD.n5213 92.5005
R6245 VDD.n5375 VDD.n5374 92.5005
R6246 VDD.n5376 VDD.n5375 92.5005
R6247 VDD.n5212 VDD.n5211 92.5005
R6248 VDD.n5377 VDD.n5212 92.5005
R6249 VDD.n5380 VDD.n5379 92.5005
R6250 VDD.n5379 VDD.n5378 92.5005
R6251 VDD.n5381 VDD.n5210 92.5005
R6252 VDD.n5210 VDD.n5209 92.5005
R6253 VDD.n5383 VDD.n5382 92.5005
R6254 VDD.n5384 VDD.n5383 92.5005
R6255 VDD.n5208 VDD.n5207 92.5005
R6256 VDD.n5385 VDD.n5208 92.5005
R6257 VDD.n5388 VDD.n5387 92.5005
R6258 VDD.n5387 VDD.n5386 92.5005
R6259 VDD.n5389 VDD.n5206 92.5005
R6260 VDD.n5206 VDD.n5205 92.5005
R6261 VDD.n5392 VDD.n5391 92.5005
R6262 VDD.n5393 VDD.n5392 92.5005
R6263 VDD.n5390 VDD.n5203 92.5005
R6264 VDD.n5394 VDD.n5203 92.5005
R6265 VDD.n5397 VDD.n5204 92.5005
R6266 VDD.n5397 VDD.n5396 92.5005
R6267 VDD.n5246 VDD.n5245 92.5005
R6268 VDD.n5306 VDD.n5246 92.5005
R6269 VDD.n5309 VDD.n5308 92.5005
R6270 VDD.n5308 VDD.n5307 92.5005
R6271 VDD.n5310 VDD.n5244 92.5005
R6272 VDD.n5244 VDD.n5243 92.5005
R6273 VDD.n5312 VDD.n5311 92.5005
R6274 VDD.n5313 VDD.n5312 92.5005
R6275 VDD.n5242 VDD.n5241 92.5005
R6276 VDD.n5314 VDD.n5242 92.5005
R6277 VDD.n5317 VDD.n5316 92.5005
R6278 VDD.n5316 VDD.n5315 92.5005
R6279 VDD.n5318 VDD.n5240 92.5005
R6280 VDD.n5240 VDD.n5239 92.5005
R6281 VDD.n5320 VDD.n5319 92.5005
R6282 VDD.n5321 VDD.n5320 92.5005
R6283 VDD.n5238 VDD.n5237 92.5005
R6284 VDD.n5322 VDD.n5238 92.5005
R6285 VDD.n5325 VDD.n5324 92.5005
R6286 VDD.n5324 VDD.n5323 92.5005
R6287 VDD.n5326 VDD.n5236 92.5005
R6288 VDD.n5236 VDD.n5235 92.5005
R6289 VDD.n5328 VDD.n5327 92.5005
R6290 VDD.n5329 VDD.n5328 92.5005
R6291 VDD.n5234 VDD.n5233 92.5005
R6292 VDD.n5330 VDD.n5234 92.5005
R6293 VDD.n5333 VDD.n5332 92.5005
R6294 VDD.n5332 VDD.n5331 92.5005
R6295 VDD.n5334 VDD.n5232 92.5005
R6296 VDD.n5232 VDD.n5231 92.5005
R6297 VDD.n5336 VDD.n5335 92.5005
R6298 VDD.n5337 VDD.n5336 92.5005
R6299 VDD.n5230 VDD.n5229 92.5005
R6300 VDD.n5338 VDD.n5230 92.5005
R6301 VDD.n5341 VDD.n5340 92.5005
R6302 VDD.n5340 VDD.n5339 92.5005
R6303 VDD.n5342 VDD.n5228 92.5005
R6304 VDD.n5228 VDD.n5227 92.5005
R6305 VDD.n5344 VDD.n5343 92.5005
R6306 VDD.n5345 VDD.n5344 92.5005
R6307 VDD.n5226 VDD.n5225 92.5005
R6308 VDD.n5346 VDD.n5226 92.5005
R6309 VDD.n5349 VDD.n5348 92.5005
R6310 VDD.n5348 VDD.n5347 92.5005
R6311 VDD.n5350 VDD.n5224 92.5005
R6312 VDD.n5224 VDD.n5223 92.5005
R6313 VDD.n5353 VDD.n5352 92.5005
R6314 VDD.n5354 VDD.n5353 92.5005
R6315 VDD.n5351 VDD.n5221 92.5005
R6316 VDD.n5355 VDD.n5221 92.5005
R6317 VDD.n5357 VDD.n5222 92.5005
R6318 VDD.n5357 VDD.n5356 92.5005
R6319 VDD.n5301 VDD.n5300 92.5005
R6320 VDD.n5248 VDD.n5247 92.5005
R6321 VDD.n5305 VDD.n5304 92.5005
R6322 VDD.n5045 VDD.n5044 92.5005
R6323 VDD.n5267 VDD.n5044 92.5005
R6324 VDD.n5270 VDD.n5269 92.5005
R6325 VDD.n5269 VDD.n5268 92.5005
R6326 VDD.n5272 VDD.n5271 92.5005
R6327 VDD.n5273 VDD.n5272 92.5005
R6328 VDD.n5266 VDD.n5265 92.5005
R6329 VDD.n5274 VDD.n5266 92.5005
R6330 VDD.n5277 VDD.n5276 92.5005
R6331 VDD.n5276 VDD.n5275 92.5005
R6332 VDD.n5278 VDD.n5264 92.5005
R6333 VDD.n5264 VDD.n5263 92.5005
R6334 VDD.n5280 VDD.n5279 92.5005
R6335 VDD.n5281 VDD.n5280 92.5005
R6336 VDD.n5262 VDD.n5261 92.5005
R6337 VDD.n5282 VDD.n5262 92.5005
R6338 VDD.n5285 VDD.n5284 92.5005
R6339 VDD.n5284 VDD.n5283 92.5005
R6340 VDD.n5286 VDD.n5260 92.5005
R6341 VDD.n5260 VDD.n5259 92.5005
R6342 VDD.n5288 VDD.n5287 92.5005
R6343 VDD.n5289 VDD.n5288 92.5005
R6344 VDD.n5257 VDD.n5256 92.5005
R6345 VDD.n5290 VDD.n5257 92.5005
R6346 VDD.n5293 VDD.n5292 92.5005
R6347 VDD.n5292 VDD.n5291 92.5005
R6348 VDD.n5294 VDD.n5254 92.5005
R6349 VDD.n5258 VDD.n5254 92.5005
R6350 VDD.n5296 VDD.n5295 92.5005
R6351 VDD.n5255 VDD.n5253 92.5005
R6352 VDD.n5250 VDD.n5249 92.5005
R6353 VDD.n5540 VDD.n5539 92.5005
R6354 VDD.n5121 VDD.n5024 92.5005
R6355 VDD.n5123 VDD.n5122 92.5005
R6356 VDD.n5120 VDD.n5119 92.5005
R6357 VDD.n5090 VDD.n5089 92.5005
R6358 VDD.n5114 VDD.n5113 92.5005
R6359 VDD.n5092 VDD.n5091 92.5005
R6360 VDD.n5108 VDD.n5107 92.5005
R6361 VDD.n5104 VDD.n5103 92.5005
R6362 VDD.n5102 VDD.n5101 92.5005
R6363 VDD.n5515 VDD.n5514 92.5005
R6364 VDD.n5519 VDD.n5518 92.5005
R6365 VDD.n5522 VDD.n5521 92.5005
R6366 VDD.n5059 VDD.n5058 92.5005
R6367 VDD.n5048 VDD.n5047 92.5005
R6368 VDD.n5531 VDD.n5530 92.5005
R6369 VDD.n5532 VDD.n5043 92.5005
R6370 VDD.n5535 VDD.n5534 92.5005
R6371 VDD.n5529 VDD.n5528 92.5005
R6372 VDD.n5057 VDD.n5050 92.5005
R6373 VDD.n5524 VDD.n5523 92.5005
R6374 VDD.n5520 VDD.n5056 92.5005
R6375 VDD.n5517 VDD.n5516 92.5005
R6376 VDD.n5060 VDD.n5036 92.5005
R6377 VDD.n5537 VDD.n5036 92.5005
R6378 VDD.n5513 VDD.n5512 92.5005
R6379 VDD.n5096 VDD.n5095 92.5005
R6380 VDD.n5098 VDD.n5097 92.5005
R6381 VDD.n5100 VDD.n5099 92.5005
R6382 VDD.n5106 VDD.n5105 92.5005
R6383 VDD.n5125 VDD.n5124 92.5005
R6384 VDD.n5118 VDD.n5117 92.5005
R6385 VDD.n5116 VDD.n5115 92.5005
R6386 VDD.n5112 VDD.n5111 92.5005
R6387 VDD.n5110 VDD.n5109 92.5005
R6388 VDD.n4936 VDD.n4928 92.5005
R6389 VDD.n5693 VDD.n5692 92.5005
R6390 VDD.n5691 VDD.n5690 92.5005
R6391 VDD.n5691 VDD.n4937 92.5005
R6392 VDD.n5683 VDD.n5682 92.5005
R6393 VDD.n5681 VDD.n5680 92.5005
R6394 VDD.n4952 VDD.n4948 92.5005
R6395 VDD.n5674 VDD.n5673 92.5005
R6396 VDD.n5671 VDD.n5670 92.5005
R6397 VDD.n4944 VDD.n4939 92.5005
R6398 VDD.n5455 VDD.n5454 92.5005
R6399 VDD.n5457 VDD.n5456 92.5005
R6400 VDD.n5459 VDD.n5458 92.5005
R6401 VDD.n5461 VDD.n5460 92.5005
R6402 VDD.n5449 VDD.n5448 92.5005
R6403 VDD.n5466 VDD.n5465 92.5005
R6404 VDD.n4935 VDD.n4934 92.5005
R6405 VDD.n4937 VDD.n4935 92.5005
R6406 VDD.n5695 VDD.n5694 92.5005
R6407 VDD.n5694 VDD.n5693 92.5005
R6408 VDD.n5696 VDD.n4932 92.5005
R6409 VDD.n4936 VDD.n4932 92.5005
R6410 VDD.n5698 VDD.n5697 92.5005
R6411 VDD.n5699 VDD.n5698 92.5005
R6412 VDD.n5441 VDD.n5440 92.5005
R6413 VDD.n5440 VDD.n5191 92.5005
R6414 VDD.n5443 VDD.n5442 92.5005
R6415 VDD.n5444 VDD.n5443 92.5005
R6416 VDD.n5151 VDD.n5150 92.5005
R6417 VDD.n5168 VDD.n5151 92.5005
R6418 VDD.n5485 VDD.n5484 92.5005
R6419 VDD.n5484 VDD.n5483 92.5005
R6420 VDD.n5486 VDD.n5088 92.5005
R6421 VDD.n5152 VDD.n5088 92.5005
R6422 VDD.n5488 VDD.n5487 92.5005
R6423 VDD.n5489 VDD.n5488 92.5005
R6424 VDD.n5132 VDD.n5131 92.5005
R6425 VDD.n5131 VDD.n5070 92.5005
R6426 VDD.n5130 VDD.n5129 92.5005
R6427 VDD.n5130 VDD.n5069 92.5005
R6428 VDD.n5128 VDD.n5064 92.5005
R6429 VDD.n5509 VDD.n5064 92.5005
R6430 VDD.n5127 VDD.n5126 92.5005
R6431 VDD.n5126 VDD.n5051 92.5005
R6432 VDD.n5148 VDD.n5147 92.5005
R6433 VDD.n5145 VDD.n5133 92.5005
R6434 VDD.n5143 VDD.n5142 92.5005
R6435 VDD.n5141 VDD.n5140 92.5005
R6436 VDD.n5138 VDD.n5135 92.5005
R6437 VDD.n5136 VDD.n5080 92.5005
R6438 VDD.n5093 VDD.n5065 92.5005
R6439 VDD.n5065 VDD.n5051 92.5005
R6440 VDD.n5508 VDD.n5507 92.5005
R6441 VDD.n5509 VDD.n5508 92.5005
R6442 VDD.n5505 VDD.n5066 92.5005
R6443 VDD.n5069 VDD.n5066 92.5005
R6444 VDD.n5082 VDD.n5067 92.5005
R6445 VDD.n5082 VDD.n5070 92.5005
R6446 VDD.n5491 VDD.n5490 92.5005
R6447 VDD.n5490 VDD.n5489 92.5005
R6448 VDD.n5155 VDD.n5084 92.5005
R6449 VDD.n5152 VDD.n5084 92.5005
R6450 VDD.n5482 VDD.n5481 92.5005
R6451 VDD.n5483 VDD.n5482 92.5005
R6452 VDD.n5166 VDD.n5154 92.5005
R6453 VDD.n5168 VDD.n5154 92.5005
R6454 VDD.n5445 VDD.n5438 92.5005
R6455 VDD.n5445 VDD.n5444 92.5005
R6456 VDD.n5447 VDD.n5446 92.5005
R6457 VDD.n5446 VDD.n5191 92.5005
R6458 VDD.n5701 VDD.n5700 92.5005
R6459 VDD.n5700 VDD.n5699 92.5005
R6460 VDD.n5506 VDD.n5061 92.5005
R6461 VDD.n5063 VDD.n5061 92.5005
R6462 VDD.n5504 VDD.n5503 92.5005
R6463 VDD.n5503 VDD.n5502 92.5005
R6464 VDD.n5079 VDD.n5068 92.5005
R6465 VDD.n5076 VDD.n5068 92.5005
R6466 VDD.n5495 VDD.n5494 92.5005
R6467 VDD.n5496 VDD.n5495 92.5005
R6468 VDD.n5492 VDD.n5078 92.5005
R6469 VDD.n5085 VDD.n5078 92.5005
R6470 VDD.n5480 VDD.n5479 92.5005
R6471 VDD.n5479 VDD.n5153 92.5005
R6472 VDD.n5478 VDD.n5167 92.5005
R6473 VDD.n5478 VDD.n5477 92.5005
R6474 VDD.n5437 VDD.n5165 92.5005
R6475 VDD.n5439 VDD.n5165 92.5005
R6476 VDD.n5470 VDD.n5469 92.5005
R6477 VDD.n5471 VDD.n5470 92.5005
R6478 VDD.n5468 VDD.n5436 92.5005
R6479 VDD.n5450 VDD.n5436 92.5005
R6480 VDD.n5435 VDD.n4926 92.5005
R6481 VDD.n5435 VDD.n4929 92.5005
R6482 VDD.n5511 VDD.n5062 92.5005
R6483 VDD.n5511 VDD.n5510 92.5005
R6484 VDD.n4263 VDD.n4260 92.5005
R6485 VDD.n4724 VDD.n4263 92.5005
R6486 VDD.n4618 VDD.n4617 92.5005
R6487 VDD.n4618 VDD.n4143 92.5005
R6488 VDD.n4404 VDD.n4403 92.5005
R6489 VDD.n4664 VDD.n4404 92.5005
R6490 VDD.n4687 VDD.n4686 92.5005
R6491 VDD.n4686 VDD.n4685 92.5005
R6492 VDD.n4688 VDD.n4384 92.5005
R6493 VDD.n4653 VDD.n4384 92.5005
R6494 VDD.n4690 VDD.n4689 92.5005
R6495 VDD.n4691 VDD.n4690 92.5005
R6496 VDD.n4402 VDD.n4383 92.5005
R6497 VDD.n4383 VDD.n4367 92.5005
R6498 VDD.n4397 VDD.n4385 92.5005
R6499 VDD.n4396 VDD.n4395 92.5005
R6500 VDD.n4394 VDD.n4393 92.5005
R6501 VDD.n4392 VDD.n4388 92.5005
R6502 VDD.n4390 VDD.n4389 92.5005
R6503 VDD.n4400 VDD.n4399 92.5005
R6504 VDD.n4289 VDD.n4288 92.5005
R6505 VDD.n4299 VDD.n4289 92.5005
R6506 VDD.n4712 VDD.n4711 92.5005
R6507 VDD.n4711 VDD.n4710 92.5005
R6508 VDD.n4713 VDD.n4286 92.5005
R6509 VDD.n4290 VDD.n4286 92.5005
R6510 VDD.n4715 VDD.n4714 92.5005
R6511 VDD.n4716 VDD.n4715 92.5005
R6512 VDD.n4287 VDD.n4285 92.5005
R6513 VDD.n4285 VDD.n4277 92.5005
R6514 VDD.n4755 VDD.n4236 92.5005
R6515 VDD.n4236 VDD.n4235 92.5005
R6516 VDD.n4778 VDD.n4777 92.5005
R6517 VDD.n4777 VDD.n4776 92.5005
R6518 VDD.n4226 VDD.n4225 92.5005
R6519 VDD.n4775 VDD.n4226 92.5005
R6520 VDD.n4773 VDD.n4772 92.5005
R6521 VDD.n4774 VDD.n4773 92.5005
R6522 VDD.n4771 VDD.n4228 92.5005
R6523 VDD.n4228 VDD.n4227 92.5005
R6524 VDD.n4770 VDD.n4769 92.5005
R6525 VDD.n4769 VDD.n4768 92.5005
R6526 VDD.n4230 VDD.n4229 92.5005
R6527 VDD.n4767 VDD.n4230 92.5005
R6528 VDD.n4765 VDD.n4764 92.5005
R6529 VDD.n4766 VDD.n4765 92.5005
R6530 VDD.n4763 VDD.n4232 92.5005
R6531 VDD.n4232 VDD.n4231 92.5005
R6532 VDD.n4762 VDD.n4761 92.5005
R6533 VDD.n4761 VDD.n4760 92.5005
R6534 VDD.n4234 VDD.n4233 92.5005
R6535 VDD.n4759 VDD.n4234 92.5005
R6536 VDD.n4757 VDD.n4756 92.5005
R6537 VDD.n4758 VDD.n4757 92.5005
R6538 VDD.n4779 VDD.n4223 92.5005
R6539 VDD.n4223 VDD.n4222 92.5005
R6540 VDD.n4782 VDD.n4781 92.5005
R6541 VDD.n4783 VDD.n4782 92.5005
R6542 VDD.n4780 VDD.n4224 92.5005
R6543 VDD.n4220 VDD.n4219 92.5005
R6544 VDD.n4787 VDD.n4786 92.5005
R6545 VDD.n4786 VDD.n4785 92.5005
R6546 VDD.n4790 VDD.n4789 92.5005
R6547 VDD.n4791 VDD.n4790 92.5005
R6548 VDD.n4216 VDD.n4215 92.5005
R6549 VDD.n4792 VDD.n4216 92.5005
R6550 VDD.n4795 VDD.n4794 92.5005
R6551 VDD.n4794 VDD.n4793 92.5005
R6552 VDD.n4796 VDD.n4214 92.5005
R6553 VDD.n4214 VDD.n4213 92.5005
R6554 VDD.n4798 VDD.n4797 92.5005
R6555 VDD.n4799 VDD.n4798 92.5005
R6556 VDD.n4212 VDD.n4211 92.5005
R6557 VDD.n4800 VDD.n4212 92.5005
R6558 VDD.n4803 VDD.n4802 92.5005
R6559 VDD.n4802 VDD.n4801 92.5005
R6560 VDD.n4804 VDD.n4210 92.5005
R6561 VDD.n4210 VDD.n4209 92.5005
R6562 VDD.n4806 VDD.n4805 92.5005
R6563 VDD.n4807 VDD.n4806 92.5005
R6564 VDD.n4208 VDD.n4207 92.5005
R6565 VDD.n4808 VDD.n4208 92.5005
R6566 VDD.n4811 VDD.n4810 92.5005
R6567 VDD.n4810 VDD.n4809 92.5005
R6568 VDD.n4812 VDD.n4206 92.5005
R6569 VDD.n4206 VDD.n4205 92.5005
R6570 VDD.n4814 VDD.n4813 92.5005
R6571 VDD.n4815 VDD.n4814 92.5005
R6572 VDD.n4204 VDD.n4203 92.5005
R6573 VDD.n4816 VDD.n4204 92.5005
R6574 VDD.n4819 VDD.n4818 92.5005
R6575 VDD.n4818 VDD.n4817 92.5005
R6576 VDD.n4820 VDD.n4202 92.5005
R6577 VDD.n4202 VDD.n4201 92.5005
R6578 VDD.n4822 VDD.n4821 92.5005
R6579 VDD.n4823 VDD.n4822 92.5005
R6580 VDD.n4200 VDD.n4199 92.5005
R6581 VDD.n4824 VDD.n4200 92.5005
R6582 VDD.n4827 VDD.n4826 92.5005
R6583 VDD.n4826 VDD.n4825 92.5005
R6584 VDD.n4828 VDD.n4198 92.5005
R6585 VDD.n4198 VDD.n4197 92.5005
R6586 VDD.n4830 VDD.n4829 92.5005
R6587 VDD.n4831 VDD.n4830 92.5005
R6588 VDD.n4196 VDD.n4195 92.5005
R6589 VDD.n4832 VDD.n4196 92.5005
R6590 VDD.n4835 VDD.n4834 92.5005
R6591 VDD.n4834 VDD.n4833 92.5005
R6592 VDD.n4836 VDD.n4194 92.5005
R6593 VDD.n4194 VDD.n4193 92.5005
R6594 VDD.n4838 VDD.n4837 92.5005
R6595 VDD.n4839 VDD.n4838 92.5005
R6596 VDD.n4192 VDD.n4191 92.5005
R6597 VDD.n4840 VDD.n4192 92.5005
R6598 VDD.n4843 VDD.n4842 92.5005
R6599 VDD.n4842 VDD.n4841 92.5005
R6600 VDD.n4844 VDD.n4189 92.5005
R6601 VDD.n4189 VDD.n4186 92.5005
R6602 VDD.n4788 VDD.n4218 92.5005
R6603 VDD.n4218 VDD.n4217 92.5005
R6604 VDD.n4181 VDD.n4180 92.5005
R6605 VDD.n4856 VDD.n4181 92.5005
R6606 VDD.n4859 VDD.n4858 92.5005
R6607 VDD.n4858 VDD.n4857 92.5005
R6608 VDD.n4860 VDD.n4179 92.5005
R6609 VDD.n4179 VDD.n4178 92.5005
R6610 VDD.n4862 VDD.n4861 92.5005
R6611 VDD.n4863 VDD.n4862 92.5005
R6612 VDD.n4177 VDD.n4176 92.5005
R6613 VDD.n4864 VDD.n4177 92.5005
R6614 VDD.n4867 VDD.n4866 92.5005
R6615 VDD.n4866 VDD.n4865 92.5005
R6616 VDD.n4868 VDD.n4175 92.5005
R6617 VDD.n4175 VDD.n4174 92.5005
R6618 VDD.n4870 VDD.n4869 92.5005
R6619 VDD.n4871 VDD.n4870 92.5005
R6620 VDD.n4172 VDD.n4171 92.5005
R6621 VDD.n4872 VDD.n4172 92.5005
R6622 VDD.n4875 VDD.n4874 92.5005
R6623 VDD.n4874 VDD.n4873 92.5005
R6624 VDD.n4876 VDD.n4170 92.5005
R6625 VDD.n4173 VDD.n4170 92.5005
R6626 VDD.n4852 VDD.n4183 92.5005
R6627 VDD.n4183 VDD.n4182 92.5005
R6628 VDD.n4851 VDD.n4850 92.5005
R6629 VDD.n4850 VDD.n4849 92.5005
R6630 VDD.n4185 VDD.n4184 92.5005
R6631 VDD.n4190 VDD.n4188 92.5005
R6632 VDD.n4846 VDD.n4845 92.5005
R6633 VDD.n4847 VDD.n4846 92.5005
R6634 VDD.n4854 VDD.n4853 92.5005
R6635 VDD.n4855 VDD.n4854 92.5005
R6636 VDD.n4879 VDD.n4878 92.5005
R6637 VDD.n4900 VDD.n4154 92.5005
R6638 VDD.n4899 VDD.n4898 92.5005
R6639 VDD.n4163 VDD.n4159 92.5005
R6640 VDD.n4893 VDD.n4892 92.5005
R6641 VDD.n4890 VDD.n4889 92.5005
R6642 VDD.n4165 VDD.n4164 92.5005
R6643 VDD.n4883 VDD.n4882 92.5005
R6644 VDD.n4881 VDD.n4168 92.5005
R6645 VDD.n4903 VDD.n4902 92.5005
R6646 VDD.n4640 VDD.n4139 92.5005
R6647 VDD.n4642 VDD.n4138 92.5005
R6648 VDD.n4414 VDD.n4413 92.5005
R6649 VDD.n4624 VDD.n4623 92.5005
R6650 VDD.n4628 VDD.n4627 92.5005
R6651 VDD.n4626 VDD.n4410 92.5005
R6652 VDD.n4637 VDD.n4636 92.5005
R6653 VDD.n4638 VDD.n4407 92.5005
R6654 VDD.n4635 VDD.n4406 92.5005
R6655 VDD.n4634 VDD.n4633 92.5005
R6656 VDD.n4630 VDD.n4629 92.5005
R6657 VDD.n4619 VDD.n4412 92.5005
R6658 VDD.n4622 VDD.n4621 92.5005
R6659 VDD.n4612 VDD.n4415 92.5005
R6660 VDD.n4615 VDD.n4614 92.5005
R6661 VDD.n4648 VDD.n4647 92.5005
R6662 VDD.n4648 VDD.n4144 92.5005
R6663 VDD.n4646 VDD.n4645 92.5005
R6664 VDD.n4644 VDD.n4408 92.5005
R6665 VDD.n4572 VDD.n4431 92.5005
R6666 VDD.n4574 VDD.n4573 92.5005
R6667 VDD.n4576 VDD.n4575 92.5005
R6668 VDD.n4577 VDD.n4433 92.5005
R6669 VDD.n4579 VDD.n4578 92.5005
R6670 VDD.n4430 VDD.n4429 92.5005
R6671 VDD.n4583 VDD.n4430 92.5005
R6672 VDD.n4586 VDD.n4585 92.5005
R6673 VDD.n4585 VDD.n4584 92.5005
R6674 VDD.n4587 VDD.n4428 92.5005
R6675 VDD.n4428 VDD.n4427 92.5005
R6676 VDD.n4589 VDD.n4588 92.5005
R6677 VDD.n4590 VDD.n4589 92.5005
R6678 VDD.n4426 VDD.n4425 92.5005
R6679 VDD.n4591 VDD.n4426 92.5005
R6680 VDD.n4594 VDD.n4593 92.5005
R6681 VDD.n4593 VDD.n4592 92.5005
R6682 VDD.n4595 VDD.n4424 92.5005
R6683 VDD.n4424 VDD.n4423 92.5005
R6684 VDD.n4597 VDD.n4596 92.5005
R6685 VDD.n4598 VDD.n4597 92.5005
R6686 VDD.n4422 VDD.n4421 92.5005
R6687 VDD.n4599 VDD.n4422 92.5005
R6688 VDD.n4602 VDD.n4601 92.5005
R6689 VDD.n4601 VDD.n4600 92.5005
R6690 VDD.n4603 VDD.n4420 92.5005
R6691 VDD.n4420 VDD.n4419 92.5005
R6692 VDD.n4606 VDD.n4605 92.5005
R6693 VDD.n4607 VDD.n4606 92.5005
R6694 VDD.n4604 VDD.n4417 92.5005
R6695 VDD.n4608 VDD.n4417 92.5005
R6696 VDD.n4611 VDD.n4418 92.5005
R6697 VDD.n4611 VDD.n4610 92.5005
R6698 VDD.n4460 VDD.n4459 92.5005
R6699 VDD.n4520 VDD.n4460 92.5005
R6700 VDD.n4523 VDD.n4522 92.5005
R6701 VDD.n4522 VDD.n4521 92.5005
R6702 VDD.n4524 VDD.n4458 92.5005
R6703 VDD.n4458 VDD.n4457 92.5005
R6704 VDD.n4526 VDD.n4525 92.5005
R6705 VDD.n4527 VDD.n4526 92.5005
R6706 VDD.n4456 VDD.n4455 92.5005
R6707 VDD.n4528 VDD.n4456 92.5005
R6708 VDD.n4531 VDD.n4530 92.5005
R6709 VDD.n4530 VDD.n4529 92.5005
R6710 VDD.n4532 VDD.n4454 92.5005
R6711 VDD.n4454 VDD.n4453 92.5005
R6712 VDD.n4534 VDD.n4533 92.5005
R6713 VDD.n4535 VDD.n4534 92.5005
R6714 VDD.n4452 VDD.n4451 92.5005
R6715 VDD.n4536 VDD.n4452 92.5005
R6716 VDD.n4539 VDD.n4538 92.5005
R6717 VDD.n4538 VDD.n4537 92.5005
R6718 VDD.n4540 VDD.n4450 92.5005
R6719 VDD.n4450 VDD.n4449 92.5005
R6720 VDD.n4542 VDD.n4541 92.5005
R6721 VDD.n4543 VDD.n4542 92.5005
R6722 VDD.n4448 VDD.n4447 92.5005
R6723 VDD.n4544 VDD.n4448 92.5005
R6724 VDD.n4547 VDD.n4546 92.5005
R6725 VDD.n4546 VDD.n4545 92.5005
R6726 VDD.n4548 VDD.n4446 92.5005
R6727 VDD.n4446 VDD.n4445 92.5005
R6728 VDD.n4550 VDD.n4549 92.5005
R6729 VDD.n4551 VDD.n4550 92.5005
R6730 VDD.n4444 VDD.n4443 92.5005
R6731 VDD.n4552 VDD.n4444 92.5005
R6732 VDD.n4555 VDD.n4554 92.5005
R6733 VDD.n4554 VDD.n4553 92.5005
R6734 VDD.n4556 VDD.n4442 92.5005
R6735 VDD.n4442 VDD.n4441 92.5005
R6736 VDD.n4558 VDD.n4557 92.5005
R6737 VDD.n4559 VDD.n4558 92.5005
R6738 VDD.n4440 VDD.n4439 92.5005
R6739 VDD.n4560 VDD.n4440 92.5005
R6740 VDD.n4563 VDD.n4562 92.5005
R6741 VDD.n4562 VDD.n4561 92.5005
R6742 VDD.n4564 VDD.n4438 92.5005
R6743 VDD.n4438 VDD.n4437 92.5005
R6744 VDD.n4567 VDD.n4566 92.5005
R6745 VDD.n4568 VDD.n4567 92.5005
R6746 VDD.n4565 VDD.n4435 92.5005
R6747 VDD.n4569 VDD.n4435 92.5005
R6748 VDD.n4571 VDD.n4436 92.5005
R6749 VDD.n4571 VDD.n4570 92.5005
R6750 VDD.n4515 VDD.n4514 92.5005
R6751 VDD.n4462 VDD.n4461 92.5005
R6752 VDD.n4519 VDD.n4518 92.5005
R6753 VDD.n4259 VDD.n4258 92.5005
R6754 VDD.n4481 VDD.n4258 92.5005
R6755 VDD.n4484 VDD.n4483 92.5005
R6756 VDD.n4483 VDD.n4482 92.5005
R6757 VDD.n4486 VDD.n4485 92.5005
R6758 VDD.n4487 VDD.n4486 92.5005
R6759 VDD.n4480 VDD.n4479 92.5005
R6760 VDD.n4488 VDD.n4480 92.5005
R6761 VDD.n4491 VDD.n4490 92.5005
R6762 VDD.n4490 VDD.n4489 92.5005
R6763 VDD.n4492 VDD.n4478 92.5005
R6764 VDD.n4478 VDD.n4477 92.5005
R6765 VDD.n4494 VDD.n4493 92.5005
R6766 VDD.n4495 VDD.n4494 92.5005
R6767 VDD.n4476 VDD.n4475 92.5005
R6768 VDD.n4496 VDD.n4476 92.5005
R6769 VDD.n4499 VDD.n4498 92.5005
R6770 VDD.n4498 VDD.n4497 92.5005
R6771 VDD.n4500 VDD.n4474 92.5005
R6772 VDD.n4474 VDD.n4473 92.5005
R6773 VDD.n4502 VDD.n4501 92.5005
R6774 VDD.n4503 VDD.n4502 92.5005
R6775 VDD.n4471 VDD.n4470 92.5005
R6776 VDD.n4504 VDD.n4471 92.5005
R6777 VDD.n4507 VDD.n4506 92.5005
R6778 VDD.n4506 VDD.n4505 92.5005
R6779 VDD.n4508 VDD.n4468 92.5005
R6780 VDD.n4472 VDD.n4468 92.5005
R6781 VDD.n4510 VDD.n4509 92.5005
R6782 VDD.n4469 VDD.n4467 92.5005
R6783 VDD.n4464 VDD.n4463 92.5005
R6784 VDD.n4754 VDD.n4753 92.5005
R6785 VDD.n4335 VDD.n4238 92.5005
R6786 VDD.n4337 VDD.n4336 92.5005
R6787 VDD.n4334 VDD.n4333 92.5005
R6788 VDD.n4304 VDD.n4303 92.5005
R6789 VDD.n4328 VDD.n4327 92.5005
R6790 VDD.n4306 VDD.n4305 92.5005
R6791 VDD.n4322 VDD.n4321 92.5005
R6792 VDD.n4318 VDD.n4317 92.5005
R6793 VDD.n4316 VDD.n4315 92.5005
R6794 VDD.n4729 VDD.n4728 92.5005
R6795 VDD.n4733 VDD.n4732 92.5005
R6796 VDD.n4736 VDD.n4735 92.5005
R6797 VDD.n4273 VDD.n4272 92.5005
R6798 VDD.n4262 VDD.n4261 92.5005
R6799 VDD.n4745 VDD.n4744 92.5005
R6800 VDD.n4746 VDD.n4257 92.5005
R6801 VDD.n4749 VDD.n4748 92.5005
R6802 VDD.n4743 VDD.n4742 92.5005
R6803 VDD.n4271 VDD.n4264 92.5005
R6804 VDD.n4738 VDD.n4737 92.5005
R6805 VDD.n4734 VDD.n4270 92.5005
R6806 VDD.n4731 VDD.n4730 92.5005
R6807 VDD.n4274 VDD.n4250 92.5005
R6808 VDD.n4751 VDD.n4250 92.5005
R6809 VDD.n4727 VDD.n4726 92.5005
R6810 VDD.n4310 VDD.n4309 92.5005
R6811 VDD.n4312 VDD.n4311 92.5005
R6812 VDD.n4314 VDD.n4313 92.5005
R6813 VDD.n4320 VDD.n4319 92.5005
R6814 VDD.n4339 VDD.n4338 92.5005
R6815 VDD.n4332 VDD.n4331 92.5005
R6816 VDD.n4330 VDD.n4329 92.5005
R6817 VDD.n4326 VDD.n4325 92.5005
R6818 VDD.n4324 VDD.n4323 92.5005
R6819 VDD.n4150 VDD.n4142 92.5005
R6820 VDD.n4907 VDD.n4906 92.5005
R6821 VDD.n4905 VDD.n4904 92.5005
R6822 VDD.n4905 VDD.n4151 92.5005
R6823 VDD.n4897 VDD.n4896 92.5005
R6824 VDD.n4895 VDD.n4894 92.5005
R6825 VDD.n4166 VDD.n4162 92.5005
R6826 VDD.n4888 VDD.n4887 92.5005
R6827 VDD.n4885 VDD.n4884 92.5005
R6828 VDD.n4158 VDD.n4153 92.5005
R6829 VDD.n4669 VDD.n4668 92.5005
R6830 VDD.n4671 VDD.n4670 92.5005
R6831 VDD.n4673 VDD.n4672 92.5005
R6832 VDD.n4675 VDD.n4674 92.5005
R6833 VDD.n4663 VDD.n4662 92.5005
R6834 VDD.n4680 VDD.n4679 92.5005
R6835 VDD.n4149 VDD.n4148 92.5005
R6836 VDD.n4151 VDD.n4149 92.5005
R6837 VDD.n4909 VDD.n4908 92.5005
R6838 VDD.n4908 VDD.n4907 92.5005
R6839 VDD.n4910 VDD.n4146 92.5005
R6840 VDD.n4150 VDD.n4146 92.5005
R6841 VDD.n4912 VDD.n4911 92.5005
R6842 VDD.n4913 VDD.n4912 92.5005
R6843 VDD.n4655 VDD.n4654 92.5005
R6844 VDD.n4654 VDD.n4405 92.5005
R6845 VDD.n4657 VDD.n4656 92.5005
R6846 VDD.n4658 VDD.n4657 92.5005
R6847 VDD.n4365 VDD.n4364 92.5005
R6848 VDD.n4382 VDD.n4365 92.5005
R6849 VDD.n4699 VDD.n4698 92.5005
R6850 VDD.n4698 VDD.n4697 92.5005
R6851 VDD.n4700 VDD.n4302 92.5005
R6852 VDD.n4366 VDD.n4302 92.5005
R6853 VDD.n4702 VDD.n4701 92.5005
R6854 VDD.n4703 VDD.n4702 92.5005
R6855 VDD.n4346 VDD.n4345 92.5005
R6856 VDD.n4345 VDD.n4284 92.5005
R6857 VDD.n4344 VDD.n4343 92.5005
R6858 VDD.n4344 VDD.n4283 92.5005
R6859 VDD.n4342 VDD.n4278 92.5005
R6860 VDD.n4723 VDD.n4278 92.5005
R6861 VDD.n4341 VDD.n4340 92.5005
R6862 VDD.n4340 VDD.n4265 92.5005
R6863 VDD.n4362 VDD.n4361 92.5005
R6864 VDD.n4359 VDD.n4347 92.5005
R6865 VDD.n4357 VDD.n4356 92.5005
R6866 VDD.n4355 VDD.n4354 92.5005
R6867 VDD.n4352 VDD.n4349 92.5005
R6868 VDD.n4350 VDD.n4294 92.5005
R6869 VDD.n4307 VDD.n4279 92.5005
R6870 VDD.n4279 VDD.n4265 92.5005
R6871 VDD.n4722 VDD.n4721 92.5005
R6872 VDD.n4723 VDD.n4722 92.5005
R6873 VDD.n4719 VDD.n4280 92.5005
R6874 VDD.n4283 VDD.n4280 92.5005
R6875 VDD.n4296 VDD.n4281 92.5005
R6876 VDD.n4296 VDD.n4284 92.5005
R6877 VDD.n4705 VDD.n4704 92.5005
R6878 VDD.n4704 VDD.n4703 92.5005
R6879 VDD.n4369 VDD.n4298 92.5005
R6880 VDD.n4366 VDD.n4298 92.5005
R6881 VDD.n4696 VDD.n4695 92.5005
R6882 VDD.n4697 VDD.n4696 92.5005
R6883 VDD.n4380 VDD.n4368 92.5005
R6884 VDD.n4382 VDD.n4368 92.5005
R6885 VDD.n4659 VDD.n4652 92.5005
R6886 VDD.n4659 VDD.n4658 92.5005
R6887 VDD.n4661 VDD.n4660 92.5005
R6888 VDD.n4660 VDD.n4405 92.5005
R6889 VDD.n4915 VDD.n4914 92.5005
R6890 VDD.n4914 VDD.n4913 92.5005
R6891 VDD.n4720 VDD.n4275 92.5005
R6892 VDD.n4277 VDD.n4275 92.5005
R6893 VDD.n4718 VDD.n4717 92.5005
R6894 VDD.n4717 VDD.n4716 92.5005
R6895 VDD.n4293 VDD.n4282 92.5005
R6896 VDD.n4290 VDD.n4282 92.5005
R6897 VDD.n4709 VDD.n4708 92.5005
R6898 VDD.n4710 VDD.n4709 92.5005
R6899 VDD.n4706 VDD.n4292 92.5005
R6900 VDD.n4299 VDD.n4292 92.5005
R6901 VDD.n4694 VDD.n4693 92.5005
R6902 VDD.n4693 VDD.n4367 92.5005
R6903 VDD.n4692 VDD.n4381 92.5005
R6904 VDD.n4692 VDD.n4691 92.5005
R6905 VDD.n4651 VDD.n4379 92.5005
R6906 VDD.n4653 VDD.n4379 92.5005
R6907 VDD.n4684 VDD.n4683 92.5005
R6908 VDD.n4685 VDD.n4684 92.5005
R6909 VDD.n4682 VDD.n4650 92.5005
R6910 VDD.n4664 VDD.n4650 92.5005
R6911 VDD.n4649 VDD.n4140 92.5005
R6912 VDD.n4649 VDD.n4143 92.5005
R6913 VDD.n4725 VDD.n4276 92.5005
R6914 VDD.n4725 VDD.n4724 92.5005
R6915 VDD.n3409 VDD.n3406 92.5005
R6916 VDD.n3870 VDD.n3409 92.5005
R6917 VDD.n3764 VDD.n3763 92.5005
R6918 VDD.n3764 VDD.n3289 92.5005
R6919 VDD.n3550 VDD.n3549 92.5005
R6920 VDD.n3810 VDD.n3550 92.5005
R6921 VDD.n3833 VDD.n3832 92.5005
R6922 VDD.n3832 VDD.n3831 92.5005
R6923 VDD.n3834 VDD.n3530 92.5005
R6924 VDD.n3799 VDD.n3530 92.5005
R6925 VDD.n3836 VDD.n3835 92.5005
R6926 VDD.n3837 VDD.n3836 92.5005
R6927 VDD.n3548 VDD.n3529 92.5005
R6928 VDD.n3529 VDD.n3513 92.5005
R6929 VDD.n3543 VDD.n3531 92.5005
R6930 VDD.n3542 VDD.n3541 92.5005
R6931 VDD.n3540 VDD.n3539 92.5005
R6932 VDD.n3538 VDD.n3534 92.5005
R6933 VDD.n3536 VDD.n3535 92.5005
R6934 VDD.n3546 VDD.n3545 92.5005
R6935 VDD.n3435 VDD.n3434 92.5005
R6936 VDD.n3445 VDD.n3435 92.5005
R6937 VDD.n3858 VDD.n3857 92.5005
R6938 VDD.n3857 VDD.n3856 92.5005
R6939 VDD.n3859 VDD.n3432 92.5005
R6940 VDD.n3436 VDD.n3432 92.5005
R6941 VDD.n3861 VDD.n3860 92.5005
R6942 VDD.n3862 VDD.n3861 92.5005
R6943 VDD.n3433 VDD.n3431 92.5005
R6944 VDD.n3431 VDD.n3423 92.5005
R6945 VDD.n3901 VDD.n3382 92.5005
R6946 VDD.n3382 VDD.n3381 92.5005
R6947 VDD.n3924 VDD.n3923 92.5005
R6948 VDD.n3923 VDD.n3922 92.5005
R6949 VDD.n3372 VDD.n3371 92.5005
R6950 VDD.n3921 VDD.n3372 92.5005
R6951 VDD.n3919 VDD.n3918 92.5005
R6952 VDD.n3920 VDD.n3919 92.5005
R6953 VDD.n3917 VDD.n3374 92.5005
R6954 VDD.n3374 VDD.n3373 92.5005
R6955 VDD.n3916 VDD.n3915 92.5005
R6956 VDD.n3915 VDD.n3914 92.5005
R6957 VDD.n3376 VDD.n3375 92.5005
R6958 VDD.n3913 VDD.n3376 92.5005
R6959 VDD.n3911 VDD.n3910 92.5005
R6960 VDD.n3912 VDD.n3911 92.5005
R6961 VDD.n3909 VDD.n3378 92.5005
R6962 VDD.n3378 VDD.n3377 92.5005
R6963 VDD.n3908 VDD.n3907 92.5005
R6964 VDD.n3907 VDD.n3906 92.5005
R6965 VDD.n3380 VDD.n3379 92.5005
R6966 VDD.n3905 VDD.n3380 92.5005
R6967 VDD.n3903 VDD.n3902 92.5005
R6968 VDD.n3904 VDD.n3903 92.5005
R6969 VDD.n3925 VDD.n3369 92.5005
R6970 VDD.n3369 VDD.n3368 92.5005
R6971 VDD.n3928 VDD.n3927 92.5005
R6972 VDD.n3929 VDD.n3928 92.5005
R6973 VDD.n3926 VDD.n3370 92.5005
R6974 VDD.n3366 VDD.n3365 92.5005
R6975 VDD.n3933 VDD.n3932 92.5005
R6976 VDD.n3932 VDD.n3931 92.5005
R6977 VDD.n3936 VDD.n3935 92.5005
R6978 VDD.n3937 VDD.n3936 92.5005
R6979 VDD.n3362 VDD.n3361 92.5005
R6980 VDD.n3938 VDD.n3362 92.5005
R6981 VDD.n3941 VDD.n3940 92.5005
R6982 VDD.n3940 VDD.n3939 92.5005
R6983 VDD.n3942 VDD.n3360 92.5005
R6984 VDD.n3360 VDD.n3359 92.5005
R6985 VDD.n3944 VDD.n3943 92.5005
R6986 VDD.n3945 VDD.n3944 92.5005
R6987 VDD.n3358 VDD.n3357 92.5005
R6988 VDD.n3946 VDD.n3358 92.5005
R6989 VDD.n3949 VDD.n3948 92.5005
R6990 VDD.n3948 VDD.n3947 92.5005
R6991 VDD.n3950 VDD.n3356 92.5005
R6992 VDD.n3356 VDD.n3355 92.5005
R6993 VDD.n3952 VDD.n3951 92.5005
R6994 VDD.n3953 VDD.n3952 92.5005
R6995 VDD.n3354 VDD.n3353 92.5005
R6996 VDD.n3954 VDD.n3354 92.5005
R6997 VDD.n3957 VDD.n3956 92.5005
R6998 VDD.n3956 VDD.n3955 92.5005
R6999 VDD.n3958 VDD.n3352 92.5005
R7000 VDD.n3352 VDD.n3351 92.5005
R7001 VDD.n3960 VDD.n3959 92.5005
R7002 VDD.n3961 VDD.n3960 92.5005
R7003 VDD.n3350 VDD.n3349 92.5005
R7004 VDD.n3962 VDD.n3350 92.5005
R7005 VDD.n3965 VDD.n3964 92.5005
R7006 VDD.n3964 VDD.n3963 92.5005
R7007 VDD.n3966 VDD.n3348 92.5005
R7008 VDD.n3348 VDD.n3347 92.5005
R7009 VDD.n3968 VDD.n3967 92.5005
R7010 VDD.n3969 VDD.n3968 92.5005
R7011 VDD.n3346 VDD.n3345 92.5005
R7012 VDD.n3970 VDD.n3346 92.5005
R7013 VDD.n3973 VDD.n3972 92.5005
R7014 VDD.n3972 VDD.n3971 92.5005
R7015 VDD.n3974 VDD.n3344 92.5005
R7016 VDD.n3344 VDD.n3343 92.5005
R7017 VDD.n3976 VDD.n3975 92.5005
R7018 VDD.n3977 VDD.n3976 92.5005
R7019 VDD.n3342 VDD.n3341 92.5005
R7020 VDD.n3978 VDD.n3342 92.5005
R7021 VDD.n3981 VDD.n3980 92.5005
R7022 VDD.n3980 VDD.n3979 92.5005
R7023 VDD.n3982 VDD.n3340 92.5005
R7024 VDD.n3340 VDD.n3339 92.5005
R7025 VDD.n3984 VDD.n3983 92.5005
R7026 VDD.n3985 VDD.n3984 92.5005
R7027 VDD.n3338 VDD.n3337 92.5005
R7028 VDD.n3986 VDD.n3338 92.5005
R7029 VDD.n3989 VDD.n3988 92.5005
R7030 VDD.n3988 VDD.n3987 92.5005
R7031 VDD.n3990 VDD.n3335 92.5005
R7032 VDD.n3335 VDD.n3332 92.5005
R7033 VDD.n3934 VDD.n3364 92.5005
R7034 VDD.n3364 VDD.n3363 92.5005
R7035 VDD.n3327 VDD.n3326 92.5005
R7036 VDD.n4002 VDD.n3327 92.5005
R7037 VDD.n4005 VDD.n4004 92.5005
R7038 VDD.n4004 VDD.n4003 92.5005
R7039 VDD.n4006 VDD.n3325 92.5005
R7040 VDD.n3325 VDD.n3324 92.5005
R7041 VDD.n4008 VDD.n4007 92.5005
R7042 VDD.n4009 VDD.n4008 92.5005
R7043 VDD.n3323 VDD.n3322 92.5005
R7044 VDD.n4010 VDD.n3323 92.5005
R7045 VDD.n4013 VDD.n4012 92.5005
R7046 VDD.n4012 VDD.n4011 92.5005
R7047 VDD.n4014 VDD.n3321 92.5005
R7048 VDD.n3321 VDD.n3320 92.5005
R7049 VDD.n4016 VDD.n4015 92.5005
R7050 VDD.n4017 VDD.n4016 92.5005
R7051 VDD.n3318 VDD.n3317 92.5005
R7052 VDD.n4018 VDD.n3318 92.5005
R7053 VDD.n4021 VDD.n4020 92.5005
R7054 VDD.n4020 VDD.n4019 92.5005
R7055 VDD.n4022 VDD.n3316 92.5005
R7056 VDD.n3319 VDD.n3316 92.5005
R7057 VDD.n3998 VDD.n3329 92.5005
R7058 VDD.n3329 VDD.n3328 92.5005
R7059 VDD.n3997 VDD.n3996 92.5005
R7060 VDD.n3996 VDD.n3995 92.5005
R7061 VDD.n3331 VDD.n3330 92.5005
R7062 VDD.n3336 VDD.n3334 92.5005
R7063 VDD.n3992 VDD.n3991 92.5005
R7064 VDD.n3993 VDD.n3992 92.5005
R7065 VDD.n4000 VDD.n3999 92.5005
R7066 VDD.n4001 VDD.n4000 92.5005
R7067 VDD.n4025 VDD.n4024 92.5005
R7068 VDD.n4046 VDD.n3300 92.5005
R7069 VDD.n4045 VDD.n4044 92.5005
R7070 VDD.n3309 VDD.n3305 92.5005
R7071 VDD.n4039 VDD.n4038 92.5005
R7072 VDD.n4036 VDD.n4035 92.5005
R7073 VDD.n3311 VDD.n3310 92.5005
R7074 VDD.n4029 VDD.n4028 92.5005
R7075 VDD.n4027 VDD.n3314 92.5005
R7076 VDD.n4049 VDD.n4048 92.5005
R7077 VDD.n3786 VDD.n3285 92.5005
R7078 VDD.n3788 VDD.n3284 92.5005
R7079 VDD.n3560 VDD.n3559 92.5005
R7080 VDD.n3770 VDD.n3769 92.5005
R7081 VDD.n3774 VDD.n3773 92.5005
R7082 VDD.n3772 VDD.n3556 92.5005
R7083 VDD.n3783 VDD.n3782 92.5005
R7084 VDD.n3784 VDD.n3553 92.5005
R7085 VDD.n3781 VDD.n3552 92.5005
R7086 VDD.n3780 VDD.n3779 92.5005
R7087 VDD.n3776 VDD.n3775 92.5005
R7088 VDD.n3765 VDD.n3558 92.5005
R7089 VDD.n3768 VDD.n3767 92.5005
R7090 VDD.n3758 VDD.n3561 92.5005
R7091 VDD.n3761 VDD.n3760 92.5005
R7092 VDD.n3794 VDD.n3793 92.5005
R7093 VDD.n3794 VDD.n3290 92.5005
R7094 VDD.n3792 VDD.n3791 92.5005
R7095 VDD.n3790 VDD.n3554 92.5005
R7096 VDD.n3718 VDD.n3577 92.5005
R7097 VDD.n3720 VDD.n3719 92.5005
R7098 VDD.n3722 VDD.n3721 92.5005
R7099 VDD.n3723 VDD.n3579 92.5005
R7100 VDD.n3725 VDD.n3724 92.5005
R7101 VDD.n3576 VDD.n3575 92.5005
R7102 VDD.n3729 VDD.n3576 92.5005
R7103 VDD.n3732 VDD.n3731 92.5005
R7104 VDD.n3731 VDD.n3730 92.5005
R7105 VDD.n3733 VDD.n3574 92.5005
R7106 VDD.n3574 VDD.n3573 92.5005
R7107 VDD.n3735 VDD.n3734 92.5005
R7108 VDD.n3736 VDD.n3735 92.5005
R7109 VDD.n3572 VDD.n3571 92.5005
R7110 VDD.n3737 VDD.n3572 92.5005
R7111 VDD.n3740 VDD.n3739 92.5005
R7112 VDD.n3739 VDD.n3738 92.5005
R7113 VDD.n3741 VDD.n3570 92.5005
R7114 VDD.n3570 VDD.n3569 92.5005
R7115 VDD.n3743 VDD.n3742 92.5005
R7116 VDD.n3744 VDD.n3743 92.5005
R7117 VDD.n3568 VDD.n3567 92.5005
R7118 VDD.n3745 VDD.n3568 92.5005
R7119 VDD.n3748 VDD.n3747 92.5005
R7120 VDD.n3747 VDD.n3746 92.5005
R7121 VDD.n3749 VDD.n3566 92.5005
R7122 VDD.n3566 VDD.n3565 92.5005
R7123 VDD.n3752 VDD.n3751 92.5005
R7124 VDD.n3753 VDD.n3752 92.5005
R7125 VDD.n3750 VDD.n3563 92.5005
R7126 VDD.n3754 VDD.n3563 92.5005
R7127 VDD.n3757 VDD.n3564 92.5005
R7128 VDD.n3757 VDD.n3756 92.5005
R7129 VDD.n3606 VDD.n3605 92.5005
R7130 VDD.n3666 VDD.n3606 92.5005
R7131 VDD.n3669 VDD.n3668 92.5005
R7132 VDD.n3668 VDD.n3667 92.5005
R7133 VDD.n3670 VDD.n3604 92.5005
R7134 VDD.n3604 VDD.n3603 92.5005
R7135 VDD.n3672 VDD.n3671 92.5005
R7136 VDD.n3673 VDD.n3672 92.5005
R7137 VDD.n3602 VDD.n3601 92.5005
R7138 VDD.n3674 VDD.n3602 92.5005
R7139 VDD.n3677 VDD.n3676 92.5005
R7140 VDD.n3676 VDD.n3675 92.5005
R7141 VDD.n3678 VDD.n3600 92.5005
R7142 VDD.n3600 VDD.n3599 92.5005
R7143 VDD.n3680 VDD.n3679 92.5005
R7144 VDD.n3681 VDD.n3680 92.5005
R7145 VDD.n3598 VDD.n3597 92.5005
R7146 VDD.n3682 VDD.n3598 92.5005
R7147 VDD.n3685 VDD.n3684 92.5005
R7148 VDD.n3684 VDD.n3683 92.5005
R7149 VDD.n3686 VDD.n3596 92.5005
R7150 VDD.n3596 VDD.n3595 92.5005
R7151 VDD.n3688 VDD.n3687 92.5005
R7152 VDD.n3689 VDD.n3688 92.5005
R7153 VDD.n3594 VDD.n3593 92.5005
R7154 VDD.n3690 VDD.n3594 92.5005
R7155 VDD.n3693 VDD.n3692 92.5005
R7156 VDD.n3692 VDD.n3691 92.5005
R7157 VDD.n3694 VDD.n3592 92.5005
R7158 VDD.n3592 VDD.n3591 92.5005
R7159 VDD.n3696 VDD.n3695 92.5005
R7160 VDD.n3697 VDD.n3696 92.5005
R7161 VDD.n3590 VDD.n3589 92.5005
R7162 VDD.n3698 VDD.n3590 92.5005
R7163 VDD.n3701 VDD.n3700 92.5005
R7164 VDD.n3700 VDD.n3699 92.5005
R7165 VDD.n3702 VDD.n3588 92.5005
R7166 VDD.n3588 VDD.n3587 92.5005
R7167 VDD.n3704 VDD.n3703 92.5005
R7168 VDD.n3705 VDD.n3704 92.5005
R7169 VDD.n3586 VDD.n3585 92.5005
R7170 VDD.n3706 VDD.n3586 92.5005
R7171 VDD.n3709 VDD.n3708 92.5005
R7172 VDD.n3708 VDD.n3707 92.5005
R7173 VDD.n3710 VDD.n3584 92.5005
R7174 VDD.n3584 VDD.n3583 92.5005
R7175 VDD.n3713 VDD.n3712 92.5005
R7176 VDD.n3714 VDD.n3713 92.5005
R7177 VDD.n3711 VDD.n3581 92.5005
R7178 VDD.n3715 VDD.n3581 92.5005
R7179 VDD.n3717 VDD.n3582 92.5005
R7180 VDD.n3717 VDD.n3716 92.5005
R7181 VDD.n3661 VDD.n3660 92.5005
R7182 VDD.n3608 VDD.n3607 92.5005
R7183 VDD.n3665 VDD.n3664 92.5005
R7184 VDD.n3405 VDD.n3404 92.5005
R7185 VDD.n3627 VDD.n3404 92.5005
R7186 VDD.n3630 VDD.n3629 92.5005
R7187 VDD.n3629 VDD.n3628 92.5005
R7188 VDD.n3632 VDD.n3631 92.5005
R7189 VDD.n3633 VDD.n3632 92.5005
R7190 VDD.n3626 VDD.n3625 92.5005
R7191 VDD.n3634 VDD.n3626 92.5005
R7192 VDD.n3637 VDD.n3636 92.5005
R7193 VDD.n3636 VDD.n3635 92.5005
R7194 VDD.n3638 VDD.n3624 92.5005
R7195 VDD.n3624 VDD.n3623 92.5005
R7196 VDD.n3640 VDD.n3639 92.5005
R7197 VDD.n3641 VDD.n3640 92.5005
R7198 VDD.n3622 VDD.n3621 92.5005
R7199 VDD.n3642 VDD.n3622 92.5005
R7200 VDD.n3645 VDD.n3644 92.5005
R7201 VDD.n3644 VDD.n3643 92.5005
R7202 VDD.n3646 VDD.n3620 92.5005
R7203 VDD.n3620 VDD.n3619 92.5005
R7204 VDD.n3648 VDD.n3647 92.5005
R7205 VDD.n3649 VDD.n3648 92.5005
R7206 VDD.n3617 VDD.n3616 92.5005
R7207 VDD.n3650 VDD.n3617 92.5005
R7208 VDD.n3653 VDD.n3652 92.5005
R7209 VDD.n3652 VDD.n3651 92.5005
R7210 VDD.n3654 VDD.n3614 92.5005
R7211 VDD.n3618 VDD.n3614 92.5005
R7212 VDD.n3656 VDD.n3655 92.5005
R7213 VDD.n3615 VDD.n3613 92.5005
R7214 VDD.n3610 VDD.n3609 92.5005
R7215 VDD.n3900 VDD.n3899 92.5005
R7216 VDD.n3481 VDD.n3384 92.5005
R7217 VDD.n3483 VDD.n3482 92.5005
R7218 VDD.n3480 VDD.n3479 92.5005
R7219 VDD.n3450 VDD.n3449 92.5005
R7220 VDD.n3474 VDD.n3473 92.5005
R7221 VDD.n3452 VDD.n3451 92.5005
R7222 VDD.n3468 VDD.n3467 92.5005
R7223 VDD.n3464 VDD.n3463 92.5005
R7224 VDD.n3462 VDD.n3461 92.5005
R7225 VDD.n3875 VDD.n3874 92.5005
R7226 VDD.n3879 VDD.n3878 92.5005
R7227 VDD.n3882 VDD.n3881 92.5005
R7228 VDD.n3419 VDD.n3418 92.5005
R7229 VDD.n3408 VDD.n3407 92.5005
R7230 VDD.n3891 VDD.n3890 92.5005
R7231 VDD.n3892 VDD.n3403 92.5005
R7232 VDD.n3895 VDD.n3894 92.5005
R7233 VDD.n3889 VDD.n3888 92.5005
R7234 VDD.n3417 VDD.n3410 92.5005
R7235 VDD.n3884 VDD.n3883 92.5005
R7236 VDD.n3880 VDD.n3416 92.5005
R7237 VDD.n3877 VDD.n3876 92.5005
R7238 VDD.n3420 VDD.n3396 92.5005
R7239 VDD.n3897 VDD.n3396 92.5005
R7240 VDD.n3873 VDD.n3872 92.5005
R7241 VDD.n3456 VDD.n3455 92.5005
R7242 VDD.n3458 VDD.n3457 92.5005
R7243 VDD.n3460 VDD.n3459 92.5005
R7244 VDD.n3466 VDD.n3465 92.5005
R7245 VDD.n3485 VDD.n3484 92.5005
R7246 VDD.n3478 VDD.n3477 92.5005
R7247 VDD.n3476 VDD.n3475 92.5005
R7248 VDD.n3472 VDD.n3471 92.5005
R7249 VDD.n3470 VDD.n3469 92.5005
R7250 VDD.n3296 VDD.n3288 92.5005
R7251 VDD.n4053 VDD.n4052 92.5005
R7252 VDD.n4051 VDD.n4050 92.5005
R7253 VDD.n4051 VDD.n3297 92.5005
R7254 VDD.n4043 VDD.n4042 92.5005
R7255 VDD.n4041 VDD.n4040 92.5005
R7256 VDD.n3312 VDD.n3308 92.5005
R7257 VDD.n4034 VDD.n4033 92.5005
R7258 VDD.n4031 VDD.n4030 92.5005
R7259 VDD.n3304 VDD.n3299 92.5005
R7260 VDD.n3815 VDD.n3814 92.5005
R7261 VDD.n3817 VDD.n3816 92.5005
R7262 VDD.n3819 VDD.n3818 92.5005
R7263 VDD.n3821 VDD.n3820 92.5005
R7264 VDD.n3809 VDD.n3808 92.5005
R7265 VDD.n3826 VDD.n3825 92.5005
R7266 VDD.n3295 VDD.n3294 92.5005
R7267 VDD.n3297 VDD.n3295 92.5005
R7268 VDD.n4055 VDD.n4054 92.5005
R7269 VDD.n4054 VDD.n4053 92.5005
R7270 VDD.n4056 VDD.n3292 92.5005
R7271 VDD.n3296 VDD.n3292 92.5005
R7272 VDD.n4058 VDD.n4057 92.5005
R7273 VDD.n4059 VDD.n4058 92.5005
R7274 VDD.n3801 VDD.n3800 92.5005
R7275 VDD.n3800 VDD.n3551 92.5005
R7276 VDD.n3803 VDD.n3802 92.5005
R7277 VDD.n3804 VDD.n3803 92.5005
R7278 VDD.n3511 VDD.n3510 92.5005
R7279 VDD.n3528 VDD.n3511 92.5005
R7280 VDD.n3845 VDD.n3844 92.5005
R7281 VDD.n3844 VDD.n3843 92.5005
R7282 VDD.n3846 VDD.n3448 92.5005
R7283 VDD.n3512 VDD.n3448 92.5005
R7284 VDD.n3848 VDD.n3847 92.5005
R7285 VDD.n3849 VDD.n3848 92.5005
R7286 VDD.n3492 VDD.n3491 92.5005
R7287 VDD.n3491 VDD.n3430 92.5005
R7288 VDD.n3490 VDD.n3489 92.5005
R7289 VDD.n3490 VDD.n3429 92.5005
R7290 VDD.n3488 VDD.n3424 92.5005
R7291 VDD.n3869 VDD.n3424 92.5005
R7292 VDD.n3487 VDD.n3486 92.5005
R7293 VDD.n3486 VDD.n3411 92.5005
R7294 VDD.n3508 VDD.n3507 92.5005
R7295 VDD.n3505 VDD.n3493 92.5005
R7296 VDD.n3503 VDD.n3502 92.5005
R7297 VDD.n3501 VDD.n3500 92.5005
R7298 VDD.n3498 VDD.n3495 92.5005
R7299 VDD.n3496 VDD.n3440 92.5005
R7300 VDD.n3453 VDD.n3425 92.5005
R7301 VDD.n3425 VDD.n3411 92.5005
R7302 VDD.n3868 VDD.n3867 92.5005
R7303 VDD.n3869 VDD.n3868 92.5005
R7304 VDD.n3865 VDD.n3426 92.5005
R7305 VDD.n3429 VDD.n3426 92.5005
R7306 VDD.n3442 VDD.n3427 92.5005
R7307 VDD.n3442 VDD.n3430 92.5005
R7308 VDD.n3851 VDD.n3850 92.5005
R7309 VDD.n3850 VDD.n3849 92.5005
R7310 VDD.n3515 VDD.n3444 92.5005
R7311 VDD.n3512 VDD.n3444 92.5005
R7312 VDD.n3842 VDD.n3841 92.5005
R7313 VDD.n3843 VDD.n3842 92.5005
R7314 VDD.n3526 VDD.n3514 92.5005
R7315 VDD.n3528 VDD.n3514 92.5005
R7316 VDD.n3805 VDD.n3798 92.5005
R7317 VDD.n3805 VDD.n3804 92.5005
R7318 VDD.n3807 VDD.n3806 92.5005
R7319 VDD.n3806 VDD.n3551 92.5005
R7320 VDD.n4061 VDD.n4060 92.5005
R7321 VDD.n4060 VDD.n4059 92.5005
R7322 VDD.n3866 VDD.n3421 92.5005
R7323 VDD.n3423 VDD.n3421 92.5005
R7324 VDD.n3864 VDD.n3863 92.5005
R7325 VDD.n3863 VDD.n3862 92.5005
R7326 VDD.n3439 VDD.n3428 92.5005
R7327 VDD.n3436 VDD.n3428 92.5005
R7328 VDD.n3855 VDD.n3854 92.5005
R7329 VDD.n3856 VDD.n3855 92.5005
R7330 VDD.n3852 VDD.n3438 92.5005
R7331 VDD.n3445 VDD.n3438 92.5005
R7332 VDD.n3840 VDD.n3839 92.5005
R7333 VDD.n3839 VDD.n3513 92.5005
R7334 VDD.n3838 VDD.n3527 92.5005
R7335 VDD.n3838 VDD.n3837 92.5005
R7336 VDD.n3797 VDD.n3525 92.5005
R7337 VDD.n3799 VDD.n3525 92.5005
R7338 VDD.n3830 VDD.n3829 92.5005
R7339 VDD.n3831 VDD.n3830 92.5005
R7340 VDD.n3828 VDD.n3796 92.5005
R7341 VDD.n3810 VDD.n3796 92.5005
R7342 VDD.n3795 VDD.n3286 92.5005
R7343 VDD.n3795 VDD.n3289 92.5005
R7344 VDD.n3871 VDD.n3422 92.5005
R7345 VDD.n3871 VDD.n3870 92.5005
R7346 VDD.n2623 VDD.n2620 92.5005
R7347 VDD.n3084 VDD.n2623 92.5005
R7348 VDD.n2978 VDD.n2977 92.5005
R7349 VDD.n2978 VDD.n2503 92.5005
R7350 VDD.n2764 VDD.n2763 92.5005
R7351 VDD.n3024 VDD.n2764 92.5005
R7352 VDD.n3047 VDD.n3046 92.5005
R7353 VDD.n3046 VDD.n3045 92.5005
R7354 VDD.n3048 VDD.n2744 92.5005
R7355 VDD.n3013 VDD.n2744 92.5005
R7356 VDD.n3050 VDD.n3049 92.5005
R7357 VDD.n3051 VDD.n3050 92.5005
R7358 VDD.n2762 VDD.n2743 92.5005
R7359 VDD.n2743 VDD.n2727 92.5005
R7360 VDD.n2757 VDD.n2745 92.5005
R7361 VDD.n2756 VDD.n2755 92.5005
R7362 VDD.n2754 VDD.n2753 92.5005
R7363 VDD.n2752 VDD.n2748 92.5005
R7364 VDD.n2750 VDD.n2749 92.5005
R7365 VDD.n2760 VDD.n2759 92.5005
R7366 VDD.n2649 VDD.n2648 92.5005
R7367 VDD.n2659 VDD.n2649 92.5005
R7368 VDD.n3072 VDD.n3071 92.5005
R7369 VDD.n3071 VDD.n3070 92.5005
R7370 VDD.n3073 VDD.n2646 92.5005
R7371 VDD.n2650 VDD.n2646 92.5005
R7372 VDD.n3075 VDD.n3074 92.5005
R7373 VDD.n3076 VDD.n3075 92.5005
R7374 VDD.n2647 VDD.n2645 92.5005
R7375 VDD.n2645 VDD.n2637 92.5005
R7376 VDD.n3115 VDD.n2596 92.5005
R7377 VDD.n2596 VDD.n2595 92.5005
R7378 VDD.n3138 VDD.n3137 92.5005
R7379 VDD.n3137 VDD.n3136 92.5005
R7380 VDD.n2586 VDD.n2585 92.5005
R7381 VDD.n3135 VDD.n2586 92.5005
R7382 VDD.n3133 VDD.n3132 92.5005
R7383 VDD.n3134 VDD.n3133 92.5005
R7384 VDD.n3131 VDD.n2588 92.5005
R7385 VDD.n2588 VDD.n2587 92.5005
R7386 VDD.n3130 VDD.n3129 92.5005
R7387 VDD.n3129 VDD.n3128 92.5005
R7388 VDD.n2590 VDD.n2589 92.5005
R7389 VDD.n3127 VDD.n2590 92.5005
R7390 VDD.n3125 VDD.n3124 92.5005
R7391 VDD.n3126 VDD.n3125 92.5005
R7392 VDD.n3123 VDD.n2592 92.5005
R7393 VDD.n2592 VDD.n2591 92.5005
R7394 VDD.n3122 VDD.n3121 92.5005
R7395 VDD.n3121 VDD.n3120 92.5005
R7396 VDD.n2594 VDD.n2593 92.5005
R7397 VDD.n3119 VDD.n2594 92.5005
R7398 VDD.n3117 VDD.n3116 92.5005
R7399 VDD.n3118 VDD.n3117 92.5005
R7400 VDD.n3139 VDD.n2583 92.5005
R7401 VDD.n2583 VDD.n2582 92.5005
R7402 VDD.n3142 VDD.n3141 92.5005
R7403 VDD.n3143 VDD.n3142 92.5005
R7404 VDD.n3140 VDD.n2584 92.5005
R7405 VDD.n2580 VDD.n2579 92.5005
R7406 VDD.n3147 VDD.n3146 92.5005
R7407 VDD.n3146 VDD.n3145 92.5005
R7408 VDD.n3150 VDD.n3149 92.5005
R7409 VDD.n3151 VDD.n3150 92.5005
R7410 VDD.n2576 VDD.n2575 92.5005
R7411 VDD.n3152 VDD.n2576 92.5005
R7412 VDD.n3155 VDD.n3154 92.5005
R7413 VDD.n3154 VDD.n3153 92.5005
R7414 VDD.n3156 VDD.n2574 92.5005
R7415 VDD.n2574 VDD.n2573 92.5005
R7416 VDD.n3158 VDD.n3157 92.5005
R7417 VDD.n3159 VDD.n3158 92.5005
R7418 VDD.n2572 VDD.n2571 92.5005
R7419 VDD.n3160 VDD.n2572 92.5005
R7420 VDD.n3163 VDD.n3162 92.5005
R7421 VDD.n3162 VDD.n3161 92.5005
R7422 VDD.n3164 VDD.n2570 92.5005
R7423 VDD.n2570 VDD.n2569 92.5005
R7424 VDD.n3166 VDD.n3165 92.5005
R7425 VDD.n3167 VDD.n3166 92.5005
R7426 VDD.n2568 VDD.n2567 92.5005
R7427 VDD.n3168 VDD.n2568 92.5005
R7428 VDD.n3171 VDD.n3170 92.5005
R7429 VDD.n3170 VDD.n3169 92.5005
R7430 VDD.n3172 VDD.n2566 92.5005
R7431 VDD.n2566 VDD.n2565 92.5005
R7432 VDD.n3174 VDD.n3173 92.5005
R7433 VDD.n3175 VDD.n3174 92.5005
R7434 VDD.n2564 VDD.n2563 92.5005
R7435 VDD.n3176 VDD.n2564 92.5005
R7436 VDD.n3179 VDD.n3178 92.5005
R7437 VDD.n3178 VDD.n3177 92.5005
R7438 VDD.n3180 VDD.n2562 92.5005
R7439 VDD.n2562 VDD.n2561 92.5005
R7440 VDD.n3182 VDD.n3181 92.5005
R7441 VDD.n3183 VDD.n3182 92.5005
R7442 VDD.n2560 VDD.n2559 92.5005
R7443 VDD.n3184 VDD.n2560 92.5005
R7444 VDD.n3187 VDD.n3186 92.5005
R7445 VDD.n3186 VDD.n3185 92.5005
R7446 VDD.n3188 VDD.n2558 92.5005
R7447 VDD.n2558 VDD.n2557 92.5005
R7448 VDD.n3190 VDD.n3189 92.5005
R7449 VDD.n3191 VDD.n3190 92.5005
R7450 VDD.n2556 VDD.n2555 92.5005
R7451 VDD.n3192 VDD.n2556 92.5005
R7452 VDD.n3195 VDD.n3194 92.5005
R7453 VDD.n3194 VDD.n3193 92.5005
R7454 VDD.n3196 VDD.n2554 92.5005
R7455 VDD.n2554 VDD.n2553 92.5005
R7456 VDD.n3198 VDD.n3197 92.5005
R7457 VDD.n3199 VDD.n3198 92.5005
R7458 VDD.n2552 VDD.n2551 92.5005
R7459 VDD.n3200 VDD.n2552 92.5005
R7460 VDD.n3203 VDD.n3202 92.5005
R7461 VDD.n3202 VDD.n3201 92.5005
R7462 VDD.n3204 VDD.n2549 92.5005
R7463 VDD.n2549 VDD.n2546 92.5005
R7464 VDD.n3148 VDD.n2578 92.5005
R7465 VDD.n2578 VDD.n2577 92.5005
R7466 VDD.n2541 VDD.n2540 92.5005
R7467 VDD.n3216 VDD.n2541 92.5005
R7468 VDD.n3219 VDD.n3218 92.5005
R7469 VDD.n3218 VDD.n3217 92.5005
R7470 VDD.n3220 VDD.n2539 92.5005
R7471 VDD.n2539 VDD.n2538 92.5005
R7472 VDD.n3222 VDD.n3221 92.5005
R7473 VDD.n3223 VDD.n3222 92.5005
R7474 VDD.n2537 VDD.n2536 92.5005
R7475 VDD.n3224 VDD.n2537 92.5005
R7476 VDD.n3227 VDD.n3226 92.5005
R7477 VDD.n3226 VDD.n3225 92.5005
R7478 VDD.n3228 VDD.n2535 92.5005
R7479 VDD.n2535 VDD.n2534 92.5005
R7480 VDD.n3230 VDD.n3229 92.5005
R7481 VDD.n3231 VDD.n3230 92.5005
R7482 VDD.n2532 VDD.n2531 92.5005
R7483 VDD.n3232 VDD.n2532 92.5005
R7484 VDD.n3235 VDD.n3234 92.5005
R7485 VDD.n3234 VDD.n3233 92.5005
R7486 VDD.n3236 VDD.n2530 92.5005
R7487 VDD.n2533 VDD.n2530 92.5005
R7488 VDD.n3212 VDD.n2543 92.5005
R7489 VDD.n2543 VDD.n2542 92.5005
R7490 VDD.n3211 VDD.n3210 92.5005
R7491 VDD.n3210 VDD.n3209 92.5005
R7492 VDD.n2545 VDD.n2544 92.5005
R7493 VDD.n2550 VDD.n2548 92.5005
R7494 VDD.n3206 VDD.n3205 92.5005
R7495 VDD.n3207 VDD.n3206 92.5005
R7496 VDD.n3214 VDD.n3213 92.5005
R7497 VDD.n3215 VDD.n3214 92.5005
R7498 VDD.n3239 VDD.n3238 92.5005
R7499 VDD.n3260 VDD.n2514 92.5005
R7500 VDD.n3259 VDD.n3258 92.5005
R7501 VDD.n2523 VDD.n2519 92.5005
R7502 VDD.n3253 VDD.n3252 92.5005
R7503 VDD.n3250 VDD.n3249 92.5005
R7504 VDD.n2525 VDD.n2524 92.5005
R7505 VDD.n3243 VDD.n3242 92.5005
R7506 VDD.n3241 VDD.n2528 92.5005
R7507 VDD.n3263 VDD.n3262 92.5005
R7508 VDD.n3000 VDD.n2499 92.5005
R7509 VDD.n3002 VDD.n2498 92.5005
R7510 VDD.n2774 VDD.n2773 92.5005
R7511 VDD.n2984 VDD.n2983 92.5005
R7512 VDD.n2988 VDD.n2987 92.5005
R7513 VDD.n2986 VDD.n2770 92.5005
R7514 VDD.n2997 VDD.n2996 92.5005
R7515 VDD.n2998 VDD.n2767 92.5005
R7516 VDD.n2995 VDD.n2766 92.5005
R7517 VDD.n2994 VDD.n2993 92.5005
R7518 VDD.n2990 VDD.n2989 92.5005
R7519 VDD.n2979 VDD.n2772 92.5005
R7520 VDD.n2982 VDD.n2981 92.5005
R7521 VDD.n2972 VDD.n2775 92.5005
R7522 VDD.n2975 VDD.n2974 92.5005
R7523 VDD.n3008 VDD.n3007 92.5005
R7524 VDD.n3008 VDD.n2504 92.5005
R7525 VDD.n3006 VDD.n3005 92.5005
R7526 VDD.n3004 VDD.n2768 92.5005
R7527 VDD.n2932 VDD.n2791 92.5005
R7528 VDD.n2934 VDD.n2933 92.5005
R7529 VDD.n2936 VDD.n2935 92.5005
R7530 VDD.n2937 VDD.n2793 92.5005
R7531 VDD.n2939 VDD.n2938 92.5005
R7532 VDD.n2790 VDD.n2789 92.5005
R7533 VDD.n2943 VDD.n2790 92.5005
R7534 VDD.n2946 VDD.n2945 92.5005
R7535 VDD.n2945 VDD.n2944 92.5005
R7536 VDD.n2947 VDD.n2788 92.5005
R7537 VDD.n2788 VDD.n2787 92.5005
R7538 VDD.n2949 VDD.n2948 92.5005
R7539 VDD.n2950 VDD.n2949 92.5005
R7540 VDD.n2786 VDD.n2785 92.5005
R7541 VDD.n2951 VDD.n2786 92.5005
R7542 VDD.n2954 VDD.n2953 92.5005
R7543 VDD.n2953 VDD.n2952 92.5005
R7544 VDD.n2955 VDD.n2784 92.5005
R7545 VDD.n2784 VDD.n2783 92.5005
R7546 VDD.n2957 VDD.n2956 92.5005
R7547 VDD.n2958 VDD.n2957 92.5005
R7548 VDD.n2782 VDD.n2781 92.5005
R7549 VDD.n2959 VDD.n2782 92.5005
R7550 VDD.n2962 VDD.n2961 92.5005
R7551 VDD.n2961 VDD.n2960 92.5005
R7552 VDD.n2963 VDD.n2780 92.5005
R7553 VDD.n2780 VDD.n2779 92.5005
R7554 VDD.n2966 VDD.n2965 92.5005
R7555 VDD.n2967 VDD.n2966 92.5005
R7556 VDD.n2964 VDD.n2777 92.5005
R7557 VDD.n2968 VDD.n2777 92.5005
R7558 VDD.n2971 VDD.n2778 92.5005
R7559 VDD.n2971 VDD.n2970 92.5005
R7560 VDD.n2820 VDD.n2819 92.5005
R7561 VDD.n2880 VDD.n2820 92.5005
R7562 VDD.n2883 VDD.n2882 92.5005
R7563 VDD.n2882 VDD.n2881 92.5005
R7564 VDD.n2884 VDD.n2818 92.5005
R7565 VDD.n2818 VDD.n2817 92.5005
R7566 VDD.n2886 VDD.n2885 92.5005
R7567 VDD.n2887 VDD.n2886 92.5005
R7568 VDD.n2816 VDD.n2815 92.5005
R7569 VDD.n2888 VDD.n2816 92.5005
R7570 VDD.n2891 VDD.n2890 92.5005
R7571 VDD.n2890 VDD.n2889 92.5005
R7572 VDD.n2892 VDD.n2814 92.5005
R7573 VDD.n2814 VDD.n2813 92.5005
R7574 VDD.n2894 VDD.n2893 92.5005
R7575 VDD.n2895 VDD.n2894 92.5005
R7576 VDD.n2812 VDD.n2811 92.5005
R7577 VDD.n2896 VDD.n2812 92.5005
R7578 VDD.n2899 VDD.n2898 92.5005
R7579 VDD.n2898 VDD.n2897 92.5005
R7580 VDD.n2900 VDD.n2810 92.5005
R7581 VDD.n2810 VDD.n2809 92.5005
R7582 VDD.n2902 VDD.n2901 92.5005
R7583 VDD.n2903 VDD.n2902 92.5005
R7584 VDD.n2808 VDD.n2807 92.5005
R7585 VDD.n2904 VDD.n2808 92.5005
R7586 VDD.n2907 VDD.n2906 92.5005
R7587 VDD.n2906 VDD.n2905 92.5005
R7588 VDD.n2908 VDD.n2806 92.5005
R7589 VDD.n2806 VDD.n2805 92.5005
R7590 VDD.n2910 VDD.n2909 92.5005
R7591 VDD.n2911 VDD.n2910 92.5005
R7592 VDD.n2804 VDD.n2803 92.5005
R7593 VDD.n2912 VDD.n2804 92.5005
R7594 VDD.n2915 VDD.n2914 92.5005
R7595 VDD.n2914 VDD.n2913 92.5005
R7596 VDD.n2916 VDD.n2802 92.5005
R7597 VDD.n2802 VDD.n2801 92.5005
R7598 VDD.n2918 VDD.n2917 92.5005
R7599 VDD.n2919 VDD.n2918 92.5005
R7600 VDD.n2800 VDD.n2799 92.5005
R7601 VDD.n2920 VDD.n2800 92.5005
R7602 VDD.n2923 VDD.n2922 92.5005
R7603 VDD.n2922 VDD.n2921 92.5005
R7604 VDD.n2924 VDD.n2798 92.5005
R7605 VDD.n2798 VDD.n2797 92.5005
R7606 VDD.n2927 VDD.n2926 92.5005
R7607 VDD.n2928 VDD.n2927 92.5005
R7608 VDD.n2925 VDD.n2795 92.5005
R7609 VDD.n2929 VDD.n2795 92.5005
R7610 VDD.n2931 VDD.n2796 92.5005
R7611 VDD.n2931 VDD.n2930 92.5005
R7612 VDD.n2875 VDD.n2874 92.5005
R7613 VDD.n2822 VDD.n2821 92.5005
R7614 VDD.n2879 VDD.n2878 92.5005
R7615 VDD.n2619 VDD.n2618 92.5005
R7616 VDD.n2841 VDD.n2618 92.5005
R7617 VDD.n2844 VDD.n2843 92.5005
R7618 VDD.n2843 VDD.n2842 92.5005
R7619 VDD.n2846 VDD.n2845 92.5005
R7620 VDD.n2847 VDD.n2846 92.5005
R7621 VDD.n2840 VDD.n2839 92.5005
R7622 VDD.n2848 VDD.n2840 92.5005
R7623 VDD.n2851 VDD.n2850 92.5005
R7624 VDD.n2850 VDD.n2849 92.5005
R7625 VDD.n2852 VDD.n2838 92.5005
R7626 VDD.n2838 VDD.n2837 92.5005
R7627 VDD.n2854 VDD.n2853 92.5005
R7628 VDD.n2855 VDD.n2854 92.5005
R7629 VDD.n2836 VDD.n2835 92.5005
R7630 VDD.n2856 VDD.n2836 92.5005
R7631 VDD.n2859 VDD.n2858 92.5005
R7632 VDD.n2858 VDD.n2857 92.5005
R7633 VDD.n2860 VDD.n2834 92.5005
R7634 VDD.n2834 VDD.n2833 92.5005
R7635 VDD.n2862 VDD.n2861 92.5005
R7636 VDD.n2863 VDD.n2862 92.5005
R7637 VDD.n2831 VDD.n2830 92.5005
R7638 VDD.n2864 VDD.n2831 92.5005
R7639 VDD.n2867 VDD.n2866 92.5005
R7640 VDD.n2866 VDD.n2865 92.5005
R7641 VDD.n2868 VDD.n2828 92.5005
R7642 VDD.n2832 VDD.n2828 92.5005
R7643 VDD.n2870 VDD.n2869 92.5005
R7644 VDD.n2829 VDD.n2827 92.5005
R7645 VDD.n2824 VDD.n2823 92.5005
R7646 VDD.n3114 VDD.n3113 92.5005
R7647 VDD.n2695 VDD.n2598 92.5005
R7648 VDD.n2697 VDD.n2696 92.5005
R7649 VDD.n2694 VDD.n2693 92.5005
R7650 VDD.n2664 VDD.n2663 92.5005
R7651 VDD.n2688 VDD.n2687 92.5005
R7652 VDD.n2666 VDD.n2665 92.5005
R7653 VDD.n2682 VDD.n2681 92.5005
R7654 VDD.n2678 VDD.n2677 92.5005
R7655 VDD.n2676 VDD.n2675 92.5005
R7656 VDD.n3089 VDD.n3088 92.5005
R7657 VDD.n3093 VDD.n3092 92.5005
R7658 VDD.n3096 VDD.n3095 92.5005
R7659 VDD.n2633 VDD.n2632 92.5005
R7660 VDD.n2622 VDD.n2621 92.5005
R7661 VDD.n3105 VDD.n3104 92.5005
R7662 VDD.n3106 VDD.n2617 92.5005
R7663 VDD.n3109 VDD.n3108 92.5005
R7664 VDD.n3103 VDD.n3102 92.5005
R7665 VDD.n2631 VDD.n2624 92.5005
R7666 VDD.n3098 VDD.n3097 92.5005
R7667 VDD.n3094 VDD.n2630 92.5005
R7668 VDD.n3091 VDD.n3090 92.5005
R7669 VDD.n2634 VDD.n2610 92.5005
R7670 VDD.n3111 VDD.n2610 92.5005
R7671 VDD.n3087 VDD.n3086 92.5005
R7672 VDD.n2670 VDD.n2669 92.5005
R7673 VDD.n2672 VDD.n2671 92.5005
R7674 VDD.n2674 VDD.n2673 92.5005
R7675 VDD.n2680 VDD.n2679 92.5005
R7676 VDD.n2699 VDD.n2698 92.5005
R7677 VDD.n2692 VDD.n2691 92.5005
R7678 VDD.n2690 VDD.n2689 92.5005
R7679 VDD.n2686 VDD.n2685 92.5005
R7680 VDD.n2684 VDD.n2683 92.5005
R7681 VDD.n2510 VDD.n2502 92.5005
R7682 VDD.n3267 VDD.n3266 92.5005
R7683 VDD.n3265 VDD.n3264 92.5005
R7684 VDD.n3265 VDD.n2511 92.5005
R7685 VDD.n3257 VDD.n3256 92.5005
R7686 VDD.n3255 VDD.n3254 92.5005
R7687 VDD.n2526 VDD.n2522 92.5005
R7688 VDD.n3248 VDD.n3247 92.5005
R7689 VDD.n3245 VDD.n3244 92.5005
R7690 VDD.n2518 VDD.n2513 92.5005
R7691 VDD.n3029 VDD.n3028 92.5005
R7692 VDD.n3031 VDD.n3030 92.5005
R7693 VDD.n3033 VDD.n3032 92.5005
R7694 VDD.n3035 VDD.n3034 92.5005
R7695 VDD.n3023 VDD.n3022 92.5005
R7696 VDD.n3040 VDD.n3039 92.5005
R7697 VDD.n2509 VDD.n2508 92.5005
R7698 VDD.n2511 VDD.n2509 92.5005
R7699 VDD.n3269 VDD.n3268 92.5005
R7700 VDD.n3268 VDD.n3267 92.5005
R7701 VDD.n3270 VDD.n2506 92.5005
R7702 VDD.n2510 VDD.n2506 92.5005
R7703 VDD.n3272 VDD.n3271 92.5005
R7704 VDD.n3273 VDD.n3272 92.5005
R7705 VDD.n3015 VDD.n3014 92.5005
R7706 VDD.n3014 VDD.n2765 92.5005
R7707 VDD.n3017 VDD.n3016 92.5005
R7708 VDD.n3018 VDD.n3017 92.5005
R7709 VDD.n2725 VDD.n2724 92.5005
R7710 VDD.n2742 VDD.n2725 92.5005
R7711 VDD.n3059 VDD.n3058 92.5005
R7712 VDD.n3058 VDD.n3057 92.5005
R7713 VDD.n3060 VDD.n2662 92.5005
R7714 VDD.n2726 VDD.n2662 92.5005
R7715 VDD.n3062 VDD.n3061 92.5005
R7716 VDD.n3063 VDD.n3062 92.5005
R7717 VDD.n2706 VDD.n2705 92.5005
R7718 VDD.n2705 VDD.n2644 92.5005
R7719 VDD.n2704 VDD.n2703 92.5005
R7720 VDD.n2704 VDD.n2643 92.5005
R7721 VDD.n2702 VDD.n2638 92.5005
R7722 VDD.n3083 VDD.n2638 92.5005
R7723 VDD.n2701 VDD.n2700 92.5005
R7724 VDD.n2700 VDD.n2625 92.5005
R7725 VDD.n2722 VDD.n2721 92.5005
R7726 VDD.n2719 VDD.n2707 92.5005
R7727 VDD.n2717 VDD.n2716 92.5005
R7728 VDD.n2715 VDD.n2714 92.5005
R7729 VDD.n2712 VDD.n2709 92.5005
R7730 VDD.n2710 VDD.n2654 92.5005
R7731 VDD.n2667 VDD.n2639 92.5005
R7732 VDD.n2639 VDD.n2625 92.5005
R7733 VDD.n3082 VDD.n3081 92.5005
R7734 VDD.n3083 VDD.n3082 92.5005
R7735 VDD.n3079 VDD.n2640 92.5005
R7736 VDD.n2643 VDD.n2640 92.5005
R7737 VDD.n2656 VDD.n2641 92.5005
R7738 VDD.n2656 VDD.n2644 92.5005
R7739 VDD.n3065 VDD.n3064 92.5005
R7740 VDD.n3064 VDD.n3063 92.5005
R7741 VDD.n2729 VDD.n2658 92.5005
R7742 VDD.n2726 VDD.n2658 92.5005
R7743 VDD.n3056 VDD.n3055 92.5005
R7744 VDD.n3057 VDD.n3056 92.5005
R7745 VDD.n2740 VDD.n2728 92.5005
R7746 VDD.n2742 VDD.n2728 92.5005
R7747 VDD.n3019 VDD.n3012 92.5005
R7748 VDD.n3019 VDD.n3018 92.5005
R7749 VDD.n3021 VDD.n3020 92.5005
R7750 VDD.n3020 VDD.n2765 92.5005
R7751 VDD.n3275 VDD.n3274 92.5005
R7752 VDD.n3274 VDD.n3273 92.5005
R7753 VDD.n3080 VDD.n2635 92.5005
R7754 VDD.n2637 VDD.n2635 92.5005
R7755 VDD.n3078 VDD.n3077 92.5005
R7756 VDD.n3077 VDD.n3076 92.5005
R7757 VDD.n2653 VDD.n2642 92.5005
R7758 VDD.n2650 VDD.n2642 92.5005
R7759 VDD.n3069 VDD.n3068 92.5005
R7760 VDD.n3070 VDD.n3069 92.5005
R7761 VDD.n3066 VDD.n2652 92.5005
R7762 VDD.n2659 VDD.n2652 92.5005
R7763 VDD.n3054 VDD.n3053 92.5005
R7764 VDD.n3053 VDD.n2727 92.5005
R7765 VDD.n3052 VDD.n2741 92.5005
R7766 VDD.n3052 VDD.n3051 92.5005
R7767 VDD.n3011 VDD.n2739 92.5005
R7768 VDD.n3013 VDD.n2739 92.5005
R7769 VDD.n3044 VDD.n3043 92.5005
R7770 VDD.n3045 VDD.n3044 92.5005
R7771 VDD.n3042 VDD.n3010 92.5005
R7772 VDD.n3024 VDD.n3010 92.5005
R7773 VDD.n3009 VDD.n2500 92.5005
R7774 VDD.n3009 VDD.n2503 92.5005
R7775 VDD.n3085 VDD.n2636 92.5005
R7776 VDD.n3085 VDD.n3084 92.5005
R7777 VDD.n1768 VDD.n1765 92.5005
R7778 VDD.n2229 VDD.n1768 92.5005
R7779 VDD.n2123 VDD.n2122 92.5005
R7780 VDD.n2123 VDD.n1648 92.5005
R7781 VDD.n1909 VDD.n1908 92.5005
R7782 VDD.n2169 VDD.n1909 92.5005
R7783 VDD.n2192 VDD.n2191 92.5005
R7784 VDD.n2191 VDD.n2190 92.5005
R7785 VDD.n2193 VDD.n1889 92.5005
R7786 VDD.n2158 VDD.n1889 92.5005
R7787 VDD.n2195 VDD.n2194 92.5005
R7788 VDD.n2196 VDD.n2195 92.5005
R7789 VDD.n1907 VDD.n1888 92.5005
R7790 VDD.n1888 VDD.n1872 92.5005
R7791 VDD.n1902 VDD.n1890 92.5005
R7792 VDD.n1901 VDD.n1900 92.5005
R7793 VDD.n1899 VDD.n1898 92.5005
R7794 VDD.n1897 VDD.n1893 92.5005
R7795 VDD.n1895 VDD.n1894 92.5005
R7796 VDD.n1905 VDD.n1904 92.5005
R7797 VDD.n1794 VDD.n1793 92.5005
R7798 VDD.n1804 VDD.n1794 92.5005
R7799 VDD.n2217 VDD.n2216 92.5005
R7800 VDD.n2216 VDD.n2215 92.5005
R7801 VDD.n2218 VDD.n1791 92.5005
R7802 VDD.n1795 VDD.n1791 92.5005
R7803 VDD.n2220 VDD.n2219 92.5005
R7804 VDD.n2221 VDD.n2220 92.5005
R7805 VDD.n1792 VDD.n1790 92.5005
R7806 VDD.n1790 VDD.n1782 92.5005
R7807 VDD.n2260 VDD.n1741 92.5005
R7808 VDD.n1741 VDD.n1740 92.5005
R7809 VDD.n2283 VDD.n2282 92.5005
R7810 VDD.n2282 VDD.n2281 92.5005
R7811 VDD.n1731 VDD.n1730 92.5005
R7812 VDD.n2280 VDD.n1731 92.5005
R7813 VDD.n2278 VDD.n2277 92.5005
R7814 VDD.n2279 VDD.n2278 92.5005
R7815 VDD.n2276 VDD.n1733 92.5005
R7816 VDD.n1733 VDD.n1732 92.5005
R7817 VDD.n2275 VDD.n2274 92.5005
R7818 VDD.n2274 VDD.n2273 92.5005
R7819 VDD.n1735 VDD.n1734 92.5005
R7820 VDD.n2272 VDD.n1735 92.5005
R7821 VDD.n2270 VDD.n2269 92.5005
R7822 VDD.n2271 VDD.n2270 92.5005
R7823 VDD.n2268 VDD.n1737 92.5005
R7824 VDD.n1737 VDD.n1736 92.5005
R7825 VDD.n2267 VDD.n2266 92.5005
R7826 VDD.n2266 VDD.n2265 92.5005
R7827 VDD.n1739 VDD.n1738 92.5005
R7828 VDD.n2264 VDD.n1739 92.5005
R7829 VDD.n2262 VDD.n2261 92.5005
R7830 VDD.n2263 VDD.n2262 92.5005
R7831 VDD.n2284 VDD.n1728 92.5005
R7832 VDD.n1728 VDD.n1727 92.5005
R7833 VDD.n2287 VDD.n2286 92.5005
R7834 VDD.n2288 VDD.n2287 92.5005
R7835 VDD.n2285 VDD.n1729 92.5005
R7836 VDD.n1725 VDD.n1724 92.5005
R7837 VDD.n2292 VDD.n2291 92.5005
R7838 VDD.n2291 VDD.n2290 92.5005
R7839 VDD.n2295 VDD.n2294 92.5005
R7840 VDD.n2296 VDD.n2295 92.5005
R7841 VDD.n1721 VDD.n1720 92.5005
R7842 VDD.n2297 VDD.n1721 92.5005
R7843 VDD.n2300 VDD.n2299 92.5005
R7844 VDD.n2299 VDD.n2298 92.5005
R7845 VDD.n2301 VDD.n1719 92.5005
R7846 VDD.n1719 VDD.n1718 92.5005
R7847 VDD.n2303 VDD.n2302 92.5005
R7848 VDD.n2304 VDD.n2303 92.5005
R7849 VDD.n1717 VDD.n1716 92.5005
R7850 VDD.n2305 VDD.n1717 92.5005
R7851 VDD.n2308 VDD.n2307 92.5005
R7852 VDD.n2307 VDD.n2306 92.5005
R7853 VDD.n2309 VDD.n1715 92.5005
R7854 VDD.n1715 VDD.n1714 92.5005
R7855 VDD.n2311 VDD.n2310 92.5005
R7856 VDD.n2312 VDD.n2311 92.5005
R7857 VDD.n1713 VDD.n1712 92.5005
R7858 VDD.n2313 VDD.n1713 92.5005
R7859 VDD.n2316 VDD.n2315 92.5005
R7860 VDD.n2315 VDD.n2314 92.5005
R7861 VDD.n2317 VDD.n1711 92.5005
R7862 VDD.n1711 VDD.n1710 92.5005
R7863 VDD.n2319 VDD.n2318 92.5005
R7864 VDD.n2320 VDD.n2319 92.5005
R7865 VDD.n1709 VDD.n1708 92.5005
R7866 VDD.n2321 VDD.n1709 92.5005
R7867 VDD.n2324 VDD.n2323 92.5005
R7868 VDD.n2323 VDD.n2322 92.5005
R7869 VDD.n2325 VDD.n1707 92.5005
R7870 VDD.n1707 VDD.n1706 92.5005
R7871 VDD.n2327 VDD.n2326 92.5005
R7872 VDD.n2328 VDD.n2327 92.5005
R7873 VDD.n1705 VDD.n1704 92.5005
R7874 VDD.n2329 VDD.n1705 92.5005
R7875 VDD.n2332 VDD.n2331 92.5005
R7876 VDD.n2331 VDD.n2330 92.5005
R7877 VDD.n2333 VDD.n1703 92.5005
R7878 VDD.n1703 VDD.n1702 92.5005
R7879 VDD.n2335 VDD.n2334 92.5005
R7880 VDD.n2336 VDD.n2335 92.5005
R7881 VDD.n1701 VDD.n1700 92.5005
R7882 VDD.n2337 VDD.n1701 92.5005
R7883 VDD.n2340 VDD.n2339 92.5005
R7884 VDD.n2339 VDD.n2338 92.5005
R7885 VDD.n2341 VDD.n1699 92.5005
R7886 VDD.n1699 VDD.n1698 92.5005
R7887 VDD.n2343 VDD.n2342 92.5005
R7888 VDD.n2344 VDD.n2343 92.5005
R7889 VDD.n1697 VDD.n1696 92.5005
R7890 VDD.n2345 VDD.n1697 92.5005
R7891 VDD.n2348 VDD.n2347 92.5005
R7892 VDD.n2347 VDD.n2346 92.5005
R7893 VDD.n2349 VDD.n1694 92.5005
R7894 VDD.n1694 VDD.n1691 92.5005
R7895 VDD.n2293 VDD.n1723 92.5005
R7896 VDD.n1723 VDD.n1722 92.5005
R7897 VDD.n1686 VDD.n1685 92.5005
R7898 VDD.n2361 VDD.n1686 92.5005
R7899 VDD.n2364 VDD.n2363 92.5005
R7900 VDD.n2363 VDD.n2362 92.5005
R7901 VDD.n2365 VDD.n1684 92.5005
R7902 VDD.n1684 VDD.n1683 92.5005
R7903 VDD.n2367 VDD.n2366 92.5005
R7904 VDD.n2368 VDD.n2367 92.5005
R7905 VDD.n1682 VDD.n1681 92.5005
R7906 VDD.n2369 VDD.n1682 92.5005
R7907 VDD.n2372 VDD.n2371 92.5005
R7908 VDD.n2371 VDD.n2370 92.5005
R7909 VDD.n2373 VDD.n1680 92.5005
R7910 VDD.n1680 VDD.n1679 92.5005
R7911 VDD.n2375 VDD.n2374 92.5005
R7912 VDD.n2376 VDD.n2375 92.5005
R7913 VDD.n1677 VDD.n1676 92.5005
R7914 VDD.n2377 VDD.n1677 92.5005
R7915 VDD.n2380 VDD.n2379 92.5005
R7916 VDD.n2379 VDD.n2378 92.5005
R7917 VDD.n2381 VDD.n1675 92.5005
R7918 VDD.n1678 VDD.n1675 92.5005
R7919 VDD.n2357 VDD.n1688 92.5005
R7920 VDD.n1688 VDD.n1687 92.5005
R7921 VDD.n2356 VDD.n2355 92.5005
R7922 VDD.n2355 VDD.n2354 92.5005
R7923 VDD.n1690 VDD.n1689 92.5005
R7924 VDD.n1695 VDD.n1693 92.5005
R7925 VDD.n2351 VDD.n2350 92.5005
R7926 VDD.n2352 VDD.n2351 92.5005
R7927 VDD.n2359 VDD.n2358 92.5005
R7928 VDD.n2360 VDD.n2359 92.5005
R7929 VDD.n2384 VDD.n2383 92.5005
R7930 VDD.n2405 VDD.n1659 92.5005
R7931 VDD.n2404 VDD.n2403 92.5005
R7932 VDD.n1668 VDD.n1664 92.5005
R7933 VDD.n2398 VDD.n2397 92.5005
R7934 VDD.n2395 VDD.n2394 92.5005
R7935 VDD.n1670 VDD.n1669 92.5005
R7936 VDD.n2388 VDD.n2387 92.5005
R7937 VDD.n2386 VDD.n1673 92.5005
R7938 VDD.n2408 VDD.n2407 92.5005
R7939 VDD.n2145 VDD.n1644 92.5005
R7940 VDD.n2147 VDD.n1643 92.5005
R7941 VDD.n1919 VDD.n1918 92.5005
R7942 VDD.n2129 VDD.n2128 92.5005
R7943 VDD.n2133 VDD.n2132 92.5005
R7944 VDD.n2131 VDD.n1915 92.5005
R7945 VDD.n2142 VDD.n2141 92.5005
R7946 VDD.n2143 VDD.n1912 92.5005
R7947 VDD.n2140 VDD.n1911 92.5005
R7948 VDD.n2139 VDD.n2138 92.5005
R7949 VDD.n2135 VDD.n2134 92.5005
R7950 VDD.n2124 VDD.n1917 92.5005
R7951 VDD.n2127 VDD.n2126 92.5005
R7952 VDD.n2117 VDD.n1920 92.5005
R7953 VDD.n2120 VDD.n2119 92.5005
R7954 VDD.n2153 VDD.n2152 92.5005
R7955 VDD.n2153 VDD.n1649 92.5005
R7956 VDD.n2151 VDD.n2150 92.5005
R7957 VDD.n2149 VDD.n1913 92.5005
R7958 VDD.n2077 VDD.n1936 92.5005
R7959 VDD.n2079 VDD.n2078 92.5005
R7960 VDD.n2081 VDD.n2080 92.5005
R7961 VDD.n2082 VDD.n1938 92.5005
R7962 VDD.n2084 VDD.n2083 92.5005
R7963 VDD.n1935 VDD.n1934 92.5005
R7964 VDD.n2088 VDD.n1935 92.5005
R7965 VDD.n2091 VDD.n2090 92.5005
R7966 VDD.n2090 VDD.n2089 92.5005
R7967 VDD.n2092 VDD.n1933 92.5005
R7968 VDD.n1933 VDD.n1932 92.5005
R7969 VDD.n2094 VDD.n2093 92.5005
R7970 VDD.n2095 VDD.n2094 92.5005
R7971 VDD.n1931 VDD.n1930 92.5005
R7972 VDD.n2096 VDD.n1931 92.5005
R7973 VDD.n2099 VDD.n2098 92.5005
R7974 VDD.n2098 VDD.n2097 92.5005
R7975 VDD.n2100 VDD.n1929 92.5005
R7976 VDD.n1929 VDD.n1928 92.5005
R7977 VDD.n2102 VDD.n2101 92.5005
R7978 VDD.n2103 VDD.n2102 92.5005
R7979 VDD.n1927 VDD.n1926 92.5005
R7980 VDD.n2104 VDD.n1927 92.5005
R7981 VDD.n2107 VDD.n2106 92.5005
R7982 VDD.n2106 VDD.n2105 92.5005
R7983 VDD.n2108 VDD.n1925 92.5005
R7984 VDD.n1925 VDD.n1924 92.5005
R7985 VDD.n2111 VDD.n2110 92.5005
R7986 VDD.n2112 VDD.n2111 92.5005
R7987 VDD.n2109 VDD.n1922 92.5005
R7988 VDD.n2113 VDD.n1922 92.5005
R7989 VDD.n2116 VDD.n1923 92.5005
R7990 VDD.n2116 VDD.n2115 92.5005
R7991 VDD.n1965 VDD.n1964 92.5005
R7992 VDD.n2025 VDD.n1965 92.5005
R7993 VDD.n2028 VDD.n2027 92.5005
R7994 VDD.n2027 VDD.n2026 92.5005
R7995 VDD.n2029 VDD.n1963 92.5005
R7996 VDD.n1963 VDD.n1962 92.5005
R7997 VDD.n2031 VDD.n2030 92.5005
R7998 VDD.n2032 VDD.n2031 92.5005
R7999 VDD.n1961 VDD.n1960 92.5005
R8000 VDD.n2033 VDD.n1961 92.5005
R8001 VDD.n2036 VDD.n2035 92.5005
R8002 VDD.n2035 VDD.n2034 92.5005
R8003 VDD.n2037 VDD.n1959 92.5005
R8004 VDD.n1959 VDD.n1958 92.5005
R8005 VDD.n2039 VDD.n2038 92.5005
R8006 VDD.n2040 VDD.n2039 92.5005
R8007 VDD.n1957 VDD.n1956 92.5005
R8008 VDD.n2041 VDD.n1957 92.5005
R8009 VDD.n2044 VDD.n2043 92.5005
R8010 VDD.n2043 VDD.n2042 92.5005
R8011 VDD.n2045 VDD.n1955 92.5005
R8012 VDD.n1955 VDD.n1954 92.5005
R8013 VDD.n2047 VDD.n2046 92.5005
R8014 VDD.n2048 VDD.n2047 92.5005
R8015 VDD.n1953 VDD.n1952 92.5005
R8016 VDD.n2049 VDD.n1953 92.5005
R8017 VDD.n2052 VDD.n2051 92.5005
R8018 VDD.n2051 VDD.n2050 92.5005
R8019 VDD.n2053 VDD.n1951 92.5005
R8020 VDD.n1951 VDD.n1950 92.5005
R8021 VDD.n2055 VDD.n2054 92.5005
R8022 VDD.n2056 VDD.n2055 92.5005
R8023 VDD.n1949 VDD.n1948 92.5005
R8024 VDD.n2057 VDD.n1949 92.5005
R8025 VDD.n2060 VDD.n2059 92.5005
R8026 VDD.n2059 VDD.n2058 92.5005
R8027 VDD.n2061 VDD.n1947 92.5005
R8028 VDD.n1947 VDD.n1946 92.5005
R8029 VDD.n2063 VDD.n2062 92.5005
R8030 VDD.n2064 VDD.n2063 92.5005
R8031 VDD.n1945 VDD.n1944 92.5005
R8032 VDD.n2065 VDD.n1945 92.5005
R8033 VDD.n2068 VDD.n2067 92.5005
R8034 VDD.n2067 VDD.n2066 92.5005
R8035 VDD.n2069 VDD.n1943 92.5005
R8036 VDD.n1943 VDD.n1942 92.5005
R8037 VDD.n2072 VDD.n2071 92.5005
R8038 VDD.n2073 VDD.n2072 92.5005
R8039 VDD.n2070 VDD.n1940 92.5005
R8040 VDD.n2074 VDD.n1940 92.5005
R8041 VDD.n2076 VDD.n1941 92.5005
R8042 VDD.n2076 VDD.n2075 92.5005
R8043 VDD.n2020 VDD.n2019 92.5005
R8044 VDD.n1967 VDD.n1966 92.5005
R8045 VDD.n2024 VDD.n2023 92.5005
R8046 VDD.n1764 VDD.n1763 92.5005
R8047 VDD.n1986 VDD.n1763 92.5005
R8048 VDD.n1989 VDD.n1988 92.5005
R8049 VDD.n1988 VDD.n1987 92.5005
R8050 VDD.n1991 VDD.n1990 92.5005
R8051 VDD.n1992 VDD.n1991 92.5005
R8052 VDD.n1985 VDD.n1984 92.5005
R8053 VDD.n1993 VDD.n1985 92.5005
R8054 VDD.n1996 VDD.n1995 92.5005
R8055 VDD.n1995 VDD.n1994 92.5005
R8056 VDD.n1997 VDD.n1983 92.5005
R8057 VDD.n1983 VDD.n1982 92.5005
R8058 VDD.n1999 VDD.n1998 92.5005
R8059 VDD.n2000 VDD.n1999 92.5005
R8060 VDD.n1981 VDD.n1980 92.5005
R8061 VDD.n2001 VDD.n1981 92.5005
R8062 VDD.n2004 VDD.n2003 92.5005
R8063 VDD.n2003 VDD.n2002 92.5005
R8064 VDD.n2005 VDD.n1979 92.5005
R8065 VDD.n1979 VDD.n1978 92.5005
R8066 VDD.n2007 VDD.n2006 92.5005
R8067 VDD.n2008 VDD.n2007 92.5005
R8068 VDD.n1976 VDD.n1975 92.5005
R8069 VDD.n2009 VDD.n1976 92.5005
R8070 VDD.n2012 VDD.n2011 92.5005
R8071 VDD.n2011 VDD.n2010 92.5005
R8072 VDD.n2013 VDD.n1973 92.5005
R8073 VDD.n1977 VDD.n1973 92.5005
R8074 VDD.n2015 VDD.n2014 92.5005
R8075 VDD.n1974 VDD.n1972 92.5005
R8076 VDD.n1969 VDD.n1968 92.5005
R8077 VDD.n2259 VDD.n2258 92.5005
R8078 VDD.n1840 VDD.n1743 92.5005
R8079 VDD.n1842 VDD.n1841 92.5005
R8080 VDD.n1839 VDD.n1838 92.5005
R8081 VDD.n1809 VDD.n1808 92.5005
R8082 VDD.n1833 VDD.n1832 92.5005
R8083 VDD.n1811 VDD.n1810 92.5005
R8084 VDD.n1827 VDD.n1826 92.5005
R8085 VDD.n1823 VDD.n1822 92.5005
R8086 VDD.n1821 VDD.n1820 92.5005
R8087 VDD.n2234 VDD.n2233 92.5005
R8088 VDD.n2238 VDD.n2237 92.5005
R8089 VDD.n2241 VDD.n2240 92.5005
R8090 VDD.n1778 VDD.n1777 92.5005
R8091 VDD.n1767 VDD.n1766 92.5005
R8092 VDD.n2250 VDD.n2249 92.5005
R8093 VDD.n2251 VDD.n1762 92.5005
R8094 VDD.n2254 VDD.n2253 92.5005
R8095 VDD.n2248 VDD.n2247 92.5005
R8096 VDD.n1776 VDD.n1769 92.5005
R8097 VDD.n2243 VDD.n2242 92.5005
R8098 VDD.n2239 VDD.n1775 92.5005
R8099 VDD.n2236 VDD.n2235 92.5005
R8100 VDD.n1779 VDD.n1755 92.5005
R8101 VDD.n2256 VDD.n1755 92.5005
R8102 VDD.n2232 VDD.n2231 92.5005
R8103 VDD.n1815 VDD.n1814 92.5005
R8104 VDD.n1817 VDD.n1816 92.5005
R8105 VDD.n1819 VDD.n1818 92.5005
R8106 VDD.n1825 VDD.n1824 92.5005
R8107 VDD.n1844 VDD.n1843 92.5005
R8108 VDD.n1837 VDD.n1836 92.5005
R8109 VDD.n1835 VDD.n1834 92.5005
R8110 VDD.n1831 VDD.n1830 92.5005
R8111 VDD.n1829 VDD.n1828 92.5005
R8112 VDD.n1655 VDD.n1647 92.5005
R8113 VDD.n2412 VDD.n2411 92.5005
R8114 VDD.n2410 VDD.n2409 92.5005
R8115 VDD.n2410 VDD.n1656 92.5005
R8116 VDD.n2402 VDD.n2401 92.5005
R8117 VDD.n2400 VDD.n2399 92.5005
R8118 VDD.n1671 VDD.n1667 92.5005
R8119 VDD.n2393 VDD.n2392 92.5005
R8120 VDD.n2390 VDD.n2389 92.5005
R8121 VDD.n1663 VDD.n1658 92.5005
R8122 VDD.n2174 VDD.n2173 92.5005
R8123 VDD.n2176 VDD.n2175 92.5005
R8124 VDD.n2178 VDD.n2177 92.5005
R8125 VDD.n2180 VDD.n2179 92.5005
R8126 VDD.n2168 VDD.n2167 92.5005
R8127 VDD.n2185 VDD.n2184 92.5005
R8128 VDD.n1654 VDD.n1653 92.5005
R8129 VDD.n1656 VDD.n1654 92.5005
R8130 VDD.n2414 VDD.n2413 92.5005
R8131 VDD.n2413 VDD.n2412 92.5005
R8132 VDD.n2415 VDD.n1651 92.5005
R8133 VDD.n1655 VDD.n1651 92.5005
R8134 VDD.n2417 VDD.n2416 92.5005
R8135 VDD.n2418 VDD.n2417 92.5005
R8136 VDD.n2160 VDD.n2159 92.5005
R8137 VDD.n2159 VDD.n1910 92.5005
R8138 VDD.n2162 VDD.n2161 92.5005
R8139 VDD.n2163 VDD.n2162 92.5005
R8140 VDD.n1870 VDD.n1869 92.5005
R8141 VDD.n1887 VDD.n1870 92.5005
R8142 VDD.n2204 VDD.n2203 92.5005
R8143 VDD.n2203 VDD.n2202 92.5005
R8144 VDD.n2205 VDD.n1807 92.5005
R8145 VDD.n1871 VDD.n1807 92.5005
R8146 VDD.n2207 VDD.n2206 92.5005
R8147 VDD.n2208 VDD.n2207 92.5005
R8148 VDD.n1851 VDD.n1850 92.5005
R8149 VDD.n1850 VDD.n1789 92.5005
R8150 VDD.n1849 VDD.n1848 92.5005
R8151 VDD.n1849 VDD.n1788 92.5005
R8152 VDD.n1847 VDD.n1783 92.5005
R8153 VDD.n2228 VDD.n1783 92.5005
R8154 VDD.n1846 VDD.n1845 92.5005
R8155 VDD.n1845 VDD.n1770 92.5005
R8156 VDD.n1867 VDD.n1866 92.5005
R8157 VDD.n1864 VDD.n1852 92.5005
R8158 VDD.n1862 VDD.n1861 92.5005
R8159 VDD.n1860 VDD.n1859 92.5005
R8160 VDD.n1857 VDD.n1854 92.5005
R8161 VDD.n1855 VDD.n1799 92.5005
R8162 VDD.n1812 VDD.n1784 92.5005
R8163 VDD.n1784 VDD.n1770 92.5005
R8164 VDD.n2227 VDD.n2226 92.5005
R8165 VDD.n2228 VDD.n2227 92.5005
R8166 VDD.n2224 VDD.n1785 92.5005
R8167 VDD.n1788 VDD.n1785 92.5005
R8168 VDD.n1801 VDD.n1786 92.5005
R8169 VDD.n1801 VDD.n1789 92.5005
R8170 VDD.n2210 VDD.n2209 92.5005
R8171 VDD.n2209 VDD.n2208 92.5005
R8172 VDD.n1874 VDD.n1803 92.5005
R8173 VDD.n1871 VDD.n1803 92.5005
R8174 VDD.n2201 VDD.n2200 92.5005
R8175 VDD.n2202 VDD.n2201 92.5005
R8176 VDD.n1885 VDD.n1873 92.5005
R8177 VDD.n1887 VDD.n1873 92.5005
R8178 VDD.n2164 VDD.n2157 92.5005
R8179 VDD.n2164 VDD.n2163 92.5005
R8180 VDD.n2166 VDD.n2165 92.5005
R8181 VDD.n2165 VDD.n1910 92.5005
R8182 VDD.n2420 VDD.n2419 92.5005
R8183 VDD.n2419 VDD.n2418 92.5005
R8184 VDD.n2225 VDD.n1780 92.5005
R8185 VDD.n1782 VDD.n1780 92.5005
R8186 VDD.n2223 VDD.n2222 92.5005
R8187 VDD.n2222 VDD.n2221 92.5005
R8188 VDD.n1798 VDD.n1787 92.5005
R8189 VDD.n1795 VDD.n1787 92.5005
R8190 VDD.n2214 VDD.n2213 92.5005
R8191 VDD.n2215 VDD.n2214 92.5005
R8192 VDD.n2211 VDD.n1797 92.5005
R8193 VDD.n1804 VDD.n1797 92.5005
R8194 VDD.n2199 VDD.n2198 92.5005
R8195 VDD.n2198 VDD.n1872 92.5005
R8196 VDD.n2197 VDD.n1886 92.5005
R8197 VDD.n2197 VDD.n2196 92.5005
R8198 VDD.n2156 VDD.n1884 92.5005
R8199 VDD.n2158 VDD.n1884 92.5005
R8200 VDD.n2189 VDD.n2188 92.5005
R8201 VDD.n2190 VDD.n2189 92.5005
R8202 VDD.n2187 VDD.n2155 92.5005
R8203 VDD.n2169 VDD.n2155 92.5005
R8204 VDD.n2154 VDD.n1645 92.5005
R8205 VDD.n2154 VDD.n1648 92.5005
R8206 VDD.n2230 VDD.n1781 92.5005
R8207 VDD.n2230 VDD.n2229 92.5005
R8208 VDD.n1268 VDD.n1267 92.5005
R8209 VDD.n878 VDD.n877 92.5005
R8210 VDD.n876 VDD.n875 92.5005
R8211 VDD.n874 VDD.n873 92.5005
R8212 VDD.n872 VDD.n871 92.5005
R8213 VDD.n870 VDD.n869 92.5005
R8214 VDD.n868 VDD.n867 92.5005
R8215 VDD.n858 VDD.n857 92.5005
R8216 VDD.n1232 VDD.n1231 92.5005
R8217 VDD.n1235 VDD.n1234 92.5005
R8218 VDD.n1237 VDD.n1236 92.5005
R8219 VDD.n1243 VDD.n1242 92.5005
R8220 VDD.n861 VDD.n860 92.5005
R8221 VDD.n865 VDD.n864 92.5005
R8222 VDD.n863 VDD.n862 92.5005
R8223 VDD.n1262 VDD.n1261 92.5005
R8224 VDD.n1264 VDD.n1263 92.5005
R8225 VDD.n1266 VDD.n1265 92.5005
R8226 VDD.n1507 VDD.n1506 92.5005
R8227 VDD.n1506 VDD.n1505 92.5005
R8228 VDD.n1474 VDD.n1473 92.5005
R8229 VDD.n1473 VDD.n1472 92.5005
R8230 VDD.n1477 VDD.n1476 92.5005
R8231 VDD.n1476 VDD.n1475 92.5005
R8232 VDD.n1480 VDD.n1479 92.5005
R8233 VDD.n1479 VDD.n1478 92.5005
R8234 VDD.n1483 VDD.n1482 92.5005
R8235 VDD.n1482 VDD.n1481 92.5005
R8236 VDD.n1486 VDD.n1485 92.5005
R8237 VDD.n1485 VDD.n1484 92.5005
R8238 VDD.n1489 VDD.n1488 92.5005
R8239 VDD.n1488 VDD.n1487 92.5005
R8240 VDD.n1492 VDD.n1491 92.5005
R8241 VDD.n1491 VDD.n1490 92.5005
R8242 VDD.n1495 VDD.n1494 92.5005
R8243 VDD.n1494 VDD.n1493 92.5005
R8244 VDD.n1498 VDD.n1497 92.5005
R8245 VDD.n1497 VDD.n1496 92.5005
R8246 VDD.n1501 VDD.n1500 92.5005
R8247 VDD.n1500 VDD.n1499 92.5005
R8248 VDD.n1504 VDD.n1503 92.5005
R8249 VDD.n1503 VDD.n1502 92.5005
R8250 VDD.n1471 VDD.n1470 92.5005
R8251 VDD.n1470 VDD.n1469 92.5005
R8252 VDD.n1468 VDD.n1467 92.5005
R8253 VDD.n1467 VDD.n1466 92.5005
R8254 VDD.n1465 VDD.n1464 92.5005
R8255 VDD.n1461 VDD.n1460 92.5005
R8256 VDD.n1459 VDD.n1458 92.5005
R8257 VDD.n1453 VDD.n1452 92.5005
R8258 VDD.n1452 VDD.n1451 92.5005
R8259 VDD.n1450 VDD.n1449 92.5005
R8260 VDD.n1449 VDD.n1448 92.5005
R8261 VDD.n1447 VDD.n1446 92.5005
R8262 VDD.n1446 VDD.n1445 92.5005
R8263 VDD.n1444 VDD.n1443 92.5005
R8264 VDD.n1443 VDD.n1442 92.5005
R8265 VDD.n1441 VDD.n1440 92.5005
R8266 VDD.n1440 VDD.n1439 92.5005
R8267 VDD.n1438 VDD.n1437 92.5005
R8268 VDD.n1437 VDD.n1436 92.5005
R8269 VDD.n1435 VDD.n1434 92.5005
R8270 VDD.n1434 VDD.n1433 92.5005
R8271 VDD.n1432 VDD.n1431 92.5005
R8272 VDD.n1431 VDD.n1430 92.5005
R8273 VDD.n1429 VDD.n1428 92.5005
R8274 VDD.n1428 VDD.n1427 92.5005
R8275 VDD.n1426 VDD.n1425 92.5005
R8276 VDD.n1425 VDD.n1424 92.5005
R8277 VDD.n1423 VDD.n1422 92.5005
R8278 VDD.n1422 VDD.n1421 92.5005
R8279 VDD.n1420 VDD.n1419 92.5005
R8280 VDD.n1419 VDD.n1418 92.5005
R8281 VDD.n1417 VDD.n1416 92.5005
R8282 VDD.n1416 VDD.n1415 92.5005
R8283 VDD.n1029 VDD.n1028 92.5005
R8284 VDD.n1028 VDD.n1027 92.5005
R8285 VDD.n1032 VDD.n1031 92.5005
R8286 VDD.n1031 VDD.n1030 92.5005
R8287 VDD.n1035 VDD.n1034 92.5005
R8288 VDD.n1034 VDD.n1033 92.5005
R8289 VDD.n1038 VDD.n1037 92.5005
R8290 VDD.n1037 VDD.n1036 92.5005
R8291 VDD.n1041 VDD.n1040 92.5005
R8292 VDD.n1040 VDD.n1039 92.5005
R8293 VDD.n1044 VDD.n1043 92.5005
R8294 VDD.n1043 VDD.n1042 92.5005
R8295 VDD.n1047 VDD.n1046 92.5005
R8296 VDD.n1046 VDD.n1045 92.5005
R8297 VDD.n1050 VDD.n1049 92.5005
R8298 VDD.n1049 VDD.n1048 92.5005
R8299 VDD.n1053 VDD.n1052 92.5005
R8300 VDD.n1052 VDD.n1051 92.5005
R8301 VDD.n1056 VDD.n1055 92.5005
R8302 VDD.n1055 VDD.n1054 92.5005
R8303 VDD.n1059 VDD.n1058 92.5005
R8304 VDD.n1058 VDD.n1057 92.5005
R8305 VDD.n1062 VDD.n1061 92.5005
R8306 VDD.n1061 VDD.n1060 92.5005
R8307 VDD.n1065 VDD.n1064 92.5005
R8308 VDD.n1064 VDD.n1063 92.5005
R8309 VDD.n1068 VDD.n1067 92.5005
R8310 VDD.n1067 VDD.n1066 92.5005
R8311 VDD.n1072 VDD.n1071 92.5005
R8312 VDD.n1071 VDD.n1070 92.5005
R8313 VDD.n1457 VDD.n1456 92.5005
R8314 VDD.n1456 VDD.n1455 92.5005
R8315 VDD.n1092 VDD.n1091 92.5005
R8316 VDD.n1091 VDD.n1090 92.5005
R8317 VDD.n1095 VDD.n1094 92.5005
R8318 VDD.n1094 VDD.n1093 92.5005
R8319 VDD.n1098 VDD.n1097 92.5005
R8320 VDD.n1097 VDD.n1096 92.5005
R8321 VDD.n1101 VDD.n1100 92.5005
R8322 VDD.n1100 VDD.n1099 92.5005
R8323 VDD.n1104 VDD.n1103 92.5005
R8324 VDD.n1103 VDD.n1102 92.5005
R8325 VDD.n1107 VDD.n1106 92.5005
R8326 VDD.n1106 VDD.n1105 92.5005
R8327 VDD.n1110 VDD.n1109 92.5005
R8328 VDD.n1109 VDD.n1108 92.5005
R8329 VDD.n1113 VDD.n1112 92.5005
R8330 VDD.n1112 VDD.n1111 92.5005
R8331 VDD.n1116 VDD.n1115 92.5005
R8332 VDD.n1115 VDD.n1114 92.5005
R8333 VDD.n1119 VDD.n1118 92.5005
R8334 VDD.n1118 VDD.n1117 92.5005
R8335 VDD.n1122 VDD.n1121 92.5005
R8336 VDD.n1121 VDD.n1120 92.5005
R8337 VDD.n1086 VDD.n1085 92.5005
R8338 VDD.n1085 VDD.n1084 92.5005
R8339 VDD.n1083 VDD.n1082 92.5005
R8340 VDD.n1082 VDD.n1081 92.5005
R8341 VDD.n1080 VDD.n1079 92.5005
R8342 VDD.n1076 VDD.n1075 92.5005
R8343 VDD.n1074 VDD.n1073 92.5005
R8344 VDD.n1089 VDD.n1088 92.5005
R8345 VDD.n1088 VDD.n1087 92.5005
R8346 VDD.n1124 VDD.n1123 92.5005
R8347 VDD.n1187 VDD.n1186 92.5005
R8348 VDD.n1180 VDD.n1179 92.5005
R8349 VDD.n1175 VDD.n1174 92.5005
R8350 VDD.n1170 VDD.n1169 92.5005
R8351 VDD.n1165 VDD.n1164 92.5005
R8352 VDD.n1160 VDD.n1159 92.5005
R8353 VDD.n1155 VDD.n1154 92.5005
R8354 VDD.n1153 VDD.n1152 92.5005
R8355 VDD.n1189 VDD.n1188 92.5005
R8356 VDD.n1200 VDD.n1199 92.5005
R8357 VDD.n1026 VDD.n1025 92.5005
R8358 VDD.n986 VDD.n985 92.5005
R8359 VDD.n991 VDD.n990 92.5005
R8360 VDD.n996 VDD.n995 92.5005
R8361 VDD.n1001 VDD.n1000 92.5005
R8362 VDD.n1007 VDD.n1006 92.5005
R8363 VDD.n1013 VDD.n1012 92.5005
R8364 VDD.n1011 VDD.n1010 92.5005
R8365 VDD.n1004 VDD.n1003 92.5005
R8366 VDD.n999 VDD.n998 92.5005
R8367 VDD.n993 VDD.n992 92.5005
R8368 VDD.n989 VDD.n988 92.5005
R8369 VDD.n980 VDD.n979 92.5005
R8370 VDD.n983 VDD.n982 92.5005
R8371 VDD.n1015 VDD.n1014 92.5005
R8372 VDD.n1020 VDD.n1019 92.5005
R8373 VDD.n1023 VDD.n1022 92.5005
R8374 VDD.n881 VDD.n880 92.5005
R8375 VDD.n926 VDD.n925 92.5005
R8376 VDD.n929 VDD.n928 92.5005
R8377 VDD.n931 VDD.n930 92.5005
R8378 VDD.n935 VDD.n934 92.5005
R8379 VDD.n938 VDD.n937 92.5005
R8380 VDD.n937 VDD.n936 92.5005
R8381 VDD.n941 VDD.n940 92.5005
R8382 VDD.n940 VDD.n939 92.5005
R8383 VDD.n944 VDD.n943 92.5005
R8384 VDD.n943 VDD.n942 92.5005
R8385 VDD.n947 VDD.n946 92.5005
R8386 VDD.n946 VDD.n945 92.5005
R8387 VDD.n950 VDD.n949 92.5005
R8388 VDD.n949 VDD.n948 92.5005
R8389 VDD.n953 VDD.n952 92.5005
R8390 VDD.n952 VDD.n951 92.5005
R8391 VDD.n956 VDD.n955 92.5005
R8392 VDD.n955 VDD.n954 92.5005
R8393 VDD.n959 VDD.n958 92.5005
R8394 VDD.n958 VDD.n957 92.5005
R8395 VDD.n962 VDD.n961 92.5005
R8396 VDD.n961 VDD.n960 92.5005
R8397 VDD.n965 VDD.n964 92.5005
R8398 VDD.n964 VDD.n963 92.5005
R8399 VDD.n968 VDD.n967 92.5005
R8400 VDD.n967 VDD.n966 92.5005
R8401 VDD.n971 VDD.n970 92.5005
R8402 VDD.n970 VDD.n969 92.5005
R8403 VDD.n974 VDD.n973 92.5005
R8404 VDD.n973 VDD.n972 92.5005
R8405 VDD.n977 VDD.n976 92.5005
R8406 VDD.n976 VDD.n975 92.5005
R8407 VDD.n1304 VDD.n1303 92.5005
R8408 VDD.n1303 VDD.n1302 92.5005
R8409 VDD.n1301 VDD.n1300 92.5005
R8410 VDD.n1300 VDD.n1299 92.5005
R8411 VDD.n1298 VDD.n1297 92.5005
R8412 VDD.n1297 VDD.n1296 92.5005
R8413 VDD.n1295 VDD.n1294 92.5005
R8414 VDD.n1294 VDD.n1293 92.5005
R8415 VDD.n1292 VDD.n1291 92.5005
R8416 VDD.n1291 VDD.n1290 92.5005
R8417 VDD.n1289 VDD.n1288 92.5005
R8418 VDD.n1288 VDD.n1287 92.5005
R8419 VDD.n1286 VDD.n1285 92.5005
R8420 VDD.n1285 VDD.n1284 92.5005
R8421 VDD.n1283 VDD.n1282 92.5005
R8422 VDD.n1282 VDD.n1281 92.5005
R8423 VDD.n1280 VDD.n1279 92.5005
R8424 VDD.n1279 VDD.n1278 92.5005
R8425 VDD.n1277 VDD.n1276 92.5005
R8426 VDD.n1276 VDD.n1275 92.5005
R8427 VDD.n1274 VDD.n1273 92.5005
R8428 VDD.n1273 VDD.n1272 92.5005
R8429 VDD.n1271 VDD.n1270 92.5005
R8430 VDD.n1270 VDD.n1269 92.5005
R8431 VDD.n884 VDD.n883 92.5005
R8432 VDD.n883 VDD.n882 92.5005
R8433 VDD.n887 VDD.n886 92.5005
R8434 VDD.n886 VDD.n885 92.5005
R8435 VDD.n890 VDD.n889 92.5005
R8436 VDD.n889 VDD.n888 92.5005
R8437 VDD.n893 VDD.n892 92.5005
R8438 VDD.n892 VDD.n891 92.5005
R8439 VDD.n896 VDD.n895 92.5005
R8440 VDD.n895 VDD.n894 92.5005
R8441 VDD.n899 VDD.n898 92.5005
R8442 VDD.n898 VDD.n897 92.5005
R8443 VDD.n902 VDD.n901 92.5005
R8444 VDD.n901 VDD.n900 92.5005
R8445 VDD.n905 VDD.n904 92.5005
R8446 VDD.n904 VDD.n903 92.5005
R8447 VDD.n908 VDD.n907 92.5005
R8448 VDD.n907 VDD.n906 92.5005
R8449 VDD.n911 VDD.n910 92.5005
R8450 VDD.n910 VDD.n909 92.5005
R8451 VDD.n914 VDD.n913 92.5005
R8452 VDD.n913 VDD.n912 92.5005
R8453 VDD.n917 VDD.n916 92.5005
R8454 VDD.n916 VDD.n915 92.5005
R8455 VDD.n920 VDD.n919 92.5005
R8456 VDD.n919 VDD.n918 92.5005
R8457 VDD.n923 VDD.n922 92.5005
R8458 VDD.n922 VDD.n921 92.5005
R8459 VDD.n1314 VDD.n1313 92.5005
R8460 VDD.n1307 VDD.n1306 92.5005
R8461 VDD.n1309 VDD.n1308 92.5005
R8462 VDD.n1365 VDD.n1364 92.5005
R8463 VDD.n1364 VDD.n1363 92.5005
R8464 VDD.n1362 VDD.n1361 92.5005
R8465 VDD.n1361 VDD.n1360 92.5005
R8466 VDD.n1359 VDD.n1358 92.5005
R8467 VDD.n1358 VDD.n1357 92.5005
R8468 VDD.n1356 VDD.n1355 92.5005
R8469 VDD.n1355 VDD.n1354 92.5005
R8470 VDD.n1353 VDD.n1352 92.5005
R8471 VDD.n1352 VDD.n1351 92.5005
R8472 VDD.n1350 VDD.n1349 92.5005
R8473 VDD.n1349 VDD.n1348 92.5005
R8474 VDD.n1347 VDD.n1346 92.5005
R8475 VDD.n1346 VDD.n1345 92.5005
R8476 VDD.n1344 VDD.n1343 92.5005
R8477 VDD.n1343 VDD.n1342 92.5005
R8478 VDD.n1341 VDD.n1340 92.5005
R8479 VDD.n1340 VDD.n1339 92.5005
R8480 VDD.n1338 VDD.n1337 92.5005
R8481 VDD.n1337 VDD.n1336 92.5005
R8482 VDD.n1335 VDD.n1334 92.5005
R8483 VDD.n1334 VDD.n1333 92.5005
R8484 VDD.n1332 VDD.n1331 92.5005
R8485 VDD.n1331 VDD.n1330 92.5005
R8486 VDD.n1329 VDD.n1328 92.5005
R8487 VDD.n1328 VDD.n1327 92.5005
R8488 VDD.n1326 VDD.n1325 92.5005
R8489 VDD.n1325 VDD.n1324 92.5005
R8490 VDD.n1323 VDD.n1322 92.5005
R8491 VDD.n1319 VDD.n1318 92.5005
R8492 VDD.n1316 VDD.n1315 92.5005
R8493 VDD.n1510 VDD.n1509 92.5005
R8494 VDD.n1527 VDD.n1526 92.5005
R8495 VDD.n1530 VDD.n1529 92.5005
R8496 VDD.n1535 VDD.n1534 92.5005
R8497 VDD.n1541 VDD.n1540 92.5005
R8498 VDD.n1546 VDD.n1545 92.5005
R8499 VDD.n1552 VDD.n1551 92.5005
R8500 VDD.n1557 VDD.n1556 92.5005
R8501 VDD.n1563 VDD.n1562 92.5005
R8502 VDD.n1566 VDD.n1565 92.5005
R8503 VDD.n1401 VDD.n1400 92.5005
R8504 VDD.n1396 VDD.n1395 92.5005
R8505 VDD.n1390 VDD.n1389 92.5005
R8506 VDD.n1385 VDD.n1384 92.5005
R8507 VDD.n1379 VDD.n1378 92.5005
R8508 VDD.n1374 VDD.n1373 92.5005
R8509 VDD.n1371 VDD.n1370 92.5005
R8510 VDD.n1368 VDD.n1367 92.5005
R8511 VDD.n1376 VDD.n1375 92.5005
R8512 VDD.n1382 VDD.n1381 92.5005
R8513 VDD.n1387 VDD.n1386 92.5005
R8514 VDD.n1393 VDD.n1392 92.5005
R8515 VDD.n1398 VDD.n1397 92.5005
R8516 VDD.n1407 VDD.n1406 92.5005
R8517 VDD.n1405 VDD.n1404 92.5005
R8518 VDD.n1409 VDD.n1408 92.5005
R8519 VDD.n1414 VDD.n1413 92.5005
R8520 VDD.n1569 VDD.n1568 92.5005
R8521 VDD.n1560 VDD.n1559 92.5005
R8522 VDD.n1532 VDD.n1531 92.5005
R8523 VDD.n1538 VDD.n1537 92.5005
R8524 VDD.n1543 VDD.n1542 92.5005
R8525 VDD.n1549 VDD.n1548 92.5005
R8526 VDD.n1554 VDD.n1553 92.5005
R8527 VDD.n1191 VDD.n1190 92.5005
R8528 VDD.n1193 VDD.n1192 92.5005
R8529 VDD.n1197 VDD.n1196 92.5005
R8530 VDD.n1196 VDD.n1195 92.5005
R8531 VDD.n1177 VDD.n1176 92.5005
R8532 VDD.n1173 VDD.n1172 92.5005
R8533 VDD.n1167 VDD.n1166 92.5005
R8534 VDD.n1163 VDD.n1162 92.5005
R8535 VDD.n1157 VDD.n1156 92.5005
R8536 VDD.n1184 VDD.n1183 92.5005
R8537 VDD.n1130 VDD.n1129 92.5005
R8538 VDD.n1126 VDD.n1125 92.5005
R8539 VDD.n1203 VDD.n1202 92.5005
R8540 VDD.n1206 VDD.n1205 92.5005
R8541 VDD.n1209 VDD.n1208 92.5005
R8542 VDD.n1214 VDD.n1213 92.5005
R8543 VDD.n1149 VDD.n1148 92.5005
R8544 VDD.n1147 VDD.n1146 92.5005
R8545 VDD.n1145 VDD.n1144 92.5005
R8546 VDD.n1143 VDD.n1142 92.5005
R8547 VDD.n1140 VDD.n1139 92.5005
R8548 VDD.n1138 VDD.n1137 92.5005
R8549 VDD.n1136 VDD.n1135 92.5005
R8550 VDD.n1134 VDD.n1133 92.5005
R8551 VDD.n1132 VDD.n1131 92.5005
R8552 VDD.n1512 VDD.n1511 92.5005
R8553 VDD.n1518 VDD.n1517 92.5005
R8554 VDD.n1520 VDD.n1519 92.5005
R8555 VDD.n1522 VDD.n1521 92.5005
R8556 VDD.n1524 VDD.n1523 92.5005
R8557 VDD.n1515 VDD.n1514 92.5005
R8558 VDD.n1245 VDD.n1244 92.5005
R8559 VDD.n1248 VDD.n1247 92.5005
R8560 VDD.n1251 VDD.n1250 92.5005
R8561 VDD.n1254 VDD.n1253 92.5005
R8562 VDD.n1260 VDD.n1259 92.5005
R8563 VDD.n1573 VDD.n1572 92.5005
R8564 VDD.n1572 VDD.n1571 92.5005
R8565 VDD.n1579 VDD.n1578 92.5005
R8566 VDD.n1578 VDD.n1577 92.5005
R8567 VDD.n1585 VDD.n1584 92.5005
R8568 VDD.n1584 VDD.n1583 92.5005
R8569 VDD.n1591 VDD.n1590 92.5005
R8570 VDD.n1590 VDD.n1589 92.5005
R8571 VDD.n1604 VDD.n1603 92.5005
R8572 VDD.n1603 VDD.n1602 92.5005
R8573 VDD.n1608 VDD.n1607 92.5005
R8574 VDD.n1607 VDD.n1606 92.5005
R8575 VDD.n1613 VDD.n1612 92.5005
R8576 VDD.n1612 VDD.n1611 92.5005
R8577 VDD.n1634 VDD.n1633 92.5005
R8578 VDD.n1633 VDD.n1632 92.5005
R8579 VDD.n1628 VDD.n1627 92.5005
R8580 VDD.n1627 VDD.n1626 92.5005
R8581 VDD.n1622 VDD.n1621 92.5005
R8582 VDD.n1621 VDD.n1620 92.5005
R8583 VDD.n1224 VDD.n1223 92.5005
R8584 VDD.n1223 VDD.n1222 92.5005
R8585 VDD.n1582 VDD.n1581 92.5005
R8586 VDD.n1581 VDD.n1580 92.5005
R8587 VDD.n1588 VDD.n1587 92.5005
R8588 VDD.n1587 VDD.n1586 92.5005
R8589 VDD.n1594 VDD.n1593 92.5005
R8590 VDD.n1593 VDD.n1592 92.5005
R8591 VDD.n1597 VDD.n1596 92.5005
R8592 VDD.n1596 VDD.n1595 92.5005
R8593 VDD.n1601 VDD.n1600 92.5005
R8594 VDD.n1600 VDD.n1599 92.5005
R8595 VDD.n1616 VDD.n1615 92.5005
R8596 VDD.n1615 VDD.n1614 92.5005
R8597 VDD.n1631 VDD.n1630 92.5005
R8598 VDD.n1630 VDD.n1629 92.5005
R8599 VDD.n1625 VDD.n1624 92.5005
R8600 VDD.n1624 VDD.n1623 92.5005
R8601 VDD.n1619 VDD.n1618 92.5005
R8602 VDD.n1618 VDD.n1617 92.5005
R8603 VDD.n1217 VDD.n1216 92.5005
R8604 VDD.n1216 VDD.n1215 92.5005
R8605 VDD.n1221 VDD.n1220 92.5005
R8606 VDD.n1220 VDD.n1219 92.5005
R8607 VDD.n1576 VDD.n1575 92.5005
R8608 VDD.n1575 VDD.n1574 92.5005
R8609 VDD.n40 VDD.n39 92.5005
R8610 VDD.n432 VDD.n431 92.5005
R8611 VDD.n430 VDD.n429 92.5005
R8612 VDD.n428 VDD.n427 92.5005
R8613 VDD.n426 VDD.n425 92.5005
R8614 VDD.n424 VDD.n423 92.5005
R8615 VDD.n422 VDD.n421 92.5005
R8616 VDD.n412 VDD.n411 92.5005
R8617 VDD.n4 VDD.n3 92.5005
R8618 VDD.n7 VDD.n6 92.5005
R8619 VDD.n9 VDD.n8 92.5005
R8620 VDD.n15 VDD.n14 92.5005
R8621 VDD.n415 VDD.n414 92.5005
R8622 VDD.n419 VDD.n418 92.5005
R8623 VDD.n417 VDD.n416 92.5005
R8624 VDD.n34 VDD.n33 92.5005
R8625 VDD.n36 VDD.n35 92.5005
R8626 VDD.n38 VDD.n37 92.5005
R8627 VDD.n279 VDD.n278 92.5005
R8628 VDD.n278 VDD.n277 92.5005
R8629 VDD.n246 VDD.n245 92.5005
R8630 VDD.n245 VDD.n244 92.5005
R8631 VDD.n249 VDD.n248 92.5005
R8632 VDD.n248 VDD.n247 92.5005
R8633 VDD.n252 VDD.n251 92.5005
R8634 VDD.n251 VDD.n250 92.5005
R8635 VDD.n255 VDD.n254 92.5005
R8636 VDD.n254 VDD.n253 92.5005
R8637 VDD.n258 VDD.n257 92.5005
R8638 VDD.n257 VDD.n256 92.5005
R8639 VDD.n261 VDD.n260 92.5005
R8640 VDD.n260 VDD.n259 92.5005
R8641 VDD.n264 VDD.n263 92.5005
R8642 VDD.n263 VDD.n262 92.5005
R8643 VDD.n267 VDD.n266 92.5005
R8644 VDD.n266 VDD.n265 92.5005
R8645 VDD.n270 VDD.n269 92.5005
R8646 VDD.n269 VDD.n268 92.5005
R8647 VDD.n273 VDD.n272 92.5005
R8648 VDD.n272 VDD.n271 92.5005
R8649 VDD.n276 VDD.n275 92.5005
R8650 VDD.n275 VDD.n274 92.5005
R8651 VDD.n243 VDD.n242 92.5005
R8652 VDD.n242 VDD.n241 92.5005
R8653 VDD.n240 VDD.n239 92.5005
R8654 VDD.n239 VDD.n238 92.5005
R8655 VDD.n237 VDD.n236 92.5005
R8656 VDD.n233 VDD.n232 92.5005
R8657 VDD.n231 VDD.n230 92.5005
R8658 VDD.n225 VDD.n224 92.5005
R8659 VDD.n224 VDD.n223 92.5005
R8660 VDD.n222 VDD.n221 92.5005
R8661 VDD.n221 VDD.n220 92.5005
R8662 VDD.n219 VDD.n218 92.5005
R8663 VDD.n218 VDD.n217 92.5005
R8664 VDD.n216 VDD.n215 92.5005
R8665 VDD.n215 VDD.n214 92.5005
R8666 VDD.n213 VDD.n212 92.5005
R8667 VDD.n212 VDD.n211 92.5005
R8668 VDD.n210 VDD.n209 92.5005
R8669 VDD.n209 VDD.n208 92.5005
R8670 VDD.n207 VDD.n206 92.5005
R8671 VDD.n206 VDD.n205 92.5005
R8672 VDD.n204 VDD.n203 92.5005
R8673 VDD.n203 VDD.n202 92.5005
R8674 VDD.n201 VDD.n200 92.5005
R8675 VDD.n200 VDD.n199 92.5005
R8676 VDD.n198 VDD.n197 92.5005
R8677 VDD.n197 VDD.n196 92.5005
R8678 VDD.n195 VDD.n194 92.5005
R8679 VDD.n194 VDD.n193 92.5005
R8680 VDD.n192 VDD.n191 92.5005
R8681 VDD.n191 VDD.n190 92.5005
R8682 VDD.n189 VDD.n188 92.5005
R8683 VDD.n188 VDD.n187 92.5005
R8684 VDD.n583 VDD.n582 92.5005
R8685 VDD.n582 VDD.n581 92.5005
R8686 VDD.n586 VDD.n585 92.5005
R8687 VDD.n585 VDD.n584 92.5005
R8688 VDD.n589 VDD.n588 92.5005
R8689 VDD.n588 VDD.n587 92.5005
R8690 VDD.n592 VDD.n591 92.5005
R8691 VDD.n591 VDD.n590 92.5005
R8692 VDD.n595 VDD.n594 92.5005
R8693 VDD.n594 VDD.n593 92.5005
R8694 VDD.n598 VDD.n597 92.5005
R8695 VDD.n597 VDD.n596 92.5005
R8696 VDD.n601 VDD.n600 92.5005
R8697 VDD.n600 VDD.n599 92.5005
R8698 VDD.n604 VDD.n603 92.5005
R8699 VDD.n603 VDD.n602 92.5005
R8700 VDD.n607 VDD.n606 92.5005
R8701 VDD.n606 VDD.n605 92.5005
R8702 VDD.n610 VDD.n609 92.5005
R8703 VDD.n609 VDD.n608 92.5005
R8704 VDD.n613 VDD.n612 92.5005
R8705 VDD.n612 VDD.n611 92.5005
R8706 VDD.n616 VDD.n615 92.5005
R8707 VDD.n615 VDD.n614 92.5005
R8708 VDD.n619 VDD.n618 92.5005
R8709 VDD.n618 VDD.n617 92.5005
R8710 VDD.n622 VDD.n621 92.5005
R8711 VDD.n621 VDD.n620 92.5005
R8712 VDD.n626 VDD.n625 92.5005
R8713 VDD.n625 VDD.n624 92.5005
R8714 VDD.n229 VDD.n228 92.5005
R8715 VDD.n228 VDD.n227 92.5005
R8716 VDD.n646 VDD.n645 92.5005
R8717 VDD.n645 VDD.n644 92.5005
R8718 VDD.n649 VDD.n648 92.5005
R8719 VDD.n648 VDD.n647 92.5005
R8720 VDD.n652 VDD.n651 92.5005
R8721 VDD.n651 VDD.n650 92.5005
R8722 VDD.n655 VDD.n654 92.5005
R8723 VDD.n654 VDD.n653 92.5005
R8724 VDD.n658 VDD.n657 92.5005
R8725 VDD.n657 VDD.n656 92.5005
R8726 VDD.n661 VDD.n660 92.5005
R8727 VDD.n660 VDD.n659 92.5005
R8728 VDD.n664 VDD.n663 92.5005
R8729 VDD.n663 VDD.n662 92.5005
R8730 VDD.n667 VDD.n666 92.5005
R8731 VDD.n666 VDD.n665 92.5005
R8732 VDD.n670 VDD.n669 92.5005
R8733 VDD.n669 VDD.n668 92.5005
R8734 VDD.n673 VDD.n672 92.5005
R8735 VDD.n672 VDD.n671 92.5005
R8736 VDD.n676 VDD.n675 92.5005
R8737 VDD.n675 VDD.n674 92.5005
R8738 VDD.n640 VDD.n639 92.5005
R8739 VDD.n639 VDD.n638 92.5005
R8740 VDD.n637 VDD.n636 92.5005
R8741 VDD.n636 VDD.n635 92.5005
R8742 VDD.n634 VDD.n633 92.5005
R8743 VDD.n630 VDD.n629 92.5005
R8744 VDD.n628 VDD.n627 92.5005
R8745 VDD.n643 VDD.n642 92.5005
R8746 VDD.n642 VDD.n641 92.5005
R8747 VDD.n678 VDD.n677 92.5005
R8748 VDD.n741 VDD.n740 92.5005
R8749 VDD.n734 VDD.n733 92.5005
R8750 VDD.n729 VDD.n728 92.5005
R8751 VDD.n724 VDD.n723 92.5005
R8752 VDD.n719 VDD.n718 92.5005
R8753 VDD.n714 VDD.n713 92.5005
R8754 VDD.n709 VDD.n708 92.5005
R8755 VDD.n707 VDD.n706 92.5005
R8756 VDD.n743 VDD.n742 92.5005
R8757 VDD.n754 VDD.n753 92.5005
R8758 VDD.n580 VDD.n579 92.5005
R8759 VDD.n540 VDD.n539 92.5005
R8760 VDD.n545 VDD.n544 92.5005
R8761 VDD.n550 VDD.n549 92.5005
R8762 VDD.n555 VDD.n554 92.5005
R8763 VDD.n561 VDD.n560 92.5005
R8764 VDD.n567 VDD.n566 92.5005
R8765 VDD.n565 VDD.n564 92.5005
R8766 VDD.n558 VDD.n557 92.5005
R8767 VDD.n553 VDD.n552 92.5005
R8768 VDD.n547 VDD.n546 92.5005
R8769 VDD.n543 VDD.n542 92.5005
R8770 VDD.n534 VDD.n533 92.5005
R8771 VDD.n537 VDD.n536 92.5005
R8772 VDD.n569 VDD.n568 92.5005
R8773 VDD.n574 VDD.n573 92.5005
R8774 VDD.n577 VDD.n576 92.5005
R8775 VDD.n435 VDD.n434 92.5005
R8776 VDD.n480 VDD.n479 92.5005
R8777 VDD.n483 VDD.n482 92.5005
R8778 VDD.n485 VDD.n484 92.5005
R8779 VDD.n489 VDD.n488 92.5005
R8780 VDD.n492 VDD.n491 92.5005
R8781 VDD.n491 VDD.n490 92.5005
R8782 VDD.n495 VDD.n494 92.5005
R8783 VDD.n494 VDD.n493 92.5005
R8784 VDD.n498 VDD.n497 92.5005
R8785 VDD.n497 VDD.n496 92.5005
R8786 VDD.n501 VDD.n500 92.5005
R8787 VDD.n500 VDD.n499 92.5005
R8788 VDD.n504 VDD.n503 92.5005
R8789 VDD.n503 VDD.n502 92.5005
R8790 VDD.n507 VDD.n506 92.5005
R8791 VDD.n506 VDD.n505 92.5005
R8792 VDD.n510 VDD.n509 92.5005
R8793 VDD.n509 VDD.n508 92.5005
R8794 VDD.n513 VDD.n512 92.5005
R8795 VDD.n512 VDD.n511 92.5005
R8796 VDD.n516 VDD.n515 92.5005
R8797 VDD.n515 VDD.n514 92.5005
R8798 VDD.n519 VDD.n518 92.5005
R8799 VDD.n518 VDD.n517 92.5005
R8800 VDD.n522 VDD.n521 92.5005
R8801 VDD.n521 VDD.n520 92.5005
R8802 VDD.n525 VDD.n524 92.5005
R8803 VDD.n524 VDD.n523 92.5005
R8804 VDD.n528 VDD.n527 92.5005
R8805 VDD.n527 VDD.n526 92.5005
R8806 VDD.n531 VDD.n530 92.5005
R8807 VDD.n530 VDD.n529 92.5005
R8808 VDD.n76 VDD.n75 92.5005
R8809 VDD.n75 VDD.n74 92.5005
R8810 VDD.n73 VDD.n72 92.5005
R8811 VDD.n72 VDD.n71 92.5005
R8812 VDD.n70 VDD.n69 92.5005
R8813 VDD.n69 VDD.n68 92.5005
R8814 VDD.n67 VDD.n66 92.5005
R8815 VDD.n66 VDD.n65 92.5005
R8816 VDD.n64 VDD.n63 92.5005
R8817 VDD.n63 VDD.n62 92.5005
R8818 VDD.n61 VDD.n60 92.5005
R8819 VDD.n60 VDD.n59 92.5005
R8820 VDD.n58 VDD.n57 92.5005
R8821 VDD.n57 VDD.n56 92.5005
R8822 VDD.n55 VDD.n54 92.5005
R8823 VDD.n54 VDD.n53 92.5005
R8824 VDD.n52 VDD.n51 92.5005
R8825 VDD.n51 VDD.n50 92.5005
R8826 VDD.n49 VDD.n48 92.5005
R8827 VDD.n48 VDD.n47 92.5005
R8828 VDD.n46 VDD.n45 92.5005
R8829 VDD.n45 VDD.n44 92.5005
R8830 VDD.n43 VDD.n42 92.5005
R8831 VDD.n42 VDD.n41 92.5005
R8832 VDD.n438 VDD.n437 92.5005
R8833 VDD.n437 VDD.n436 92.5005
R8834 VDD.n441 VDD.n440 92.5005
R8835 VDD.n440 VDD.n439 92.5005
R8836 VDD.n444 VDD.n443 92.5005
R8837 VDD.n443 VDD.n442 92.5005
R8838 VDD.n447 VDD.n446 92.5005
R8839 VDD.n446 VDD.n445 92.5005
R8840 VDD.n450 VDD.n449 92.5005
R8841 VDD.n449 VDD.n448 92.5005
R8842 VDD.n453 VDD.n452 92.5005
R8843 VDD.n452 VDD.n451 92.5005
R8844 VDD.n456 VDD.n455 92.5005
R8845 VDD.n455 VDD.n454 92.5005
R8846 VDD.n459 VDD.n458 92.5005
R8847 VDD.n458 VDD.n457 92.5005
R8848 VDD.n462 VDD.n461 92.5005
R8849 VDD.n461 VDD.n460 92.5005
R8850 VDD.n465 VDD.n464 92.5005
R8851 VDD.n464 VDD.n463 92.5005
R8852 VDD.n468 VDD.n467 92.5005
R8853 VDD.n467 VDD.n466 92.5005
R8854 VDD.n471 VDD.n470 92.5005
R8855 VDD.n470 VDD.n469 92.5005
R8856 VDD.n474 VDD.n473 92.5005
R8857 VDD.n473 VDD.n472 92.5005
R8858 VDD.n477 VDD.n476 92.5005
R8859 VDD.n476 VDD.n475 92.5005
R8860 VDD.n86 VDD.n85 92.5005
R8861 VDD.n79 VDD.n78 92.5005
R8862 VDD.n81 VDD.n80 92.5005
R8863 VDD.n137 VDD.n136 92.5005
R8864 VDD.n136 VDD.n135 92.5005
R8865 VDD.n134 VDD.n133 92.5005
R8866 VDD.n133 VDD.n132 92.5005
R8867 VDD.n131 VDD.n130 92.5005
R8868 VDD.n130 VDD.n129 92.5005
R8869 VDD.n128 VDD.n127 92.5005
R8870 VDD.n127 VDD.n126 92.5005
R8871 VDD.n125 VDD.n124 92.5005
R8872 VDD.n124 VDD.n123 92.5005
R8873 VDD.n122 VDD.n121 92.5005
R8874 VDD.n121 VDD.n120 92.5005
R8875 VDD.n119 VDD.n118 92.5005
R8876 VDD.n118 VDD.n117 92.5005
R8877 VDD.n116 VDD.n115 92.5005
R8878 VDD.n115 VDD.n114 92.5005
R8879 VDD.n113 VDD.n112 92.5005
R8880 VDD.n112 VDD.n111 92.5005
R8881 VDD.n110 VDD.n109 92.5005
R8882 VDD.n109 VDD.n108 92.5005
R8883 VDD.n107 VDD.n106 92.5005
R8884 VDD.n106 VDD.n105 92.5005
R8885 VDD.n104 VDD.n103 92.5005
R8886 VDD.n103 VDD.n102 92.5005
R8887 VDD.n101 VDD.n100 92.5005
R8888 VDD.n100 VDD.n99 92.5005
R8889 VDD.n98 VDD.n97 92.5005
R8890 VDD.n97 VDD.n96 92.5005
R8891 VDD.n95 VDD.n94 92.5005
R8892 VDD.n91 VDD.n90 92.5005
R8893 VDD.n88 VDD.n87 92.5005
R8894 VDD.n282 VDD.n281 92.5005
R8895 VDD.n299 VDD.n298 92.5005
R8896 VDD.n302 VDD.n301 92.5005
R8897 VDD.n307 VDD.n306 92.5005
R8898 VDD.n313 VDD.n312 92.5005
R8899 VDD.n318 VDD.n317 92.5005
R8900 VDD.n324 VDD.n323 92.5005
R8901 VDD.n329 VDD.n328 92.5005
R8902 VDD.n335 VDD.n334 92.5005
R8903 VDD.n338 VDD.n337 92.5005
R8904 VDD.n173 VDD.n172 92.5005
R8905 VDD.n168 VDD.n167 92.5005
R8906 VDD.n162 VDD.n161 92.5005
R8907 VDD.n157 VDD.n156 92.5005
R8908 VDD.n151 VDD.n150 92.5005
R8909 VDD.n146 VDD.n145 92.5005
R8910 VDD.n143 VDD.n142 92.5005
R8911 VDD.n140 VDD.n139 92.5005
R8912 VDD.n148 VDD.n147 92.5005
R8913 VDD.n154 VDD.n153 92.5005
R8914 VDD.n159 VDD.n158 92.5005
R8915 VDD.n165 VDD.n164 92.5005
R8916 VDD.n170 VDD.n169 92.5005
R8917 VDD.n179 VDD.n178 92.5005
R8918 VDD.n177 VDD.n176 92.5005
R8919 VDD.n181 VDD.n180 92.5005
R8920 VDD.n186 VDD.n185 92.5005
R8921 VDD.n341 VDD.n340 92.5005
R8922 VDD.n332 VDD.n331 92.5005
R8923 VDD.n304 VDD.n303 92.5005
R8924 VDD.n310 VDD.n309 92.5005
R8925 VDD.n315 VDD.n314 92.5005
R8926 VDD.n321 VDD.n320 92.5005
R8927 VDD.n326 VDD.n325 92.5005
R8928 VDD.n745 VDD.n744 92.5005
R8929 VDD.n747 VDD.n746 92.5005
R8930 VDD.n751 VDD.n750 92.5005
R8931 VDD.n750 VDD.n749 92.5005
R8932 VDD.n731 VDD.n730 92.5005
R8933 VDD.n727 VDD.n726 92.5005
R8934 VDD.n721 VDD.n720 92.5005
R8935 VDD.n717 VDD.n716 92.5005
R8936 VDD.n711 VDD.n710 92.5005
R8937 VDD.n738 VDD.n737 92.5005
R8938 VDD.n684 VDD.n683 92.5005
R8939 VDD.n680 VDD.n679 92.5005
R8940 VDD.n757 VDD.n756 92.5005
R8941 VDD.n760 VDD.n759 92.5005
R8942 VDD.n763 VDD.n762 92.5005
R8943 VDD.n768 VDD.n767 92.5005
R8944 VDD.n703 VDD.n702 92.5005
R8945 VDD.n701 VDD.n700 92.5005
R8946 VDD.n699 VDD.n698 92.5005
R8947 VDD.n697 VDD.n696 92.5005
R8948 VDD.n694 VDD.n693 92.5005
R8949 VDD.n692 VDD.n691 92.5005
R8950 VDD.n690 VDD.n689 92.5005
R8951 VDD.n688 VDD.n687 92.5005
R8952 VDD.n686 VDD.n685 92.5005
R8953 VDD.n284 VDD.n283 92.5005
R8954 VDD.n290 VDD.n289 92.5005
R8955 VDD.n292 VDD.n291 92.5005
R8956 VDD.n294 VDD.n293 92.5005
R8957 VDD.n296 VDD.n295 92.5005
R8958 VDD.n287 VDD.n286 92.5005
R8959 VDD.n17 VDD.n16 92.5005
R8960 VDD.n20 VDD.n19 92.5005
R8961 VDD.n23 VDD.n22 92.5005
R8962 VDD.n26 VDD.n25 92.5005
R8963 VDD.n32 VDD.n31 92.5005
R8964 VDD.n345 VDD.n344 92.5005
R8965 VDD.n344 VDD.n343 92.5005
R8966 VDD.n351 VDD.n350 92.5005
R8967 VDD.n350 VDD.n349 92.5005
R8968 VDD.n357 VDD.n356 92.5005
R8969 VDD.n356 VDD.n355 92.5005
R8970 VDD.n363 VDD.n362 92.5005
R8971 VDD.n362 VDD.n361 92.5005
R8972 VDD.n376 VDD.n375 92.5005
R8973 VDD.n375 VDD.n374 92.5005
R8974 VDD.n380 VDD.n379 92.5005
R8975 VDD.n379 VDD.n378 92.5005
R8976 VDD.n385 VDD.n384 92.5005
R8977 VDD.n384 VDD.n383 92.5005
R8978 VDD.n406 VDD.n405 92.5005
R8979 VDD.n405 VDD.n404 92.5005
R8980 VDD.n400 VDD.n399 92.5005
R8981 VDD.n399 VDD.n398 92.5005
R8982 VDD.n394 VDD.n393 92.5005
R8983 VDD.n393 VDD.n392 92.5005
R8984 VDD.n778 VDD.n777 92.5005
R8985 VDD.n777 VDD.n776 92.5005
R8986 VDD.n354 VDD.n353 92.5005
R8987 VDD.n353 VDD.n352 92.5005
R8988 VDD.n360 VDD.n359 92.5005
R8989 VDD.n359 VDD.n358 92.5005
R8990 VDD.n366 VDD.n365 92.5005
R8991 VDD.n365 VDD.n364 92.5005
R8992 VDD.n369 VDD.n368 92.5005
R8993 VDD.n368 VDD.n367 92.5005
R8994 VDD.n373 VDD.n372 92.5005
R8995 VDD.n372 VDD.n371 92.5005
R8996 VDD.n388 VDD.n387 92.5005
R8997 VDD.n387 VDD.n386 92.5005
R8998 VDD.n403 VDD.n402 92.5005
R8999 VDD.n402 VDD.n401 92.5005
R9000 VDD.n397 VDD.n396 92.5005
R9001 VDD.n396 VDD.n395 92.5005
R9002 VDD.n391 VDD.n390 92.5005
R9003 VDD.n390 VDD.n389 92.5005
R9004 VDD.n771 VDD.n770 92.5005
R9005 VDD.n770 VDD.n769 92.5005
R9006 VDD.n775 VDD.n774 92.5005
R9007 VDD.n774 VDD.n773 92.5005
R9008 VDD.n348 VDD.n347 92.5005
R9009 VDD.n347 VDD.n346 92.5005
R9010 VDD.n5750 VDD.t188 91.8719
R9011 VDD.n4110 VDD.t74 91.8719
R9012 VDD.n2469 VDD.t165 91.8719
R9013 VDD.n829 VDD.t205 91.8719
R9014 VDD.n12093 VDD.n7371 90.4767
R9015 VDD.n12678 VDD.n6717 88.8476
R9016 VDD.n6743 VDD.n6742 88.8476
R9017 VDD.n12446 VDD.n12426 87.8351
R9018 VDD.n12436 VDD.n12426 86.0979
R9019 VDD.n9978 VDD.n9973 86.0424
R9020 VDD.n12433 VDD.n12426 85.2548
R9021 VDD.n5764 VDD.t14 84.4681
R9022 VDD.n4124 VDD.t12 84.4681
R9023 VDD.n2484 VDD.t162 84.4681
R9024 VDD.n844 VDD.t30 84.4681
R9025 VDD.n8196 VDD.n8103 83.4438
R9026 VDD.n6635 VDD.n6634 83.4438
R9027 VDD.n8147 VDD.n8093 83.4431
R9028 VDD.n12716 VDD.n6595 83.4431
R9029 VDD.n5750 VDD.n5749 83.1021
R9030 VDD.n4110 VDD.n4109 83.1021
R9031 VDD.n2469 VDD.n2468 83.1021
R9032 VDD.n829 VDD.n828 83.1021
R9033 VDD.n9952 VDD.n9951 82.6643
R9034 VDD.n9190 VDD.n9189 80.7889
R9035 VDD.n5739 VDD.t10 78.5582
R9036 VDD.n4099 VDD.t111 78.5582
R9037 VDD.n2458 VDD.t138 78.5582
R9038 VDD.n818 VDD.t170 78.5582
R9039 VDD.n12094 VDD.n12093 78.4132
R9040 VDD.n6250 VDD.n6249 78.4132
R9041 VDD.n6121 VDD.n5879 78.4132
R9042 VDD.n5396 VDD.n5395 78.4132
R9043 VDD.n5267 VDD.n5025 78.4132
R9044 VDD.n4610 VDD.n4609 78.4132
R9045 VDD.n4481 VDD.n4239 78.4132
R9046 VDD.n3756 VDD.n3755 78.4132
R9047 VDD.n3627 VDD.n3385 78.4132
R9048 VDD.n2970 VDD.n2969 78.4132
R9049 VDD.n2841 VDD.n2599 78.4132
R9050 VDD.n2115 VDD.n2114 78.4132
R9051 VDD.n1986 VDD.n1744 78.4132
R9052 VDD.n9220 VDD.t6 75.5912
R9053 VDD.t160 VDD.n9220 75.5912
R9054 VDD.n12248 VDD.n7070 74.6009
R9055 VDD.n7861 VDD.n7749 72.0905
R9056 VDD.n7909 VDD.n7749 72.0905
R9057 VDD.n7860 VDD.n7749 72.0905
R9058 VDD.n7855 VDD.n7749 72.0905
R9059 VDD.n7918 VDD.n7749 72.0905
R9060 VDD.n7854 VDD.n7749 72.0905
R9061 VDD.n7849 VDD.n7749 72.0905
R9062 VDD.n7927 VDD.n7749 72.0905
R9063 VDD.n7955 VDD.n7749 72.0905
R9064 VDD.n7829 VDD.n7749 72.0905
R9065 VDD.n7824 VDD.n7749 72.0905
R9066 VDD.n7964 VDD.n7749 72.0905
R9067 VDD.n7823 VDD.n7749 72.0905
R9068 VDD.n7818 VDD.n7749 72.0905
R9069 VDD.n7973 VDD.n7749 72.0905
R9070 VDD.n7817 VDD.n7749 72.0905
R9071 VDD.n5796 VDD.n5795 72.0905
R9072 VDD.n6281 VDD.n5796 72.0905
R9073 VDD.n6152 VDD.n6105 72.0905
R9074 VDD.n6391 VDD.n5880 72.0905
R9075 VDD.n6391 VDD.n5881 72.0905
R9076 VDD.n6391 VDD.n5882 72.0905
R9077 VDD.n6391 VDD.n5883 72.0905
R9078 VDD.n6391 VDD.n5884 72.0905
R9079 VDD.n6391 VDD.n5885 72.0905
R9080 VDD.n6391 VDD.n5886 72.0905
R9081 VDD.n6391 VDD.n5887 72.0905
R9082 VDD.n6391 VDD.n5892 72.0905
R9083 VDD.n6391 VDD.n5893 72.0905
R9084 VDD.n6391 VDD.n5894 72.0905
R9085 VDD.n6391 VDD.n5895 72.0905
R9086 VDD.n6391 VDD.n5896 72.0905
R9087 VDD.n4942 VDD.n4941 72.0905
R9088 VDD.n5427 VDD.n4942 72.0905
R9089 VDD.n5298 VDD.n5251 72.0905
R9090 VDD.n5537 VDD.n5026 72.0905
R9091 VDD.n5537 VDD.n5027 72.0905
R9092 VDD.n5537 VDD.n5028 72.0905
R9093 VDD.n5537 VDD.n5029 72.0905
R9094 VDD.n5537 VDD.n5030 72.0905
R9095 VDD.n5537 VDD.n5031 72.0905
R9096 VDD.n5537 VDD.n5032 72.0905
R9097 VDD.n5537 VDD.n5033 72.0905
R9098 VDD.n5537 VDD.n5038 72.0905
R9099 VDD.n5537 VDD.n5039 72.0905
R9100 VDD.n5537 VDD.n5040 72.0905
R9101 VDD.n5537 VDD.n5041 72.0905
R9102 VDD.n5537 VDD.n5042 72.0905
R9103 VDD.n4156 VDD.n4155 72.0905
R9104 VDD.n4641 VDD.n4156 72.0905
R9105 VDD.n4512 VDD.n4465 72.0905
R9106 VDD.n4751 VDD.n4240 72.0905
R9107 VDD.n4751 VDD.n4241 72.0905
R9108 VDD.n4751 VDD.n4242 72.0905
R9109 VDD.n4751 VDD.n4243 72.0905
R9110 VDD.n4751 VDD.n4244 72.0905
R9111 VDD.n4751 VDD.n4245 72.0905
R9112 VDD.n4751 VDD.n4246 72.0905
R9113 VDD.n4751 VDD.n4247 72.0905
R9114 VDD.n4751 VDD.n4252 72.0905
R9115 VDD.n4751 VDD.n4253 72.0905
R9116 VDD.n4751 VDD.n4254 72.0905
R9117 VDD.n4751 VDD.n4255 72.0905
R9118 VDD.n4751 VDD.n4256 72.0905
R9119 VDD.n3302 VDD.n3301 72.0905
R9120 VDD.n3787 VDD.n3302 72.0905
R9121 VDD.n3658 VDD.n3611 72.0905
R9122 VDD.n3897 VDD.n3386 72.0905
R9123 VDD.n3897 VDD.n3387 72.0905
R9124 VDD.n3897 VDD.n3388 72.0905
R9125 VDD.n3897 VDD.n3389 72.0905
R9126 VDD.n3897 VDD.n3390 72.0905
R9127 VDD.n3897 VDD.n3391 72.0905
R9128 VDD.n3897 VDD.n3392 72.0905
R9129 VDD.n3897 VDD.n3393 72.0905
R9130 VDD.n3897 VDD.n3398 72.0905
R9131 VDD.n3897 VDD.n3399 72.0905
R9132 VDD.n3897 VDD.n3400 72.0905
R9133 VDD.n3897 VDD.n3401 72.0905
R9134 VDD.n3897 VDD.n3402 72.0905
R9135 VDD.n2516 VDD.n2515 72.0905
R9136 VDD.n3001 VDD.n2516 72.0905
R9137 VDD.n2872 VDD.n2825 72.0905
R9138 VDD.n3111 VDD.n2600 72.0905
R9139 VDD.n3111 VDD.n2601 72.0905
R9140 VDD.n3111 VDD.n2602 72.0905
R9141 VDD.n3111 VDD.n2603 72.0905
R9142 VDD.n3111 VDD.n2604 72.0905
R9143 VDD.n3111 VDD.n2605 72.0905
R9144 VDD.n3111 VDD.n2606 72.0905
R9145 VDD.n3111 VDD.n2607 72.0905
R9146 VDD.n3111 VDD.n2612 72.0905
R9147 VDD.n3111 VDD.n2613 72.0905
R9148 VDD.n3111 VDD.n2614 72.0905
R9149 VDD.n3111 VDD.n2615 72.0905
R9150 VDD.n3111 VDD.n2616 72.0905
R9151 VDD.n1661 VDD.n1660 72.0905
R9152 VDD.n2146 VDD.n1661 72.0905
R9153 VDD.n2017 VDD.n1970 72.0905
R9154 VDD.n2256 VDD.n1745 72.0905
R9155 VDD.n2256 VDD.n1746 72.0905
R9156 VDD.n2256 VDD.n1747 72.0905
R9157 VDD.n2256 VDD.n1748 72.0905
R9158 VDD.n2256 VDD.n1749 72.0905
R9159 VDD.n2256 VDD.n1750 72.0905
R9160 VDD.n2256 VDD.n1751 72.0905
R9161 VDD.n2256 VDD.n1752 72.0905
R9162 VDD.n2256 VDD.n1757 72.0905
R9163 VDD.n2256 VDD.n1758 72.0905
R9164 VDD.n2256 VDD.n1759 72.0905
R9165 VDD.n2256 VDD.n1760 72.0905
R9166 VDD.n2256 VDD.n1761 72.0905
R9167 VDD.n6380 VDD.n5905 71.1543
R9168 VDD.n5807 VDD.n5791 71.1543
R9169 VDD.n5526 VDD.n5051 71.1543
R9170 VDD.n4953 VDD.n4937 71.1543
R9171 VDD.n4740 VDD.n4265 71.1543
R9172 VDD.n4167 VDD.n4151 71.1543
R9173 VDD.n3886 VDD.n3411 71.1543
R9174 VDD.n3313 VDD.n3297 71.1543
R9175 VDD.n3100 VDD.n2625 71.1543
R9176 VDD.n2527 VDD.n2511 71.1543
R9177 VDD.n2245 VDD.n1770 71.1543
R9178 VDD.n1672 VDD.n1656 71.1543
R9179 VDD.n12474 VDD.n12473 70.7591
R9180 VDD.n6638 VDD.n6631 70.5361
R9181 VDD.n6640 VDD.n6639 70.5361
R9182 VDD.n6642 VDD.n6641 70.5361
R9183 VDD.n6645 VDD.n6629 70.5361
R9184 VDD.n6647 VDD.n6646 70.5361
R9185 VDD.n6649 VDD.n6648 70.5361
R9186 VDD.n6652 VDD.n6627 70.5361
R9187 VDD.n6654 VDD.n6653 70.5361
R9188 VDD.n6656 VDD.n6655 70.5361
R9189 VDD.n6659 VDD.n6625 70.5361
R9190 VDD.n6661 VDD.n6660 70.5361
R9191 VDD.n6697 VDD.n6662 70.5361
R9192 VDD.n6696 VDD.n6695 70.5361
R9193 VDD.n6694 VDD.n6693 70.5361
R9194 VDD.n6690 VDD.n6663 70.5361
R9195 VDD.n6689 VDD.n6688 70.5361
R9196 VDD.n6687 VDD.n6686 70.5361
R9197 VDD.n6683 VDD.n6665 70.5361
R9198 VDD.n6682 VDD.n6681 70.5361
R9199 VDD.n6680 VDD.n6679 70.5361
R9200 VDD.n6676 VDD.n6667 70.5361
R9201 VDD.n6675 VDD.n6674 70.5361
R9202 VDD.n6673 VDD.n6672 70.5361
R9203 VDD.n6670 VDD.n6669 70.5361
R9204 VDD.n12769 VDD.n6579 70.5361
R9205 VDD.n12768 VDD.n12767 70.5361
R9206 VDD.n12766 VDD.n12765 70.5361
R9207 VDD.n12762 VDD.n6581 70.5361
R9208 VDD.n12761 VDD.n12760 70.5361
R9209 VDD.n12759 VDD.n12758 70.5361
R9210 VDD.n12755 VDD.n6583 70.5361
R9211 VDD.n12754 VDD.n12753 70.5361
R9212 VDD.n12752 VDD.n12751 70.5361
R9213 VDD.n12748 VDD.n6585 70.5361
R9214 VDD.n12747 VDD.n12746 70.5361
R9215 VDD.n12745 VDD.n12744 70.5361
R9216 VDD.n12741 VDD.n6587 70.5361
R9217 VDD.n12740 VDD.n12739 70.5361
R9218 VDD.n12738 VDD.n12737 70.5361
R9219 VDD.n12734 VDD.n6589 70.5361
R9220 VDD.n12733 VDD.n12732 70.5361
R9221 VDD.n12731 VDD.n12730 70.5361
R9222 VDD.n12727 VDD.n6591 70.5361
R9223 VDD.n12726 VDD.n12725 70.5361
R9224 VDD.n12724 VDD.n12723 70.5361
R9225 VDD.n12720 VDD.n6593 70.5361
R9226 VDD.n12719 VDD.n12718 70.5361
R9227 VDD.n12717 VDD.n12716 70.5361
R9228 VDD.n8109 VDD.n8102 70.5361
R9229 VDD.n8183 VDD.n8101 70.5361
R9230 VDD.n8130 VDD.n8100 70.5361
R9231 VDD.n8132 VDD.n8099 70.5361
R9232 VDD.n8173 VDD.n8098 70.5361
R9233 VDD.n8139 VDD.n8097 70.5361
R9234 VDD.n8141 VDD.n8096 70.5361
R9235 VDD.n8162 VDD.n8095 70.5361
R9236 VDD.n8147 VDD.n8094 70.5361
R9237 VDD.n8162 VDD.n8094 70.5361
R9238 VDD.n8141 VDD.n8095 70.5361
R9239 VDD.n8139 VDD.n8096 70.5361
R9240 VDD.n8173 VDD.n8097 70.5361
R9241 VDD.n8132 VDD.n8098 70.5361
R9242 VDD.n8130 VDD.n8099 70.5361
R9243 VDD.n8183 VDD.n8100 70.5361
R9244 VDD.n8109 VDD.n8101 70.5361
R9245 VDD.n8103 VDD.n8102 70.5361
R9246 VDD.n12718 VDD.n12717 70.5361
R9247 VDD.n12720 VDD.n12719 70.5361
R9248 VDD.n12723 VDD.n6593 70.5361
R9249 VDD.n12725 VDD.n12724 70.5361
R9250 VDD.n12727 VDD.n12726 70.5361
R9251 VDD.n12730 VDD.n6591 70.5361
R9252 VDD.n12732 VDD.n12731 70.5361
R9253 VDD.n12734 VDD.n12733 70.5361
R9254 VDD.n12737 VDD.n6589 70.5361
R9255 VDD.n12739 VDD.n12738 70.5361
R9256 VDD.n12741 VDD.n12740 70.5361
R9257 VDD.n12744 VDD.n6587 70.5361
R9258 VDD.n12746 VDD.n12745 70.5361
R9259 VDD.n12748 VDD.n12747 70.5361
R9260 VDD.n12751 VDD.n6585 70.5361
R9261 VDD.n12753 VDD.n12752 70.5361
R9262 VDD.n12755 VDD.n12754 70.5361
R9263 VDD.n12758 VDD.n6583 70.5361
R9264 VDD.n12760 VDD.n12759 70.5361
R9265 VDD.n12762 VDD.n12761 70.5361
R9266 VDD.n12765 VDD.n6581 70.5361
R9267 VDD.n12767 VDD.n12766 70.5361
R9268 VDD.n12769 VDD.n12768 70.5361
R9269 VDD.n6669 VDD.n6579 70.5361
R9270 VDD.n6672 VDD.n6670 70.5361
R9271 VDD.n6674 VDD.n6673 70.5361
R9272 VDD.n6676 VDD.n6675 70.5361
R9273 VDD.n6679 VDD.n6667 70.5361
R9274 VDD.n6681 VDD.n6680 70.5361
R9275 VDD.n6683 VDD.n6682 70.5361
R9276 VDD.n6686 VDD.n6665 70.5361
R9277 VDD.n6688 VDD.n6687 70.5361
R9278 VDD.n6690 VDD.n6689 70.5361
R9279 VDD.n6693 VDD.n6663 70.5361
R9280 VDD.n6695 VDD.n6694 70.5361
R9281 VDD.n6697 VDD.n6696 70.5361
R9282 VDD.n6662 VDD.n6661 70.5361
R9283 VDD.n6660 VDD.n6659 70.5361
R9284 VDD.n6656 VDD.n6625 70.5361
R9285 VDD.n6655 VDD.n6654 70.5361
R9286 VDD.n6653 VDD.n6652 70.5361
R9287 VDD.n6649 VDD.n6627 70.5361
R9288 VDD.n6648 VDD.n6647 70.5361
R9289 VDD.n6646 VDD.n6645 70.5361
R9290 VDD.n6642 VDD.n6629 70.5361
R9291 VDD.n6641 VDD.n6640 70.5361
R9292 VDD.n6639 VDD.n6638 70.5361
R9293 VDD.n6635 VDD.n6631 70.5361
R9294 VDD.n10965 VDD.n10964 69.0092
R9295 VDD.n10993 VDD.n10992 69.0092
R9296 VDD.n6271 VDD.n5784 67.9542
R9297 VDD.n6051 VDD.n5784 67.9542
R9298 VDD.n6317 VDD.n6306 67.9542
R9299 VDD.n6317 VDD.n6307 67.9542
R9300 VDD.n6317 VDD.n6316 67.9542
R9301 VDD.n5998 VDD.n5931 67.9542
R9302 VDD.n5988 VDD.n5931 67.9542
R9303 VDD.n5993 VDD.n5931 67.9542
R9304 VDD.n5417 VDD.n4930 67.9542
R9305 VDD.n5197 VDD.n4930 67.9542
R9306 VDD.n5463 VDD.n5452 67.9542
R9307 VDD.n5463 VDD.n5453 67.9542
R9308 VDD.n5463 VDD.n5462 67.9542
R9309 VDD.n5144 VDD.n5077 67.9542
R9310 VDD.n5134 VDD.n5077 67.9542
R9311 VDD.n5139 VDD.n5077 67.9542
R9312 VDD.n4631 VDD.n4144 67.9542
R9313 VDD.n4411 VDD.n4144 67.9542
R9314 VDD.n4677 VDD.n4666 67.9542
R9315 VDD.n4677 VDD.n4667 67.9542
R9316 VDD.n4677 VDD.n4676 67.9542
R9317 VDD.n4358 VDD.n4291 67.9542
R9318 VDD.n4348 VDD.n4291 67.9542
R9319 VDD.n4353 VDD.n4291 67.9542
R9320 VDD.n3777 VDD.n3290 67.9542
R9321 VDD.n3557 VDD.n3290 67.9542
R9322 VDD.n3823 VDD.n3812 67.9542
R9323 VDD.n3823 VDD.n3813 67.9542
R9324 VDD.n3823 VDD.n3822 67.9542
R9325 VDD.n3504 VDD.n3437 67.9542
R9326 VDD.n3494 VDD.n3437 67.9542
R9327 VDD.n3499 VDD.n3437 67.9542
R9328 VDD.n2991 VDD.n2504 67.9542
R9329 VDD.n2771 VDD.n2504 67.9542
R9330 VDD.n3037 VDD.n3026 67.9542
R9331 VDD.n3037 VDD.n3027 67.9542
R9332 VDD.n3037 VDD.n3036 67.9542
R9333 VDD.n2718 VDD.n2651 67.9542
R9334 VDD.n2708 VDD.n2651 67.9542
R9335 VDD.n2713 VDD.n2651 67.9542
R9336 VDD.n2136 VDD.n1649 67.9542
R9337 VDD.n1916 VDD.n1649 67.9542
R9338 VDD.n2182 VDD.n2171 67.9542
R9339 VDD.n2182 VDD.n2172 67.9542
R9340 VDD.n2182 VDD.n2181 67.9542
R9341 VDD.n1863 VDD.n1796 67.9542
R9342 VDD.n1853 VDD.n1796 67.9542
R9343 VDD.n1858 VDD.n1796 67.9542
R9344 VDD.n6619 VDD.n6618 66.8858
R9345 VDD.n6617 VDD.n6616 66.8858
R9346 VDD.n6615 VDD.n6613 66.8858
R9347 VDD.n8124 VDD.n8123 66.8856
R9348 VDD.n6618 VDD.n6617 66.8854
R9349 VDD.n6616 VDD.n6615 66.8854
R9350 VDD.n12480 VDD.n12479 64.5694
R9351 VDD.n12463 VDD.n12462 64.5694
R9352 VDD.n9209 VDD.n9207 64.4031
R9353 VDD.n12497 VDD.n12496 60.3019
R9354 VDD.n12450 VDD.n6901 60.3019
R9355 VDD.n9651 VDD.t33 60.2505
R9356 VDD.n9663 VDD.t54 60.2505
R9357 VDD.n10794 VDD.t51 60.2505
R9358 VDD.n10806 VDD.t36 60.2505
R9359 VDD.n8963 VDD.t59 60.2505
R9360 VDD.n8870 VDD.t40 60.2505
R9361 VDD.n9002 VDD.t48 60.2505
R9362 VDD.n8989 VDD.t42 60.2505
R9363 VDD.n9277 VDD.t57 60.2505
R9364 VDD.n9407 VDD.t45 60.2505
R9365 VDD.n6260 VDD.n6259 60.14
R9366 VDD.n6318 VDD.n6303 60.14
R9367 VDD.n5992 VDD.n5991 60.14
R9368 VDD.n5406 VDD.n5405 60.14
R9369 VDD.n5464 VDD.n5449 60.14
R9370 VDD.n5138 VDD.n5137 60.14
R9371 VDD.n4620 VDD.n4619 60.14
R9372 VDD.n4678 VDD.n4663 60.14
R9373 VDD.n4352 VDD.n4351 60.14
R9374 VDD.n3766 VDD.n3765 60.14
R9375 VDD.n3824 VDD.n3809 60.14
R9376 VDD.n3498 VDD.n3497 60.14
R9377 VDD.n2980 VDD.n2979 60.14
R9378 VDD.n3038 VDD.n3023 60.14
R9379 VDD.n2712 VDD.n2711 60.14
R9380 VDD.n2125 VDD.n2124 60.14
R9381 VDD.n2183 VDD.n2168 60.14
R9382 VDD.n1857 VDD.n1856 60.14
R9383 VDD.n6273 VDD.n6272 60.1394
R9384 VDD.n6310 VDD.n6305 60.1394
R9385 VDD.n6000 VDD.n5999 60.1394
R9386 VDD.n5419 VDD.n5418 60.1394
R9387 VDD.n5456 VDD.n5451 60.1394
R9388 VDD.n5146 VDD.n5145 60.1394
R9389 VDD.n4633 VDD.n4632 60.1394
R9390 VDD.n4670 VDD.n4665 60.1394
R9391 VDD.n4360 VDD.n4359 60.1394
R9392 VDD.n3779 VDD.n3778 60.1394
R9393 VDD.n3816 VDD.n3811 60.1394
R9394 VDD.n3506 VDD.n3505 60.1394
R9395 VDD.n2993 VDD.n2992 60.1394
R9396 VDD.n3030 VDD.n3025 60.1394
R9397 VDD.n2720 VDD.n2719 60.1394
R9398 VDD.n2138 VDD.n2137 60.1394
R9399 VDD.n2175 VDD.n2170 60.1394
R9400 VDD.n1865 VDD.n1864 60.1394
R9401 VDD.n9196 VDD.n9195 60.1048
R9402 VDD.n10983 VDD.n9196 60.1048
R9403 VDD.n10044 VDD.t149 59.2764
R9404 VDD.n10603 VDD.t151 59.2764
R9405 VDD.n10542 VDD.t29 59.2764
R9406 VDD.t35 VDD.n9561 59.2764
R9407 VDD.t39 VDD.n10732 59.2764
R9408 VDD.t41 VDD.n8915 59.2764
R9409 VDD.t47 VDD.n9368 59.2764
R9410 VDD.n8197 VDD.n8094 57.2334
R9411 VDD.n8197 VDD.n8095 57.2334
R9412 VDD.n8197 VDD.n8096 57.2334
R9413 VDD.n8197 VDD.n8097 57.2334
R9414 VDD.n8197 VDD.n8098 57.2334
R9415 VDD.n8197 VDD.n8099 57.2334
R9416 VDD.n8197 VDD.n8100 57.2334
R9417 VDD.n8197 VDD.n8101 57.2334
R9418 VDD.n8197 VDD.n8102 57.2334
R9419 VDD.n12717 VDD.n6580 57.2334
R9420 VDD.n12719 VDD.n6580 57.2334
R9421 VDD.n6593 VDD.n6580 57.2334
R9422 VDD.n12724 VDD.n6580 57.2334
R9423 VDD.n12726 VDD.n6580 57.2334
R9424 VDD.n6591 VDD.n6580 57.2334
R9425 VDD.n12731 VDD.n6580 57.2334
R9426 VDD.n12733 VDD.n6580 57.2334
R9427 VDD.n6589 VDD.n6580 57.2334
R9428 VDD.n12738 VDD.n6580 57.2334
R9429 VDD.n12740 VDD.n6580 57.2334
R9430 VDD.n6587 VDD.n6580 57.2334
R9431 VDD.n12745 VDD.n6580 57.2334
R9432 VDD.n12747 VDD.n6580 57.2334
R9433 VDD.n6585 VDD.n6580 57.2334
R9434 VDD.n12752 VDD.n6580 57.2334
R9435 VDD.n12754 VDD.n6580 57.2334
R9436 VDD.n6583 VDD.n6580 57.2334
R9437 VDD.n12759 VDD.n6580 57.2334
R9438 VDD.n12761 VDD.n6580 57.2334
R9439 VDD.n6581 VDD.n6580 57.2334
R9440 VDD.n12766 VDD.n6580 57.2334
R9441 VDD.n12768 VDD.n6580 57.2334
R9442 VDD.n6580 VDD.n6579 57.2334
R9443 VDD.n6670 VDD.n6580 57.2334
R9444 VDD.n6673 VDD.n6580 57.2334
R9445 VDD.n6675 VDD.n6580 57.2334
R9446 VDD.n6667 VDD.n6580 57.2334
R9447 VDD.n6680 VDD.n6580 57.2334
R9448 VDD.n6682 VDD.n6580 57.2334
R9449 VDD.n6665 VDD.n6580 57.2334
R9450 VDD.n6687 VDD.n6580 57.2334
R9451 VDD.n6689 VDD.n6580 57.2334
R9452 VDD.n6663 VDD.n6580 57.2334
R9453 VDD.n6694 VDD.n6580 57.2334
R9454 VDD.n6696 VDD.n6580 57.2334
R9455 VDD.n6662 VDD.n6580 57.2334
R9456 VDD.n6660 VDD.n6580 57.2334
R9457 VDD.n6625 VDD.n6580 57.2334
R9458 VDD.n6655 VDD.n6580 57.2334
R9459 VDD.n6653 VDD.n6580 57.2334
R9460 VDD.n6627 VDD.n6580 57.2334
R9461 VDD.n6648 VDD.n6580 57.2334
R9462 VDD.n6646 VDD.n6580 57.2334
R9463 VDD.n6629 VDD.n6580 57.2334
R9464 VDD.n6641 VDD.n6580 57.2334
R9465 VDD.n6639 VDD.n6580 57.2334
R9466 VDD.n6631 VDD.n6580 57.2334
R9467 VDD.n10962 VDD.n9219 57.2295
R9468 VDD.n10990 VDD.n10987 57.2295
R9469 VDD.n6343 VDD.n5939 55.1287
R9470 VDD.n5489 VDD.n5085 55.1287
R9471 VDD.n4703 VDD.n4299 55.1287
R9472 VDD.n3849 VDD.n3445 55.1287
R9473 VDD.n3063 VDD.n2659 55.1287
R9474 VDD.n2208 VDD.n1804 55.1287
R9475 VDD.n8125 VDD.n8114 54.6255
R9476 VDD.n9976 VDD.n9973 54.3813
R9477 VDD.n11641 VDD.n7611 54.2862
R9478 VDD.n8114 VDD.n8092 53.8338
R9479 VDD.n8567 VDD.n7754 53.8338
R9480 VDD.n8557 VDD.n7755 53.8338
R9481 VDD.n8557 VDD.n8556 53.8338
R9482 VDD.n8556 VDD.n8555 53.8338
R9483 VDD.n8555 VDD.n7773 53.8338
R9484 VDD.n8546 VDD.n7773 53.8338
R9485 VDD.n8546 VDD.n8545 53.8338
R9486 VDD.n8545 VDD.n8544 53.8338
R9487 VDD.n8544 VDD.n7782 53.8338
R9488 VDD.n10045 VDD.n10044 52.6902
R9489 VDD.n10604 VDD.n10603 52.6902
R9490 VDD.n10543 VDD.n10542 52.6902
R9491 VDD.n9632 VDD.n9561 52.6902
R9492 VDD.n10732 VDD.n10726 52.6902
R9493 VDD.n8915 VDD.n8888 52.6902
R9494 VDD.n9368 VDD.n9364 52.6902
R9495 VDD.n8570 VDD.n7756 51.067
R9496 VDD.n8574 VDD.n7757 51.067
R9497 VDD.n8578 VDD.n7758 51.067
R9498 VDD.n8582 VDD.n7759 51.067
R9499 VDD.n8589 VDD.n7760 51.067
R9500 VDD.n8591 VDD.n7753 51.067
R9501 VDD.n8573 VDD.n7756 51.0665
R9502 VDD.n8577 VDD.n7757 51.0665
R9503 VDD.n8581 VDD.n7758 51.0665
R9504 VDD.n8584 VDD.n7759 51.0665
R9505 VDD.n8589 VDD.n8588 51.0665
R9506 VDD.n8592 VDD.n8591 51.0665
R9507 VDD.n7928 VDD.n7848 50.7006
R9508 VDD.n7816 VDD.n7815 50.7006
R9509 VDD.n6283 VDD.n6282 50.7006
R9510 VDD.n6390 VDD.n5897 50.7006
R9511 VDD.n5955 VDD.n5888 50.7006
R9512 VDD.n5429 VDD.n5428 50.7006
R9513 VDD.n5536 VDD.n5043 50.7006
R9514 VDD.n5101 VDD.n5034 50.7006
R9515 VDD.n4643 VDD.n4642 50.7006
R9516 VDD.n4750 VDD.n4257 50.7006
R9517 VDD.n4315 VDD.n4248 50.7006
R9518 VDD.n3789 VDD.n3788 50.7006
R9519 VDD.n3896 VDD.n3403 50.7006
R9520 VDD.n3461 VDD.n3394 50.7006
R9521 VDD.n3003 VDD.n3002 50.7006
R9522 VDD.n3110 VDD.n2617 50.7006
R9523 VDD.n2675 VDD.n2608 50.7006
R9524 VDD.n2148 VDD.n2147 50.7006
R9525 VDD.n2255 VDD.n1762 50.7006
R9526 VDD.n1820 VDD.n1753 50.7006
R9527 VDD.n7954 VDD.n7830 50.6999
R9528 VDD.n7865 VDD.n7864 50.6999
R9529 VDD.n6542 VDD.n6541 50.6999
R9530 VDD.n6254 VDD.n6056 50.6999
R9531 VDD.n6254 VDD.n6253 50.6999
R9532 VDD.n6153 VDD.n6104 50.6999
R9533 VDD.n6151 VDD.n6107 50.6999
R9534 VDD.n6392 VDD.n5878 50.6999
R9535 VDD.n6372 VDD.n5891 50.6999
R9536 VDD.n5688 VDD.n5687 50.6999
R9537 VDD.n5400 VDD.n5202 50.6999
R9538 VDD.n5400 VDD.n5399 50.6999
R9539 VDD.n5299 VDD.n5250 50.6999
R9540 VDD.n5297 VDD.n5253 50.6999
R9541 VDD.n5538 VDD.n5024 50.6999
R9542 VDD.n5518 VDD.n5037 50.6999
R9543 VDD.n4902 VDD.n4901 50.6999
R9544 VDD.n4614 VDD.n4416 50.6999
R9545 VDD.n4614 VDD.n4613 50.6999
R9546 VDD.n4513 VDD.n4464 50.6999
R9547 VDD.n4511 VDD.n4467 50.6999
R9548 VDD.n4752 VDD.n4238 50.6999
R9549 VDD.n4732 VDD.n4251 50.6999
R9550 VDD.n4048 VDD.n4047 50.6999
R9551 VDD.n3760 VDD.n3562 50.6999
R9552 VDD.n3760 VDD.n3759 50.6999
R9553 VDD.n3659 VDD.n3610 50.6999
R9554 VDD.n3657 VDD.n3613 50.6999
R9555 VDD.n3898 VDD.n3384 50.6999
R9556 VDD.n3878 VDD.n3397 50.6999
R9557 VDD.n3262 VDD.n3261 50.6999
R9558 VDD.n2974 VDD.n2776 50.6999
R9559 VDD.n2974 VDD.n2973 50.6999
R9560 VDD.n2873 VDD.n2824 50.6999
R9561 VDD.n2871 VDD.n2827 50.6999
R9562 VDD.n3112 VDD.n2598 50.6999
R9563 VDD.n3092 VDD.n2611 50.6999
R9564 VDD.n2407 VDD.n2406 50.6999
R9565 VDD.n2119 VDD.n1921 50.6999
R9566 VDD.n2119 VDD.n2118 50.6999
R9567 VDD.n2018 VDD.n1969 50.6999
R9568 VDD.n2016 VDD.n1972 50.6999
R9569 VDD.n2257 VDD.n1743 50.6999
R9570 VDD.n2237 VDD.n1756 50.6999
R9571 VDD.n7785 VDD.n7782 50.6672
R9572 VDD.n5994 VDD.n5993 49.0945
R9573 VDD.n5997 VDD.n5988 49.0945
R9574 VDD.n5999 VDD.n5998 49.0945
R9575 VDD.n6270 VDD.n6051 49.0945
R9576 VDD.n6273 VDD.n6271 49.0945
R9577 VDD.n6271 VDD.n6270 49.0945
R9578 VDD.n6259 VDD.n6051 49.0945
R9579 VDD.n6316 VDD.n6315 49.0945
R9580 VDD.n6312 VDD.n6307 49.0945
R9581 VDD.n6310 VDD.n6306 49.0945
R9582 VDD.n6312 VDD.n6306 49.0945
R9583 VDD.n6315 VDD.n6307 49.0945
R9584 VDD.n6316 VDD.n6303 49.0945
R9585 VDD.n5998 VDD.n5997 49.0945
R9586 VDD.n5994 VDD.n5988 49.0945
R9587 VDD.n5993 VDD.n5992 49.0945
R9588 VDD.n5140 VDD.n5139 49.0945
R9589 VDD.n5143 VDD.n5134 49.0945
R9590 VDD.n5145 VDD.n5144 49.0945
R9591 VDD.n5416 VDD.n5197 49.0945
R9592 VDD.n5419 VDD.n5417 49.0945
R9593 VDD.n5417 VDD.n5416 49.0945
R9594 VDD.n5405 VDD.n5197 49.0945
R9595 VDD.n5462 VDD.n5461 49.0945
R9596 VDD.n5458 VDD.n5453 49.0945
R9597 VDD.n5456 VDD.n5452 49.0945
R9598 VDD.n5458 VDD.n5452 49.0945
R9599 VDD.n5461 VDD.n5453 49.0945
R9600 VDD.n5462 VDD.n5449 49.0945
R9601 VDD.n5144 VDD.n5143 49.0945
R9602 VDD.n5140 VDD.n5134 49.0945
R9603 VDD.n5139 VDD.n5138 49.0945
R9604 VDD.n4354 VDD.n4353 49.0945
R9605 VDD.n4357 VDD.n4348 49.0945
R9606 VDD.n4359 VDD.n4358 49.0945
R9607 VDD.n4630 VDD.n4411 49.0945
R9608 VDD.n4633 VDD.n4631 49.0945
R9609 VDD.n4631 VDD.n4630 49.0945
R9610 VDD.n4619 VDD.n4411 49.0945
R9611 VDD.n4676 VDD.n4675 49.0945
R9612 VDD.n4672 VDD.n4667 49.0945
R9613 VDD.n4670 VDD.n4666 49.0945
R9614 VDD.n4672 VDD.n4666 49.0945
R9615 VDD.n4675 VDD.n4667 49.0945
R9616 VDD.n4676 VDD.n4663 49.0945
R9617 VDD.n4358 VDD.n4357 49.0945
R9618 VDD.n4354 VDD.n4348 49.0945
R9619 VDD.n4353 VDD.n4352 49.0945
R9620 VDD.n3500 VDD.n3499 49.0945
R9621 VDD.n3503 VDD.n3494 49.0945
R9622 VDD.n3505 VDD.n3504 49.0945
R9623 VDD.n3776 VDD.n3557 49.0945
R9624 VDD.n3779 VDD.n3777 49.0945
R9625 VDD.n3777 VDD.n3776 49.0945
R9626 VDD.n3765 VDD.n3557 49.0945
R9627 VDD.n3822 VDD.n3821 49.0945
R9628 VDD.n3818 VDD.n3813 49.0945
R9629 VDD.n3816 VDD.n3812 49.0945
R9630 VDD.n3818 VDD.n3812 49.0945
R9631 VDD.n3821 VDD.n3813 49.0945
R9632 VDD.n3822 VDD.n3809 49.0945
R9633 VDD.n3504 VDD.n3503 49.0945
R9634 VDD.n3500 VDD.n3494 49.0945
R9635 VDD.n3499 VDD.n3498 49.0945
R9636 VDD.n2714 VDD.n2713 49.0945
R9637 VDD.n2717 VDD.n2708 49.0945
R9638 VDD.n2719 VDD.n2718 49.0945
R9639 VDD.n2990 VDD.n2771 49.0945
R9640 VDD.n2993 VDD.n2991 49.0945
R9641 VDD.n2991 VDD.n2990 49.0945
R9642 VDD.n2979 VDD.n2771 49.0945
R9643 VDD.n3036 VDD.n3035 49.0945
R9644 VDD.n3032 VDD.n3027 49.0945
R9645 VDD.n3030 VDD.n3026 49.0945
R9646 VDD.n3032 VDD.n3026 49.0945
R9647 VDD.n3035 VDD.n3027 49.0945
R9648 VDD.n3036 VDD.n3023 49.0945
R9649 VDD.n2718 VDD.n2717 49.0945
R9650 VDD.n2714 VDD.n2708 49.0945
R9651 VDD.n2713 VDD.n2712 49.0945
R9652 VDD.n1859 VDD.n1858 49.0945
R9653 VDD.n1862 VDD.n1853 49.0945
R9654 VDD.n1864 VDD.n1863 49.0945
R9655 VDD.n2135 VDD.n1916 49.0945
R9656 VDD.n2138 VDD.n2136 49.0945
R9657 VDD.n2136 VDD.n2135 49.0945
R9658 VDD.n2124 VDD.n1916 49.0945
R9659 VDD.n2181 VDD.n2180 49.0945
R9660 VDD.n2177 VDD.n2172 49.0945
R9661 VDD.n2175 VDD.n2171 49.0945
R9662 VDD.n2177 VDD.n2171 49.0945
R9663 VDD.n2180 VDD.n2172 49.0945
R9664 VDD.n2181 VDD.n2168 49.0945
R9665 VDD.n1863 VDD.n1862 49.0945
R9666 VDD.n1859 VDD.n1853 49.0945
R9667 VDD.n1858 VDD.n1857 49.0945
R9668 VDD.n998 VDD.n997 49.0945
R9669 VDD.n1003 VDD.n1002 49.0945
R9670 VDD.n1202 VDD.n1201 49.0945
R9671 VDD.n1205 VDD.n1204 49.0945
R9672 VDD.n1208 VDD.n1207 49.0945
R9673 VDD.n1247 VDD.n1246 49.0945
R9674 VDD.n1250 VDD.n1249 49.0945
R9675 VDD.n1253 VDD.n1252 49.0945
R9676 VDD.n552 VDD.n551 49.0945
R9677 VDD.n557 VDD.n556 49.0945
R9678 VDD.n756 VDD.n755 49.0945
R9679 VDD.n759 VDD.n758 49.0945
R9680 VDD.n762 VDD.n761 49.0945
R9681 VDD.n19 VDD.n18 49.0945
R9682 VDD.n22 VDD.n21 49.0945
R9683 VDD.n25 VDD.n24 49.0945
R9684 VDD.n8198 VDD.n8087 49.0838
R9685 VDD.n8203 VDD.n8201 49.0838
R9686 VDD.n8202 VDD.n8081 49.0838
R9687 VDD.n8214 VDD.n8213 49.0838
R9688 VDD.n8217 VDD.n8076 49.0838
R9689 VDD.n8219 VDD.n8218 49.0838
R9690 VDD.n8229 VDD.n8070 49.0838
R9691 VDD.n8230 VDD.n8065 49.0838
R9692 VDD.n8235 VDD.n8233 49.0838
R9693 VDD.n8234 VDD.n8059 49.0838
R9694 VDD.n8247 VDD.n8245 49.0838
R9695 VDD.n8246 VDD.n8053 49.0838
R9696 VDD.n8258 VDD.n8257 49.0838
R9697 VDD.n8261 VDD.n8048 49.0838
R9698 VDD.n8263 VDD.n8262 49.0838
R9699 VDD.n8273 VDD.n8042 49.0838
R9700 VDD.n8274 VDD.n8037 49.0838
R9701 VDD.n8279 VDD.n8277 49.0838
R9702 VDD.n8278 VDD.n8030 49.0838
R9703 VDD.n8289 VDD.n8288 49.0838
R9704 VDD.n8292 VDD.n8025 49.0838
R9705 VDD.n8294 VDD.n8293 49.0838
R9706 VDD.n8304 VDD.n8019 49.0838
R9707 VDD.n8305 VDD.n8014 49.0838
R9708 VDD.n8310 VDD.n8308 49.0838
R9709 VDD.n8309 VDD.n8008 49.0838
R9710 VDD.n8322 VDD.n8320 49.0838
R9711 VDD.n8321 VDD.n8002 49.0838
R9712 VDD.n8334 VDD.n8332 49.0838
R9713 VDD.n8333 VDD.n7988 49.0838
R9714 VDD.n8497 VDD.n7989 49.0838
R9715 VDD.n8488 VDD.n8339 49.0838
R9716 VDD.n8487 VDD.n8340 49.0838
R9717 VDD.n8484 VDD.n8483 49.0838
R9718 VDD.n8354 VDD.n8345 49.0838
R9719 VDD.n8473 VDD.n8355 49.0838
R9720 VDD.n8472 VDD.n8356 49.0838
R9721 VDD.n8469 VDD.n8468 49.0838
R9722 VDD.n8370 VDD.n8362 49.0838
R9723 VDD.n8459 VDD.n8371 49.0838
R9724 VDD.n8458 VDD.n8372 49.0838
R9725 VDD.n8455 VDD.n8454 49.0838
R9726 VDD.n8387 VDD.n8378 49.0838
R9727 VDD.n8444 VDD.n8388 49.0838
R9728 VDD.n8443 VDD.n8389 49.0838
R9729 VDD.n8440 VDD.n8439 49.0838
R9730 VDD.n8404 VDD.n8395 49.0838
R9731 VDD.n8429 VDD.n8405 49.0838
R9732 VDD.n8428 VDD.n8406 49.0838
R9733 VDD.n8425 VDD.n8424 49.0838
R9734 VDD.n8413 VDD.n8412 49.0838
R9735 VDD.n8568 VDD.n7764 49.0838
R9736 VDD.n9980 VDD.n9973 48.3613
R9737 VDD.n6553 VDD.n5783 48.0774
R9738 VDD.n5699 VDD.n4929 48.0774
R9739 VDD.n4913 VDD.n4143 48.0774
R9740 VDD.n4059 VDD.n3289 48.0774
R9741 VDD.n3273 VDD.n2503 48.0774
R9742 VDD.n2418 VDD.n1648 48.0774
R9743 VDD.n6598 VDD.n6596 46.4193
R9744 VDD.n10041 VDD.n10032 46.104
R9745 VDD.n10600 VDD.n10591 46.104
R9746 VDD.n10552 VDD.n10551 46.104
R9747 VDD.n9630 VDD.n9564 46.104
R9748 VDD.n10738 VDD.n10737 46.104
R9749 VDD.n8910 VDD.n8891 46.104
R9750 VDD.n9375 VDD.n9362 46.104
R9751 VDD.n9593 VDD.n9589 44.9671
R9752 VDD.n10764 VDD.n10699 44.9671
R9753 VDD.n7848 VDD.n7749 44.7682
R9754 VDD.n7815 VDD.n7749 44.7682
R9755 VDD.n6283 VDD.n5796 44.7682
R9756 VDD.n6391 VDD.n5888 44.7682
R9757 VDD.n6391 VDD.n6390 44.7682
R9758 VDD.n5429 VDD.n4942 44.7682
R9759 VDD.n5537 VDD.n5034 44.7682
R9760 VDD.n5537 VDD.n5536 44.7682
R9761 VDD.n4643 VDD.n4156 44.7682
R9762 VDD.n4751 VDD.n4248 44.7682
R9763 VDD.n4751 VDD.n4750 44.7682
R9764 VDD.n3789 VDD.n3302 44.7682
R9765 VDD.n3897 VDD.n3394 44.7682
R9766 VDD.n3897 VDD.n3896 44.7682
R9767 VDD.n3003 VDD.n2516 44.7682
R9768 VDD.n3111 VDD.n2608 44.7682
R9769 VDD.n3111 VDD.n3110 44.7682
R9770 VDD.n2148 VDD.n1661 44.7682
R9771 VDD.n2256 VDD.n1753 44.7682
R9772 VDD.n2256 VDD.n2255 44.7682
R9773 VDD.n7865 VDD.n7749 44.768
R9774 VDD.n7830 VDD.n7749 44.768
R9775 VDD.n6541 VDD.n5796 44.768
R9776 VDD.n6056 VDD.n5796 44.768
R9777 VDD.n6253 VDD.n5796 44.768
R9778 VDD.n6153 VDD.n6152 44.768
R9779 VDD.n6152 VDD.n6151 44.768
R9780 VDD.n6392 VDD.n6391 44.768
R9781 VDD.n6391 VDD.n5891 44.768
R9782 VDD.n5687 VDD.n4942 44.768
R9783 VDD.n5202 VDD.n4942 44.768
R9784 VDD.n5399 VDD.n4942 44.768
R9785 VDD.n5299 VDD.n5298 44.768
R9786 VDD.n5298 VDD.n5297 44.768
R9787 VDD.n5538 VDD.n5537 44.768
R9788 VDD.n5537 VDD.n5037 44.768
R9789 VDD.n4901 VDD.n4156 44.768
R9790 VDD.n4416 VDD.n4156 44.768
R9791 VDD.n4613 VDD.n4156 44.768
R9792 VDD.n4513 VDD.n4512 44.768
R9793 VDD.n4512 VDD.n4511 44.768
R9794 VDD.n4752 VDD.n4751 44.768
R9795 VDD.n4751 VDD.n4251 44.768
R9796 VDD.n4047 VDD.n3302 44.768
R9797 VDD.n3562 VDD.n3302 44.768
R9798 VDD.n3759 VDD.n3302 44.768
R9799 VDD.n3659 VDD.n3658 44.768
R9800 VDD.n3658 VDD.n3657 44.768
R9801 VDD.n3898 VDD.n3897 44.768
R9802 VDD.n3897 VDD.n3397 44.768
R9803 VDD.n3261 VDD.n2516 44.768
R9804 VDD.n2776 VDD.n2516 44.768
R9805 VDD.n2973 VDD.n2516 44.768
R9806 VDD.n2873 VDD.n2872 44.768
R9807 VDD.n2872 VDD.n2871 44.768
R9808 VDD.n3112 VDD.n3111 44.768
R9809 VDD.n3111 VDD.n2611 44.768
R9810 VDD.n2406 VDD.n1661 44.768
R9811 VDD.n1921 VDD.n1661 44.768
R9812 VDD.n2118 VDD.n1661 44.768
R9813 VDD.n2018 VDD.n2017 44.768
R9814 VDD.n2017 VDD.n2016 44.768
R9815 VDD.n2257 VDD.n2256 44.768
R9816 VDD.n2256 VDD.n1756 44.768
R9817 VDD.n1321 VDD.n1320 44.768
R9818 VDD.n93 VDD.n92 44.768
R9819 VDD.n11025 VDD.n8732 44.4161
R9820 VDD.n9182 VDD.n9173 44.4161
R9821 VDD.n6547 VDD.n5791 43.5902
R9822 VDD.n5693 VDD.n4937 43.5902
R9823 VDD.n4907 VDD.n4151 43.5902
R9824 VDD.n4053 VDD.n3297 43.5902
R9825 VDD.n3267 VDD.n2511 43.5902
R9826 VDD.n2412 VDD.n1656 43.5902
R9827 VDD.n6485 VDD.n6484 41.7887
R9828 VDD.n6428 VDD.n6427 41.7887
R9829 VDD.n5631 VDD.n5630 41.7887
R9830 VDD.n5574 VDD.n5573 41.7887
R9831 VDD.n4845 VDD.n4844 41.7887
R9832 VDD.n4788 VDD.n4787 41.7887
R9833 VDD.n3991 VDD.n3990 41.7887
R9834 VDD.n3934 VDD.n3933 41.7887
R9835 VDD.n3205 VDD.n3204 41.7887
R9836 VDD.n3148 VDD.n3147 41.7887
R9837 VDD.n2350 VDD.n2349 41.7887
R9838 VDD.n2293 VDD.n2292 41.7887
R9839 VDD.n1074 VDD.n1072 41.7887
R9840 VDD.n1459 VDD.n1457 41.7887
R9841 VDD.n628 VDD.n626 41.7887
R9842 VDD.n231 VDD.n229 41.7887
R9843 VDD.n8196 VDD.n8195 41.7222
R9844 VDD.n6634 VDD.n6602 41.7222
R9845 VDD.n12713 VDD.n6595 41.7221
R9846 VDD.n8150 VDD.n8093 41.7221
R9847 VDD.n6260 VDD.n5784 41.6217
R9848 VDD.n6318 VDD.n6317 41.6217
R9849 VDD.n5991 VDD.n5931 41.6217
R9850 VDD.n5406 VDD.n4930 41.6217
R9851 VDD.n5464 VDD.n5463 41.6217
R9852 VDD.n5137 VDD.n5077 41.6217
R9853 VDD.n4620 VDD.n4144 41.6217
R9854 VDD.n4678 VDD.n4677 41.6217
R9855 VDD.n4351 VDD.n4291 41.6217
R9856 VDD.n3766 VDD.n3290 41.6217
R9857 VDD.n3824 VDD.n3823 41.6217
R9858 VDD.n3497 VDD.n3437 41.6217
R9859 VDD.n2980 VDD.n2504 41.6217
R9860 VDD.n3038 VDD.n3037 41.6217
R9861 VDD.n2711 VDD.n2651 41.6217
R9862 VDD.n2125 VDD.n1649 41.6217
R9863 VDD.n2183 VDD.n2182 41.6217
R9864 VDD.n1856 VDD.n1796 41.6217
R9865 VDD.n1212 VDD.n1211 41.6217
R9866 VDD.n1258 VDD.n1257 41.6217
R9867 VDD.n766 VDD.n765 41.6217
R9868 VDD.n30 VDD.n29 41.6217
R9869 VDD.n6272 VDD.n5784 41.6215
R9870 VDD.n6317 VDD.n6305 41.6215
R9871 VDD.n6000 VDD.n5931 41.6215
R9872 VDD.n5418 VDD.n4930 41.6215
R9873 VDD.n5463 VDD.n5451 41.6215
R9874 VDD.n5146 VDD.n5077 41.6215
R9875 VDD.n4632 VDD.n4144 41.6215
R9876 VDD.n4677 VDD.n4665 41.6215
R9877 VDD.n4360 VDD.n4291 41.6215
R9878 VDD.n3778 VDD.n3290 41.6215
R9879 VDD.n3823 VDD.n3811 41.6215
R9880 VDD.n3506 VDD.n3437 41.6215
R9881 VDD.n2992 VDD.n2504 41.6215
R9882 VDD.n3037 VDD.n3025 41.6215
R9883 VDD.n2720 VDD.n2651 41.6215
R9884 VDD.n2137 VDD.n1649 41.6215
R9885 VDD.n2182 VDD.n2170 41.6215
R9886 VDD.n1865 VDD.n1796 41.6215
R9887 VDD.n1009 VDD.n1008 41.6215
R9888 VDD.n1257 VDD.n1256 41.6215
R9889 VDD.n563 VDD.n562 41.6215
R9890 VDD.n29 VDD.n28 41.6215
R9891 VDD.n8590 VDD.n7754 41.1672
R9892 VDD.n9657 VDD.n9645 40.9783
R9893 VDD.n9668 VDD.n9659 40.9783
R9894 VDD.n10800 VDD.n10788 40.9783
R9895 VDD.n10811 VDD.n10802 40.9783
R9896 VDD.n8876 VDD.n8864 40.9783
R9897 VDD.n8954 VDD.n8861 40.9783
R9898 VDD.n8974 VDD.n8857 40.9783
R9899 VDD.n9007 VDD.n8998 40.9783
R9900 VDD.n8977 VDD.n8834 40.9783
R9901 VDD.n8996 VDD.n8829 40.9783
R9902 VDD.n9287 VDD.n9275 40.9783
R9903 VDD.n9417 VDD.n9405 40.9783
R9904 VDD.n7974 VDD.n7817 40.8219
R9905 VDD.n7973 VDD.n7972 40.8219
R9906 VDD.n7822 VDD.n7818 40.8219
R9907 VDD.n7965 VDD.n7823 40.8219
R9908 VDD.n7964 VDD.n7963 40.8219
R9909 VDD.n7828 VDD.n7824 40.8219
R9910 VDD.n7956 VDD.n7829 40.8219
R9911 VDD.n7955 VDD.n7954 40.8219
R9912 VDD.n7927 VDD.n7926 40.8219
R9913 VDD.n7853 VDD.n7849 40.8219
R9914 VDD.n7919 VDD.n7854 40.8219
R9915 VDD.n7918 VDD.n7917 40.8219
R9916 VDD.n7859 VDD.n7855 40.8219
R9917 VDD.n7910 VDD.n7860 40.8219
R9918 VDD.n7909 VDD.n7908 40.8219
R9919 VDD.n7864 VDD.n7861 40.8219
R9920 VDD.n7817 VDD.n7816 40.8219
R9921 VDD.n7974 VDD.n7973 40.8219
R9922 VDD.n7972 VDD.n7818 40.8219
R9923 VDD.n7823 VDD.n7822 40.8219
R9924 VDD.n7965 VDD.n7964 40.8219
R9925 VDD.n7963 VDD.n7824 40.8219
R9926 VDD.n7829 VDD.n7828 40.8219
R9927 VDD.n7956 VDD.n7955 40.8219
R9928 VDD.n7928 VDD.n7927 40.8219
R9929 VDD.n7926 VDD.n7849 40.8219
R9930 VDD.n7854 VDD.n7853 40.8219
R9931 VDD.n7919 VDD.n7918 40.8219
R9932 VDD.n7917 VDD.n7855 40.8219
R9933 VDD.n7860 VDD.n7859 40.8219
R9934 VDD.n7910 VDD.n7909 40.8219
R9935 VDD.n7908 VDD.n7861 40.8219
R9936 VDD.n6107 VDD.n6105 40.8219
R9937 VDD.n6384 VDD.n5896 40.8219
R9938 VDD.n5901 VDD.n5895 40.8219
R9939 VDD.n5912 VDD.n5894 40.8219
R9940 VDD.n6375 VDD.n5893 40.8219
R9941 VDD.n6372 VDD.n5892 40.8219
R9942 VDD.n5957 VDD.n5887 40.8219
R9943 VDD.n5961 VDD.n5886 40.8219
R9944 VDD.n5945 VDD.n5885 40.8219
R9945 VDD.n5967 VDD.n5884 40.8219
R9946 VDD.n5943 VDD.n5883 40.8219
R9947 VDD.n5973 VDD.n5882 40.8219
R9948 VDD.n5976 VDD.n5881 40.8219
R9949 VDD.n5880 VDD.n5878 40.8219
R9950 VDD.n6281 VDD.n6280 40.8219
R9951 VDD.n6542 VDD.n5795 40.8219
R9952 VDD.n6280 VDD.n5795 40.8219
R9953 VDD.n6282 VDD.n6281 40.8219
R9954 VDD.n6105 VDD.n6104 40.8219
R9955 VDD.n5955 VDD.n5887 40.8219
R9956 VDD.n5957 VDD.n5886 40.8219
R9957 VDD.n5961 VDD.n5885 40.8219
R9958 VDD.n5945 VDD.n5884 40.8219
R9959 VDD.n5967 VDD.n5883 40.8219
R9960 VDD.n5943 VDD.n5882 40.8219
R9961 VDD.n5973 VDD.n5881 40.8219
R9962 VDD.n5976 VDD.n5880 40.8219
R9963 VDD.n5897 VDD.n5896 40.8219
R9964 VDD.n6384 VDD.n5895 40.8219
R9965 VDD.n5901 VDD.n5894 40.8219
R9966 VDD.n5912 VDD.n5893 40.8219
R9967 VDD.n6375 VDD.n5892 40.8219
R9968 VDD.n5253 VDD.n5251 40.8219
R9969 VDD.n5530 VDD.n5042 40.8219
R9970 VDD.n5047 VDD.n5041 40.8219
R9971 VDD.n5058 VDD.n5040 40.8219
R9972 VDD.n5521 VDD.n5039 40.8219
R9973 VDD.n5518 VDD.n5038 40.8219
R9974 VDD.n5103 VDD.n5033 40.8219
R9975 VDD.n5107 VDD.n5032 40.8219
R9976 VDD.n5091 VDD.n5031 40.8219
R9977 VDD.n5113 VDD.n5030 40.8219
R9978 VDD.n5089 VDD.n5029 40.8219
R9979 VDD.n5119 VDD.n5028 40.8219
R9980 VDD.n5122 VDD.n5027 40.8219
R9981 VDD.n5026 VDD.n5024 40.8219
R9982 VDD.n5427 VDD.n5426 40.8219
R9983 VDD.n5688 VDD.n4941 40.8219
R9984 VDD.n5426 VDD.n4941 40.8219
R9985 VDD.n5428 VDD.n5427 40.8219
R9986 VDD.n5251 VDD.n5250 40.8219
R9987 VDD.n5101 VDD.n5033 40.8219
R9988 VDD.n5103 VDD.n5032 40.8219
R9989 VDD.n5107 VDD.n5031 40.8219
R9990 VDD.n5091 VDD.n5030 40.8219
R9991 VDD.n5113 VDD.n5029 40.8219
R9992 VDD.n5089 VDD.n5028 40.8219
R9993 VDD.n5119 VDD.n5027 40.8219
R9994 VDD.n5122 VDD.n5026 40.8219
R9995 VDD.n5043 VDD.n5042 40.8219
R9996 VDD.n5530 VDD.n5041 40.8219
R9997 VDD.n5047 VDD.n5040 40.8219
R9998 VDD.n5058 VDD.n5039 40.8219
R9999 VDD.n5521 VDD.n5038 40.8219
R10000 VDD.n4467 VDD.n4465 40.8219
R10001 VDD.n4744 VDD.n4256 40.8219
R10002 VDD.n4261 VDD.n4255 40.8219
R10003 VDD.n4272 VDD.n4254 40.8219
R10004 VDD.n4735 VDD.n4253 40.8219
R10005 VDD.n4732 VDD.n4252 40.8219
R10006 VDD.n4317 VDD.n4247 40.8219
R10007 VDD.n4321 VDD.n4246 40.8219
R10008 VDD.n4305 VDD.n4245 40.8219
R10009 VDD.n4327 VDD.n4244 40.8219
R10010 VDD.n4303 VDD.n4243 40.8219
R10011 VDD.n4333 VDD.n4242 40.8219
R10012 VDD.n4336 VDD.n4241 40.8219
R10013 VDD.n4240 VDD.n4238 40.8219
R10014 VDD.n4641 VDD.n4640 40.8219
R10015 VDD.n4902 VDD.n4155 40.8219
R10016 VDD.n4640 VDD.n4155 40.8219
R10017 VDD.n4642 VDD.n4641 40.8219
R10018 VDD.n4465 VDD.n4464 40.8219
R10019 VDD.n4315 VDD.n4247 40.8219
R10020 VDD.n4317 VDD.n4246 40.8219
R10021 VDD.n4321 VDD.n4245 40.8219
R10022 VDD.n4305 VDD.n4244 40.8219
R10023 VDD.n4327 VDD.n4243 40.8219
R10024 VDD.n4303 VDD.n4242 40.8219
R10025 VDD.n4333 VDD.n4241 40.8219
R10026 VDD.n4336 VDD.n4240 40.8219
R10027 VDD.n4257 VDD.n4256 40.8219
R10028 VDD.n4744 VDD.n4255 40.8219
R10029 VDD.n4261 VDD.n4254 40.8219
R10030 VDD.n4272 VDD.n4253 40.8219
R10031 VDD.n4735 VDD.n4252 40.8219
R10032 VDD.n3613 VDD.n3611 40.8219
R10033 VDD.n3890 VDD.n3402 40.8219
R10034 VDD.n3407 VDD.n3401 40.8219
R10035 VDD.n3418 VDD.n3400 40.8219
R10036 VDD.n3881 VDD.n3399 40.8219
R10037 VDD.n3878 VDD.n3398 40.8219
R10038 VDD.n3463 VDD.n3393 40.8219
R10039 VDD.n3467 VDD.n3392 40.8219
R10040 VDD.n3451 VDD.n3391 40.8219
R10041 VDD.n3473 VDD.n3390 40.8219
R10042 VDD.n3449 VDD.n3389 40.8219
R10043 VDD.n3479 VDD.n3388 40.8219
R10044 VDD.n3482 VDD.n3387 40.8219
R10045 VDD.n3386 VDD.n3384 40.8219
R10046 VDD.n3787 VDD.n3786 40.8219
R10047 VDD.n4048 VDD.n3301 40.8219
R10048 VDD.n3786 VDD.n3301 40.8219
R10049 VDD.n3788 VDD.n3787 40.8219
R10050 VDD.n3611 VDD.n3610 40.8219
R10051 VDD.n3461 VDD.n3393 40.8219
R10052 VDD.n3463 VDD.n3392 40.8219
R10053 VDD.n3467 VDD.n3391 40.8219
R10054 VDD.n3451 VDD.n3390 40.8219
R10055 VDD.n3473 VDD.n3389 40.8219
R10056 VDD.n3449 VDD.n3388 40.8219
R10057 VDD.n3479 VDD.n3387 40.8219
R10058 VDD.n3482 VDD.n3386 40.8219
R10059 VDD.n3403 VDD.n3402 40.8219
R10060 VDD.n3890 VDD.n3401 40.8219
R10061 VDD.n3407 VDD.n3400 40.8219
R10062 VDD.n3418 VDD.n3399 40.8219
R10063 VDD.n3881 VDD.n3398 40.8219
R10064 VDD.n2827 VDD.n2825 40.8219
R10065 VDD.n3104 VDD.n2616 40.8219
R10066 VDD.n2621 VDD.n2615 40.8219
R10067 VDD.n2632 VDD.n2614 40.8219
R10068 VDD.n3095 VDD.n2613 40.8219
R10069 VDD.n3092 VDD.n2612 40.8219
R10070 VDD.n2677 VDD.n2607 40.8219
R10071 VDD.n2681 VDD.n2606 40.8219
R10072 VDD.n2665 VDD.n2605 40.8219
R10073 VDD.n2687 VDD.n2604 40.8219
R10074 VDD.n2663 VDD.n2603 40.8219
R10075 VDD.n2693 VDD.n2602 40.8219
R10076 VDD.n2696 VDD.n2601 40.8219
R10077 VDD.n2600 VDD.n2598 40.8219
R10078 VDD.n3001 VDD.n3000 40.8219
R10079 VDD.n3262 VDD.n2515 40.8219
R10080 VDD.n3000 VDD.n2515 40.8219
R10081 VDD.n3002 VDD.n3001 40.8219
R10082 VDD.n2825 VDD.n2824 40.8219
R10083 VDD.n2675 VDD.n2607 40.8219
R10084 VDD.n2677 VDD.n2606 40.8219
R10085 VDD.n2681 VDD.n2605 40.8219
R10086 VDD.n2665 VDD.n2604 40.8219
R10087 VDD.n2687 VDD.n2603 40.8219
R10088 VDD.n2663 VDD.n2602 40.8219
R10089 VDD.n2693 VDD.n2601 40.8219
R10090 VDD.n2696 VDD.n2600 40.8219
R10091 VDD.n2617 VDD.n2616 40.8219
R10092 VDD.n3104 VDD.n2615 40.8219
R10093 VDD.n2621 VDD.n2614 40.8219
R10094 VDD.n2632 VDD.n2613 40.8219
R10095 VDD.n3095 VDD.n2612 40.8219
R10096 VDD.n1972 VDD.n1970 40.8219
R10097 VDD.n2249 VDD.n1761 40.8219
R10098 VDD.n1766 VDD.n1760 40.8219
R10099 VDD.n1777 VDD.n1759 40.8219
R10100 VDD.n2240 VDD.n1758 40.8219
R10101 VDD.n2237 VDD.n1757 40.8219
R10102 VDD.n1822 VDD.n1752 40.8219
R10103 VDD.n1826 VDD.n1751 40.8219
R10104 VDD.n1810 VDD.n1750 40.8219
R10105 VDD.n1832 VDD.n1749 40.8219
R10106 VDD.n1808 VDD.n1748 40.8219
R10107 VDD.n1838 VDD.n1747 40.8219
R10108 VDD.n1841 VDD.n1746 40.8219
R10109 VDD.n1745 VDD.n1743 40.8219
R10110 VDD.n2146 VDD.n2145 40.8219
R10111 VDD.n2407 VDD.n1660 40.8219
R10112 VDD.n2145 VDD.n1660 40.8219
R10113 VDD.n2147 VDD.n2146 40.8219
R10114 VDD.n1970 VDD.n1969 40.8219
R10115 VDD.n1820 VDD.n1752 40.8219
R10116 VDD.n1822 VDD.n1751 40.8219
R10117 VDD.n1826 VDD.n1750 40.8219
R10118 VDD.n1810 VDD.n1749 40.8219
R10119 VDD.n1832 VDD.n1748 40.8219
R10120 VDD.n1808 VDD.n1747 40.8219
R10121 VDD.n1838 VDD.n1746 40.8219
R10122 VDD.n1841 VDD.n1745 40.8219
R10123 VDD.n1762 VDD.n1761 40.8219
R10124 VDD.n2249 VDD.n1760 40.8219
R10125 VDD.n1766 VDD.n1759 40.8219
R10126 VDD.n1777 VDD.n1758 40.8219
R10127 VDD.n2240 VDD.n1757 40.8219
R10128 VDD.n1318 VDD.n1317 40.8219
R10129 VDD.n1373 VDD.n1372 40.8219
R10130 VDD.n1378 VDD.n1377 40.8219
R10131 VDD.n1384 VDD.n1383 40.8219
R10132 VDD.n1389 VDD.n1388 40.8219
R10133 VDD.n1395 VDD.n1394 40.8219
R10134 VDD.n1199 VDD.n1198 40.8219
R10135 VDD.n1025 VDD.n1024 40.8219
R10136 VDD.n1565 VDD.n1564 40.8219
R10137 VDD.n1562 VDD.n1561 40.8219
R10138 VDD.n1556 VDD.n1555 40.8219
R10139 VDD.n1551 VDD.n1550 40.8219
R10140 VDD.n1545 VDD.n1544 40.8219
R10141 VDD.n1540 VDD.n1539 40.8219
R10142 VDD.n1534 VDD.n1533 40.8219
R10143 VDD.n1529 VDD.n1528 40.8219
R10144 VDD.n90 VDD.n89 40.8219
R10145 VDD.n145 VDD.n144 40.8219
R10146 VDD.n150 VDD.n149 40.8219
R10147 VDD.n156 VDD.n155 40.8219
R10148 VDD.n161 VDD.n160 40.8219
R10149 VDD.n167 VDD.n166 40.8219
R10150 VDD.n753 VDD.n752 40.8219
R10151 VDD.n579 VDD.n578 40.8219
R10152 VDD.n337 VDD.n336 40.8219
R10153 VDD.n334 VDD.n333 40.8219
R10154 VDD.n328 VDD.n327 40.8219
R10155 VDD.n323 VDD.n322 40.8219
R10156 VDD.n317 VDD.n316 40.8219
R10157 VDD.n312 VDD.n311 40.8219
R10158 VDD.n306 VDD.n305 40.8219
R10159 VDD.n301 VDD.n300 40.8219
R10160 VDD.n8198 VDD.n8197 39.5838
R10161 VDD.n10054 VDD.n10028 39.5177
R10162 VDD.n10613 VDD.n10588 39.5177
R10163 VDD.n10537 VDD.n10503 39.5177
R10164 VDD.n9622 VDD.n9569 39.5177
R10165 VDD.n10747 VDD.n10746 39.5177
R10166 VDD.n8904 VDD.n8765 39.5177
R10167 VDD.n9385 VDD.n9361 39.5177
R10168 VDD.n11449 VDD.n11448 39.2068
R10169 VDD.n6729 VDD.n6728 38.7994
R10170 VDD.n6733 VDD.n6732 38.7994
R10171 VDD.n6735 VDD.n6726 38.7994
R10172 VDD.n6740 VDD.n6739 38.7994
R10173 VDD.n6038 VDD.n6037 38.7994
R10174 VDD.n6036 VDD.n6027 38.7994
R10175 VDD.n6032 VDD.n6031 38.7994
R10176 VDD.n6382 VDD.n6381 38.7994
R10177 VDD.n5792 VDD.n5782 38.7994
R10178 VDD.n6536 VDD.n5800 38.7994
R10179 VDD.n6535 VDD.n5801 38.7994
R10180 VDD.n6527 VDD.n6526 38.7994
R10181 VDD.n5184 VDD.n5183 38.7994
R10182 VDD.n5182 VDD.n5173 38.7994
R10183 VDD.n5178 VDD.n5177 38.7994
R10184 VDD.n5528 VDD.n5527 38.7994
R10185 VDD.n4938 VDD.n4928 38.7994
R10186 VDD.n5682 VDD.n4946 38.7994
R10187 VDD.n5681 VDD.n4947 38.7994
R10188 VDD.n5673 VDD.n5672 38.7994
R10189 VDD.n4398 VDD.n4397 38.7994
R10190 VDD.n4396 VDD.n4387 38.7994
R10191 VDD.n4392 VDD.n4391 38.7994
R10192 VDD.n4742 VDD.n4741 38.7994
R10193 VDD.n4152 VDD.n4142 38.7994
R10194 VDD.n4896 VDD.n4160 38.7994
R10195 VDD.n4895 VDD.n4161 38.7994
R10196 VDD.n4887 VDD.n4886 38.7994
R10197 VDD.n3544 VDD.n3543 38.7994
R10198 VDD.n3542 VDD.n3533 38.7994
R10199 VDD.n3538 VDD.n3537 38.7994
R10200 VDD.n3888 VDD.n3887 38.7994
R10201 VDD.n3298 VDD.n3288 38.7994
R10202 VDD.n4042 VDD.n3306 38.7994
R10203 VDD.n4041 VDD.n3307 38.7994
R10204 VDD.n4033 VDD.n4032 38.7994
R10205 VDD.n2758 VDD.n2757 38.7994
R10206 VDD.n2756 VDD.n2747 38.7994
R10207 VDD.n2752 VDD.n2751 38.7994
R10208 VDD.n3102 VDD.n3101 38.7994
R10209 VDD.n2512 VDD.n2502 38.7994
R10210 VDD.n3256 VDD.n2520 38.7994
R10211 VDD.n3255 VDD.n2521 38.7994
R10212 VDD.n3247 VDD.n3246 38.7994
R10213 VDD.n1903 VDD.n1902 38.7994
R10214 VDD.n1901 VDD.n1892 38.7994
R10215 VDD.n1897 VDD.n1896 38.7994
R10216 VDD.n2247 VDD.n2246 38.7994
R10217 VDD.n1657 VDD.n1647 38.7994
R10218 VDD.n2401 VDD.n1665 38.7994
R10219 VDD.n2400 VDD.n1666 38.7994
R10220 VDD.n2392 VDD.n2391 38.7994
R10221 VDD.n1194 VDD.n1191 38.7994
R10222 VDD.n1172 VDD.n1171 38.7994
R10223 VDD.n1162 VDD.n1161 38.7994
R10224 VDD.n748 VDD.n745 38.7994
R10225 VDD.n726 VDD.n725 38.7994
R10226 VDD.n716 VDD.n715 38.7994
R10227 VDD.n6734 VDD.n6733 38.7989
R10228 VDD.n6738 VDD.n6726 38.7989
R10229 VDD.n6741 VDD.n6740 38.7989
R10230 VDD.n6728 VDD.n6715 38.7989
R10231 VDD.n6033 VDD.n6027 38.7989
R10232 VDD.n6031 VDD.n6030 38.7989
R10233 VDD.n6039 VDD.n6038 38.7989
R10234 VDD.n6381 VDD.n5904 38.7989
R10235 VDD.n6546 VDD.n5792 38.7989
R10236 VDD.n6526 VDD.n6525 38.7989
R10237 VDD.n5806 VDD.n5801 38.7989
R10238 VDD.n5800 VDD.n5793 38.7989
R10239 VDD.n5179 VDD.n5173 38.7989
R10240 VDD.n5177 VDD.n5176 38.7989
R10241 VDD.n5185 VDD.n5184 38.7989
R10242 VDD.n5527 VDD.n5050 38.7989
R10243 VDD.n5692 VDD.n4938 38.7989
R10244 VDD.n5672 VDD.n5671 38.7989
R10245 VDD.n4952 VDD.n4947 38.7989
R10246 VDD.n4946 VDD.n4939 38.7989
R10247 VDD.n4393 VDD.n4387 38.7989
R10248 VDD.n4391 VDD.n4390 38.7989
R10249 VDD.n4399 VDD.n4398 38.7989
R10250 VDD.n4741 VDD.n4264 38.7989
R10251 VDD.n4906 VDD.n4152 38.7989
R10252 VDD.n4886 VDD.n4885 38.7989
R10253 VDD.n4166 VDD.n4161 38.7989
R10254 VDD.n4160 VDD.n4153 38.7989
R10255 VDD.n3539 VDD.n3533 38.7989
R10256 VDD.n3537 VDD.n3536 38.7989
R10257 VDD.n3545 VDD.n3544 38.7989
R10258 VDD.n3887 VDD.n3410 38.7989
R10259 VDD.n4052 VDD.n3298 38.7989
R10260 VDD.n4032 VDD.n4031 38.7989
R10261 VDD.n3312 VDD.n3307 38.7989
R10262 VDD.n3306 VDD.n3299 38.7989
R10263 VDD.n2753 VDD.n2747 38.7989
R10264 VDD.n2751 VDD.n2750 38.7989
R10265 VDD.n2759 VDD.n2758 38.7989
R10266 VDD.n3101 VDD.n2624 38.7989
R10267 VDD.n3266 VDD.n2512 38.7989
R10268 VDD.n3246 VDD.n3245 38.7989
R10269 VDD.n2526 VDD.n2521 38.7989
R10270 VDD.n2520 VDD.n2513 38.7989
R10271 VDD.n1898 VDD.n1892 38.7989
R10272 VDD.n1896 VDD.n1895 38.7989
R10273 VDD.n1904 VDD.n1903 38.7989
R10274 VDD.n2246 VDD.n1769 38.7989
R10275 VDD.n2411 VDD.n1657 38.7989
R10276 VDD.n2391 VDD.n2390 38.7989
R10277 VDD.n1671 VDD.n1666 38.7989
R10278 VDD.n1665 VDD.n1658 38.7989
R10279 VDD.n1234 VDD.n1233 38.7989
R10280 VDD.n1242 VDD.n1240 38.7989
R10281 VDD.n1381 VDD.n1380 38.7989
R10282 VDD.n1194 VDD.n1193 38.7989
R10283 VDD.n1183 VDD.n1182 38.7989
R10284 VDD.n6 VDD.n5 38.7989
R10285 VDD.n14 VDD.n12 38.7989
R10286 VDD.n153 VDD.n152 38.7989
R10287 VDD.n748 VDD.n747 38.7989
R10288 VDD.n737 VDD.n736 38.7989
R10289 VDD.n6379 VDD.n5910 38.7987
R10290 VDD.n6366 VDD.n5909 38.7987
R10291 VDD.n6379 VDD.n6378 38.7987
R10292 VDD.n6370 VDD.n5909 38.7987
R10293 VDD.n5964 VDD.n5908 38.7987
R10294 VDD.n5970 VDD.n5907 38.7987
R10295 VDD.n5979 VDD.n5906 38.7987
R10296 VDD.n5971 VDD.n5906 38.7987
R10297 VDD.n5965 VDD.n5907 38.7987
R10298 VDD.n5959 VDD.n5908 38.7987
R10299 VDD.n5525 VDD.n5056 38.7987
R10300 VDD.n5512 VDD.n5055 38.7987
R10301 VDD.n5525 VDD.n5524 38.7987
R10302 VDD.n5516 VDD.n5055 38.7987
R10303 VDD.n5110 VDD.n5054 38.7987
R10304 VDD.n5116 VDD.n5053 38.7987
R10305 VDD.n5125 VDD.n5052 38.7987
R10306 VDD.n5117 VDD.n5052 38.7987
R10307 VDD.n5111 VDD.n5053 38.7987
R10308 VDD.n5105 VDD.n5054 38.7987
R10309 VDD.n4739 VDD.n4270 38.7987
R10310 VDD.n4726 VDD.n4269 38.7987
R10311 VDD.n4739 VDD.n4738 38.7987
R10312 VDD.n4730 VDD.n4269 38.7987
R10313 VDD.n4324 VDD.n4268 38.7987
R10314 VDD.n4330 VDD.n4267 38.7987
R10315 VDD.n4339 VDD.n4266 38.7987
R10316 VDD.n4331 VDD.n4266 38.7987
R10317 VDD.n4325 VDD.n4267 38.7987
R10318 VDD.n4319 VDD.n4268 38.7987
R10319 VDD.n3885 VDD.n3416 38.7987
R10320 VDD.n3872 VDD.n3415 38.7987
R10321 VDD.n3885 VDD.n3884 38.7987
R10322 VDD.n3876 VDD.n3415 38.7987
R10323 VDD.n3470 VDD.n3414 38.7987
R10324 VDD.n3476 VDD.n3413 38.7987
R10325 VDD.n3485 VDD.n3412 38.7987
R10326 VDD.n3477 VDD.n3412 38.7987
R10327 VDD.n3471 VDD.n3413 38.7987
R10328 VDD.n3465 VDD.n3414 38.7987
R10329 VDD.n3099 VDD.n2630 38.7987
R10330 VDD.n3086 VDD.n2629 38.7987
R10331 VDD.n3099 VDD.n3098 38.7987
R10332 VDD.n3090 VDD.n2629 38.7987
R10333 VDD.n2684 VDD.n2628 38.7987
R10334 VDD.n2690 VDD.n2627 38.7987
R10335 VDD.n2699 VDD.n2626 38.7987
R10336 VDD.n2691 VDD.n2626 38.7987
R10337 VDD.n2685 VDD.n2627 38.7987
R10338 VDD.n2679 VDD.n2628 38.7987
R10339 VDD.n2244 VDD.n1775 38.7987
R10340 VDD.n2231 VDD.n1774 38.7987
R10341 VDD.n2244 VDD.n2243 38.7987
R10342 VDD.n2235 VDD.n1774 38.7987
R10343 VDD.n1829 VDD.n1773 38.7987
R10344 VDD.n1835 VDD.n1772 38.7987
R10345 VDD.n1844 VDD.n1771 38.7987
R10346 VDD.n1836 VDD.n1771 38.7987
R10347 VDD.n1830 VDD.n1772 38.7987
R10348 VDD.n1824 VDD.n1773 38.7987
R10349 VDD.n1392 VDD.n1391 38.7987
R10350 VDD.n1404 VDD.n1403 38.7987
R10351 VDD.n1537 VDD.n1536 38.7987
R10352 VDD.n1548 VDD.n1547 38.7987
R10353 VDD.n1559 VDD.n1558 38.7987
R10354 VDD.n164 VDD.n163 38.7987
R10355 VDD.n176 VDD.n175 38.7987
R10356 VDD.n309 VDD.n308 38.7987
R10357 VDD.n320 VDD.n319 38.7987
R10358 VDD.n331 VDD.n330 38.7987
R10359 VDD.n8571 VDD.n7761 38.777
R10360 VDD.n10429 VDD.n10427 38.4005
R10361 VDD.n6364 VDD.n6363 36.539
R10362 VDD.n6356 VDD.n5924 36.539
R10363 VDD.n5510 VDD.n5509 36.539
R10364 VDD.n5502 VDD.n5070 36.539
R10365 VDD.n4724 VDD.n4723 36.539
R10366 VDD.n4716 VDD.n4284 36.539
R10367 VDD.n3870 VDD.n3869 36.539
R10368 VDD.n3862 VDD.n3430 36.539
R10369 VDD.n3084 VDD.n3083 36.539
R10370 VDD.n3076 VDD.n2644 36.539
R10371 VDD.n2229 VDD.n2228 36.539
R10372 VDD.n2221 VDD.n1789 36.539
R10373 VDD.n9423 VDD.n9403 36.2246
R10374 VDD.n10430 VDD.n10429 36.2136
R10375 VDD.n9968 VDD.n9967 36.1417
R10376 VDD.n9967 VDD.n9908 36.1417
R10377 VDD.n9959 VDD.n9908 36.1417
R10378 VDD.n9960 VDD.n9959 36.1417
R10379 VDD.n9945 VDD.n9913 36.1417
R10380 VDD.n9945 VDD.n9915 36.1417
R10381 VDD.n9920 VDD.n9915 36.1417
R10382 VDD.n9938 VDD.n9920 36.1417
R10383 VDD.n9938 VDD.n9921 36.1417
R10384 VDD.n9933 VDD.n9921 36.1417
R10385 VDD.n9933 VDD.n9931 36.1417
R10386 VDD.n5760 VDD.n5744 36.1417
R10387 VDD.n5760 VDD.n5759 36.1417
R10388 VDD.n5759 VDD.n5748 36.1417
R10389 VDD.n5755 VDD.n5748 36.1417
R10390 VDD.n5725 VDD.n5717 36.1417
R10391 VDD.n5736 VDD.n5717 36.1417
R10392 VDD.n5736 VDD.n5713 36.1417
R10393 VDD.n5767 VDD.n5713 36.1417
R10394 VDD.n4120 VDD.n4104 36.1417
R10395 VDD.n4120 VDD.n4119 36.1417
R10396 VDD.n4119 VDD.n4108 36.1417
R10397 VDD.n4115 VDD.n4108 36.1417
R10398 VDD.n4085 VDD.n4077 36.1417
R10399 VDD.n4096 VDD.n4077 36.1417
R10400 VDD.n4096 VDD.n4073 36.1417
R10401 VDD.n4127 VDD.n4073 36.1417
R10402 VDD.n2480 VDD.n2463 36.1417
R10403 VDD.n2480 VDD.n2479 36.1417
R10404 VDD.n2479 VDD.n2467 36.1417
R10405 VDD.n2475 VDD.n2467 36.1417
R10406 VDD.n2444 VDD.n2436 36.1417
R10407 VDD.n2455 VDD.n2436 36.1417
R10408 VDD.n2455 VDD.n2432 36.1417
R10409 VDD.n2487 VDD.n2432 36.1417
R10410 VDD.n840 VDD.n823 36.1417
R10411 VDD.n840 VDD.n839 36.1417
R10412 VDD.n839 VDD.n827 36.1417
R10413 VDD.n835 VDD.n827 36.1417
R10414 VDD.n804 VDD.n796 36.1417
R10415 VDD.n815 VDD.n796 36.1417
R10416 VDD.n815 VDD.n792 36.1417
R10417 VDD.n847 VDD.n792 36.1417
R10418 VDD.n6488 VDD.n5826 35.9626
R10419 VDD.n5634 VDD.n4972 35.9626
R10420 VDD.n4848 VDD.n4186 35.9626
R10421 VDD.n3994 VDD.n3332 35.9626
R10422 VDD.n3208 VDD.n2546 35.9626
R10423 VDD.n2353 VDD.n1691 35.9626
R10424 VDD.n1070 VDD.n1069 35.9626
R10425 VDD.n624 VDD.n623 35.9626
R10426 VDD.n6391 VDD.n5879 35.2569
R10427 VDD.n5537 VDD.n5025 35.2569
R10428 VDD.n4751 VDD.n4239 35.2569
R10429 VDD.n3897 VDD.n3385 35.2569
R10430 VDD.n3111 VDD.n2599 35.2569
R10431 VDD.n2256 VDD.n1744 35.2569
R10432 VDD.n1411 VDD.n1410 35.2569
R10433 VDD.n183 VDD.n182 35.2569
R10434 VDD.n12407 VDD.n6934 34.6359
R10435 VDD.n6249 VDD.n5796 34.6159
R10436 VDD.n5395 VDD.n4942 34.6159
R10437 VDD.n4609 VDD.n4156 34.6159
R10438 VDD.n3755 VDD.n3302 34.6159
R10439 VDD.n2969 VDD.n2516 34.6159
R10440 VDD.n2114 VDD.n1661 34.6159
R10441 VDD.n1017 VDD.n1016 34.6159
R10442 VDD.n571 VDD.n570 34.6159
R10443 VDD.n11648 VDD.n11647 34.3808
R10444 VDD.n12090 VDD.n12089 34.3388
R10445 VDD.n8542 VDD.n8541 34.2989
R10446 VDD.n8123 VDD.n8122 33.9026
R10447 VDD.n8197 VDD.n8196 33.8538
R10448 VDD.n6634 VDD.n6580 33.8538
R10449 VDD.n8197 VDD.n8093 33.8536
R10450 VDD.n6595 VDD.n6580 33.8536
R10451 VDD.n8124 VDD.n8116 33.4435
R10452 VDD.n8115 VDD.n8113 33.4435
R10453 VDD.n8188 VDD.n8187 33.4435
R10454 VDD.n8134 VDD.n8126 33.4435
R10455 VDD.n8176 VDD.n8135 33.4435
R10456 VDD.n8167 VDD.n8166 33.4435
R10457 VDD.n8152 VDD.n8144 33.4435
R10458 VDD.n6934 VDD.n6933 33.4435
R10459 VDD.n12412 VDD.n12411 33.4435
R10460 VDD.n7127 VDD.n7069 33.4435
R10461 VDD.n12090 VDD.n7372 33.4435
R10462 VDD.n11644 VDD.n11643 33.4435
R10463 VDD.n11648 VDD.n7610 33.4435
R10464 VDD.n8542 VDD.n7783 33.4435
R10465 VDD.n8538 VDD.n8537 33.4435
R10466 VDD.n8535 VDD.n7786 33.4435
R10467 VDD.n8528 VDD.n8527 33.4435
R10468 VDD.n7797 VDD.n7793 33.4435
R10469 VDD.n8518 VDD.n8517 33.4435
R10470 VDD.n7803 VDD.n7798 33.4435
R10471 VDD.n8508 VDD.n7804 33.4435
R10472 VDD.n8123 VDD.n8112 33.4435
R10473 VDD.n11219 VDD.n11217 33.4435
R10474 VDD.n5864 VDD.n5861 33.4435
R10475 VDD.n5827 VDD.n5825 33.4435
R10476 VDD.n6520 VDD.n6519 33.4435
R10477 VDD.n6539 VDD.n5797 33.4435
R10478 VDD.n6532 VDD.n6531 33.4435
R10479 VDD.n5809 VDD.n5804 33.4435
R10480 VDD.n6265 VDD.n6264 33.4435
R10481 VDD.n6266 VDD.n6049 33.4435
R10482 VDD.n6279 VDD.n6278 33.4435
R10483 VDD.n6213 VDD.n6072 33.4435
R10484 VDD.n6220 VDD.n6073 33.4435
R10485 VDD.n6157 VDD.n6102 33.4435
R10486 VDD.n5010 VDD.n5007 33.4435
R10487 VDD.n4973 VDD.n4971 33.4435
R10488 VDD.n5666 VDD.n5665 33.4435
R10489 VDD.n5685 VDD.n4943 33.4435
R10490 VDD.n5678 VDD.n5677 33.4435
R10491 VDD.n4955 VDD.n4950 33.4435
R10492 VDD.n5411 VDD.n5410 33.4435
R10493 VDD.n5412 VDD.n5195 33.4435
R10494 VDD.n5425 VDD.n5424 33.4435
R10495 VDD.n5359 VDD.n5218 33.4435
R10496 VDD.n5366 VDD.n5219 33.4435
R10497 VDD.n5303 VDD.n5248 33.4435
R10498 VDD.n4224 VDD.n4221 33.4435
R10499 VDD.n4187 VDD.n4185 33.4435
R10500 VDD.n4880 VDD.n4879 33.4435
R10501 VDD.n4899 VDD.n4157 33.4435
R10502 VDD.n4892 VDD.n4891 33.4435
R10503 VDD.n4169 VDD.n4164 33.4435
R10504 VDD.n4625 VDD.n4624 33.4435
R10505 VDD.n4626 VDD.n4409 33.4435
R10506 VDD.n4639 VDD.n4638 33.4435
R10507 VDD.n4573 VDD.n4432 33.4435
R10508 VDD.n4580 VDD.n4433 33.4435
R10509 VDD.n4517 VDD.n4462 33.4435
R10510 VDD.n3370 VDD.n3367 33.4435
R10511 VDD.n3333 VDD.n3331 33.4435
R10512 VDD.n4026 VDD.n4025 33.4435
R10513 VDD.n4045 VDD.n3303 33.4435
R10514 VDD.n4038 VDD.n4037 33.4435
R10515 VDD.n3315 VDD.n3310 33.4435
R10516 VDD.n3771 VDD.n3770 33.4435
R10517 VDD.n3772 VDD.n3555 33.4435
R10518 VDD.n3785 VDD.n3784 33.4435
R10519 VDD.n3719 VDD.n3578 33.4435
R10520 VDD.n3726 VDD.n3579 33.4435
R10521 VDD.n3663 VDD.n3608 33.4435
R10522 VDD.n2584 VDD.n2581 33.4435
R10523 VDD.n2547 VDD.n2545 33.4435
R10524 VDD.n3240 VDD.n3239 33.4435
R10525 VDD.n3259 VDD.n2517 33.4435
R10526 VDD.n3252 VDD.n3251 33.4435
R10527 VDD.n2529 VDD.n2524 33.4435
R10528 VDD.n2985 VDD.n2984 33.4435
R10529 VDD.n2986 VDD.n2769 33.4435
R10530 VDD.n2999 VDD.n2998 33.4435
R10531 VDD.n2933 VDD.n2792 33.4435
R10532 VDD.n2940 VDD.n2793 33.4435
R10533 VDD.n2877 VDD.n2822 33.4435
R10534 VDD.n1729 VDD.n1726 33.4435
R10535 VDD.n1692 VDD.n1690 33.4435
R10536 VDD.n2385 VDD.n2384 33.4435
R10537 VDD.n2404 VDD.n1662 33.4435
R10538 VDD.n2397 VDD.n2396 33.4435
R10539 VDD.n1674 VDD.n1669 33.4435
R10540 VDD.n2130 VDD.n2129 33.4435
R10541 VDD.n2131 VDD.n1914 33.4435
R10542 VDD.n2144 VDD.n2143 33.4435
R10543 VDD.n2078 VDD.n1937 33.4435
R10544 VDD.n2085 VDD.n1938 33.4435
R10545 VDD.n2022 VDD.n1967 33.4435
R10546 VDD.n1464 VDD.n1463 33.4435
R10547 VDD.n1079 VDD.n1078 33.4435
R10548 VDD.n1179 VDD.n1178 33.4435
R10549 VDD.n1169 VDD.n1168 33.4435
R10550 VDD.n1159 VDD.n1158 33.4435
R10551 VDD.n1310 VDD.n1307 33.4435
R10552 VDD.n236 VDD.n235 33.4435
R10553 VDD.n633 VDD.n632 33.4435
R10554 VDD.n733 VDD.n732 33.4435
R10555 VDD.n723 VDD.n722 33.4435
R10556 VDD.n713 VDD.n712 33.4435
R10557 VDD.n82 VDD.n79 33.4435
R10558 VDD.n8113 VDD.n8111 33.4431
R10559 VDD.n8187 VDD.n8186 33.4431
R10560 VDD.n8177 VDD.n8134 33.4431
R10561 VDD.n8143 VDD.n8135 33.4431
R10562 VDD.n8166 VDD.n8165 33.4431
R10563 VDD.n8153 VDD.n8152 33.4431
R10564 VDD.n12411 VDD.n12410 33.4431
R10565 VDD.n6936 VDD.n6934 33.4431
R10566 VDD.n7132 VDD.n7127 33.4431
R10567 VDD.n12091 VDD.n12090 33.4431
R10568 VDD.n11649 VDD.n11648 33.4431
R10569 VDD.n11643 VDD.n7612 33.4431
R10570 VDD.n7808 VDD.n7804 33.4431
R10571 VDD.n8509 VDD.n7803 33.4431
R10572 VDD.n8517 VDD.n8516 33.4431
R10573 VDD.n8519 VDD.n7797 33.4431
R10574 VDD.n8527 VDD.n8526 33.4431
R10575 VDD.n7792 VDD.n7786 33.4431
R10576 VDD.n8537 VDD.n8536 33.4431
R10577 VDD.n8543 VDD.n8542 33.4431
R10578 VDD.n11217 VDD.n11216 33.4431
R10579 VDD.n12696 VDD.n6613 33.4431
R10580 VDD.n5861 VDD.n5860 33.4431
R10581 VDD.n5828 VDD.n5827 33.4431
R10582 VDD.n6521 VDD.n6520 33.4431
R10583 VDD.n6522 VDD.n5809 33.4431
R10584 VDD.n6531 VDD.n6530 33.4431
R10585 VDD.n5803 VDD.n5797 33.4431
R10586 VDD.n6285 VDD.n6279 33.4431
R10587 VDD.n6277 VDD.n6049 33.4431
R10588 VDD.n6267 VDD.n6265 33.4431
R10589 VDD.n6220 VDD.n6219 33.4431
R10590 VDD.n6215 VDD.n6072 33.4431
R10591 VDD.n6158 VDD.n6157 33.4431
R10592 VDD.n5007 VDD.n5006 33.4431
R10593 VDD.n4974 VDD.n4973 33.4431
R10594 VDD.n5667 VDD.n5666 33.4431
R10595 VDD.n5668 VDD.n4955 33.4431
R10596 VDD.n5677 VDD.n5676 33.4431
R10597 VDD.n4949 VDD.n4943 33.4431
R10598 VDD.n5431 VDD.n5425 33.4431
R10599 VDD.n5423 VDD.n5195 33.4431
R10600 VDD.n5413 VDD.n5411 33.4431
R10601 VDD.n5366 VDD.n5365 33.4431
R10602 VDD.n5361 VDD.n5218 33.4431
R10603 VDD.n5304 VDD.n5303 33.4431
R10604 VDD.n4221 VDD.n4220 33.4431
R10605 VDD.n4188 VDD.n4187 33.4431
R10606 VDD.n4881 VDD.n4880 33.4431
R10607 VDD.n4882 VDD.n4169 33.4431
R10608 VDD.n4891 VDD.n4890 33.4431
R10609 VDD.n4163 VDD.n4157 33.4431
R10610 VDD.n4645 VDD.n4639 33.4431
R10611 VDD.n4637 VDD.n4409 33.4431
R10612 VDD.n4627 VDD.n4625 33.4431
R10613 VDD.n4580 VDD.n4579 33.4431
R10614 VDD.n4575 VDD.n4432 33.4431
R10615 VDD.n4518 VDD.n4517 33.4431
R10616 VDD.n3367 VDD.n3366 33.4431
R10617 VDD.n3334 VDD.n3333 33.4431
R10618 VDD.n4027 VDD.n4026 33.4431
R10619 VDD.n4028 VDD.n3315 33.4431
R10620 VDD.n4037 VDD.n4036 33.4431
R10621 VDD.n3309 VDD.n3303 33.4431
R10622 VDD.n3791 VDD.n3785 33.4431
R10623 VDD.n3783 VDD.n3555 33.4431
R10624 VDD.n3773 VDD.n3771 33.4431
R10625 VDD.n3726 VDD.n3725 33.4431
R10626 VDD.n3721 VDD.n3578 33.4431
R10627 VDD.n3664 VDD.n3663 33.4431
R10628 VDD.n2581 VDD.n2580 33.4431
R10629 VDD.n2548 VDD.n2547 33.4431
R10630 VDD.n3241 VDD.n3240 33.4431
R10631 VDD.n3242 VDD.n2529 33.4431
R10632 VDD.n3251 VDD.n3250 33.4431
R10633 VDD.n2523 VDD.n2517 33.4431
R10634 VDD.n3005 VDD.n2999 33.4431
R10635 VDD.n2997 VDD.n2769 33.4431
R10636 VDD.n2987 VDD.n2985 33.4431
R10637 VDD.n2940 VDD.n2939 33.4431
R10638 VDD.n2935 VDD.n2792 33.4431
R10639 VDD.n2878 VDD.n2877 33.4431
R10640 VDD.n1726 VDD.n1725 33.4431
R10641 VDD.n1693 VDD.n1692 33.4431
R10642 VDD.n2386 VDD.n2385 33.4431
R10643 VDD.n2387 VDD.n1674 33.4431
R10644 VDD.n2396 VDD.n2395 33.4431
R10645 VDD.n1668 VDD.n1662 33.4431
R10646 VDD.n2150 VDD.n2144 33.4431
R10647 VDD.n2142 VDD.n1914 33.4431
R10648 VDD.n2132 VDD.n2130 33.4431
R10649 VDD.n2085 VDD.n2084 33.4431
R10650 VDD.n2080 VDD.n1937 33.4431
R10651 VDD.n2023 VDD.n2022 33.4431
R10652 VDD.n1152 VDD.n1151 33.4431
R10653 VDD.n1019 VDD.n1018 33.4431
R10654 VDD.n1006 VDD.n1005 33.4431
R10655 VDD.n995 VDD.n994 33.4431
R10656 VDD.n934 VDD.n933 33.4431
R10657 VDD.n928 VDD.n927 33.4431
R10658 VDD.n1310 VDD.n1309 33.4431
R10659 VDD.n706 VDD.n705 33.4431
R10660 VDD.n573 VDD.n572 33.4431
R10661 VDD.n560 VDD.n559 33.4431
R10662 VDD.n549 VDD.n548 33.4431
R10663 VDD.n488 VDD.n487 33.4431
R10664 VDD.n482 VDD.n481 33.4431
R10665 VDD.n82 VDD.n81 33.4431
R10666 VDD.n7133 VDD.n7123 33.4428
R10667 VDD.n7144 VDD.n7142 33.4428
R10668 VDD.n7151 VDD.n7119 33.4428
R10669 VDD.n7152 VDD.n7115 33.4428
R10670 VDD.n7163 VDD.n7162 33.4428
R10671 VDD.n7164 VDD.n7111 33.4428
R10672 VDD.n7175 VDD.n7173 33.4428
R10673 VDD.n7182 VDD.n7107 33.4428
R10674 VDD.n7183 VDD.n7103 33.4428
R10675 VDD.n7194 VDD.n7192 33.4428
R10676 VDD.n7201 VDD.n7099 33.4428
R10677 VDD.n7202 VDD.n7095 33.4428
R10678 VDD.n7214 VDD.n7211 33.4428
R10679 VDD.n7212 VDD.n7091 33.4428
R10680 VDD.n7225 VDD.n7223 33.4428
R10681 VDD.n7232 VDD.n7087 33.4428
R10682 VDD.n7233 VDD.n7083 33.4428
R10683 VDD.n7244 VDD.n7242 33.4428
R10684 VDD.n7251 VDD.n7079 33.4428
R10685 VDD.n7252 VDD.n7073 33.4428
R10686 VDD.n7946 VDD.n7945 33.4428
R10687 VDD.n7938 VDD.n7840 33.4428
R10688 VDD.n7936 VDD.n7935 33.4428
R10689 VDD.n7900 VDD.n7899 33.4428
R10690 VDD.n7892 VDD.n7872 33.4428
R10691 VDD.n7890 VDD.n7889 33.4428
R10692 VDD.n7882 VDD.n7881 33.4428
R10693 VDD.n7134 VDD.n7133 33.4428
R10694 VDD.n7142 VDD.n7141 33.4428
R10695 VDD.n7143 VDD.n7119 33.4428
R10696 VDD.n7153 VDD.n7152 33.4428
R10697 VDD.n7162 VDD.n7161 33.4428
R10698 VDD.n7165 VDD.n7164 33.4428
R10699 VDD.n7173 VDD.n7172 33.4428
R10700 VDD.n7174 VDD.n7107 33.4428
R10701 VDD.n7184 VDD.n7183 33.4428
R10702 VDD.n7192 VDD.n7191 33.4428
R10703 VDD.n7193 VDD.n7099 33.4428
R10704 VDD.n7203 VDD.n7202 33.4428
R10705 VDD.n7211 VDD.n7210 33.4428
R10706 VDD.n7213 VDD.n7212 33.4428
R10707 VDD.n7223 VDD.n7222 33.4428
R10708 VDD.n7224 VDD.n7087 33.4428
R10709 VDD.n7234 VDD.n7233 33.4428
R10710 VDD.n7242 VDD.n7241 33.4428
R10711 VDD.n7243 VDD.n7079 33.4428
R10712 VDD.n7253 VDD.n7252 33.4428
R10713 VDD.n7947 VDD.n7946 33.4428
R10714 VDD.n7840 VDD.n7836 33.4428
R10715 VDD.n7937 VDD.n7936 33.4428
R10716 VDD.n7901 VDD.n7900 33.4428
R10717 VDD.n7872 VDD.n7868 33.4428
R10718 VDD.n7891 VDD.n7890 33.4428
R10719 VDD.n7881 VDD.n7874 33.4428
R10720 VDD.n6620 VDD.n6619 33.4428
R10721 VDD.n5952 VDD.n5889 33.4428
R10722 VDD.n5949 VDD.n5889 33.4428
R10723 VDD.n5098 VDD.n5035 33.4428
R10724 VDD.n5095 VDD.n5035 33.4428
R10725 VDD.n4312 VDD.n4249 33.4428
R10726 VDD.n4309 VDD.n4249 33.4428
R10727 VDD.n3458 VDD.n3395 33.4428
R10728 VDD.n3455 VDD.n3395 33.4428
R10729 VDD.n2672 VDD.n2609 33.4428
R10730 VDD.n2669 VDD.n2609 33.4428
R10731 VDD.n1817 VDD.n1754 33.4428
R10732 VDD.n1814 VDD.n1754 33.4428
R10733 VDD.n1413 VDD.n1412 33.4428
R10734 VDD.n185 VDD.n184 33.4428
R10735 VDD.n6424 VDD.n5857 32.9658
R10736 VDD.n5570 VDD.n5003 32.9658
R10737 VDD.n4784 VDD.n4217 32.9658
R10738 VDD.n3930 VDD.n3363 32.9658
R10739 VDD.n3144 VDD.n2577 32.9658
R10740 VDD.n2289 VDD.n1722 32.9658
R10741 VDD.n1455 VDD.n1454 32.9658
R10742 VDD.n227 VDD.n226 32.9658
R10743 VDD.n10066 VDD.n10063 32.9315
R10744 VDD.n10625 VDD.n10624 32.9315
R10745 VDD.n10564 VDD.n10563 32.9315
R10746 VDD.n9615 VDD.n9573 32.9315
R10747 VDD.n10721 VDD.n10720 32.9315
R10748 VDD.n9441 VDD.n9440 32.9315
R10749 VDD.n6157 VDD.n6156 32.6607
R10750 VDD.n5303 VDD.n5302 32.6607
R10751 VDD.n4517 VDD.n4516 32.6607
R10752 VDD.n3663 VDD.n3662 32.6607
R10753 VDD.n2877 VDD.n2876 32.6607
R10754 VDD.n2022 VDD.n2021 32.6607
R10755 VDD.n1311 VDD.n1310 32.6607
R10756 VDD.n83 VDD.n82 32.6607
R10757 VDD.n12473 VDD.n12472 31.4488
R10758 VDD.n6553 VDD.n5784 30.1287
R10759 VDD.n5699 VDD.n4930 30.1287
R10760 VDD.n4913 VDD.n4144 30.1287
R10761 VDD.n4059 VDD.n3290 30.1287
R10762 VDD.n3273 VDD.n2504 30.1287
R10763 VDD.n2418 VDD.n1649 30.1287
R10764 VDD.n6041 VDD.n6040 30.1181
R10765 VDD.n6321 VDD.n6320 30.1181
R10766 VDD.n6309 VDD.n5787 30.1181
R10767 VDD.n6347 VDD.n5934 30.1181
R10768 VDD.n6003 VDD.n6002 30.1181
R10769 VDD.n5187 VDD.n5186 30.1181
R10770 VDD.n5467 VDD.n5466 30.1181
R10771 VDD.n5455 VDD.n4933 30.1181
R10772 VDD.n5493 VDD.n5080 30.1181
R10773 VDD.n5149 VDD.n5148 30.1181
R10774 VDD.n4401 VDD.n4400 30.1181
R10775 VDD.n4681 VDD.n4680 30.1181
R10776 VDD.n4669 VDD.n4147 30.1181
R10777 VDD.n4707 VDD.n4294 30.1181
R10778 VDD.n4363 VDD.n4362 30.1181
R10779 VDD.n3547 VDD.n3546 30.1181
R10780 VDD.n3827 VDD.n3826 30.1181
R10781 VDD.n3815 VDD.n3293 30.1181
R10782 VDD.n3853 VDD.n3440 30.1181
R10783 VDD.n3509 VDD.n3508 30.1181
R10784 VDD.n2761 VDD.n2760 30.1181
R10785 VDD.n3041 VDD.n3040 30.1181
R10786 VDD.n3029 VDD.n2507 30.1181
R10787 VDD.n3067 VDD.n2654 30.1181
R10788 VDD.n2723 VDD.n2722 30.1181
R10789 VDD.n1906 VDD.n1905 30.1181
R10790 VDD.n2186 VDD.n2185 30.1181
R10791 VDD.n2174 VDD.n1652 30.1181
R10792 VDD.n2212 VDD.n1799 30.1181
R10793 VDD.n1868 VDD.n1867 30.1181
R10794 VDD.n866 VDD.n861 30.1181
R10795 VDD.n1218 VDD.n1214 30.1181
R10796 VDD.n1141 VDD.n1130 30.1181
R10797 VDD.n1598 VDD.n1260 30.1181
R10798 VDD.n1516 VDD.n1515 30.1181
R10799 VDD.n420 VDD.n415 30.1181
R10800 VDD.n772 VDD.n768 30.1181
R10801 VDD.n695 VDD.n684 30.1181
R10802 VDD.n370 VDD.n32 30.1181
R10803 VDD.n288 VDD.n287 30.1181
R10804 VDD.n6261 VDD.n6260 30.0704
R10805 VDD.n6319 VDD.n6318 30.0704
R10806 VDD.n5991 VDD.n5990 30.0704
R10807 VDD.n5407 VDD.n5406 30.0704
R10808 VDD.n5465 VDD.n5464 30.0704
R10809 VDD.n5137 VDD.n5136 30.0704
R10810 VDD.n4621 VDD.n4620 30.0704
R10811 VDD.n4679 VDD.n4678 30.0704
R10812 VDD.n4351 VDD.n4350 30.0704
R10813 VDD.n3767 VDD.n3766 30.0704
R10814 VDD.n3825 VDD.n3824 30.0704
R10815 VDD.n3497 VDD.n3496 30.0704
R10816 VDD.n2981 VDD.n2980 30.0704
R10817 VDD.n3039 VDD.n3038 30.0704
R10818 VDD.n2711 VDD.n2710 30.0704
R10819 VDD.n2126 VDD.n2125 30.0704
R10820 VDD.n2184 VDD.n2183 30.0704
R10821 VDD.n1856 VDD.n1855 30.0704
R10822 VDD.n988 VDD.n987 30.0704
R10823 VDD.n1213 VDD.n1212 30.0704
R10824 VDD.n1259 VDD.n1258 30.0704
R10825 VDD.n542 VDD.n541 30.0704
R10826 VDD.n767 VDD.n766 30.0704
R10827 VDD.n31 VDD.n30 30.0704
R10828 VDD.n6001 VDD.n6000 30.0702
R10829 VDD.n6272 VDD.n6046 30.0702
R10830 VDD.n6308 VDD.n6305 30.0702
R10831 VDD.n5147 VDD.n5146 30.0702
R10832 VDD.n5418 VDD.n5192 30.0702
R10833 VDD.n5454 VDD.n5451 30.0702
R10834 VDD.n4361 VDD.n4360 30.0702
R10835 VDD.n4632 VDD.n4406 30.0702
R10836 VDD.n4668 VDD.n4665 30.0702
R10837 VDD.n3507 VDD.n3506 30.0702
R10838 VDD.n3778 VDD.n3552 30.0702
R10839 VDD.n3814 VDD.n3811 30.0702
R10840 VDD.n2721 VDD.n2720 30.0702
R10841 VDD.n2992 VDD.n2766 30.0702
R10842 VDD.n3028 VDD.n3025 30.0702
R10843 VDD.n1866 VDD.n1865 30.0702
R10844 VDD.n2137 VDD.n1911 30.0702
R10845 VDD.n2173 VDD.n2170 30.0702
R10846 VDD.n1010 VDD.n1009 30.0702
R10847 VDD.n1129 VDD.n1127 30.0702
R10848 VDD.n564 VDD.n563 30.0702
R10849 VDD.n683 VDD.n681 30.0702
R10850 VDD.n10076 VDD.n10075 29.6384
R10851 VDD.n10636 VDD.n10635 29.6384
R10852 VDD.n10528 VDD.n10515 29.6384
R10853 VDD.n9606 VDD.n9605 29.6384
R10854 VDD.n10762 VDD.n10702 29.6384
R10855 VDD.n9431 VDD.n9430 29.6384
R10856 VDD.n8125 VDD.n8113 29.5303
R10857 VDD.n8187 VDD.n8125 29.5303
R10858 VDD.n8134 VDD.n8125 29.5303
R10859 VDD.n8135 VDD.n8125 29.5303
R10860 VDD.n8166 VDD.n8125 29.5303
R10861 VDD.n8152 VDD.n8125 29.5303
R10862 VDD.n12411 VDD.n6932 29.5303
R10863 VDD.n7127 VDD.n7071 29.5303
R10864 VDD.n8537 VDD.n7785 29.5303
R10865 VDD.n7786 VDD.n7785 29.5303
R10866 VDD.n8527 VDD.n7785 29.5303
R10867 VDD.n7797 VDD.n7785 29.5303
R10868 VDD.n8517 VDD.n7785 29.5303
R10869 VDD.n7803 VDD.n7785 29.5303
R10870 VDD.n7804 VDD.n7785 29.5303
R10871 VDD.n8125 VDD.n8124 29.5303
R10872 VDD.n11217 VDD.n6607 29.5303
R10873 VDD.n12694 VDD.n6618 29.5303
R10874 VDD.n12694 VDD.n6616 29.5303
R10875 VDD.n12694 VDD.n6613 29.5303
R10876 VDD.n6425 VDD.n5861 29.5303
R10877 VDD.n6487 VDD.n5827 29.5303
R10878 VDD.n5797 VDD.n5796 29.5303
R10879 VDD.n6531 VDD.n5796 29.5303
R10880 VDD.n5809 VDD.n5796 29.5303
R10881 VDD.n6520 VDD.n5796 29.5303
R10882 VDD.n6265 VDD.n5796 29.5303
R10883 VDD.n6049 VDD.n5796 29.5303
R10884 VDD.n6279 VDD.n5796 29.5303
R10885 VDD.n6221 VDD.n6072 29.5303
R10886 VDD.n6221 VDD.n6220 29.5303
R10887 VDD.n5571 VDD.n5007 29.5303
R10888 VDD.n5633 VDD.n4973 29.5303
R10889 VDD.n4943 VDD.n4942 29.5303
R10890 VDD.n5677 VDD.n4942 29.5303
R10891 VDD.n4955 VDD.n4942 29.5303
R10892 VDD.n5666 VDD.n4942 29.5303
R10893 VDD.n5411 VDD.n4942 29.5303
R10894 VDD.n5195 VDD.n4942 29.5303
R10895 VDD.n5425 VDD.n4942 29.5303
R10896 VDD.n5367 VDD.n5218 29.5303
R10897 VDD.n5367 VDD.n5366 29.5303
R10898 VDD.n4785 VDD.n4221 29.5303
R10899 VDD.n4847 VDD.n4187 29.5303
R10900 VDD.n4157 VDD.n4156 29.5303
R10901 VDD.n4891 VDD.n4156 29.5303
R10902 VDD.n4169 VDD.n4156 29.5303
R10903 VDD.n4880 VDD.n4156 29.5303
R10904 VDD.n4625 VDD.n4156 29.5303
R10905 VDD.n4409 VDD.n4156 29.5303
R10906 VDD.n4639 VDD.n4156 29.5303
R10907 VDD.n4581 VDD.n4432 29.5303
R10908 VDD.n4581 VDD.n4580 29.5303
R10909 VDD.n3931 VDD.n3367 29.5303
R10910 VDD.n3993 VDD.n3333 29.5303
R10911 VDD.n3303 VDD.n3302 29.5303
R10912 VDD.n4037 VDD.n3302 29.5303
R10913 VDD.n3315 VDD.n3302 29.5303
R10914 VDD.n4026 VDD.n3302 29.5303
R10915 VDD.n3771 VDD.n3302 29.5303
R10916 VDD.n3555 VDD.n3302 29.5303
R10917 VDD.n3785 VDD.n3302 29.5303
R10918 VDD.n3727 VDD.n3578 29.5303
R10919 VDD.n3727 VDD.n3726 29.5303
R10920 VDD.n3145 VDD.n2581 29.5303
R10921 VDD.n3207 VDD.n2547 29.5303
R10922 VDD.n2517 VDD.n2516 29.5303
R10923 VDD.n3251 VDD.n2516 29.5303
R10924 VDD.n2529 VDD.n2516 29.5303
R10925 VDD.n3240 VDD.n2516 29.5303
R10926 VDD.n2985 VDD.n2516 29.5303
R10927 VDD.n2769 VDD.n2516 29.5303
R10928 VDD.n2999 VDD.n2516 29.5303
R10929 VDD.n2941 VDD.n2792 29.5303
R10930 VDD.n2941 VDD.n2940 29.5303
R10931 VDD.n2290 VDD.n1726 29.5303
R10932 VDD.n2352 VDD.n1692 29.5303
R10933 VDD.n1662 VDD.n1661 29.5303
R10934 VDD.n2396 VDD.n1661 29.5303
R10935 VDD.n1674 VDD.n1661 29.5303
R10936 VDD.n2385 VDD.n1661 29.5303
R10937 VDD.n2130 VDD.n1661 29.5303
R10938 VDD.n1914 VDD.n1661 29.5303
R10939 VDD.n2144 VDD.n1661 29.5303
R10940 VDD.n2086 VDD.n1937 29.5303
R10941 VDD.n2086 VDD.n2085 29.5303
R10942 VDD.n1463 VDD.n1462 29.5303
R10943 VDD.n1078 VDD.n1077 29.5303
R10944 VDD.n1018 VDD.n1017 29.5303
R10945 VDD.n933 VDD.n932 29.5303
R10946 VDD.n235 VDD.n234 29.5303
R10947 VDD.n632 VDD.n631 29.5303
R10948 VDD.n572 VDD.n571 29.5303
R10949 VDD.n487 VDD.n486 29.5303
R10950 VDD.n7133 VDD.n7071 29.5301
R10951 VDD.n7142 VDD.n7071 29.5301
R10952 VDD.n7119 VDD.n7071 29.5301
R10953 VDD.n7152 VDD.n7071 29.5301
R10954 VDD.n7162 VDD.n7071 29.5301
R10955 VDD.n7164 VDD.n7071 29.5301
R10956 VDD.n7173 VDD.n7071 29.5301
R10957 VDD.n7107 VDD.n7071 29.5301
R10958 VDD.n7183 VDD.n7071 29.5301
R10959 VDD.n7192 VDD.n7071 29.5301
R10960 VDD.n7099 VDD.n7071 29.5301
R10961 VDD.n7202 VDD.n7071 29.5301
R10962 VDD.n7211 VDD.n7071 29.5301
R10963 VDD.n7212 VDD.n7071 29.5301
R10964 VDD.n7223 VDD.n7071 29.5301
R10965 VDD.n7087 VDD.n7071 29.5301
R10966 VDD.n7233 VDD.n7071 29.5301
R10967 VDD.n7242 VDD.n7071 29.5301
R10968 VDD.n7079 VDD.n7071 29.5301
R10969 VDD.n7252 VDD.n7071 29.5301
R10970 VDD.n7946 VDD.n7749 29.5301
R10971 VDD.n7840 VDD.n7749 29.5301
R10972 VDD.n7936 VDD.n7749 29.5301
R10973 VDD.n7900 VDD.n7749 29.5301
R10974 VDD.n7872 VDD.n7749 29.5301
R10975 VDD.n7890 VDD.n7749 29.5301
R10976 VDD.n7881 VDD.n7749 29.5301
R10977 VDD.n6619 VDD.n6607 29.5301
R10978 VDD.n6617 VDD.n6607 29.5301
R10979 VDD.n6615 VDD.n6607 29.5301
R10980 VDD.n6391 VDD.n5889 29.5301
R10981 VDD.n5537 VDD.n5035 29.5301
R10982 VDD.n4751 VDD.n4249 29.5301
R10983 VDD.n3897 VDD.n3395 29.5301
R10984 VDD.n3111 VDD.n2609 29.5301
R10985 VDD.n2256 VDD.n1754 29.5301
R10986 VDD.n1412 VDD.n1411 29.5301
R10987 VDD.n184 VDD.n183 29.5301
R10988 VDD.n6022 VDD.n6007 29.4877
R10989 VDD.n6293 VDD.n6045 29.4877
R10990 VDD.n5168 VDD.n5153 29.4877
R10991 VDD.n5439 VDD.n5191 29.4877
R10992 VDD.n4382 VDD.n4367 29.4877
R10993 VDD.n4653 VDD.n4405 29.4877
R10994 VDD.n3528 VDD.n3513 29.4877
R10995 VDD.n3799 VDD.n3551 29.4877
R10996 VDD.n2742 VDD.n2727 29.4877
R10997 VDD.n3013 VDD.n2765 29.4877
R10998 VDD.n1887 VDD.n1872 29.4877
R10999 VDD.n2158 VDD.n1910 29.4877
R11000 VDD.n9180 VDD.n9179 29.4133
R11001 VDD.n9179 VDD.n8734 29.4133
R11002 VDD.t105 VDD.n5930 28.8467
R11003 VDD.n6337 VDD.t100 28.8467
R11004 VDD.n6325 VDD.t174 28.8467
R11005 VDD.t103 VDD.n5076 28.8467
R11006 VDD.n5483 VDD.t146 28.8467
R11007 VDD.n5471 VDD.t158 28.8467
R11008 VDD.t122 VDD.n4290 28.8467
R11009 VDD.n4697 VDD.t186 28.8467
R11010 VDD.n4685 VDD.t180 28.8467
R11011 VDD.t120 VDD.n3436 28.8467
R11012 VDD.n3843 VDD.t125 28.8467
R11013 VDD.n3831 VDD.t7 28.8467
R11014 VDD.t98 VDD.n2650 28.8467
R11015 VDD.n3057 VDD.t82 28.8467
R11016 VDD.n3045 VDD.t177 28.8467
R11017 VDD.t94 VDD.n1795 28.8467
R11018 VDD.n2202 VDD.t20 28.8467
R11019 VDD.n2190 VDD.t101 28.8467
R11020 VDD.n5764 VDD.t187 28.1564
R11021 VDD.n4124 VDD.t73 28.1564
R11022 VDD.n2484 VDD.t164 28.1564
R11023 VDD.n844 VDD.t204 28.1564
R11024 VDD.n6222 VDD.n6071 28.0793
R11025 VDD.n5368 VDD.n5217 28.0793
R11026 VDD.n4582 VDD.n4431 28.0793
R11027 VDD.n3728 VDD.n3577 28.0793
R11028 VDD.n2942 VDD.n2791 28.0793
R11029 VDD.n2087 VDD.n1936 28.0793
R11030 VDD.n880 VDD.n879 28.0793
R11031 VDD.n434 VDD.n433 28.0793
R11032 VDD.n6010 VDD.t108 27.6955
R11033 VDD.n6010 VDD.t106 27.6955
R11034 VDD.n6014 VDD.t70 27.6955
R11035 VDD.n6014 VDD.t175 27.6955
R11036 VDD.n5156 VDD.t107 27.6955
R11037 VDD.n5156 VDD.t104 27.6955
R11038 VDD.n5160 VDD.t197 27.6955
R11039 VDD.n5160 VDD.t159 27.6955
R11040 VDD.n4370 VDD.t119 27.6955
R11041 VDD.n4370 VDD.t123 27.6955
R11042 VDD.n4374 VDD.t81 27.6955
R11043 VDD.n4374 VDD.t181 27.6955
R11044 VDD.n3516 VDD.t117 27.6955
R11045 VDD.n3516 VDD.t121 27.6955
R11046 VDD.n3520 VDD.t66 27.6955
R11047 VDD.n3520 VDD.t8 27.6955
R11048 VDD.n2730 VDD.t97 27.6955
R11049 VDD.n2730 VDD.t99 27.6955
R11050 VDD.n2734 VDD.t62 27.6955
R11051 VDD.n2734 VDD.t178 27.6955
R11052 VDD.n1875 VDD.t93 27.6955
R11053 VDD.n1875 VDD.t95 27.6955
R11054 VDD.n1879 VDD.t19 27.6955
R11055 VDD.n1879 VDD.t102 27.6955
R11056 VDD.n1229 VDD.t87 27.6955
R11057 VDD.n1229 VDD.t89 27.6955
R11058 VDD.n1228 VDD.t64 27.6955
R11059 VDD.n1228 VDD.t78 27.6955
R11060 VDD.n1 VDD.t91 27.6955
R11061 VDD.n1 VDD.t86 27.6955
R11062 VDD.n0 VDD.t202 27.6955
R11063 VDD.n0 VDD.t157 27.6955
R11064 VDD.n12481 VDD.n12480 27.5177
R11065 VDD.n6733 VDD.n6702 26.8524
R11066 VDD.n6726 VDD.n6702 26.8524
R11067 VDD.n6740 VDD.n6702 26.8524
R11068 VDD.n6728 VDD.n6702 26.8524
R11069 VDD.n6027 VDD.n5940 26.8524
R11070 VDD.n6031 VDD.n5940 26.8524
R11071 VDD.n6038 VDD.n5940 26.8524
R11072 VDD.n6381 VDD.n6380 26.8524
R11073 VDD.n6544 VDD.n5792 26.8524
R11074 VDD.n5807 VDD.n5801 26.8524
R11075 VDD.n6526 VDD.n5807 26.8524
R11076 VDD.n5807 VDD.n5800 26.8524
R11077 VDD.n5173 VDD.n5086 26.8524
R11078 VDD.n5177 VDD.n5086 26.8524
R11079 VDD.n5184 VDD.n5086 26.8524
R11080 VDD.n5527 VDD.n5526 26.8524
R11081 VDD.n5690 VDD.n4938 26.8524
R11082 VDD.n4953 VDD.n4947 26.8524
R11083 VDD.n5672 VDD.n4953 26.8524
R11084 VDD.n4953 VDD.n4946 26.8524
R11085 VDD.n4387 VDD.n4300 26.8524
R11086 VDD.n4391 VDD.n4300 26.8524
R11087 VDD.n4398 VDD.n4300 26.8524
R11088 VDD.n4741 VDD.n4740 26.8524
R11089 VDD.n4904 VDD.n4152 26.8524
R11090 VDD.n4167 VDD.n4161 26.8524
R11091 VDD.n4886 VDD.n4167 26.8524
R11092 VDD.n4167 VDD.n4160 26.8524
R11093 VDD.n3533 VDD.n3446 26.8524
R11094 VDD.n3537 VDD.n3446 26.8524
R11095 VDD.n3544 VDD.n3446 26.8524
R11096 VDD.n3887 VDD.n3886 26.8524
R11097 VDD.n4050 VDD.n3298 26.8524
R11098 VDD.n3313 VDD.n3307 26.8524
R11099 VDD.n4032 VDD.n3313 26.8524
R11100 VDD.n3313 VDD.n3306 26.8524
R11101 VDD.n2747 VDD.n2660 26.8524
R11102 VDD.n2751 VDD.n2660 26.8524
R11103 VDD.n2758 VDD.n2660 26.8524
R11104 VDD.n3101 VDD.n3100 26.8524
R11105 VDD.n3264 VDD.n2512 26.8524
R11106 VDD.n2527 VDD.n2521 26.8524
R11107 VDD.n3246 VDD.n2527 26.8524
R11108 VDD.n2527 VDD.n2520 26.8524
R11109 VDD.n1892 VDD.n1805 26.8524
R11110 VDD.n1896 VDD.n1805 26.8524
R11111 VDD.n1903 VDD.n1805 26.8524
R11112 VDD.n2246 VDD.n2245 26.8524
R11113 VDD.n2409 VDD.n1657 26.8524
R11114 VDD.n1672 VDD.n1666 26.8524
R11115 VDD.n2391 VDD.n1672 26.8524
R11116 VDD.n1672 VDD.n1665 26.8524
R11117 VDD.n1240 VDD.n1239 26.8524
R11118 VDD.n1239 VDD.n1238 26.8524
R11119 VDD.n1197 VDD.n1194 26.8524
R11120 VDD.n1182 VDD.n1181 26.8524
R11121 VDD.n12 VDD.n11 26.8524
R11122 VDD.n11 VDD.n10 26.8524
R11123 VDD.n751 VDD.n748 26.8524
R11124 VDD.n736 VDD.n735 26.8524
R11125 VDD.n6380 VDD.n6379 26.8521
R11126 VDD.n6380 VDD.n5909 26.8521
R11127 VDD.n6380 VDD.n5906 26.8521
R11128 VDD.n6380 VDD.n5907 26.8521
R11129 VDD.n6380 VDD.n5908 26.8521
R11130 VDD.n5526 VDD.n5525 26.8521
R11131 VDD.n5526 VDD.n5055 26.8521
R11132 VDD.n5526 VDD.n5052 26.8521
R11133 VDD.n5526 VDD.n5053 26.8521
R11134 VDD.n5526 VDD.n5054 26.8521
R11135 VDD.n4740 VDD.n4739 26.8521
R11136 VDD.n4740 VDD.n4269 26.8521
R11137 VDD.n4740 VDD.n4266 26.8521
R11138 VDD.n4740 VDD.n4267 26.8521
R11139 VDD.n4740 VDD.n4268 26.8521
R11140 VDD.n3886 VDD.n3885 26.8521
R11141 VDD.n3886 VDD.n3415 26.8521
R11142 VDD.n3886 VDD.n3412 26.8521
R11143 VDD.n3886 VDD.n3413 26.8521
R11144 VDD.n3886 VDD.n3414 26.8521
R11145 VDD.n3100 VDD.n3099 26.8521
R11146 VDD.n3100 VDD.n2629 26.8521
R11147 VDD.n3100 VDD.n2626 26.8521
R11148 VDD.n3100 VDD.n2627 26.8521
R11149 VDD.n3100 VDD.n2628 26.8521
R11150 VDD.n2245 VDD.n2244 26.8521
R11151 VDD.n2245 VDD.n1774 26.8521
R11152 VDD.n2245 VDD.n1771 26.8521
R11153 VDD.n2245 VDD.n1772 26.8521
R11154 VDD.n2245 VDD.n1773 26.8521
R11155 VDD.n1403 VDD.n1402 26.8521
R11156 VDD.n175 VDD.n174 26.8521
R11157 VDD.n10478 VDD.n6914 26.6499
R11158 VDD.n10448 VDD.n6914 26.6499
R11159 VDD.n10448 VDD.n6922 26.6499
R11160 VDD.n10481 VDD.n6922 26.6499
R11161 VDD.n10493 VDD.n10433 26.6499
R11162 VDD.n10422 VDD.n10421 26.6499
R11163 VDD.n10495 VDD.n10163 26.6499
R11164 VDD.n11025 VDD.n8733 26.6499
R11165 VDD.n8733 VDD.n8728 26.6499
R11166 VDD.n10995 VDD.n8728 26.6499
R11167 VDD.n10995 VDD.n8731 26.6499
R11168 VDD.n10988 VDD.n10986 26.6499
R11169 VDD.n10986 VDD.n8730 26.6499
R11170 VDD.n10998 VDD.n8729 26.6499
R11171 VDD.n9182 VDD.n9175 26.6499
R11172 VDD.n9184 VDD.n9171 26.6499
R11173 VDD.n9209 VDD.n9200 26.6499
R11174 VDD.n9217 VDD.n9200 26.6499
R11175 VDD.n9217 VDD.n9206 26.6499
R11176 VDD.n9218 VDD.n9206 26.6499
R11177 VDD.n10950 VDD.n9222 26.6499
R11178 VDD.n10958 VDD.n9223 26.6499
R11179 VDD.n9980 VDD.n9979 26.3534
R11180 VDD.n6029 VDD.n5935 26.3534
R11181 VDD.n5175 VDD.n5081 26.3534
R11182 VDD.n4389 VDD.n4295 26.3534
R11183 VDD.n3535 VDD.n3441 26.3534
R11184 VDD.n2749 VDD.n2655 26.3534
R11185 VDD.n1894 VDD.n1800 26.3534
R11186 VDD.n1605 VDD.n1243 26.3534
R11187 VDD.n377 VDD.n15 26.3534
R11188 VDD.n10075 VDD.n10025 26.3453
R11189 VDD.n10635 VDD.n10144 26.3453
R11190 VDD.n10520 VDD.n10515 26.3453
R11191 VDD.n9605 VDD.n9604 26.3453
R11192 VDD.n10717 VDD.n10702 26.3453
R11193 VDD.n9432 VDD.n9431 26.3453
R11194 VDD.n9651 VDD.n9650 26.3366
R11195 VDD.n9666 VDD.n9663 26.3366
R11196 VDD.n10794 VDD.n10793 26.3366
R11197 VDD.n10809 VDD.n10806 26.3366
R11198 VDD.n8870 VDD.n8869 26.3366
R11199 VDD.n8963 VDD.n8962 26.3366
R11200 VDD.n8966 VDD.n8963 26.3366
R11201 VDD.n9005 VDD.n9002 26.3366
R11202 VDD.n8989 VDD.n8985 26.3366
R11203 VDD.n8989 VDD.n8988 26.3366
R11204 VDD.n9280 VDD.n9277 26.3366
R11205 VDD.n9410 VDD.n9407 26.3366
R11206 VDD.n9977 VDD.n9976 25.9875
R11207 VDD.n6106 VDD.n6101 25.7394
R11208 VDD.n5252 VDD.n5247 25.7394
R11209 VDD.n4466 VDD.n4461 25.7394
R11210 VDD.n3612 VDD.n3607 25.7394
R11211 VDD.n2826 VDD.n2821 25.7394
R11212 VDD.n1971 VDD.n1966 25.7394
R11213 VDD.n1306 VDD.n1305 25.7394
R11214 VDD.n78 VDD.n77 25.7394
R11215 VDD.n8572 VDD.n8571 25.6005
R11216 VDD.n8575 VDD.n8572 25.6005
R11217 VDD.n8576 VDD.n8575 25.6005
R11218 VDD.n8579 VDD.n8576 25.6005
R11219 VDD.n8580 VDD.n8579 25.6005
R11220 VDD.n8583 VDD.n8580 25.6005
R11221 VDD.n8585 VDD.n8583 25.6005
R11222 VDD.n8586 VDD.n8585 25.6005
R11223 VDD.n8587 VDD.n8586 25.6005
R11224 VDD.n8587 VDD.n7752 25.6005
R11225 VDD.n8593 VDD.n7752 25.6005
R11226 VDD.n8594 VDD.n8593 25.6005
R11227 VDD.n8596 VDD.n8594 25.6005
R11228 VDD.n8596 VDD.n8595 25.6005
R11229 VDD.n8595 VDD.n7732 25.6005
R11230 VDD.n11439 VDD.n7732 25.6005
R11231 VDD.n11439 VDD.n11438 25.6005
R11232 VDD.n11438 VDD.n11437 25.6005
R11233 VDD.n11437 VDD.n7733 25.6005
R11234 VDD.n8625 VDD.n7733 25.6005
R11235 VDD.n11420 VDD.n8625 25.6005
R11236 VDD.n11420 VDD.n11419 25.6005
R11237 VDD.n11419 VDD.n11418 25.6005
R11238 VDD.n11418 VDD.n8626 25.6005
R11239 VDD.n8656 VDD.n8626 25.6005
R11240 VDD.n11401 VDD.n8656 25.6005
R11241 VDD.n11401 VDD.n11400 25.6005
R11242 VDD.n11400 VDD.n11399 25.6005
R11243 VDD.n11399 VDD.n8657 25.6005
R11244 VDD.n8694 VDD.n8657 25.6005
R11245 VDD.n8696 VDD.n8694 25.6005
R11246 VDD.n8697 VDD.n8696 25.6005
R11247 VDD.n11376 VDD.n8697 25.6005
R11248 VDD.n11376 VDD.n11375 25.6005
R11249 VDD.n11375 VDD.n11374 25.6005
R11250 VDD.n11374 VDD.n8698 25.6005
R11251 VDD.n11030 VDD.n8698 25.6005
R11252 VDD.n11357 VDD.n11030 25.6005
R11253 VDD.n11357 VDD.n11356 25.6005
R11254 VDD.n11356 VDD.n11355 25.6005
R11255 VDD.n11355 VDD.n11031 25.6005
R11256 VDD.n11060 VDD.n11031 25.6005
R11257 VDD.n11338 VDD.n11060 25.6005
R11258 VDD.n11338 VDD.n11337 25.6005
R11259 VDD.n11337 VDD.n11336 25.6005
R11260 VDD.n11336 VDD.n11061 25.6005
R11261 VDD.n11323 VDD.n11061 25.6005
R11262 VDD.n11323 VDD.n11322 25.6005
R11263 VDD.n11322 VDD.n11321 25.6005
R11264 VDD.n11321 VDD.n11078 25.6005
R11265 VDD.n11114 VDD.n11078 25.6005
R11266 VDD.n11304 VDD.n11114 25.6005
R11267 VDD.n11304 VDD.n11303 25.6005
R11268 VDD.n11303 VDD.n11302 25.6005
R11269 VDD.n11302 VDD.n11115 25.6005
R11270 VDD.n11145 VDD.n11115 25.6005
R11271 VDD.n11285 VDD.n11145 25.6005
R11272 VDD.n11285 VDD.n11284 25.6005
R11273 VDD.n11284 VDD.n11283 25.6005
R11274 VDD.n11283 VDD.n11146 25.6005
R11275 VDD.n11176 VDD.n11146 25.6005
R11276 VDD.n11266 VDD.n11176 25.6005
R11277 VDD.n11266 VDD.n11265 25.6005
R11278 VDD.n11265 VDD.n11264 25.6005
R11279 VDD.n11264 VDD.n11177 25.6005
R11280 VDD.n11235 VDD.n11177 25.6005
R11281 VDD.n11237 VDD.n11235 25.6005
R11282 VDD.n11238 VDD.n11237 25.6005
R11283 VDD.n11241 VDD.n11238 25.6005
R11284 VDD.n11241 VDD.n11240 25.6005
R11285 VDD.n11240 VDD.n11239 25.6005
R11286 VDD.n11239 VDD.n6598 25.6005
R11287 VDD.n12678 VDD.n12677 25.6005
R11288 VDD.n12677 VDD.n12676 25.6005
R11289 VDD.n12676 VDD.n6718 25.6005
R11290 VDD.n12666 VDD.n6718 25.6005
R11291 VDD.n12666 VDD.n12665 25.6005
R11292 VDD.n12665 VDD.n12664 25.6005
R11293 VDD.n12664 VDD.n6751 25.6005
R11294 VDD.n12654 VDD.n6751 25.6005
R11295 VDD.n12654 VDD.n12653 25.6005
R11296 VDD.n12653 VDD.n12652 25.6005
R11297 VDD.n12652 VDD.n6761 25.6005
R11298 VDD.n12642 VDD.n6761 25.6005
R11299 VDD.n12642 VDD.n12641 25.6005
R11300 VDD.n12641 VDD.n12640 25.6005
R11301 VDD.n12640 VDD.n6773 25.6005
R11302 VDD.n12630 VDD.n6773 25.6005
R11303 VDD.n12630 VDD.n12629 25.6005
R11304 VDD.n12629 VDD.n12628 25.6005
R11305 VDD.n12628 VDD.n6785 25.6005
R11306 VDD.n12618 VDD.n6785 25.6005
R11307 VDD.n12618 VDD.n12617 25.6005
R11308 VDD.n12617 VDD.n12616 25.6005
R11309 VDD.n12616 VDD.n6795 25.6005
R11310 VDD.n12606 VDD.n6795 25.6005
R11311 VDD.n12606 VDD.n12605 25.6005
R11312 VDD.n12605 VDD.n12604 25.6005
R11313 VDD.n12604 VDD.n6807 25.6005
R11314 VDD.n12594 VDD.n6807 25.6005
R11315 VDD.n12594 VDD.n12593 25.6005
R11316 VDD.n12593 VDD.n12592 25.6005
R11317 VDD.n12592 VDD.n6818 25.6005
R11318 VDD.n12582 VDD.n6818 25.6005
R11319 VDD.n12582 VDD.n12581 25.6005
R11320 VDD.n12581 VDD.n12580 25.6005
R11321 VDD.n12580 VDD.n6827 25.6005
R11322 VDD.n12570 VDD.n6827 25.6005
R11323 VDD.n12570 VDD.n12569 25.6005
R11324 VDD.n12569 VDD.n12568 25.6005
R11325 VDD.n12568 VDD.n6839 25.6005
R11326 VDD.n12558 VDD.n6839 25.6005
R11327 VDD.n12558 VDD.n12557 25.6005
R11328 VDD.n12557 VDD.n12556 25.6005
R11329 VDD.n12556 VDD.n6851 25.6005
R11330 VDD.n12546 VDD.n6851 25.6005
R11331 VDD.n12546 VDD.n12545 25.6005
R11332 VDD.n12545 VDD.n12544 25.6005
R11333 VDD.n12544 VDD.n6861 25.6005
R11334 VDD.n12534 VDD.n6861 25.6005
R11335 VDD.n12534 VDD.n12533 25.6005
R11336 VDD.n12533 VDD.n12532 25.6005
R11337 VDD.n12532 VDD.n6872 25.6005
R11338 VDD.n12522 VDD.n6872 25.6005
R11339 VDD.n12522 VDD.n12521 25.6005
R11340 VDD.n12521 VDD.n12520 25.6005
R11341 VDD.n12520 VDD.n6883 25.6005
R11342 VDD.n12510 VDD.n6883 25.6005
R11343 VDD.n12510 VDD.n12509 25.6005
R11344 VDD.n12509 VDD.n12508 25.6005
R11345 VDD.n12508 VDD.n6895 25.6005
R11346 VDD.n12498 VDD.n6895 25.6005
R11347 VDD.n12498 VDD.n12497 25.6005
R11348 VDD.n6730 VDD.n6717 25.6005
R11349 VDD.n6731 VDD.n6730 25.6005
R11350 VDD.n6731 VDD.n6727 25.6005
R11351 VDD.n6736 VDD.n6727 25.6005
R11352 VDD.n6737 VDD.n6736 25.6005
R11353 VDD.n6737 VDD.n6725 25.6005
R11354 VDD.n6742 VDD.n6725 25.6005
R11355 VDD.n6744 VDD.n6743 25.6005
R11356 VDD.n12672 VDD.n6744 25.6005
R11357 VDD.n12672 VDD.n12671 25.6005
R11358 VDD.n12671 VDD.n12670 25.6005
R11359 VDD.n12670 VDD.n6745 25.6005
R11360 VDD.n12660 VDD.n6745 25.6005
R11361 VDD.n12660 VDD.n12659 25.6005
R11362 VDD.n12659 VDD.n12658 25.6005
R11363 VDD.n12658 VDD.n6756 25.6005
R11364 VDD.n12648 VDD.n6756 25.6005
R11365 VDD.n12648 VDD.n12647 25.6005
R11366 VDD.n12647 VDD.n12646 25.6005
R11367 VDD.n12646 VDD.n6767 25.6005
R11368 VDD.n12636 VDD.n6767 25.6005
R11369 VDD.n12636 VDD.n12635 25.6005
R11370 VDD.n12635 VDD.n12634 25.6005
R11371 VDD.n12634 VDD.n6779 25.6005
R11372 VDD.n12624 VDD.n6779 25.6005
R11373 VDD.n12624 VDD.n12623 25.6005
R11374 VDD.n12623 VDD.n12622 25.6005
R11375 VDD.n12622 VDD.n6791 25.6005
R11376 VDD.n12612 VDD.n6791 25.6005
R11377 VDD.n12612 VDD.n12611 25.6005
R11378 VDD.n12611 VDD.n12610 25.6005
R11379 VDD.n12610 VDD.n6801 25.6005
R11380 VDD.n12600 VDD.n6801 25.6005
R11381 VDD.n12600 VDD.n12599 25.6005
R11382 VDD.n12599 VDD.n12598 25.6005
R11383 VDD.n12598 VDD.n6813 25.6005
R11384 VDD.n12588 VDD.n6813 25.6005
R11385 VDD.n12588 VDD.n12587 25.6005
R11386 VDD.n12587 VDD.n12586 25.6005
R11387 VDD.n12586 VDD.n6822 25.6005
R11388 VDD.n12576 VDD.n6822 25.6005
R11389 VDD.n12576 VDD.n12575 25.6005
R11390 VDD.n12575 VDD.n12574 25.6005
R11391 VDD.n12574 VDD.n6833 25.6005
R11392 VDD.n12564 VDD.n6833 25.6005
R11393 VDD.n12564 VDD.n12563 25.6005
R11394 VDD.n12563 VDD.n12562 25.6005
R11395 VDD.n12562 VDD.n6845 25.6005
R11396 VDD.n12552 VDD.n6845 25.6005
R11397 VDD.n12552 VDD.n12551 25.6005
R11398 VDD.n12551 VDD.n12550 25.6005
R11399 VDD.n12550 VDD.n6855 25.6005
R11400 VDD.n12540 VDD.n6855 25.6005
R11401 VDD.n12540 VDD.n12539 25.6005
R11402 VDD.n12539 VDD.n12538 25.6005
R11403 VDD.n12538 VDD.n6867 25.6005
R11404 VDD.n12528 VDD.n6867 25.6005
R11405 VDD.n12528 VDD.n12527 25.6005
R11406 VDD.n12527 VDD.n12526 25.6005
R11407 VDD.n12526 VDD.n6877 25.6005
R11408 VDD.n12516 VDD.n6877 25.6005
R11409 VDD.n12516 VDD.n12515 25.6005
R11410 VDD.n12515 VDD.n12514 25.6005
R11411 VDD.n12514 VDD.n6889 25.6005
R11412 VDD.n12504 VDD.n6889 25.6005
R11413 VDD.n12504 VDD.n12503 25.6005
R11414 VDD.n12503 VDD.n12502 25.6005
R11415 VDD.n12502 VDD.n6901 25.6005
R11416 VDD.n6040 VDD.n6025 25.6005
R11417 VDD.n6035 VDD.n6025 25.6005
R11418 VDD.n6035 VDD.n6034 25.6005
R11419 VDD.n6034 VDD.n6028 25.6005
R11420 VDD.n6029 VDD.n6028 25.6005
R11421 VDD.n6492 VDD.n6491 25.6005
R11422 VDD.n6491 VDD.n5824 25.6005
R11423 VDD.n5830 VDD.n5824 25.6005
R11424 VDD.n6485 VDD.n5830 25.6005
R11425 VDD.n6429 VDD.n6428 25.6005
R11426 VDD.n6429 VDD.n5855 25.6005
R11427 VDD.n6435 VDD.n5855 25.6005
R11428 VDD.n6436 VDD.n6435 25.6005
R11429 VDD.n6437 VDD.n6436 25.6005
R11430 VDD.n6437 VDD.n5851 25.6005
R11431 VDD.n6443 VDD.n5851 25.6005
R11432 VDD.n6444 VDD.n6443 25.6005
R11433 VDD.n6445 VDD.n6444 25.6005
R11434 VDD.n6445 VDD.n5847 25.6005
R11435 VDD.n6451 VDD.n5847 25.6005
R11436 VDD.n6452 VDD.n6451 25.6005
R11437 VDD.n6453 VDD.n6452 25.6005
R11438 VDD.n6453 VDD.n5843 25.6005
R11439 VDD.n6459 VDD.n5843 25.6005
R11440 VDD.n6460 VDD.n6459 25.6005
R11441 VDD.n6461 VDD.n6460 25.6005
R11442 VDD.n6461 VDD.n5839 25.6005
R11443 VDD.n6467 VDD.n5839 25.6005
R11444 VDD.n6468 VDD.n6467 25.6005
R11445 VDD.n6469 VDD.n6468 25.6005
R11446 VDD.n6469 VDD.n5835 25.6005
R11447 VDD.n6475 VDD.n5835 25.6005
R11448 VDD.n6476 VDD.n6475 25.6005
R11449 VDD.n6477 VDD.n6476 25.6005
R11450 VDD.n6477 VDD.n5831 25.6005
R11451 VDD.n6483 VDD.n5831 25.6005
R11452 VDD.n6484 VDD.n6483 25.6005
R11453 VDD.n6421 VDD.n6419 25.6005
R11454 VDD.n6421 VDD.n6420 25.6005
R11455 VDD.n6420 VDD.n5859 25.6005
R11456 VDD.n6427 VDD.n5859 25.6005
R11457 VDD.n6320 VDD.n6302 25.6005
R11458 VDD.n6314 VDD.n6302 25.6005
R11459 VDD.n6314 VDD.n6313 25.6005
R11460 VDD.n6313 VDD.n6311 25.6005
R11461 VDD.n6311 VDD.n6309 25.6005
R11462 VDD.n5989 VDD.n5934 25.6005
R11463 VDD.n5995 VDD.n5989 25.6005
R11464 VDD.n5996 VDD.n5995 25.6005
R11465 VDD.n5996 VDD.n5987 25.6005
R11466 VDD.n6002 VDD.n5987 25.6005
R11467 VDD.n5186 VDD.n5171 25.6005
R11468 VDD.n5181 VDD.n5171 25.6005
R11469 VDD.n5181 VDD.n5180 25.6005
R11470 VDD.n5180 VDD.n5174 25.6005
R11471 VDD.n5175 VDD.n5174 25.6005
R11472 VDD.n5638 VDD.n5637 25.6005
R11473 VDD.n5637 VDD.n4970 25.6005
R11474 VDD.n4976 VDD.n4970 25.6005
R11475 VDD.n5631 VDD.n4976 25.6005
R11476 VDD.n5575 VDD.n5574 25.6005
R11477 VDD.n5575 VDD.n5001 25.6005
R11478 VDD.n5581 VDD.n5001 25.6005
R11479 VDD.n5582 VDD.n5581 25.6005
R11480 VDD.n5583 VDD.n5582 25.6005
R11481 VDD.n5583 VDD.n4997 25.6005
R11482 VDD.n5589 VDD.n4997 25.6005
R11483 VDD.n5590 VDD.n5589 25.6005
R11484 VDD.n5591 VDD.n5590 25.6005
R11485 VDD.n5591 VDD.n4993 25.6005
R11486 VDD.n5597 VDD.n4993 25.6005
R11487 VDD.n5598 VDD.n5597 25.6005
R11488 VDD.n5599 VDD.n5598 25.6005
R11489 VDD.n5599 VDD.n4989 25.6005
R11490 VDD.n5605 VDD.n4989 25.6005
R11491 VDD.n5606 VDD.n5605 25.6005
R11492 VDD.n5607 VDD.n5606 25.6005
R11493 VDD.n5607 VDD.n4985 25.6005
R11494 VDD.n5613 VDD.n4985 25.6005
R11495 VDD.n5614 VDD.n5613 25.6005
R11496 VDD.n5615 VDD.n5614 25.6005
R11497 VDD.n5615 VDD.n4981 25.6005
R11498 VDD.n5621 VDD.n4981 25.6005
R11499 VDD.n5622 VDD.n5621 25.6005
R11500 VDD.n5623 VDD.n5622 25.6005
R11501 VDD.n5623 VDD.n4977 25.6005
R11502 VDD.n5629 VDD.n4977 25.6005
R11503 VDD.n5630 VDD.n5629 25.6005
R11504 VDD.n5567 VDD.n5565 25.6005
R11505 VDD.n5567 VDD.n5566 25.6005
R11506 VDD.n5566 VDD.n5005 25.6005
R11507 VDD.n5573 VDD.n5005 25.6005
R11508 VDD.n5466 VDD.n5448 25.6005
R11509 VDD.n5460 VDD.n5448 25.6005
R11510 VDD.n5460 VDD.n5459 25.6005
R11511 VDD.n5459 VDD.n5457 25.6005
R11512 VDD.n5457 VDD.n5455 25.6005
R11513 VDD.n5135 VDD.n5080 25.6005
R11514 VDD.n5141 VDD.n5135 25.6005
R11515 VDD.n5142 VDD.n5141 25.6005
R11516 VDD.n5142 VDD.n5133 25.6005
R11517 VDD.n5148 VDD.n5133 25.6005
R11518 VDD.n4400 VDD.n4385 25.6005
R11519 VDD.n4395 VDD.n4385 25.6005
R11520 VDD.n4395 VDD.n4394 25.6005
R11521 VDD.n4394 VDD.n4388 25.6005
R11522 VDD.n4389 VDD.n4388 25.6005
R11523 VDD.n4852 VDD.n4851 25.6005
R11524 VDD.n4851 VDD.n4184 25.6005
R11525 VDD.n4190 VDD.n4184 25.6005
R11526 VDD.n4845 VDD.n4190 25.6005
R11527 VDD.n4789 VDD.n4788 25.6005
R11528 VDD.n4789 VDD.n4215 25.6005
R11529 VDD.n4795 VDD.n4215 25.6005
R11530 VDD.n4796 VDD.n4795 25.6005
R11531 VDD.n4797 VDD.n4796 25.6005
R11532 VDD.n4797 VDD.n4211 25.6005
R11533 VDD.n4803 VDD.n4211 25.6005
R11534 VDD.n4804 VDD.n4803 25.6005
R11535 VDD.n4805 VDD.n4804 25.6005
R11536 VDD.n4805 VDD.n4207 25.6005
R11537 VDD.n4811 VDD.n4207 25.6005
R11538 VDD.n4812 VDD.n4811 25.6005
R11539 VDD.n4813 VDD.n4812 25.6005
R11540 VDD.n4813 VDD.n4203 25.6005
R11541 VDD.n4819 VDD.n4203 25.6005
R11542 VDD.n4820 VDD.n4819 25.6005
R11543 VDD.n4821 VDD.n4820 25.6005
R11544 VDD.n4821 VDD.n4199 25.6005
R11545 VDD.n4827 VDD.n4199 25.6005
R11546 VDD.n4828 VDD.n4827 25.6005
R11547 VDD.n4829 VDD.n4828 25.6005
R11548 VDD.n4829 VDD.n4195 25.6005
R11549 VDD.n4835 VDD.n4195 25.6005
R11550 VDD.n4836 VDD.n4835 25.6005
R11551 VDD.n4837 VDD.n4836 25.6005
R11552 VDD.n4837 VDD.n4191 25.6005
R11553 VDD.n4843 VDD.n4191 25.6005
R11554 VDD.n4844 VDD.n4843 25.6005
R11555 VDD.n4781 VDD.n4779 25.6005
R11556 VDD.n4781 VDD.n4780 25.6005
R11557 VDD.n4780 VDD.n4219 25.6005
R11558 VDD.n4787 VDD.n4219 25.6005
R11559 VDD.n4680 VDD.n4662 25.6005
R11560 VDD.n4674 VDD.n4662 25.6005
R11561 VDD.n4674 VDD.n4673 25.6005
R11562 VDD.n4673 VDD.n4671 25.6005
R11563 VDD.n4671 VDD.n4669 25.6005
R11564 VDD.n4349 VDD.n4294 25.6005
R11565 VDD.n4355 VDD.n4349 25.6005
R11566 VDD.n4356 VDD.n4355 25.6005
R11567 VDD.n4356 VDD.n4347 25.6005
R11568 VDD.n4362 VDD.n4347 25.6005
R11569 VDD.n3546 VDD.n3531 25.6005
R11570 VDD.n3541 VDD.n3531 25.6005
R11571 VDD.n3541 VDD.n3540 25.6005
R11572 VDD.n3540 VDD.n3534 25.6005
R11573 VDD.n3535 VDD.n3534 25.6005
R11574 VDD.n3998 VDD.n3997 25.6005
R11575 VDD.n3997 VDD.n3330 25.6005
R11576 VDD.n3336 VDD.n3330 25.6005
R11577 VDD.n3991 VDD.n3336 25.6005
R11578 VDD.n3935 VDD.n3934 25.6005
R11579 VDD.n3935 VDD.n3361 25.6005
R11580 VDD.n3941 VDD.n3361 25.6005
R11581 VDD.n3942 VDD.n3941 25.6005
R11582 VDD.n3943 VDD.n3942 25.6005
R11583 VDD.n3943 VDD.n3357 25.6005
R11584 VDD.n3949 VDD.n3357 25.6005
R11585 VDD.n3950 VDD.n3949 25.6005
R11586 VDD.n3951 VDD.n3950 25.6005
R11587 VDD.n3951 VDD.n3353 25.6005
R11588 VDD.n3957 VDD.n3353 25.6005
R11589 VDD.n3958 VDD.n3957 25.6005
R11590 VDD.n3959 VDD.n3958 25.6005
R11591 VDD.n3959 VDD.n3349 25.6005
R11592 VDD.n3965 VDD.n3349 25.6005
R11593 VDD.n3966 VDD.n3965 25.6005
R11594 VDD.n3967 VDD.n3966 25.6005
R11595 VDD.n3967 VDD.n3345 25.6005
R11596 VDD.n3973 VDD.n3345 25.6005
R11597 VDD.n3974 VDD.n3973 25.6005
R11598 VDD.n3975 VDD.n3974 25.6005
R11599 VDD.n3975 VDD.n3341 25.6005
R11600 VDD.n3981 VDD.n3341 25.6005
R11601 VDD.n3982 VDD.n3981 25.6005
R11602 VDD.n3983 VDD.n3982 25.6005
R11603 VDD.n3983 VDD.n3337 25.6005
R11604 VDD.n3989 VDD.n3337 25.6005
R11605 VDD.n3990 VDD.n3989 25.6005
R11606 VDD.n3927 VDD.n3925 25.6005
R11607 VDD.n3927 VDD.n3926 25.6005
R11608 VDD.n3926 VDD.n3365 25.6005
R11609 VDD.n3933 VDD.n3365 25.6005
R11610 VDD.n3826 VDD.n3808 25.6005
R11611 VDD.n3820 VDD.n3808 25.6005
R11612 VDD.n3820 VDD.n3819 25.6005
R11613 VDD.n3819 VDD.n3817 25.6005
R11614 VDD.n3817 VDD.n3815 25.6005
R11615 VDD.n3495 VDD.n3440 25.6005
R11616 VDD.n3501 VDD.n3495 25.6005
R11617 VDD.n3502 VDD.n3501 25.6005
R11618 VDD.n3502 VDD.n3493 25.6005
R11619 VDD.n3508 VDD.n3493 25.6005
R11620 VDD.n2760 VDD.n2745 25.6005
R11621 VDD.n2755 VDD.n2745 25.6005
R11622 VDD.n2755 VDD.n2754 25.6005
R11623 VDD.n2754 VDD.n2748 25.6005
R11624 VDD.n2749 VDD.n2748 25.6005
R11625 VDD.n3212 VDD.n3211 25.6005
R11626 VDD.n3211 VDD.n2544 25.6005
R11627 VDD.n2550 VDD.n2544 25.6005
R11628 VDD.n3205 VDD.n2550 25.6005
R11629 VDD.n3149 VDD.n3148 25.6005
R11630 VDD.n3149 VDD.n2575 25.6005
R11631 VDD.n3155 VDD.n2575 25.6005
R11632 VDD.n3156 VDD.n3155 25.6005
R11633 VDD.n3157 VDD.n3156 25.6005
R11634 VDD.n3157 VDD.n2571 25.6005
R11635 VDD.n3163 VDD.n2571 25.6005
R11636 VDD.n3164 VDD.n3163 25.6005
R11637 VDD.n3165 VDD.n3164 25.6005
R11638 VDD.n3165 VDD.n2567 25.6005
R11639 VDD.n3171 VDD.n2567 25.6005
R11640 VDD.n3172 VDD.n3171 25.6005
R11641 VDD.n3173 VDD.n3172 25.6005
R11642 VDD.n3173 VDD.n2563 25.6005
R11643 VDD.n3179 VDD.n2563 25.6005
R11644 VDD.n3180 VDD.n3179 25.6005
R11645 VDD.n3181 VDD.n3180 25.6005
R11646 VDD.n3181 VDD.n2559 25.6005
R11647 VDD.n3187 VDD.n2559 25.6005
R11648 VDD.n3188 VDD.n3187 25.6005
R11649 VDD.n3189 VDD.n3188 25.6005
R11650 VDD.n3189 VDD.n2555 25.6005
R11651 VDD.n3195 VDD.n2555 25.6005
R11652 VDD.n3196 VDD.n3195 25.6005
R11653 VDD.n3197 VDD.n3196 25.6005
R11654 VDD.n3197 VDD.n2551 25.6005
R11655 VDD.n3203 VDD.n2551 25.6005
R11656 VDD.n3204 VDD.n3203 25.6005
R11657 VDD.n3141 VDD.n3139 25.6005
R11658 VDD.n3141 VDD.n3140 25.6005
R11659 VDD.n3140 VDD.n2579 25.6005
R11660 VDD.n3147 VDD.n2579 25.6005
R11661 VDD.n3040 VDD.n3022 25.6005
R11662 VDD.n3034 VDD.n3022 25.6005
R11663 VDD.n3034 VDD.n3033 25.6005
R11664 VDD.n3033 VDD.n3031 25.6005
R11665 VDD.n3031 VDD.n3029 25.6005
R11666 VDD.n2709 VDD.n2654 25.6005
R11667 VDD.n2715 VDD.n2709 25.6005
R11668 VDD.n2716 VDD.n2715 25.6005
R11669 VDD.n2716 VDD.n2707 25.6005
R11670 VDD.n2722 VDD.n2707 25.6005
R11671 VDD.n1905 VDD.n1890 25.6005
R11672 VDD.n1900 VDD.n1890 25.6005
R11673 VDD.n1900 VDD.n1899 25.6005
R11674 VDD.n1899 VDD.n1893 25.6005
R11675 VDD.n1894 VDD.n1893 25.6005
R11676 VDD.n2357 VDD.n2356 25.6005
R11677 VDD.n2356 VDD.n1689 25.6005
R11678 VDD.n1695 VDD.n1689 25.6005
R11679 VDD.n2350 VDD.n1695 25.6005
R11680 VDD.n2294 VDD.n2293 25.6005
R11681 VDD.n2294 VDD.n1720 25.6005
R11682 VDD.n2300 VDD.n1720 25.6005
R11683 VDD.n2301 VDD.n2300 25.6005
R11684 VDD.n2302 VDD.n2301 25.6005
R11685 VDD.n2302 VDD.n1716 25.6005
R11686 VDD.n2308 VDD.n1716 25.6005
R11687 VDD.n2309 VDD.n2308 25.6005
R11688 VDD.n2310 VDD.n2309 25.6005
R11689 VDD.n2310 VDD.n1712 25.6005
R11690 VDD.n2316 VDD.n1712 25.6005
R11691 VDD.n2317 VDD.n2316 25.6005
R11692 VDD.n2318 VDD.n2317 25.6005
R11693 VDD.n2318 VDD.n1708 25.6005
R11694 VDD.n2324 VDD.n1708 25.6005
R11695 VDD.n2325 VDD.n2324 25.6005
R11696 VDD.n2326 VDD.n2325 25.6005
R11697 VDD.n2326 VDD.n1704 25.6005
R11698 VDD.n2332 VDD.n1704 25.6005
R11699 VDD.n2333 VDD.n2332 25.6005
R11700 VDD.n2334 VDD.n2333 25.6005
R11701 VDD.n2334 VDD.n1700 25.6005
R11702 VDD.n2340 VDD.n1700 25.6005
R11703 VDD.n2341 VDD.n2340 25.6005
R11704 VDD.n2342 VDD.n2341 25.6005
R11705 VDD.n2342 VDD.n1696 25.6005
R11706 VDD.n2348 VDD.n1696 25.6005
R11707 VDD.n2349 VDD.n2348 25.6005
R11708 VDD.n2286 VDD.n2284 25.6005
R11709 VDD.n2286 VDD.n2285 25.6005
R11710 VDD.n2285 VDD.n1724 25.6005
R11711 VDD.n2292 VDD.n1724 25.6005
R11712 VDD.n2185 VDD.n2167 25.6005
R11713 VDD.n2179 VDD.n2167 25.6005
R11714 VDD.n2179 VDD.n2178 25.6005
R11715 VDD.n2178 VDD.n2176 25.6005
R11716 VDD.n2176 VDD.n2174 25.6005
R11717 VDD.n1854 VDD.n1799 25.6005
R11718 VDD.n1860 VDD.n1854 25.6005
R11719 VDD.n1861 VDD.n1860 25.6005
R11720 VDD.n1861 VDD.n1852 25.6005
R11721 VDD.n1867 VDD.n1852 25.6005
R11722 VDD.n861 VDD.n858 25.6005
R11723 VDD.n1235 VDD.n1232 25.6005
R11724 VDD.n1237 VDD.n1235 25.6005
R11725 VDD.n1243 VDD.n1237 25.6005
R11726 VDD.n1086 VDD.n1083 25.6005
R11727 VDD.n1083 VDD.n1080 25.6005
R11728 VDD.n1080 VDD.n1076 25.6005
R11729 VDD.n1076 VDD.n1074 25.6005
R11730 VDD.n1457 VDD.n1453 25.6005
R11731 VDD.n1453 VDD.n1450 25.6005
R11732 VDD.n1450 VDD.n1447 25.6005
R11733 VDD.n1447 VDD.n1444 25.6005
R11734 VDD.n1444 VDD.n1441 25.6005
R11735 VDD.n1441 VDD.n1438 25.6005
R11736 VDD.n1438 VDD.n1435 25.6005
R11737 VDD.n1435 VDD.n1432 25.6005
R11738 VDD.n1432 VDD.n1429 25.6005
R11739 VDD.n1429 VDD.n1426 25.6005
R11740 VDD.n1426 VDD.n1423 25.6005
R11741 VDD.n1423 VDD.n1420 25.6005
R11742 VDD.n1420 VDD.n1417 25.6005
R11743 VDD.n1032 VDD.n1029 25.6005
R11744 VDD.n1035 VDD.n1032 25.6005
R11745 VDD.n1038 VDD.n1035 25.6005
R11746 VDD.n1041 VDD.n1038 25.6005
R11747 VDD.n1044 VDD.n1041 25.6005
R11748 VDD.n1047 VDD.n1044 25.6005
R11749 VDD.n1050 VDD.n1047 25.6005
R11750 VDD.n1053 VDD.n1050 25.6005
R11751 VDD.n1056 VDD.n1053 25.6005
R11752 VDD.n1059 VDD.n1056 25.6005
R11753 VDD.n1062 VDD.n1059 25.6005
R11754 VDD.n1065 VDD.n1062 25.6005
R11755 VDD.n1068 VDD.n1065 25.6005
R11756 VDD.n1072 VDD.n1068 25.6005
R11757 VDD.n1471 VDD.n1468 25.6005
R11758 VDD.n1468 VDD.n1465 25.6005
R11759 VDD.n1465 VDD.n1461 25.6005
R11760 VDD.n1461 VDD.n1459 25.6005
R11761 VDD.n1214 VDD.n1209 25.6005
R11762 VDD.n1209 VDD.n1206 25.6005
R11763 VDD.n1206 VDD.n1203 25.6005
R11764 VDD.n1130 VDD.n1126 25.6005
R11765 VDD.n1260 VDD.n1254 25.6005
R11766 VDD.n1254 VDD.n1251 25.6005
R11767 VDD.n1251 VDD.n1248 25.6005
R11768 VDD.n1248 VDD.n1245 25.6005
R11769 VDD.n415 VDD.n412 25.6005
R11770 VDD.n7 VDD.n4 25.6005
R11771 VDD.n9 VDD.n7 25.6005
R11772 VDD.n15 VDD.n9 25.6005
R11773 VDD.n640 VDD.n637 25.6005
R11774 VDD.n637 VDD.n634 25.6005
R11775 VDD.n634 VDD.n630 25.6005
R11776 VDD.n630 VDD.n628 25.6005
R11777 VDD.n229 VDD.n225 25.6005
R11778 VDD.n225 VDD.n222 25.6005
R11779 VDD.n222 VDD.n219 25.6005
R11780 VDD.n219 VDD.n216 25.6005
R11781 VDD.n216 VDD.n213 25.6005
R11782 VDD.n213 VDD.n210 25.6005
R11783 VDD.n210 VDD.n207 25.6005
R11784 VDD.n207 VDD.n204 25.6005
R11785 VDD.n204 VDD.n201 25.6005
R11786 VDD.n201 VDD.n198 25.6005
R11787 VDD.n198 VDD.n195 25.6005
R11788 VDD.n195 VDD.n192 25.6005
R11789 VDD.n192 VDD.n189 25.6005
R11790 VDD.n586 VDD.n583 25.6005
R11791 VDD.n589 VDD.n586 25.6005
R11792 VDD.n592 VDD.n589 25.6005
R11793 VDD.n595 VDD.n592 25.6005
R11794 VDD.n598 VDD.n595 25.6005
R11795 VDD.n601 VDD.n598 25.6005
R11796 VDD.n604 VDD.n601 25.6005
R11797 VDD.n607 VDD.n604 25.6005
R11798 VDD.n610 VDD.n607 25.6005
R11799 VDD.n613 VDD.n610 25.6005
R11800 VDD.n616 VDD.n613 25.6005
R11801 VDD.n619 VDD.n616 25.6005
R11802 VDD.n622 VDD.n619 25.6005
R11803 VDD.n626 VDD.n622 25.6005
R11804 VDD.n243 VDD.n240 25.6005
R11805 VDD.n240 VDD.n237 25.6005
R11806 VDD.n237 VDD.n233 25.6005
R11807 VDD.n233 VDD.n231 25.6005
R11808 VDD.n768 VDD.n763 25.6005
R11809 VDD.n763 VDD.n760 25.6005
R11810 VDD.n760 VDD.n757 25.6005
R11811 VDD.n684 VDD.n680 25.6005
R11812 VDD.n32 VDD.n26 25.6005
R11813 VDD.n26 VDD.n23 25.6005
R11814 VDD.n23 VDD.n20 25.6005
R11815 VDD.n20 VDD.n17 25.6005
R11816 VDD.n7815 VDD.n7809 25.3507
R11817 VDD.n7848 VDD.n7842 25.3507
R11818 VDD.n6284 VDD.n6283 25.3507
R11819 VDD.n6390 VDD.n6389 25.3507
R11820 VDD.n5953 VDD.n5888 25.3507
R11821 VDD.n5430 VDD.n5429 25.3507
R11822 VDD.n5536 VDD.n5535 25.3507
R11823 VDD.n5099 VDD.n5034 25.3507
R11824 VDD.n4644 VDD.n4643 25.3507
R11825 VDD.n4750 VDD.n4749 25.3507
R11826 VDD.n4313 VDD.n4248 25.3507
R11827 VDD.n3790 VDD.n3789 25.3507
R11828 VDD.n3896 VDD.n3895 25.3507
R11829 VDD.n3459 VDD.n3394 25.3507
R11830 VDD.n3004 VDD.n3003 25.3507
R11831 VDD.n3110 VDD.n3109 25.3507
R11832 VDD.n2673 VDD.n2608 25.3507
R11833 VDD.n2149 VDD.n2148 25.3507
R11834 VDD.n2255 VDD.n2254 25.3507
R11835 VDD.n1818 VDD.n1753 25.3507
R11836 VDD.n1022 VDD.n1021 25.3507
R11837 VDD.n1367 VDD.n1366 25.3507
R11838 VDD.n1568 VDD.n1567 25.3507
R11839 VDD.n576 VDD.n575 25.3507
R11840 VDD.n139 VDD.n138 25.3507
R11841 VDD.n340 VDD.n339 25.3507
R11842 VDD.n7831 VDD.n7830 25.3505
R11843 VDD.n7866 VDD.n7865 25.3505
R11844 VDD.n6154 VDD.n6153 25.3505
R11845 VDD.n6151 VDD.n6150 25.3505
R11846 VDD.n6368 VDD.n5891 25.3505
R11847 VDD.n6393 VDD.n6392 25.3505
R11848 VDD.n6253 VDD.n6252 25.3505
R11849 VDD.n6056 VDD.n6053 25.3505
R11850 VDD.n6541 VDD.n6540 25.3505
R11851 VDD.n5300 VDD.n5299 25.3505
R11852 VDD.n5297 VDD.n5296 25.3505
R11853 VDD.n5514 VDD.n5037 25.3505
R11854 VDD.n5539 VDD.n5538 25.3505
R11855 VDD.n5399 VDD.n5398 25.3505
R11856 VDD.n5202 VDD.n5199 25.3505
R11857 VDD.n5687 VDD.n5686 25.3505
R11858 VDD.n4514 VDD.n4513 25.3505
R11859 VDD.n4511 VDD.n4510 25.3505
R11860 VDD.n4728 VDD.n4251 25.3505
R11861 VDD.n4753 VDD.n4752 25.3505
R11862 VDD.n4613 VDD.n4612 25.3505
R11863 VDD.n4416 VDD.n4413 25.3505
R11864 VDD.n4901 VDD.n4900 25.3505
R11865 VDD.n3660 VDD.n3659 25.3505
R11866 VDD.n3657 VDD.n3656 25.3505
R11867 VDD.n3874 VDD.n3397 25.3505
R11868 VDD.n3899 VDD.n3898 25.3505
R11869 VDD.n3759 VDD.n3758 25.3505
R11870 VDD.n3562 VDD.n3559 25.3505
R11871 VDD.n4047 VDD.n4046 25.3505
R11872 VDD.n2874 VDD.n2873 25.3505
R11873 VDD.n2871 VDD.n2870 25.3505
R11874 VDD.n3088 VDD.n2611 25.3505
R11875 VDD.n3113 VDD.n3112 25.3505
R11876 VDD.n2973 VDD.n2972 25.3505
R11877 VDD.n2776 VDD.n2773 25.3505
R11878 VDD.n3261 VDD.n3260 25.3505
R11879 VDD.n2019 VDD.n2018 25.3505
R11880 VDD.n2016 VDD.n2015 25.3505
R11881 VDD.n2233 VDD.n1756 25.3505
R11882 VDD.n2258 VDD.n2257 25.3505
R11883 VDD.n2118 VDD.n2117 25.3505
R11884 VDD.n1921 VDD.n1918 25.3505
R11885 VDD.n2406 VDD.n2405 25.3505
R11886 VDD.n1313 VDD.n1312 25.3505
R11887 VDD.n1322 VDD.n1321 25.3505
R11888 VDD.n1400 VDD.n1399 25.3505
R11889 VDD.n1509 VDD.n1508 25.3505
R11890 VDD.n979 VDD.n978 25.3505
R11891 VDD.n985 VDD.n984 25.3505
R11892 VDD.n1186 VDD.n1185 25.3505
R11893 VDD.n85 VDD.n84 25.3505
R11894 VDD.n94 VDD.n93 25.3505
R11895 VDD.n172 VDD.n171 25.3505
R11896 VDD.n281 VDD.n280 25.3505
R11897 VDD.n533 VDD.n532 25.3505
R11898 VDD.n539 VDD.n538 25.3505
R11899 VDD.n740 VDD.n739 25.3505
R11900 VDD.n12489 VDD.n12488 23.5867
R11901 VDD.n12462 VDD.n12438 23.5867
R11902 VDD.n9951 VDD.t194 23.5572
R11903 VDD.n5749 VDD.t189 23.5572
R11904 VDD.n4109 VDD.t72 23.5572
R11905 VDD.n2468 VDD.t163 23.5572
R11906 VDD.n828 VDD.t203 23.5572
R11907 VDD.n9978 VDD.n9977 23.4711
R11908 VDD.n12420 VDD.n6923 23.2949
R11909 VDD.n10980 VDD.n9197 23.2817
R11910 VDD.n10983 VDD.n10982 23.2817
R11911 VDD.n5939 VDD.n5931 23.0774
R11912 VDD.n6343 VDD.n5940 23.0774
R11913 VDD.n6317 VDD.n5783 23.0774
R11914 VDD.n5085 VDD.n5077 23.0774
R11915 VDD.n5489 VDD.n5086 23.0774
R11916 VDD.n5463 VDD.n4929 23.0774
R11917 VDD.n4299 VDD.n4291 23.0774
R11918 VDD.n4703 VDD.n4300 23.0774
R11919 VDD.n4677 VDD.n4143 23.0774
R11920 VDD.n3445 VDD.n3437 23.0774
R11921 VDD.n3849 VDD.n3446 23.0774
R11922 VDD.n3823 VDD.n3289 23.0774
R11923 VDD.n2659 VDD.n2651 23.0774
R11924 VDD.n3063 VDD.n2660 23.0774
R11925 VDD.n3037 VDD.n2503 23.0774
R11926 VDD.n1804 VDD.n1796 23.0774
R11927 VDD.n2208 VDD.n1805 23.0774
R11928 VDD.n2182 VDD.n1648 23.0774
R11929 VDD.n10067 VDD.n10066 23.0522
R11930 VDD.n10625 VDD.n10587 23.0522
R11931 VDD.n10564 VDD.n10502 23.0522
R11932 VDD.n9585 VDD.n9573 23.0522
R11933 VDD.n10720 VDD.n10718 23.0522
R11934 VDD.n9440 VDD.n9392 23.0522
R11935 VDD.n8932 VDD.n8931 22.1478
R11936 VDD.n9263 VDD.n9261 22.1478
R11937 VDD.n10923 VDD.n9342 22.1478
R11938 VDD.n8788 VDD.n8787 22.1478
R11939 VDD.n8813 VDD.n8794 22.1478
R11940 VDD.n5923 VDD.t0 21.7954
R11941 VDD.t173 VDD.n5790 21.7954
R11942 VDD.n6547 VDD.t173 21.7954
R11943 VDD.n5069 VDD.t61 21.7954
R11944 VDD.t193 VDD.n4936 21.7954
R11945 VDD.n5693 VDD.t193 21.7954
R11946 VDD.n4283 VDD.t118 21.7954
R11947 VDD.t79 VDD.n4150 21.7954
R11948 VDD.n4907 VDD.t79 21.7954
R11949 VDD.n3429 VDD.t25 21.7954
R11950 VDD.t26 VDD.n3296 21.7954
R11951 VDD.n4053 VDD.t26 21.7954
R11952 VDD.n2643 VDD.t96 21.7954
R11953 VDD.t179 VDD.n2510 21.7954
R11954 VDD.n3267 VDD.t179 21.7954
R11955 VDD.n1788 VDD.t92 21.7954
R11956 VDD.t17 VDD.n1655 21.7954
R11957 VDD.n2412 VDD.t17 21.7954
R11958 VDD.n1190 VDD.t71 21.7954
R11959 VDD.n744 VDD.t201 21.7954
R11960 VDD.n10478 VDD.n6923 21.468
R11961 VDD.n10101 VDD.n10100 21.2396
R11962 VDD.n10097 VDD.n10096 21.1681
R11963 VDD.n5745 VDD.n5740 21.1346
R11964 VDD.n4105 VDD.n4100 21.1346
R11965 VDD.n2464 VDD.n2459 21.1346
R11966 VDD.n824 VDD.n819 21.1346
R11967 VDD.n9962 VDD.n9910 20.9478
R11968 VDD.n8590 VDD.n7756 20.7186
R11969 VDD.n8590 VDD.n7757 20.7186
R11970 VDD.n8590 VDD.n7758 20.7186
R11971 VDD.n8590 VDD.n7759 20.7186
R11972 VDD.n8590 VDD.n8589 20.7186
R11973 VDD.n8591 VDD.n8590 20.7186
R11974 VDD.n6493 VDD.n6492 20.6044
R11975 VDD.n5639 VDD.n5638 20.6044
R11976 VDD.n4853 VDD.n4852 20.6044
R11977 VDD.n3999 VDD.n3998 20.6044
R11978 VDD.n3213 VDD.n3212 20.6044
R11979 VDD.n2358 VDD.n2357 20.6044
R11980 VDD.n1089 VDD.n1086 20.6044
R11981 VDD.n643 VDD.n640 20.6044
R11982 VDD.n9652 VDD.n9647 20.5156
R11983 VDD.n10795 VDD.n10790 20.5156
R11984 VDD.n8871 VDD.n8866 20.5156
R11985 VDD.n9665 VDD.n9664 20.5153
R11986 VDD.n10808 VDD.n10807 20.5153
R11987 VDD.n9004 VDD.n9003 20.5153
R11988 VDD.n9282 VDD.n9281 20.5152
R11989 VDD.n9412 VDD.n9411 20.5152
R11990 VDD.n6350 VDD.n5931 20.5133
R11991 VDD.n6006 VDD.n5940 20.5133
R11992 VDD.n6317 VDD.n6304 20.5133
R11993 VDD.n5496 VDD.n5077 20.5133
R11994 VDD.n5152 VDD.n5086 20.5133
R11995 VDD.n5463 VDD.n5450 20.5133
R11996 VDD.n4710 VDD.n4291 20.5133
R11997 VDD.n4366 VDD.n4300 20.5133
R11998 VDD.n4677 VDD.n4664 20.5133
R11999 VDD.n3856 VDD.n3437 20.5133
R12000 VDD.n3512 VDD.n3446 20.5133
R12001 VDD.n3823 VDD.n3810 20.5133
R12002 VDD.n3070 VDD.n2651 20.5133
R12003 VDD.n2726 VDD.n2660 20.5133
R12004 VDD.n3037 VDD.n3024 20.5133
R12005 VDD.n2215 VDD.n1796 20.5133
R12006 VDD.n1871 VDD.n1805 20.5133
R12007 VDD.n2182 VDD.n2169 20.5133
R12008 VDD.n12691 VDD.n12690 20.3855
R12009 VDD.n10494 VDD.n10420 20.0857
R12010 VDD.n8968 VDD.n8860 19.9534
R12011 VDD.n8968 VDD.n8967 19.9534
R12012 VDD.n8990 VDD.n8832 19.9534
R12013 VDD.n8990 VDD.n8833 19.9534
R12014 VDD.n10957 VDD.n9197 19.9425
R12015 VDD.n10982 VDD.n9070 19.9425
R12016 VDD.n9695 VDD.n9642 19.7698
R12017 VDD.n9702 VDD.n9640 19.7698
R12018 VDD.n10852 VDD.n10688 19.7698
R12019 VDD.n10845 VDD.n10686 19.7698
R12020 VDD.n9593 VDD.n9584 19.7591
R12021 VDD.n10764 VDD.n10763 19.7591
R12022 VDD.n9403 VDD.n9397 19.7591
R12023 VDD.n9690 VDD.n9643 19.7549
R12024 VDD.n9707 VDD.n9639 19.7549
R12025 VDD.n10857 VDD.n10689 19.7549
R12026 VDD.n10840 VDD.n10685 19.7549
R12027 VDD.n9923 VDD.t211 19.7525
R12028 VDD.n9740 VDD.n9560 19.7383
R12029 VDD.n9712 VDD.n9638 19.7383
R12030 VDD.n10862 VDD.n10681 19.7383
R12031 VDD.n10835 VDD.n10684 19.7383
R12032 VDD.n9744 VDD.n9559 19.7199
R12033 VDD.n9717 VDD.n9637 19.7199
R12034 VDD.n9547 VDD.n9545 19.7199
R12035 VDD.n9535 VDD.n9530 19.7199
R12036 VDD.n9789 VDD.n9517 19.7199
R12037 VDD.n9802 VDD.n9503 19.7199
R12038 VDD.n9492 VDD.n9487 19.7199
R12039 VDD.n9863 VDD.n9862 19.7199
R12040 VDD.n10890 VDD.n10889 19.7199
R12041 VDD.n10868 VDD.n10691 19.7199
R12042 VDD.n10830 VDD.n10683 19.7199
R12043 VDD.n8940 VDD.n8882 19.7199
R12044 VDD.n8843 VDD.n8784 19.7199
R12045 VDD.n9026 VDD.n8798 19.7199
R12046 VDD.n9302 VDD.n9301 19.7199
R12047 VDD.n9738 VDD.n9737 19.6997
R12048 VDD.n9722 VDD.n9636 19.6997
R12049 VDD.n9762 VDD.n9761 19.6997
R12050 VDD.n9773 VDD.n9772 19.6997
R12051 VDD.n9783 VDD.n9782 19.6997
R12052 VDD.n9809 VDD.n9808 19.6997
R12053 VDD.n9820 VDD.n9819 19.6997
R12054 VDD.n9855 VDD.n9854 19.6997
R12055 VDD.n10882 VDD.n10678 19.6997
R12056 VDD.n10877 VDD.n10876 19.6997
R12057 VDD.n10825 VDD.n10682 19.6997
R12058 VDD.n8945 VDD.n8880 19.6997
R12059 VDD.n8848 VDD.n8789 19.6997
R12060 VDD.n9021 VDD.n8796 19.6997
R12061 VDD.n9296 VDD.n9264 19.6997
R12062 VDD.n9729 VDD.n9728 19.6777
R12063 VDD.n10820 VDD.n10690 19.6777
R12064 VDD.n8950 VDD.n8878 19.6777
R12065 VDD.n8853 VDD.n8790 19.6777
R12066 VDD.n9016 VDD.n8797 19.6777
R12067 VDD.n9291 VDD.n9265 19.6777
R12068 VDD.n12423 VDD.n6912 19.6557
R12069 VDD.n10043 VDD.n10042 19.3601
R12070 VDD.n10602 VDD.n10601 19.3601
R12071 VDD.n9369 VDD.n9367 19.3601
R12072 VDD.n10541 VDD.n10540 19.3599
R12073 VDD.n9635 VDD.n9634 19.3599
R12074 VDD.n10733 VDD.n10731 19.3599
R12075 VDD.n8914 VDD.n8887 19.3599
R12076 VDD.n10482 VDD.n10447 19.2933
R12077 VDD.n10024 VDD.n10021 19.131
R12078 VDD.n10143 VDD.n10142 19.131
R12079 VDD.n10529 VDD.n10514 19.131
R12080 VDD.n9657 VDD.n9656 19.0069
R12081 VDD.n9671 VDD.n9659 19.0069
R12082 VDD.n10800 VDD.n10799 19.0069
R12083 VDD.n10814 VDD.n10802 19.0069
R12084 VDD.n8876 VDD.n8875 19.0069
R12085 VDD.n8954 VDD.n8862 19.0069
R12086 VDD.n8974 VDD.n8973 19.0069
R12087 VDD.n9010 VDD.n8998 19.0069
R12088 VDD.n8977 VDD.n8835 19.0069
R12089 VDD.n8996 VDD.n8995 19.0069
R12090 VDD.n9287 VDD.n9286 19.0069
R12091 VDD.n9417 VDD.n9416 19.0069
R12092 VDD.n9341 VDD.n9340 18.986
R12093 VDD.n9422 VDD.n9421 18.9099
R12094 VDD.n6419 VDD.n6418 18.7439
R12095 VDD.n5565 VDD.n5564 18.7439
R12096 VDD.n4779 VDD.n4778 18.7439
R12097 VDD.n3925 VDD.n3924 18.7439
R12098 VDD.n3139 VDD.n3138 18.7439
R12099 VDD.n2284 VDD.n2283 18.7439
R12100 VDD.n1474 VDD.n1471 18.7439
R12101 VDD.n246 VDD.n243 18.7439
R12102 VDD.n10447 VDD.n10434 17.9019
R12103 VDD.n9951 VDD.t133 17.8272
R12104 VDD.n5749 VDD.t15 17.8272
R12105 VDD.n4109 VDD.t13 17.8272
R12106 VDD.n2468 VDD.t200 17.8272
R12107 VDD.n828 VDD.t31 17.8272
R12108 VDD.n12248 VDD.n7071 17.8254
R12109 VDD.t183 VDD.n6712 17.6875
R12110 VDD.n9060 VDD.n9059 17.6125
R12111 VDD.n9138 VDD.n9090 17.3826
R12112 VDD.n9968 VDD.n9907 17.2489
R12113 VDD.n9931 VDD.n9918 17.2489
R12114 VDD.n9916 VDD.n9913 17.2489
R12115 VDD.n5755 VDD.n5741 17.2489
R12116 VDD.n4115 VDD.n4101 17.2489
R12117 VDD.n2475 VDD.n2460 17.2489
R12118 VDD.n835 VDD.n820 17.2489
R12119 VDD.n9149 VDD.n9148 16.6542
R12120 VDD.n12680 VDD.n6713 16.4884
R12121 VDD.n6722 VDD.n6720 16.4884
R12122 VDD.n12674 VDD.n6721 16.4884
R12123 VDD.n6748 VDD.n6747 16.4884
R12124 VDD.n12668 VDD.n6749 16.4884
R12125 VDD.n6754 VDD.n6753 16.4884
R12126 VDD.n10243 VDD.n6758 16.4884
R12127 VDD.n12656 VDD.n6759 16.4884
R12128 VDD.n6764 VDD.n6763 16.4884
R12129 VDD.n12650 VDD.n6765 16.4884
R12130 VDD.n6770 VDD.n6769 16.4884
R12131 VDD.n12644 VDD.n6771 16.4884
R12132 VDD.n12638 VDD.n6777 16.4884
R12133 VDD.n6782 VDD.n6781 16.4884
R12134 VDD.n12632 VDD.n6783 16.4884
R12135 VDD.n6788 VDD.n6787 16.4884
R12136 VDD.n12626 VDD.n6789 16.4884
R12137 VDD.n10226 VDD.n10225 16.4884
R12138 VDD.n12620 VDD.n6793 16.4884
R12139 VDD.n6798 VDD.n6797 16.4884
R12140 VDD.n12614 VDD.n6799 16.4884
R12141 VDD.n6804 VDD.n6803 16.4884
R12142 VDD.n12608 VDD.n6805 16.4884
R12143 VDD.n6810 VDD.n6809 16.4884
R12144 VDD.n12602 VDD.n6811 16.4884
R12145 VDD.n6816 VDD.n6815 16.4884
R12146 VDD.n10211 VDD.n6820 16.4884
R12147 VDD.n10334 VDD.n6824 16.4884
R12148 VDD.n12584 VDD.n6825 16.4884
R12149 VDD.n6830 VDD.n6829 16.4884
R12150 VDD.n12578 VDD.n6831 16.4884
R12151 VDD.n12572 VDD.n6837 16.4884
R12152 VDD.n6842 VDD.n6841 16.4884
R12153 VDD.n12566 VDD.n6843 16.4884
R12154 VDD.n6848 VDD.n6847 16.4884
R12155 VDD.n12560 VDD.n6849 16.4884
R12156 VDD.n10193 VDD.n10192 16.4884
R12157 VDD.n12554 VDD.n6853 16.4884
R12158 VDD.n6858 VDD.n6857 16.4884
R12159 VDD.n12548 VDD.n6859 16.4884
R12160 VDD.n6864 VDD.n6863 16.4884
R12161 VDD.n12542 VDD.n6865 16.4884
R12162 VDD.n6870 VDD.n6869 16.4884
R12163 VDD.n10182 VDD.n6874 16.4884
R12164 VDD.n12530 VDD.n6875 16.4884
R12165 VDD.n6880 VDD.n6879 16.4884
R12166 VDD.n12524 VDD.n6881 16.4884
R12167 VDD.n6886 VDD.n6885 16.4884
R12168 VDD.n12518 VDD.n6887 16.4884
R12169 VDD.n6892 VDD.n6891 16.4884
R12170 VDD.n12512 VDD.n6893 16.4884
R12171 VDD.n12506 VDD.n6899 16.4884
R12172 VDD.n6904 VDD.n6903 16.4884
R12173 VDD.n12500 VDD.n6905 16.4884
R12174 VDD.n10420 VDD.n10164 16.4884
R12175 VDD.n10062 VDD.n10028 16.466
R12176 VDD.n10623 VDD.n10588 16.466
R12177 VDD.n10562 VDD.n10503 16.466
R12178 VDD.n9616 VDD.n9569 16.466
R12179 VDD.n10748 VDD.n10747 16.466
R12180 VDD.n9061 VDD.n8765 16.466
R12181 VDD.n9391 VDD.n9361 16.466
R12182 VDD.n12431 VDD.n12428 16.4319
R12183 VDD.n12467 VDD.n12435 16.4313
R12184 VDD.n12371 VDD.n6967 16.1937
R12185 VDD.n9152 VDD.n9151 15.9242
R12186 VDD.n6898 VDD.t28 15.8888
R12187 VDD.n9923 VDD.t210 15.6574
R12188 VDD.n6341 VDD.n6003 15.6165
R12189 VDD.n6295 VDD.n5787 15.6165
R12190 VDD.n5487 VDD.n5149 15.6165
R12191 VDD.n5441 VDD.n4933 15.6165
R12192 VDD.n4701 VDD.n4363 15.6165
R12193 VDD.n4655 VDD.n4147 15.6165
R12194 VDD.n3847 VDD.n3509 15.6165
R12195 VDD.n3801 VDD.n3293 15.6165
R12196 VDD.n3061 VDD.n2723 15.6165
R12197 VDD.n3015 VDD.n2507 15.6165
R12198 VDD.n2206 VDD.n1868 15.6165
R12199 VDD.n2160 VDD.n1652 15.6165
R12200 VDD.n1516 VDD.n1512 15.6165
R12201 VDD.n1141 VDD.n1140 15.6165
R12202 VDD.n288 VDD.n284 15.6165
R12203 VDD.n695 VDD.n694 15.6165
R12204 VDD.n12248 VDD.n12247 15.0799
R12205 VDD.n10099 VDD.n10006 15.056
R12206 VDD.n9190 VDD.n9075 14.8411
R12207 VDD.t0 VDD.n5917 14.7441
R12208 VDD.n6350 VDD.t105 14.7441
R12209 VDD.t100 VDD.n6006 14.7441
R12210 VDD.n6331 VDD.t69 14.7441
R12211 VDD.n6298 VDD.t69 14.7441
R12212 VDD.n6304 VDD.t174 14.7441
R12213 VDD.t61 VDD.n5063 14.7441
R12214 VDD.n5496 VDD.t103 14.7441
R12215 VDD.t146 VDD.n5152 14.7441
R12216 VDD.n5477 VDD.t147 14.7441
R12217 VDD.n5444 VDD.t147 14.7441
R12218 VDD.n5450 VDD.t158 14.7441
R12219 VDD.t118 VDD.n4277 14.7441
R12220 VDD.n4710 VDD.t122 14.7441
R12221 VDD.t186 VDD.n4366 14.7441
R12222 VDD.n4691 VDD.t80 14.7441
R12223 VDD.n4658 VDD.t80 14.7441
R12224 VDD.n4664 VDD.t180 14.7441
R12225 VDD.t25 VDD.n3423 14.7441
R12226 VDD.n3856 VDD.t120 14.7441
R12227 VDD.t125 VDD.n3512 14.7441
R12228 VDD.n3837 VDD.t65 14.7441
R12229 VDD.n3804 VDD.t65 14.7441
R12230 VDD.n3810 VDD.t7 14.7441
R12231 VDD.t96 VDD.n2637 14.7441
R12232 VDD.n3070 VDD.t98 14.7441
R12233 VDD.t82 VDD.n2726 14.7441
R12234 VDD.n3051 VDD.t32 14.7441
R12235 VDD.n3018 VDD.t32 14.7441
R12236 VDD.n3024 VDD.t177 14.7441
R12237 VDD.t92 VDD.n1782 14.7441
R12238 VDD.n2215 VDD.t94 14.7441
R12239 VDD.t20 VDD.n1871 14.7441
R12240 VDD.n2196 VDD.t18 14.7441
R12241 VDD.n2163 VDD.t18 14.7441
R12242 VDD.n2169 VDD.t101 14.7441
R12243 VDD.n1580 VDD.t9 14.7441
R12244 VDD.n1595 VDD.t88 14.7441
R12245 VDD.n1606 VDD.t172 14.7441
R12246 VDD.n1629 VDD.t63 14.7441
R12247 VDD.n1215 VDD.t77 14.7441
R12248 VDD.n352 VDD.t90 14.7441
R12249 VDD.n367 VDD.t85 14.7441
R12250 VDD.n378 VDD.t136 14.7441
R12251 VDD.n401 VDD.t137 14.7441
R12252 VDD.n769 VDD.t156 14.7441
R12253 VDD.n6836 VDD.t154 14.6897
R12254 VDD.n10109 VDD.n10108 14.6773
R12255 VDD.n12474 VDD.n12433 14.4934
R12256 VDD.n12433 VDD.n12430 14.4934
R12257 VDD.n8197 VDD.n8092 14.2505
R12258 VDD.n6003 VDD.n5986 14.2085
R12259 VDD.n6551 VDD.n5787 14.2085
R12260 VDD.n5149 VDD.n5132 14.2085
R12261 VDD.n5697 VDD.n4933 14.2085
R12262 VDD.n4363 VDD.n4346 14.2085
R12263 VDD.n4911 VDD.n4147 14.2085
R12264 VDD.n3509 VDD.n3492 14.2085
R12265 VDD.n4057 VDD.n3293 14.2085
R12266 VDD.n2723 VDD.n2706 14.2085
R12267 VDD.n3271 VDD.n2507 14.2085
R12268 VDD.n1868 VDD.n1851 14.2085
R12269 VDD.n2416 VDD.n1652 14.2085
R12270 VDD.n1518 VDD.n1516 14.2085
R12271 VDD.n1143 VDD.n1141 14.2085
R12272 VDD.n290 VDD.n288 14.2085
R12273 VDD.n697 VDD.n695 14.2085
R12274 VDD.n6337 VDD.n6007 14.1031
R12275 VDD.n6331 VDD.n6022 14.1031
R12276 VDD.n6298 VDD.n6293 14.1031
R12277 VDD.n6325 VDD.n6045 14.1031
R12278 VDD.n5483 VDD.n5153 14.1031
R12279 VDD.n5477 VDD.n5168 14.1031
R12280 VDD.n5444 VDD.n5439 14.1031
R12281 VDD.n5471 VDD.n5191 14.1031
R12282 VDD.n4697 VDD.n4367 14.1031
R12283 VDD.n4691 VDD.n4382 14.1031
R12284 VDD.n4658 VDD.n4653 14.1031
R12285 VDD.n4685 VDD.n4405 14.1031
R12286 VDD.n3843 VDD.n3513 14.1031
R12287 VDD.n3837 VDD.n3528 14.1031
R12288 VDD.n3804 VDD.n3799 14.1031
R12289 VDD.n3831 VDD.n3551 14.1031
R12290 VDD.n3057 VDD.n2727 14.1031
R12291 VDD.n3051 VDD.n2742 14.1031
R12292 VDD.n3018 VDD.n3013 14.1031
R12293 VDD.n3045 VDD.n2765 14.1031
R12294 VDD.n2202 VDD.n1872 14.1031
R12295 VDD.n2196 VDD.n1887 14.1031
R12296 VDD.n2163 VDD.n2158 14.1031
R12297 VDD.n2190 VDD.n1910 14.1031
R12298 VDD.n6712 VDD.n6702 14.0901
R12299 VDD.n12453 VDD.n12452 13.7591
R12300 VDD.n10073 VDD.n10072 13.5534
R12301 VDD.n10055 VDD.n10031 13.5534
R12302 VDD.n10049 VDD.n10038 13.5534
R12303 VDD.n10633 VDD.n10632 13.5534
R12304 VDD.n10614 VDD.n10590 13.5534
R12305 VDD.n10608 VDD.n10597 13.5534
R12306 VDD.n10521 VDD.n10519 13.5534
R12307 VDD.n10556 VDD.n10534 13.5534
R12308 VDD.n10550 VDD.n10549 13.5534
R12309 VDD.n9592 VDD.n9591 13.5534
R12310 VDD.n9603 VDD.n9602 13.5534
R12311 VDD.n9614 VDD.n9613 13.5534
R12312 VDD.n9621 VDD.n9620 13.5534
R12313 VDD.n9629 VDD.n9628 13.5534
R12314 VDD.n10704 VDD.n10701 13.5534
R12315 VDD.n10757 VDD.n10710 13.5534
R12316 VDD.n10751 VDD.n10714 13.5534
R12317 VDD.n10745 VDD.n10744 13.5534
R12318 VDD.n10727 VDD.n10725 13.5534
R12319 VDD.n8934 VDD.n8886 13.5534
R12320 VDD.n9051 VDD.n9050 13.5534
R12321 VDD.n9032 VDD.n8799 13.5534
R12322 VDD.n8909 VDD.n8896 13.5534
R12323 VDD.n9313 VDD.n9312 13.5534
R12324 VDD.n9376 VDD.n9363 13.5534
R12325 VDD.n9443 VDD.n9442 13.5534
R12326 VDD.n9434 VDD.n9433 13.5534
R12327 VDD.n9400 VDD.n9398 13.5534
R12328 VDD.n12494 VDD.n6909 13.5534
R12329 VDD.n12487 VDD.n12486 13.5534
R12330 VDD.n12475 VDD.n12432 13.5534
R12331 VDD.n12461 VDD.n12439 13.5534
R12332 VDD.n12455 VDD.n12447 13.5534
R12333 VDD.n6776 VDD.t185 13.4906
R12334 VDD.n5790 VDD.n5784 13.462
R12335 VDD.n4936 VDD.n4930 13.462
R12336 VDD.n4150 VDD.n4144 13.462
R12337 VDD.n3296 VDD.n3290 13.462
R12338 VDD.n2510 VDD.n2504 13.462
R12339 VDD.n1655 VDD.n1649 13.462
R12340 VDD.n10432 VDD.n10423 13.3252
R12341 VDD.n12468 VDD.n12436 12.8072
R12342 VDD.n12465 VDD.n12436 12.8072
R12343 VDD.n10064 VDD.n10013 12.8005
R12344 VDD.n10617 VDD.n10586 12.8005
R12345 VDD.n10506 VDD.n10501 12.8005
R12346 VDD.n8928 VDD.n8771 12.8005
R12347 VDD.n9048 VDD.n9040 12.8005
R12348 VDD.n8811 VDD.n8795 12.8005
R12349 VDD.n8903 VDD.n8902 12.8005
R12350 VDD.n9310 VDD.n9309 12.8005
R12351 VDD.n9331 VDD.n9328 12.8005
R12352 VDD.n9386 VDD.n9355 12.8005
R12353 VDD.t144 VDD.n5715 12.789
R12354 VDD.t109 VDD.n4075 12.789
R12355 VDD.t23 VDD.n2434 12.789
R12356 VDD.t126 VDD.n794 12.789
R12357 VDD.n9739 VDD.n9730 12.6901
R12358 VDD.n9763 VDD.n9548 12.6901
R12359 VDD.n9775 VDD.n9523 12.6901
R12360 VDD.n9784 VDD.n9518 12.6901
R12361 VDD.n9810 VDD.n9504 12.6901
R12362 VDD.n9822 VDD.n9480 12.6901
R12363 VDD.n10878 VDD.n10692 12.6901
R12364 VDD.n8590 VDD.n7755 12.6672
R12365 VDD.n9856 VDD.n9837 12.2367
R12366 VDD.n10883 VDD.n10680 12.2367
R12367 VDD.n12425 VDD.n12423 12.2348
R12368 VDD.n9976 VDD.n9975 12.1342
R12369 VDD.n5981 VDD.n5877 12.0325
R12370 VDD.n6517 VDD.n5788 12.0325
R12371 VDD.n5127 VDD.n5023 12.0325
R12372 VDD.n5663 VDD.n4934 12.0325
R12373 VDD.n4341 VDD.n4237 12.0325
R12374 VDD.n4877 VDD.n4148 12.0325
R12375 VDD.n3487 VDD.n3383 12.0325
R12376 VDD.n4023 VDD.n3294 12.0325
R12377 VDD.n2701 VDD.n2597 12.0325
R12378 VDD.n3237 VDD.n2508 12.0325
R12379 VDD.n1846 VDD.n1742 12.0325
R12380 VDD.n2382 VDD.n1653 12.0325
R12381 VDD.n1525 VDD.n1524 12.0325
R12382 VDD.n1150 VDD.n1149 12.0325
R12383 VDD.n297 VDD.n296 12.0325
R12384 VDD.n704 VDD.n703 12.0325
R12385 VDD.n12692 VDD.t4 11.8979
R12386 VDD.n10964 VDD.n10962 11.7802
R12387 VDD.n10992 VDD.n10990 11.7802
R12388 VDD.n9110 VDD.n9091 11.6711
R12389 VDD.n10975 VDD.n10973 11.5947
R12390 VDD.n12536 VDD.t150 11.3921
R12391 VDD.n9971 VDD.n9970 11.1178
R12392 VDD.n10978 VDD.n9199 10.8935
R12393 VDD.n10959 VDD.n9205 10.8935
R12394 VDD.n6041 VDD.n5928 10.4112
R12395 VDD.n6042 VDD.n6041 10.4112
R12396 VDD.n5187 VDD.n5074 10.4112
R12397 VDD.n5188 VDD.n5187 10.4112
R12398 VDD.n4401 VDD.n4288 10.4112
R12399 VDD.n4402 VDD.n4401 10.4112
R12400 VDD.n3547 VDD.n3434 10.4112
R12401 VDD.n3548 VDD.n3547 10.4112
R12402 VDD.n2761 VDD.n2648 10.4112
R12403 VDD.n2762 VDD.n2761 10.4112
R12404 VDD.n1906 VDD.n1793 10.4112
R12405 VDD.n1907 VDD.n1906 10.4112
R12406 VDD.n866 VDD.n865 10.4112
R12407 VDD.n868 VDD.n866 10.4112
R12408 VDD.n420 VDD.n419 10.4112
R12409 VDD.n422 VDD.n420 10.4112
R12410 VDD.n12590 VDD.t27 10.193
R12411 VDD.n10162 VDD.n6920 9.89321
R12412 VDD.n10053 VDD.n10032 9.87981
R12413 VDD.n10612 VDD.n10591 9.87981
R12414 VDD.n10553 VDD.n10552 9.87981
R12415 VDD.n9623 VDD.n9564 9.87981
R12416 VDD.n10738 VDD.n10722 9.87981
R12417 VDD.n8905 VDD.n8891 9.87981
R12418 VDD.n9384 VDD.n9362 9.87981
R12419 VDD.n10479 VDD.n6967 9.59343
R12420 VDD.n12456 VDD.n12446 9.33286
R12421 VDD.n12453 VDD.n12446 9.33286
R12422 VDD.n10048 VDD.n10037 9.3005
R12423 VDD.n10047 VDD.n10040 9.3005
R12424 VDD.n10047 VDD.n10046 9.3005
R12425 VDD.n10050 VDD.n10049 9.3005
R12426 VDD.n10052 VDD.n10051 9.3005
R12427 VDD.n10053 VDD.n10052 9.3005
R12428 VDD.n10036 VDD.n10033 9.3005
R12429 VDD.n10029 VDD.n10014 9.3005
R12430 VDD.n10023 VDD.n10022 9.3005
R12431 VDD.n10071 VDD.n10070 9.3005
R12432 VDD.n10021 VDD.n10019 9.3005
R12433 VDD.n10069 VDD.n10068 9.3005
R12434 VDD.n10068 VDD.n10067 9.3005
R12435 VDD.n10077 VDD.n10020 9.3005
R12436 VDD.n10077 VDD.n10076 9.3005
R12437 VDD.n10035 VDD.n10031 9.3005
R12438 VDD.n10061 VDD.n10060 9.3005
R12439 VDD.n10062 VDD.n10061 9.3005
R12440 VDD.n10058 VDD.n10030 9.3005
R12441 VDD.n10092 VDD.n10007 9.3005
R12442 VDD.n10105 VDD.n10103 9.3005
R12443 VDD.n10091 VDD.n10090 9.3005
R12444 VDD.n10096 VDD.n10088 9.3005
R12445 VDD.n10112 VDD.n10111 9.3005
R12446 VDD.n10111 VDD.n10110 9.3005
R12447 VDD.n10104 VDD.n10095 9.3005
R12448 VDD.n10110 VDD.n10095 9.3005
R12449 VDD.n10107 VDD.n10106 9.3005
R12450 VDD.n10094 VDD.n10093 9.3005
R12451 VDD.n10110 VDD.n10094 9.3005
R12452 VDD.n10607 VDD.n10596 9.3005
R12453 VDD.n10606 VDD.n10599 9.3005
R12454 VDD.n10606 VDD.n10605 9.3005
R12455 VDD.n10609 VDD.n10608 9.3005
R12456 VDD.n10611 VDD.n10610 9.3005
R12457 VDD.n10612 VDD.n10611 9.3005
R12458 VDD.n10595 VDD.n10592 9.3005
R12459 VDD.n10619 VDD.n10618 9.3005
R12460 VDD.n10141 VDD.n10140 9.3005
R12461 VDD.n10147 VDD.n10146 9.3005
R12462 VDD.n10142 VDD.n10138 9.3005
R12463 VDD.n10585 VDD.n10584 9.3005
R12464 VDD.n10587 VDD.n10585 9.3005
R12465 VDD.n10638 VDD.n10637 9.3005
R12466 VDD.n10637 VDD.n10636 9.3005
R12467 VDD.n10594 VDD.n10590 9.3005
R12468 VDD.n10622 VDD.n10621 9.3005
R12469 VDD.n10623 VDD.n10622 9.3005
R12470 VDD.n10620 VDD.n10589 9.3005
R12471 VDD.n10438 VDD.n10434 9.3005
R12472 VDD.n10555 VDD.n10532 9.3005
R12473 VDD.n10547 VDD.n10539 9.3005
R12474 VDD.n10554 VDD.n10536 9.3005
R12475 VDD.n10554 VDD.n10553 9.3005
R12476 VDD.n10546 VDD.n10545 9.3005
R12477 VDD.n10545 VDD.n10538 9.3005
R12478 VDD.n10549 VDD.n10548 9.3005
R12479 VDD.n10525 VDD.n10524 9.3005
R12480 VDD.n10514 VDD.n10513 9.3005
R12481 VDD.n10518 VDD.n10517 9.3005
R12482 VDD.n10509 VDD.n10504 9.3005
R12483 VDD.n10557 VDD.n10556 9.3005
R12484 VDD.n10561 VDD.n10560 9.3005
R12485 VDD.n10562 VDD.n10561 9.3005
R12486 VDD.n10508 VDD.n10507 9.3005
R12487 VDD.n10500 VDD.n10153 9.3005
R12488 VDD.n10502 VDD.n10500 9.3005
R12489 VDD.n10527 VDD.n10526 9.3005
R12490 VDD.n10528 VDD.n10527 9.3005
R12491 VDD.n9929 VDD.n9928 9.3005
R12492 VDD.n9626 VDD.n9566 9.3005
R12493 VDD.n9568 VDD.n9567 9.3005
R12494 VDD.n9613 VDD.n9612 9.3005
R12495 VDD.n9563 VDD.n9562 9.3005
R12496 VDD.n9631 VDD.n9563 9.3005
R12497 VDD.n9628 VDD.n9627 9.3005
R12498 VDD.n9625 VDD.n9624 9.3005
R12499 VDD.n9624 VDD.n9623 9.3005
R12500 VDD.n9620 VDD.n9619 9.3005
R12501 VDD.n9618 VDD.n9617 9.3005
R12502 VDD.n9617 VDD.n9616 9.3005
R12503 VDD.n9572 VDD.n9571 9.3005
R12504 VDD.n9591 VDD.n9590 9.3005
R12505 VDD.n9608 VDD.n9607 9.3005
R12506 VDD.n9607 VDD.n9606 9.3005
R12507 VDD.n9602 VDD.n9601 9.3005
R12508 VDD.n9586 VDD.n9575 9.3005
R12509 VDD.n9586 VDD.n9585 9.3005
R12510 VDD.n9596 VDD.n9595 9.3005
R12511 VDD.n9670 VDD.n9660 9.3005
R12512 VDD.n9672 VDD.n9671 9.3005
R12513 VDD.n9669 VDD.n9662 9.3005
R12514 VDD.n9669 VDD.n9668 9.3005
R12515 VDD.n9656 VDD.n9644 9.3005
R12516 VDD.n9655 VDD.n9654 9.3005
R12517 VDD.n9653 VDD.n9646 9.3005
R12518 VDD.n9646 VDD.n9645 9.3005
R12519 VDD.n9726 VDD.n9676 9.3005
R12520 VDD.n9721 VDD.n9677 9.3005
R12521 VDD.n9716 VDD.n9678 9.3005
R12522 VDD.n9711 VDD.n9679 9.3005
R12523 VDD.n9706 VDD.n9680 9.3005
R12524 VDD.n9701 VDD.n9681 9.3005
R12525 VDD.n9696 VDD.n9682 9.3005
R12526 VDD.n9691 VDD.n9683 9.3005
R12527 VDD.n9686 VDD.n9685 9.3005
R12528 VDD.n9684 VDD.n9560 9.3005
R12529 VDD.n9688 VDD.n9687 9.3005
R12530 VDD.n9690 VDD.n9689 9.3005
R12531 VDD.n9693 VDD.n9692 9.3005
R12532 VDD.n9695 VDD.n9694 9.3005
R12533 VDD.n9698 VDD.n9697 9.3005
R12534 VDD.n9700 VDD.n9699 9.3005
R12535 VDD.n9703 VDD.n9702 9.3005
R12536 VDD.n9705 VDD.n9704 9.3005
R12537 VDD.n9708 VDD.n9707 9.3005
R12538 VDD.n9710 VDD.n9709 9.3005
R12539 VDD.n9713 VDD.n9712 9.3005
R12540 VDD.n9715 VDD.n9714 9.3005
R12541 VDD.n9718 VDD.n9717 9.3005
R12542 VDD.n9720 VDD.n9719 9.3005
R12543 VDD.n9723 VDD.n9722 9.3005
R12544 VDD.n9725 VDD.n9724 9.3005
R12545 VDD.n9728 VDD.n9727 9.3005
R12546 VDD.n9737 VDD.n9736 9.3005
R12547 VDD.n9734 VDD.n9733 9.3005
R12548 VDD.n9745 VDD.n9744 9.3005
R12549 VDD.n9742 VDD.n9741 9.3005
R12550 VDD.n9732 VDD.n9731 9.3005
R12551 VDD.n9761 VDD.n9760 9.3005
R12552 VDD.n9756 VDD.n9755 9.3005
R12553 VDD.n9765 VDD.n9543 9.3005
R12554 VDD.n9753 VDD.n9545 9.3005
R12555 VDD.n9752 VDD.n9549 9.3005
R12556 VDD.n9533 VDD.n9532 9.3005
R12557 VDD.n9536 VDD.n9535 9.3005
R12558 VDD.n9529 VDD.n9526 9.3005
R12559 VDD.n9772 VDD.n9771 9.3005
R12560 VDD.n9774 VDD.n9522 9.3005
R12561 VDD.n9782 VDD.n9509 9.3005
R12562 VDD.n9516 VDD.n9512 9.3005
R12563 VDD.n9790 VDD.n9789 9.3005
R12564 VDD.n9787 VDD.n9786 9.3005
R12565 VDD.n9781 VDD.n9780 9.3005
R12566 VDD.n9808 VDD.n9807 9.3005
R12567 VDD.n9813 VDD.n9812 9.3005
R12568 VDD.n9803 VDD.n9802 9.3005
R12569 VDD.n9801 VDD.n9800 9.3005
R12570 VDD.n9798 VDD.n9505 9.3005
R12571 VDD.n9490 VDD.n9489 9.3005
R12572 VDD.n9493 VDD.n9492 9.3005
R12573 VDD.n9486 VDD.n9483 9.3005
R12574 VDD.n9819 VDD.n9818 9.3005
R12575 VDD.n9821 VDD.n9479 9.3005
R12576 VDD.n9854 VDD.n9853 9.3005
R12577 VDD.n9865 VDD.n9864 9.3005
R12578 VDD.n9862 VDD.n9861 9.3005
R12579 VDD.n9859 VDD.n9858 9.3005
R12580 VDD.n9852 VDD.n9851 9.3005
R12581 VDD.n10678 VDD.n10677 9.3005
R12582 VDD.n10892 VDD.n10891 9.3005
R12583 VDD.n10889 VDD.n10672 9.3005
R12584 VDD.n10887 VDD.n10886 9.3005
R12585 VDD.n10881 VDD.n10880 9.3005
R12586 VDD.n10813 VDD.n10803 9.3005
R12587 VDD.n10815 VDD.n10814 9.3005
R12588 VDD.n10812 VDD.n10805 9.3005
R12589 VDD.n10812 VDD.n10811 9.3005
R12590 VDD.n10799 VDD.n10787 9.3005
R12591 VDD.n10798 VDD.n10797 9.3005
R12592 VDD.n10796 VDD.n10789 9.3005
R12593 VDD.n10789 VDD.n10788 9.3005
R12594 VDD.n10821 VDD.n10786 9.3005
R12595 VDD.n10826 VDD.n10785 9.3005
R12596 VDD.n10831 VDD.n10784 9.3005
R12597 VDD.n10836 VDD.n10783 9.3005
R12598 VDD.n10841 VDD.n10782 9.3005
R12599 VDD.n10846 VDD.n10781 9.3005
R12600 VDD.n10851 VDD.n10780 9.3005
R12601 VDD.n10856 VDD.n10779 9.3005
R12602 VDD.n10861 VDD.n10778 9.3005
R12603 VDD.n10863 VDD.n10862 9.3005
R12604 VDD.n10860 VDD.n10859 9.3005
R12605 VDD.n10858 VDD.n10857 9.3005
R12606 VDD.n10855 VDD.n10854 9.3005
R12607 VDD.n10853 VDD.n10852 9.3005
R12608 VDD.n10850 VDD.n10849 9.3005
R12609 VDD.n10848 VDD.n10847 9.3005
R12610 VDD.n10845 VDD.n10844 9.3005
R12611 VDD.n10843 VDD.n10842 9.3005
R12612 VDD.n10840 VDD.n10839 9.3005
R12613 VDD.n10838 VDD.n10837 9.3005
R12614 VDD.n10835 VDD.n10834 9.3005
R12615 VDD.n10833 VDD.n10832 9.3005
R12616 VDD.n10830 VDD.n10829 9.3005
R12617 VDD.n10828 VDD.n10827 9.3005
R12618 VDD.n10825 VDD.n10824 9.3005
R12619 VDD.n10823 VDD.n10822 9.3005
R12620 VDD.n10820 VDD.n10819 9.3005
R12621 VDD.n10876 VDD.n10875 9.3005
R12622 VDD.n10872 VDD.n10871 9.3005
R12623 VDD.n10869 VDD.n10868 9.3005
R12624 VDD.n10865 VDD.n10776 9.3005
R12625 VDD.n10771 VDD.n10693 9.3005
R12626 VDD.n10750 VDD.n10713 9.3005
R12627 VDD.n10742 VDD.n10723 9.3005
R12628 VDD.n10730 VDD.n10728 9.3005
R12629 VDD.n10735 VDD.n10734 9.3005
R12630 VDD.n10736 VDD.n10735 9.3005
R12631 VDD.n10727 VDD.n10724 9.3005
R12632 VDD.n10741 VDD.n10740 9.3005
R12633 VDD.n10740 VDD.n10722 9.3005
R12634 VDD.n10744 VDD.n10743 9.3005
R12635 VDD.n10749 VDD.n10716 9.3005
R12636 VDD.n10749 VDD.n10748 9.3005
R12637 VDD.n10752 VDD.n10751 9.3005
R12638 VDD.n10704 VDD.n10703 9.3005
R12639 VDD.n10761 VDD.n10760 9.3005
R12640 VDD.n10762 VDD.n10761 9.3005
R12641 VDD.n10754 VDD.n10711 9.3005
R12642 VDD.n10718 VDD.n10711 9.3005
R12643 VDD.n10758 VDD.n10757 9.3005
R12644 VDD.n10767 VDD.n10766 9.3005
R12645 VDD.n8781 VDD.n8778 9.3005
R12646 VDD.n9037 VDD.n9034 9.3005
R12647 VDD.n9036 VDD.n9035 9.3005
R12648 VDD.n9039 VDD.n9038 9.3005
R12649 VDD.n9045 VDD.n9044 9.3005
R12650 VDD.n8842 VDD.n8838 9.3005
R12651 VDD.n8847 VDD.n8837 9.3005
R12652 VDD.n8852 VDD.n8836 9.3005
R12653 VDD.n8854 VDD.n8853 9.3005
R12654 VDD.n8851 VDD.n8850 9.3005
R12655 VDD.n8849 VDD.n8848 9.3005
R12656 VDD.n8846 VDD.n8845 9.3005
R12657 VDD.n8844 VDD.n8843 9.3005
R12658 VDD.n8841 VDD.n8840 9.3005
R12659 VDD.n8805 VDD.n8804 9.3005
R12660 VDD.n8816 VDD.n8814 9.3005
R12661 VDD.n8815 VDD.n8810 9.3005
R12662 VDD.n8818 VDD.n8817 9.3005
R12663 VDD.n8807 VDD.n8806 9.3005
R12664 VDD.n9027 VDD.n8825 9.3005
R12665 VDD.n9026 VDD.n9025 9.3005
R12666 VDD.n9017 VDD.n8827 9.3005
R12667 VDD.n9024 VDD.n9023 9.3005
R12668 VDD.n9019 VDD.n9018 9.3005
R12669 VDD.n9016 VDD.n9015 9.3005
R12670 VDD.n9021 VDD.n9020 9.3005
R12671 VDD.n9022 VDD.n8826 9.3005
R12672 VDD.n9029 VDD.n9028 9.3005
R12673 VDD.n8981 VDD.n8980 9.3005
R12674 VDD.n8994 VDD.n8993 9.3005
R12675 VDD.n8979 VDD.n8835 9.3005
R12676 VDD.n8982 VDD.n8831 9.3005
R12677 VDD.n8982 VDD.n8834 9.3005
R12678 VDD.n8992 VDD.n8830 9.3005
R12679 VDD.n8830 VDD.n8829 9.3005
R12680 VDD.n8995 VDD.n8828 9.3005
R12681 VDD.n9009 VDD.n8999 9.3005
R12682 VDD.n9011 VDD.n9010 9.3005
R12683 VDD.n9008 VDD.n9001 9.3005
R12684 VDD.n9008 VDD.n9007 9.3005
R12685 VDD.n8973 VDD.n8856 9.3005
R12686 VDD.n8956 VDD.n8862 9.3005
R12687 VDD.n8875 VDD.n8863 9.3005
R12688 VDD.n8874 VDD.n8873 9.3005
R12689 VDD.n8872 VDD.n8865 9.3005
R12690 VDD.n8865 VDD.n8864 9.3005
R12691 VDD.n8958 VDD.n8957 9.3005
R12692 VDD.n8959 VDD.n8859 9.3005
R12693 VDD.n8959 VDD.n8861 9.3005
R12694 VDD.n8972 VDD.n8971 9.3005
R12695 VDD.n8970 VDD.n8858 9.3005
R12696 VDD.n8858 VDD.n8857 9.3005
R12697 VDD.n8949 VDD.n8879 9.3005
R12698 VDD.n8944 VDD.n8881 9.3005
R12699 VDD.n8939 VDD.n8883 9.3005
R12700 VDD.n8951 VDD.n8950 9.3005
R12701 VDD.n8948 VDD.n8947 9.3005
R12702 VDD.n8946 VDD.n8945 9.3005
R12703 VDD.n8943 VDD.n8942 9.3005
R12704 VDD.n8941 VDD.n8940 9.3005
R12705 VDD.n8938 VDD.n8937 9.3005
R12706 VDD.n8918 VDD.n8917 9.3005
R12707 VDD.n8916 VDD.n8770 9.3005
R12708 VDD.n8925 VDD.n8924 9.3005
R12709 VDD.n8923 VDD.n8922 9.3005
R12710 VDD.n8920 VDD.n8919 9.3005
R12711 VDD.n8892 VDD.n8889 9.3005
R12712 VDD.n8896 VDD.n8895 9.3005
R12713 VDD.n8912 VDD.n8890 9.3005
R12714 VDD.n8912 VDD.n8911 9.3005
R12715 VDD.n8899 VDD.n8897 9.3005
R12716 VDD.n8901 VDD.n8900 9.3005
R12717 VDD.n8764 VDD.n8762 9.3005
R12718 VDD.n9063 VDD.n9062 9.3005
R12719 VDD.n9062 VDD.n9061 9.3005
R12720 VDD.n8906 VDD.n8898 9.3005
R12721 VDD.n8906 VDD.n8905 9.3005
R12722 VDD.n9285 VDD.n9284 9.3005
R12723 VDD.n9283 VDD.n9276 9.3005
R12724 VDD.n9276 VDD.n9275 9.3005
R12725 VDD.n9286 VDD.n9274 9.3005
R12726 VDD.n9272 VDD.n9267 9.3005
R12727 VDD.n9301 VDD.n9300 9.3005
R12728 VDD.n9292 VDD.n9273 9.3005
R12729 VDD.n9299 VDD.n9266 9.3005
R12730 VDD.n9294 VDD.n9293 9.3005
R12731 VDD.n9291 VDD.n9290 9.3005
R12732 VDD.n9296 VDD.n9295 9.3005
R12733 VDD.n9298 VDD.n9297 9.3005
R12734 VDD.n9271 VDD.n9270 9.3005
R12735 VDD.n9314 VDD.n9256 9.3005
R12736 VDD.n9306 VDD.n9303 9.3005
R12737 VDD.n9305 VDD.n9304 9.3005
R12738 VDD.n9308 VDD.n9307 9.3005
R12739 VDD.n9316 VDD.n9315 9.3005
R12740 VDD.n9334 VDD.n9330 9.3005
R12741 VDD.n9333 VDD.n9332 9.3005
R12742 VDD.n9339 VDD.n9338 9.3005
R12743 VDD.n9329 VDD.n9327 9.3005
R12744 VDD.n9336 VDD.n9335 9.3005
R12745 VDD.n9371 VDD.n9366 9.3005
R12746 VDD.n9373 VDD.n9372 9.3005
R12747 VDD.n9374 VDD.n9373 9.3005
R12748 VDD.n9370 VDD.n9363 9.3005
R12749 VDD.n9415 VDD.n9414 9.3005
R12750 VDD.n9413 VDD.n9406 9.3005
R12751 VDD.n9406 VDD.n9405 9.3005
R12752 VDD.n9416 VDD.n9404 9.3005
R12753 VDD.n9402 VDD.n9399 9.3005
R12754 VDD.n9428 VDD.n9427 9.3005
R12755 VDD.n9436 VDD.n9393 9.3005
R12756 VDD.n9435 VDD.n9434 9.3005
R12757 VDD.n9429 VDD.n9395 9.3005
R12758 VDD.n9430 VDD.n9429 9.3005
R12759 VDD.n9426 VDD.n9398 9.3005
R12760 VDD.n9425 VDD.n9424 9.3005
R12761 VDD.n9424 VDD.n9423 9.3005
R12762 VDD.n9421 VDD.n9420 9.3005
R12763 VDD.n9438 VDD.n9437 9.3005
R12764 VDD.n9438 VDD.n9392 9.3005
R12765 VDD.n9359 VDD.n9358 9.3005
R12766 VDD.n9381 VDD.n9380 9.3005
R12767 VDD.n9383 VDD.n9382 9.3005
R12768 VDD.n9384 VDD.n9383 9.3005
R12769 VDD.n9379 VDD.n9354 9.3005
R12770 VDD.n9390 VDD.n9389 9.3005
R12771 VDD.n9391 VDD.n9390 9.3005
R12772 VDD.n9218 VDD.n9205 9.3005
R12773 VDD.n9217 VDD.n9205 9.3005
R12774 VDD.n9209 VDD.n9205 9.3005
R12775 VDD.n10996 VDD.n8729 9.3005
R12776 VDD.n11025 VDD.n8721 9.3005
R12777 VDD.n8731 VDD.n8721 9.3005
R12778 VDD.n8728 VDD.n8721 9.3005
R12779 VDD.n9154 VDD.n9084 9.3005
R12780 VDD.n9159 VDD.n9158 9.3005
R12781 VDD.n9102 VDD.n9101 9.3005
R12782 VDD.n9099 VDD.n9088 9.3005
R12783 VDD.n9141 VDD.n9140 9.3005
R12784 VDD.n9139 VDD.n9106 9.3005
R12785 VDD.n9130 VDD.n9109 9.3005
R12786 VDD.n9132 VDD.n9131 9.3005
R12787 VDD.n9129 VDD.n9128 9.3005
R12788 VDD.n9120 VDD.n9119 9.3005
R12789 VDD.n9117 VDD.n9113 9.3005
R12790 VDD.n9116 VDD.n9115 9.3005
R12791 VDD.n9094 VDD.n9093 9.3005
R12792 VDD.n9156 VDD.n9155 9.3005
R12793 VDD.n10448 VDD.n6920 9.3005
R12794 VDD.n10481 VDD.n6920 9.3005
R12795 VDD.n10492 VDD.n10491 9.3005
R12796 VDD.n10478 VDD.n6920 9.3005
R12797 VDD.n12448 VDD.n12440 9.3005
R12798 VDD.n12443 VDD.n12442 9.3005
R12799 VDD.n12424 VDD.n6907 9.3005
R12800 VDD.n12486 VDD.n12485 9.3005
R12801 VDD.n12492 VDD.n6911 9.3005
R12802 VDD.n12492 VDD.n12491 9.3005
R12803 VDD.n12493 VDD.n6908 9.3005
R12804 VDD.n12495 VDD.n12494 9.3005
R12805 VDD.n12441 VDD.n12437 9.3005
R12806 VDD.n12464 VDD.n12437 9.3005
R12807 VDD.n12444 VDD.n12439 9.3005
R12808 VDD.n12459 VDD.n12445 9.3005
R12809 VDD.n12459 VDD.n12458 9.3005
R12810 VDD.n12449 VDD.n12447 9.3005
R12811 VDD.n12452 VDD.n12451 9.3005
R12812 VDD.n12452 VDD.n12426 9.3005
R12813 VDD.n12483 VDD.n12427 9.3005
R12814 VDD.n12470 VDD.n12469 9.3005
R12815 VDD.n12478 VDD.n12477 9.3005
R12816 VDD.n10212 VDD.t148 9.29365
R12817 VDD.n9049 VDD.n8786 9.1381
R12818 VDD.n9033 VDD.n8793 9.1381
R12819 VDD.n8933 VDD.n8921 9.1381
R12820 VDD.n9311 VDD.n9259 9.1381
R12821 VDD.n10924 VDD.n9337 9.1381
R12822 VDD.n9049 VDD.n8785 9.12656
R12823 VDD.n9033 VDD.n8792 9.12656
R12824 VDD.n8933 VDD.n8926 9.12656
R12825 VDD.n9311 VDD.n9257 9.12656
R12826 VDD.n10925 VDD.n10924 9.12656
R12827 VDD.n9049 VDD.n8783 9.11505
R12828 VDD.n9033 VDD.n8791 9.11505
R12829 VDD.n8933 VDD.n8884 9.11505
R12830 VDD.n9311 VDD.n9260 9.11505
R12831 VDD.n10432 VDD.n6919 9.01711
R12832 VDD.n11218 VDD.n6622 8.99396
R12833 VDD.n6387 VDD.n5900 8.9605
R12834 VDD.n6257 VDD.n6256 8.9605
R12835 VDD.n5533 VDD.n5046 8.9605
R12836 VDD.n5403 VDD.n5402 8.9605
R12837 VDD.n4747 VDD.n4260 8.9605
R12838 VDD.n4617 VDD.n4616 8.9605
R12839 VDD.n3893 VDD.n3406 8.9605
R12840 VDD.n3763 VDD.n3762 8.9605
R12841 VDD.n3107 VDD.n2620 8.9605
R12842 VDD.n2977 VDD.n2976 8.9605
R12843 VDD.n2252 VDD.n1765 8.9605
R12844 VDD.n2122 VDD.n2121 8.9605
R12845 VDD.n1369 VDD.n1268 8.9605
R12846 VDD.n981 VDD.n878 8.9605
R12847 VDD.n141 VDD.n40 8.9605
R12848 VDD.n535 VDD.n432 8.9605
R12849 VDD.n12490 VDD.n12489 8.9077
R12850 VDD.n12457 VDD.n12438 8.9077
R12851 VDD.n9739 VDD.n9642 8.90247
R12852 VDD.n9739 VDD.n9640 8.90247
R12853 VDD.n10878 VDD.n10688 8.90247
R12854 VDD.n10878 VDD.n10686 8.90247
R12855 VDD.n9739 VDD.n9643 8.89163
R12856 VDD.n9739 VDD.n9639 8.89163
R12857 VDD.n10878 VDD.n10689 8.89163
R12858 VDD.n10878 VDD.n10685 8.89163
R12859 VDD.n9739 VDD.n9638 8.88085
R12860 VDD.n9740 VDD.n9739 8.88085
R12861 VDD.n10878 VDD.n10684 8.88085
R12862 VDD.n10878 VDD.n10681 8.88085
R12863 VDD.n9739 VDD.n9559 8.87012
R12864 VDD.n9739 VDD.n9637 8.87012
R12865 VDD.n9763 VDD.n9547 8.87012
R12866 VDD.n9530 VDD.n9523 8.87012
R12867 VDD.n9784 VDD.n9517 8.87012
R12868 VDD.n9810 VDD.n9503 8.87012
R12869 VDD.n9487 VDD.n9480 8.87012
R12870 VDD.n9863 VDD.n9856 8.87012
R12871 VDD.n10890 VDD.n10883 8.87012
R12872 VDD.n10878 VDD.n10691 8.87012
R12873 VDD.n10878 VDD.n10683 8.87012
R12874 VDD.n9049 VDD.n8784 8.87012
R12875 VDD.n9033 VDD.n8798 8.87012
R12876 VDD.n8933 VDD.n8882 8.87012
R12877 VDD.n9311 VDD.n9302 8.87012
R12878 VDD.n9739 VDD.n9738 8.85944
R12879 VDD.n9739 VDD.n9636 8.85944
R12880 VDD.n9763 VDD.n9762 8.85944
R12881 VDD.n9773 VDD.n9523 8.85944
R12882 VDD.n9784 VDD.n9783 8.85944
R12883 VDD.n9810 VDD.n9809 8.85944
R12884 VDD.n9820 VDD.n9480 8.85944
R12885 VDD.n9856 VDD.n9855 8.85944
R12886 VDD.n10883 VDD.n10882 8.85944
R12887 VDD.n10878 VDD.n10877 8.85944
R12888 VDD.n10878 VDD.n10682 8.85944
R12889 VDD.n9049 VDD.n8789 8.85944
R12890 VDD.n9033 VDD.n8796 8.85944
R12891 VDD.n8933 VDD.n8880 8.85944
R12892 VDD.n9311 VDD.n9264 8.85944
R12893 VDD.n9959 VDD.n9909 8.85536
R12894 VDD.n9965 VDD.n9908 8.85536
R12895 VDD.n9967 VDD.n9966 8.85536
R12896 VDD.n9961 VDD.n9960 8.85536
R12897 VDD.n9945 VDD.n9944 8.85536
R12898 VDD.n9943 VDD.n9915 8.85536
R12899 VDD.n9920 VDD.n9917 8.85536
R12900 VDD.n9939 VDD.n9938 8.85536
R12901 VDD.n9921 VDD.n9919 8.85536
R12902 VDD.n9933 VDD.n9932 8.85536
R12903 VDD.n5744 VDD.n5743 8.85536
R12904 VDD.n5761 VDD.n5760 8.85536
R12905 VDD.n5759 VDD.n5742 8.85536
R12906 VDD.n5748 VDD.n5747 8.85536
R12907 VDD.n5725 VDD.n5724 8.85536
R12908 VDD.n5717 VDD.n5716 8.85536
R12909 VDD.n5716 VDD.n5715 8.85536
R12910 VDD.n5737 VDD.n5736 8.85536
R12911 VDD.n5738 VDD.n5737 8.85536
R12912 VDD.n5714 VDD.n5713 8.85536
R12913 VDD.n5739 VDD.n5714 8.85536
R12914 VDD.n5767 VDD.n5766 8.85536
R12915 VDD.n5766 VDD.n5765 8.85536
R12916 VDD.n4104 VDD.n4103 8.85536
R12917 VDD.n4121 VDD.n4120 8.85536
R12918 VDD.n4119 VDD.n4102 8.85536
R12919 VDD.n4108 VDD.n4107 8.85536
R12920 VDD.n4085 VDD.n4084 8.85536
R12921 VDD.n4077 VDD.n4076 8.85536
R12922 VDD.n4076 VDD.n4075 8.85536
R12923 VDD.n4097 VDD.n4096 8.85536
R12924 VDD.n4098 VDD.n4097 8.85536
R12925 VDD.n4074 VDD.n4073 8.85536
R12926 VDD.n4099 VDD.n4074 8.85536
R12927 VDD.n4127 VDD.n4126 8.85536
R12928 VDD.n4126 VDD.n4125 8.85536
R12929 VDD.n2463 VDD.n2462 8.85536
R12930 VDD.n2481 VDD.n2480 8.85536
R12931 VDD.n2479 VDD.n2461 8.85536
R12932 VDD.n2467 VDD.n2466 8.85536
R12933 VDD.n2444 VDD.n2443 8.85536
R12934 VDD.n2436 VDD.n2435 8.85536
R12935 VDD.n2435 VDD.n2434 8.85536
R12936 VDD.n2456 VDD.n2455 8.85536
R12937 VDD.n2457 VDD.n2456 8.85536
R12938 VDD.n2433 VDD.n2432 8.85536
R12939 VDD.n2458 VDD.n2433 8.85536
R12940 VDD.n2487 VDD.n2486 8.85536
R12941 VDD.n2486 VDD.n2485 8.85536
R12942 VDD.n823 VDD.n822 8.85536
R12943 VDD.n841 VDD.n840 8.85536
R12944 VDD.n839 VDD.n821 8.85536
R12945 VDD.n827 VDD.n826 8.85536
R12946 VDD.n804 VDD.n803 8.85536
R12947 VDD.n796 VDD.n795 8.85536
R12948 VDD.n795 VDD.n794 8.85536
R12949 VDD.n816 VDD.n815 8.85536
R12950 VDD.n817 VDD.n816 8.85536
R12951 VDD.n793 VDD.n792 8.85536
R12952 VDD.n818 VDD.n793 8.85536
R12953 VDD.n847 VDD.n846 8.85536
R12954 VDD.n846 VDD.n845 8.85536
R12955 VDD.n9151 VDD.n9150 8.85412
R12956 VDD.n9739 VDD.n9729 8.84881
R12957 VDD.n10878 VDD.n10690 8.84881
R12958 VDD.n8933 VDD.n8878 8.84881
R12959 VDD.n9049 VDD.n8790 8.84881
R12960 VDD.n9033 VDD.n8797 8.84881
R12961 VDD.n9311 VDD.n9265 8.84881
R12962 VDD.n9150 VDD.n9149 8.84352
R12963 VDD.n9150 VDD.n9090 8.83298
R12964 VDD.n10958 VDD.n9204 8.78757
R12965 VDD.n10493 VDD.n6915 8.77128
R12966 VDD.n12434 VDD.n12426 8.76719
R12967 VDD.n8990 VDD.n8989 8.76429
R12968 VDD.n8968 VDD.n8963 8.76429
R12969 VDD.n5982 VDD.n5981 8.7045
R12970 VDD.n5983 VDD.n5982 8.7045
R12971 VDD.n5986 VDD.n5983 8.7045
R12972 VDD.n6341 VDD.n6340 8.7045
R12973 VDD.n6340 VDD.n6339 8.7045
R12974 VDD.n6339 VDD.n6004 8.7045
R12975 VDD.n6296 VDD.n6004 8.7045
R12976 VDD.n6296 VDD.n6295 8.7045
R12977 VDD.n6551 VDD.n6550 8.7045
R12978 VDD.n6550 VDD.n6549 8.7045
R12979 VDD.n6549 VDD.n5788 8.7045
R12980 VDD.n5128 VDD.n5127 8.7045
R12981 VDD.n5129 VDD.n5128 8.7045
R12982 VDD.n5132 VDD.n5129 8.7045
R12983 VDD.n5487 VDD.n5486 8.7045
R12984 VDD.n5486 VDD.n5485 8.7045
R12985 VDD.n5485 VDD.n5150 8.7045
R12986 VDD.n5442 VDD.n5150 8.7045
R12987 VDD.n5442 VDD.n5441 8.7045
R12988 VDD.n5697 VDD.n5696 8.7045
R12989 VDD.n5696 VDD.n5695 8.7045
R12990 VDD.n5695 VDD.n4934 8.7045
R12991 VDD.n4342 VDD.n4341 8.7045
R12992 VDD.n4343 VDD.n4342 8.7045
R12993 VDD.n4346 VDD.n4343 8.7045
R12994 VDD.n4701 VDD.n4700 8.7045
R12995 VDD.n4700 VDD.n4699 8.7045
R12996 VDD.n4699 VDD.n4364 8.7045
R12997 VDD.n4656 VDD.n4364 8.7045
R12998 VDD.n4656 VDD.n4655 8.7045
R12999 VDD.n4911 VDD.n4910 8.7045
R13000 VDD.n4910 VDD.n4909 8.7045
R13001 VDD.n4909 VDD.n4148 8.7045
R13002 VDD.n3488 VDD.n3487 8.7045
R13003 VDD.n3489 VDD.n3488 8.7045
R13004 VDD.n3492 VDD.n3489 8.7045
R13005 VDD.n3847 VDD.n3846 8.7045
R13006 VDD.n3846 VDD.n3845 8.7045
R13007 VDD.n3845 VDD.n3510 8.7045
R13008 VDD.n3802 VDD.n3510 8.7045
R13009 VDD.n3802 VDD.n3801 8.7045
R13010 VDD.n4057 VDD.n4056 8.7045
R13011 VDD.n4056 VDD.n4055 8.7045
R13012 VDD.n4055 VDD.n3294 8.7045
R13013 VDD.n2702 VDD.n2701 8.7045
R13014 VDD.n2703 VDD.n2702 8.7045
R13015 VDD.n2706 VDD.n2703 8.7045
R13016 VDD.n3061 VDD.n3060 8.7045
R13017 VDD.n3060 VDD.n3059 8.7045
R13018 VDD.n3059 VDD.n2724 8.7045
R13019 VDD.n3016 VDD.n2724 8.7045
R13020 VDD.n3016 VDD.n3015 8.7045
R13021 VDD.n3271 VDD.n3270 8.7045
R13022 VDD.n3270 VDD.n3269 8.7045
R13023 VDD.n3269 VDD.n2508 8.7045
R13024 VDD.n1847 VDD.n1846 8.7045
R13025 VDD.n1848 VDD.n1847 8.7045
R13026 VDD.n1851 VDD.n1848 8.7045
R13027 VDD.n2206 VDD.n2205 8.7045
R13028 VDD.n2205 VDD.n2204 8.7045
R13029 VDD.n2204 VDD.n1869 8.7045
R13030 VDD.n2161 VDD.n1869 8.7045
R13031 VDD.n2161 VDD.n2160 8.7045
R13032 VDD.n2416 VDD.n2415 8.7045
R13033 VDD.n2415 VDD.n2414 8.7045
R13034 VDD.n2414 VDD.n1653 8.7045
R13035 VDD.n1524 VDD.n1522 8.7045
R13036 VDD.n1522 VDD.n1520 8.7045
R13037 VDD.n1520 VDD.n1518 8.7045
R13038 VDD.n1134 VDD.n1132 8.7045
R13039 VDD.n1136 VDD.n1134 8.7045
R13040 VDD.n1138 VDD.n1136 8.7045
R13041 VDD.n1140 VDD.n1138 8.7045
R13042 VDD.n1145 VDD.n1143 8.7045
R13043 VDD.n1147 VDD.n1145 8.7045
R13044 VDD.n1149 VDD.n1147 8.7045
R13045 VDD.n296 VDD.n294 8.7045
R13046 VDD.n294 VDD.n292 8.7045
R13047 VDD.n292 VDD.n290 8.7045
R13048 VDD.n688 VDD.n686 8.7045
R13049 VDD.n690 VDD.n688 8.7045
R13050 VDD.n692 VDD.n690 8.7045
R13051 VDD.n694 VDD.n692 8.7045
R13052 VDD.n699 VDD.n697 8.7045
R13053 VDD.n701 VDD.n699 8.7045
R13054 VDD.n703 VDD.n701 8.7045
R13055 VDD.n9182 VDD.n9174 8.65557
R13056 VDD.n10988 VDD.n8727 8.65557
R13057 VDD.n12429 VDD.n12426 8.59505
R13058 VDD.n6600 VDD.n6580 8.46493
R13059 VDD.n9189 VDD.n9076 8.45089
R13060 VDD.n10958 VDD.n10957 8.45089
R13061 VDD.n10952 VDD.n9222 8.45089
R13062 VDD.n10432 VDD.n10431 8.45089
R13063 VDD.n9185 VDD.n9184 8.45089
R13064 VDD.n9182 VDD.n9181 8.45089
R13065 VDD.n10960 VDD.n9219 8.45089
R13066 VDD.n11000 VDD.n8730 8.45089
R13067 VDD.n10988 VDD.n10987 8.45089
R13068 VDD.n9070 VDD.n8729 8.45089
R13069 VDD.n10493 VDD.n10492 8.45089
R13070 VDD.n10435 VDD.n10422 8.45089
R13071 VDD.n10496 VDD.n10495 8.45089
R13072 VDD.n12490 VDD.n12426 8.42955
R13073 VDD.n12457 VDD.n12426 8.42955
R13074 VDD.n9218 VDD.n9199 8.40959
R13075 VDD.n9217 VDD.n9199 8.40959
R13076 VDD.n9209 VDD.n9199 8.40959
R13077 VDD.n11026 VDD.n11025 8.40959
R13078 VDD.n11026 VDD.n8731 8.40959
R13079 VDD.n11026 VDD.n8728 8.40959
R13080 VDD.n10481 VDD.n6913 8.40959
R13081 VDD.n10448 VDD.n6913 8.40959
R13082 VDD.n10478 VDD.n6913 8.40959
R13083 VDD.n12662 VDD.t184 8.39432
R13084 VDD.n12426 VDD.n12421 8.39432
R13085 VDD.n9965 VDD.n9964 8.39408
R13086 VDD.n9964 VDD.n9909 8.39408
R13087 VDD.n9966 VDD.n9907 8.39408
R13088 VDD.n9962 VDD.n9961 8.39408
R13089 VDD.n9944 VDD.n9916 8.39408
R13090 VDD.n9942 VDD.n9917 8.39408
R13091 VDD.n9940 VDD.n9919 8.39408
R13092 VDD.n9943 VDD.n9942 8.39408
R13093 VDD.n9940 VDD.n9939 8.39408
R13094 VDD.n9932 VDD.n9918 8.39408
R13095 VDD.n5762 VDD.n5742 8.39408
R13096 VDD.n5762 VDD.n5761 8.39408
R13097 VDD.n5747 VDD.n5741 8.39408
R13098 VDD.n4122 VDD.n4102 8.39408
R13099 VDD.n4122 VDD.n4121 8.39408
R13100 VDD.n4107 VDD.n4101 8.39408
R13101 VDD.n2482 VDD.n2461 8.39408
R13102 VDD.n2482 VDD.n2481 8.39408
R13103 VDD.n2466 VDD.n2460 8.39408
R13104 VDD.n842 VDD.n821 8.39408
R13105 VDD.n842 VDD.n841 8.39408
R13106 VDD.n826 VDD.n820 8.39408
R13107 VDD.n5743 VDD.n5740 8.39405
R13108 VDD.n4103 VDD.n4100 8.39405
R13109 VDD.n2462 VDD.n2459 8.39405
R13110 VDD.n822 VDD.n819 8.39405
R13111 VDD.n12426 VDD.n12425 8.2703
R13112 VDD.n10244 VDD.t184 8.09454
R13113 VDD.n9161 VDD.n9082 8.08763
R13114 VDD.n10973 VDD.n10972 8.07007
R13115 VDD.n8499 VDD.n7747 8.06816
R13116 VDD.n7728 VDD.n7719 8.06816
R13117 VDD.n11441 VDD.n7729 8.06816
R13118 VDD.n11426 VDD.n8616 8.06816
R13119 VDD.n11425 VDD.n8617 8.06816
R13120 VDD.n11422 VDD.n8623 8.06816
R13121 VDD.n8629 VDD.n8628 8.06816
R13122 VDD.n11416 VDD.n8630 8.06816
R13123 VDD.n11406 VDD.n8648 8.06816
R13124 VDD.n11403 VDD.n8654 8.06816
R13125 VDD.n11397 VDD.n8660 8.06816
R13126 VDD.n11391 VDD.n8668 8.06816
R13127 VDD.n11390 VDD.n8669 8.06816
R13128 VDD.n11382 VDD.n8685 8.06816
R13129 VDD.n11381 VDD.n8686 8.06816
R13130 VDD.n11378 VDD.n8692 8.06816
R13131 VDD.n8701 VDD.n8700 8.06816
R13132 VDD.n11372 VDD.n8702 8.06816
R13133 VDD.n11359 VDD.n11028 8.06816
R13134 VDD.n11034 VDD.n11033 8.06816
R13135 VDD.n11353 VDD.n11035 8.06816
R13136 VDD.n11344 VDD.n11052 8.06816
R13137 VDD.n11343 VDD.n11053 8.06816
R13138 VDD.n11095 VDD.n11063 8.06816
R13139 VDD.n11334 VDD.n11064 8.06816
R13140 VDD.n11075 VDD.n11074 8.06816
R13141 VDD.n11325 VDD.n11076 8.06816
R13142 VDD.n11081 VDD.n11080 8.06816
R13143 VDD.n11319 VDD.n11082 8.06816
R13144 VDD.n11310 VDD.n11105 8.06816
R13145 VDD.n11309 VDD.n11106 8.06816
R13146 VDD.n11306 VDD.n11112 8.06816
R13147 VDD.n11118 VDD.n11117 8.06816
R13148 VDD.n11300 VDD.n11119 8.06816
R13149 VDD.n11291 VDD.n11136 8.06816
R13150 VDD.n11287 VDD.n11143 8.06816
R13151 VDD.n11149 VDD.n11148 8.06816
R13152 VDD.n11281 VDD.n11150 8.06816
R13153 VDD.n11272 VDD.n11167 8.06816
R13154 VDD.n11271 VDD.n11168 8.06816
R13155 VDD.n11268 VDD.n11174 8.06816
R13156 VDD.n11262 VDD.n11181 8.06816
R13157 VDD.n11256 VDD.n11189 8.06816
R13158 VDD.n11255 VDD.n11190 8.06816
R13159 VDD.n11247 VDD.n11206 8.06816
R13160 VDD.n11246 VDD.n11207 8.06816
R13161 VDD.n11243 VDD.n11213 8.06816
R13162 VDD.n11214 VDD.n6599 8.06816
R13163 VDD.n12710 VDD.n6600 8.06816
R13164 VDD.n9926 VDD.n9923 7.96135
R13165 VDD.n9116 VDD.n9091 7.52991
R13166 VDD.n9650 VDD.n9649 7.45411
R13167 VDD.n9667 VDD.n9666 7.45411
R13168 VDD.n10793 VDD.n10792 7.45411
R13169 VDD.n10810 VDD.n10809 7.45411
R13170 VDD.n8869 VDD.n8868 7.45411
R13171 VDD.n8962 VDD.n8961 7.45411
R13172 VDD.n8966 VDD.n8965 7.45411
R13173 VDD.n9006 VDD.n9005 7.45411
R13174 VDD.n8985 VDD.n8984 7.45411
R13175 VDD.n8988 VDD.n8987 7.45411
R13176 VDD.n9280 VDD.n9279 7.45411
R13177 VDD.n9410 VDD.n9409 7.45411
R13178 VDD.n9838 VDD.n9837 7.33876
R13179 VDD.n10879 VDD.n10680 7.33876
R13180 VDD.n6011 VDD.n6010 7.09014
R13181 VDD.n6015 VDD.n6014 7.09014
R13182 VDD.n5157 VDD.n5156 7.09014
R13183 VDD.n5161 VDD.n5160 7.09014
R13184 VDD.n4371 VDD.n4370 7.09014
R13185 VDD.n4375 VDD.n4374 7.09014
R13186 VDD.n3517 VDD.n3516 7.09014
R13187 VDD.n3521 VDD.n3520 7.09014
R13188 VDD.n2731 VDD.n2730 7.09014
R13189 VDD.n2735 VDD.n2734 7.09014
R13190 VDD.n1876 VDD.n1875 7.09014
R13191 VDD.n1880 VDD.n1879 7.09014
R13192 VDD.n1230 VDD.n1229 7.09014
R13193 VDD.n1637 VDD.n1228 7.09014
R13194 VDD.n2 VDD.n1 7.09014
R13195 VDD.n409 VDD.n0 7.09014
R13196 VDD.n6163 VDD.n6099 7.07692
R13197 VDD.n6164 VDD.n6163 7.07692
R13198 VDD.n6165 VDD.n6164 7.07692
R13199 VDD.n6165 VDD.n6095 7.07692
R13200 VDD.n6171 VDD.n6095 7.07692
R13201 VDD.n6172 VDD.n6171 7.07692
R13202 VDD.n6173 VDD.n6172 7.07692
R13203 VDD.n6173 VDD.n6091 7.07692
R13204 VDD.n6179 VDD.n6091 7.07692
R13205 VDD.n6180 VDD.n6179 7.07692
R13206 VDD.n6181 VDD.n6180 7.07692
R13207 VDD.n6181 VDD.n6087 7.07692
R13208 VDD.n6187 VDD.n6087 7.07692
R13209 VDD.n6188 VDD.n6187 7.07692
R13210 VDD.n6189 VDD.n6188 7.07692
R13211 VDD.n6189 VDD.n6083 7.07692
R13212 VDD.n6195 VDD.n6083 7.07692
R13213 VDD.n6196 VDD.n6195 7.07692
R13214 VDD.n6197 VDD.n6196 7.07692
R13215 VDD.n6197 VDD.n6079 7.07692
R13216 VDD.n6203 VDD.n6079 7.07692
R13217 VDD.n6204 VDD.n6203 7.07692
R13218 VDD.n6206 VDD.n6204 7.07692
R13219 VDD.n6206 VDD.n6205 7.07692
R13220 VDD.n6205 VDD.n6076 7.07692
R13221 VDD.n5309 VDD.n5245 7.07692
R13222 VDD.n5310 VDD.n5309 7.07692
R13223 VDD.n5311 VDD.n5310 7.07692
R13224 VDD.n5311 VDD.n5241 7.07692
R13225 VDD.n5317 VDD.n5241 7.07692
R13226 VDD.n5318 VDD.n5317 7.07692
R13227 VDD.n5319 VDD.n5318 7.07692
R13228 VDD.n5319 VDD.n5237 7.07692
R13229 VDD.n5325 VDD.n5237 7.07692
R13230 VDD.n5326 VDD.n5325 7.07692
R13231 VDD.n5327 VDD.n5326 7.07692
R13232 VDD.n5327 VDD.n5233 7.07692
R13233 VDD.n5333 VDD.n5233 7.07692
R13234 VDD.n5334 VDD.n5333 7.07692
R13235 VDD.n5335 VDD.n5334 7.07692
R13236 VDD.n5335 VDD.n5229 7.07692
R13237 VDD.n5341 VDD.n5229 7.07692
R13238 VDD.n5342 VDD.n5341 7.07692
R13239 VDD.n5343 VDD.n5342 7.07692
R13240 VDD.n5343 VDD.n5225 7.07692
R13241 VDD.n5349 VDD.n5225 7.07692
R13242 VDD.n5350 VDD.n5349 7.07692
R13243 VDD.n5352 VDD.n5350 7.07692
R13244 VDD.n5352 VDD.n5351 7.07692
R13245 VDD.n5351 VDD.n5222 7.07692
R13246 VDD.n4523 VDD.n4459 7.07692
R13247 VDD.n4524 VDD.n4523 7.07692
R13248 VDD.n4525 VDD.n4524 7.07692
R13249 VDD.n4525 VDD.n4455 7.07692
R13250 VDD.n4531 VDD.n4455 7.07692
R13251 VDD.n4532 VDD.n4531 7.07692
R13252 VDD.n4533 VDD.n4532 7.07692
R13253 VDD.n4533 VDD.n4451 7.07692
R13254 VDD.n4539 VDD.n4451 7.07692
R13255 VDD.n4540 VDD.n4539 7.07692
R13256 VDD.n4541 VDD.n4540 7.07692
R13257 VDD.n4541 VDD.n4447 7.07692
R13258 VDD.n4547 VDD.n4447 7.07692
R13259 VDD.n4548 VDD.n4547 7.07692
R13260 VDD.n4549 VDD.n4548 7.07692
R13261 VDD.n4549 VDD.n4443 7.07692
R13262 VDD.n4555 VDD.n4443 7.07692
R13263 VDD.n4556 VDD.n4555 7.07692
R13264 VDD.n4557 VDD.n4556 7.07692
R13265 VDD.n4557 VDD.n4439 7.07692
R13266 VDD.n4563 VDD.n4439 7.07692
R13267 VDD.n4564 VDD.n4563 7.07692
R13268 VDD.n4566 VDD.n4564 7.07692
R13269 VDD.n4566 VDD.n4565 7.07692
R13270 VDD.n4565 VDD.n4436 7.07692
R13271 VDD.n3669 VDD.n3605 7.07692
R13272 VDD.n3670 VDD.n3669 7.07692
R13273 VDD.n3671 VDD.n3670 7.07692
R13274 VDD.n3671 VDD.n3601 7.07692
R13275 VDD.n3677 VDD.n3601 7.07692
R13276 VDD.n3678 VDD.n3677 7.07692
R13277 VDD.n3679 VDD.n3678 7.07692
R13278 VDD.n3679 VDD.n3597 7.07692
R13279 VDD.n3685 VDD.n3597 7.07692
R13280 VDD.n3686 VDD.n3685 7.07692
R13281 VDD.n3687 VDD.n3686 7.07692
R13282 VDD.n3687 VDD.n3593 7.07692
R13283 VDD.n3693 VDD.n3593 7.07692
R13284 VDD.n3694 VDD.n3693 7.07692
R13285 VDD.n3695 VDD.n3694 7.07692
R13286 VDD.n3695 VDD.n3589 7.07692
R13287 VDD.n3701 VDD.n3589 7.07692
R13288 VDD.n3702 VDD.n3701 7.07692
R13289 VDD.n3703 VDD.n3702 7.07692
R13290 VDD.n3703 VDD.n3585 7.07692
R13291 VDD.n3709 VDD.n3585 7.07692
R13292 VDD.n3710 VDD.n3709 7.07692
R13293 VDD.n3712 VDD.n3710 7.07692
R13294 VDD.n3712 VDD.n3711 7.07692
R13295 VDD.n3711 VDD.n3582 7.07692
R13296 VDD.n2883 VDD.n2819 7.07692
R13297 VDD.n2884 VDD.n2883 7.07692
R13298 VDD.n2885 VDD.n2884 7.07692
R13299 VDD.n2885 VDD.n2815 7.07692
R13300 VDD.n2891 VDD.n2815 7.07692
R13301 VDD.n2892 VDD.n2891 7.07692
R13302 VDD.n2893 VDD.n2892 7.07692
R13303 VDD.n2893 VDD.n2811 7.07692
R13304 VDD.n2899 VDD.n2811 7.07692
R13305 VDD.n2900 VDD.n2899 7.07692
R13306 VDD.n2901 VDD.n2900 7.07692
R13307 VDD.n2901 VDD.n2807 7.07692
R13308 VDD.n2907 VDD.n2807 7.07692
R13309 VDD.n2908 VDD.n2907 7.07692
R13310 VDD.n2909 VDD.n2908 7.07692
R13311 VDD.n2909 VDD.n2803 7.07692
R13312 VDD.n2915 VDD.n2803 7.07692
R13313 VDD.n2916 VDD.n2915 7.07692
R13314 VDD.n2917 VDD.n2916 7.07692
R13315 VDD.n2917 VDD.n2799 7.07692
R13316 VDD.n2923 VDD.n2799 7.07692
R13317 VDD.n2924 VDD.n2923 7.07692
R13318 VDD.n2926 VDD.n2924 7.07692
R13319 VDD.n2926 VDD.n2925 7.07692
R13320 VDD.n2925 VDD.n2796 7.07692
R13321 VDD.n2028 VDD.n1964 7.07692
R13322 VDD.n2029 VDD.n2028 7.07692
R13323 VDD.n2030 VDD.n2029 7.07692
R13324 VDD.n2030 VDD.n1960 7.07692
R13325 VDD.n2036 VDD.n1960 7.07692
R13326 VDD.n2037 VDD.n2036 7.07692
R13327 VDD.n2038 VDD.n2037 7.07692
R13328 VDD.n2038 VDD.n1956 7.07692
R13329 VDD.n2044 VDD.n1956 7.07692
R13330 VDD.n2045 VDD.n2044 7.07692
R13331 VDD.n2046 VDD.n2045 7.07692
R13332 VDD.n2046 VDD.n1952 7.07692
R13333 VDD.n2052 VDD.n1952 7.07692
R13334 VDD.n2053 VDD.n2052 7.07692
R13335 VDD.n2054 VDD.n2053 7.07692
R13336 VDD.n2054 VDD.n1948 7.07692
R13337 VDD.n2060 VDD.n1948 7.07692
R13338 VDD.n2061 VDD.n2060 7.07692
R13339 VDD.n2062 VDD.n2061 7.07692
R13340 VDD.n2062 VDD.n1944 7.07692
R13341 VDD.n2068 VDD.n1944 7.07692
R13342 VDD.n2069 VDD.n2068 7.07692
R13343 VDD.n2071 VDD.n2069 7.07692
R13344 VDD.n2071 VDD.n2070 7.07692
R13345 VDD.n2070 VDD.n1941 7.07692
R13346 VDD.n1304 VDD.n1301 7.07692
R13347 VDD.n1301 VDD.n1298 7.07692
R13348 VDD.n1298 VDD.n1295 7.07692
R13349 VDD.n1295 VDD.n1292 7.07692
R13350 VDD.n1292 VDD.n1289 7.07692
R13351 VDD.n1289 VDD.n1286 7.07692
R13352 VDD.n1286 VDD.n1283 7.07692
R13353 VDD.n1283 VDD.n1280 7.07692
R13354 VDD.n1280 VDD.n1277 7.07692
R13355 VDD.n1277 VDD.n1274 7.07692
R13356 VDD.n1274 VDD.n1271 7.07692
R13357 VDD.n887 VDD.n884 7.07692
R13358 VDD.n890 VDD.n887 7.07692
R13359 VDD.n893 VDD.n890 7.07692
R13360 VDD.n896 VDD.n893 7.07692
R13361 VDD.n899 VDD.n896 7.07692
R13362 VDD.n902 VDD.n899 7.07692
R13363 VDD.n905 VDD.n902 7.07692
R13364 VDD.n908 VDD.n905 7.07692
R13365 VDD.n911 VDD.n908 7.07692
R13366 VDD.n914 VDD.n911 7.07692
R13367 VDD.n917 VDD.n914 7.07692
R13368 VDD.n920 VDD.n917 7.07692
R13369 VDD.n923 VDD.n920 7.07692
R13370 VDD.n76 VDD.n73 7.07692
R13371 VDD.n73 VDD.n70 7.07692
R13372 VDD.n70 VDD.n67 7.07692
R13373 VDD.n67 VDD.n64 7.07692
R13374 VDD.n64 VDD.n61 7.07692
R13375 VDD.n61 VDD.n58 7.07692
R13376 VDD.n58 VDD.n55 7.07692
R13377 VDD.n55 VDD.n52 7.07692
R13378 VDD.n52 VDD.n49 7.07692
R13379 VDD.n49 VDD.n46 7.07692
R13380 VDD.n46 VDD.n43 7.07692
R13381 VDD.n441 VDD.n438 7.07692
R13382 VDD.n444 VDD.n441 7.07692
R13383 VDD.n447 VDD.n444 7.07692
R13384 VDD.n450 VDD.n447 7.07692
R13385 VDD.n453 VDD.n450 7.07692
R13386 VDD.n456 VDD.n453 7.07692
R13387 VDD.n459 VDD.n456 7.07692
R13388 VDD.n462 VDD.n459 7.07692
R13389 VDD.n465 VDD.n462 7.07692
R13390 VDD.n468 VDD.n465 7.07692
R13391 VDD.n471 VDD.n468 7.07692
R13392 VDD.n474 VDD.n471 7.07692
R13393 VDD.n477 VDD.n474 7.07692
R13394 VDD.n6364 VDD.n5905 7.05178
R13395 VDD.n6363 VDD.n5917 7.05178
R13396 VDD.n6356 VDD.n5923 7.05178
R13397 VDD.n5930 VDD.n5924 7.05178
R13398 VDD.n5510 VDD.n5051 7.05178
R13399 VDD.n5509 VDD.n5063 7.05178
R13400 VDD.n5502 VDD.n5069 7.05178
R13401 VDD.n5076 VDD.n5070 7.05178
R13402 VDD.n4724 VDD.n4265 7.05178
R13403 VDD.n4723 VDD.n4277 7.05178
R13404 VDD.n4716 VDD.n4283 7.05178
R13405 VDD.n4290 VDD.n4284 7.05178
R13406 VDD.n3870 VDD.n3411 7.05178
R13407 VDD.n3869 VDD.n3423 7.05178
R13408 VDD.n3862 VDD.n3429 7.05178
R13409 VDD.n3436 VDD.n3430 7.05178
R13410 VDD.n3084 VDD.n2625 7.05178
R13411 VDD.n3083 VDD.n2637 7.05178
R13412 VDD.n3076 VDD.n2643 7.05178
R13413 VDD.n2650 VDD.n2644 7.05178
R13414 VDD.n2229 VDD.n1770 7.05178
R13415 VDD.n2228 VDD.n1782 7.05178
R13416 VDD.n2221 VDD.n1788 7.05178
R13417 VDD.n1795 VDD.n1789 7.05178
R13418 VDD.n10997 VDD.n8730 6.89484
R13419 VDD.n9184 VDD.n9167 6.89484
R13420 VDD.n9170 VDD.n9076 6.89484
R13421 VDD.n10960 VDD.n9202 6.89484
R13422 VDD.n9222 VDD.n9203 6.89484
R13423 VDD.n10422 VDD.n6916 6.89484
R13424 VDD.n10495 VDD.n6917 6.89484
R13425 VDD.n9652 VDD.n9651 6.80334
R13426 VDD.n10795 VDD.n10794 6.80334
R13427 VDD.n8871 VDD.n8870 6.80334
R13428 VDD.n9282 VDD.n9277 6.80105
R13429 VDD.n9412 VDD.n9407 6.80105
R13430 VDD.n9664 VDD.n9663 6.80104
R13431 VDD.n10807 VDD.n10806 6.80104
R13432 VDD.n9003 VDD.n9002 6.80104
R13433 VDD.n6216 VDD.n6214 6.59444
R13434 VDD.n6217 VDD.n6216 6.59444
R13435 VDD.n6218 VDD.n6217 6.59444
R13436 VDD.n6218 VDD.n6069 6.59444
R13437 VDD.n6226 VDD.n6069 6.59444
R13438 VDD.n6227 VDD.n6226 6.59444
R13439 VDD.n6228 VDD.n6227 6.59444
R13440 VDD.n6228 VDD.n6065 6.59444
R13441 VDD.n6234 VDD.n6065 6.59444
R13442 VDD.n6235 VDD.n6234 6.59444
R13443 VDD.n6236 VDD.n6235 6.59444
R13444 VDD.n6236 VDD.n6061 6.59444
R13445 VDD.n6242 VDD.n6061 6.59444
R13446 VDD.n6243 VDD.n6242 6.59444
R13447 VDD.n6245 VDD.n6243 6.59444
R13448 VDD.n6245 VDD.n6244 6.59444
R13449 VDD.n6244 VDD.n6058 6.59444
R13450 VDD.n5362 VDD.n5360 6.59444
R13451 VDD.n5363 VDD.n5362 6.59444
R13452 VDD.n5364 VDD.n5363 6.59444
R13453 VDD.n5364 VDD.n5215 6.59444
R13454 VDD.n5372 VDD.n5215 6.59444
R13455 VDD.n5373 VDD.n5372 6.59444
R13456 VDD.n5374 VDD.n5373 6.59444
R13457 VDD.n5374 VDD.n5211 6.59444
R13458 VDD.n5380 VDD.n5211 6.59444
R13459 VDD.n5381 VDD.n5380 6.59444
R13460 VDD.n5382 VDD.n5381 6.59444
R13461 VDD.n5382 VDD.n5207 6.59444
R13462 VDD.n5388 VDD.n5207 6.59444
R13463 VDD.n5389 VDD.n5388 6.59444
R13464 VDD.n5391 VDD.n5389 6.59444
R13465 VDD.n5391 VDD.n5390 6.59444
R13466 VDD.n5390 VDD.n5204 6.59444
R13467 VDD.n4576 VDD.n4574 6.59444
R13468 VDD.n4577 VDD.n4576 6.59444
R13469 VDD.n4578 VDD.n4577 6.59444
R13470 VDD.n4578 VDD.n4429 6.59444
R13471 VDD.n4586 VDD.n4429 6.59444
R13472 VDD.n4587 VDD.n4586 6.59444
R13473 VDD.n4588 VDD.n4587 6.59444
R13474 VDD.n4588 VDD.n4425 6.59444
R13475 VDD.n4594 VDD.n4425 6.59444
R13476 VDD.n4595 VDD.n4594 6.59444
R13477 VDD.n4596 VDD.n4595 6.59444
R13478 VDD.n4596 VDD.n4421 6.59444
R13479 VDD.n4602 VDD.n4421 6.59444
R13480 VDD.n4603 VDD.n4602 6.59444
R13481 VDD.n4605 VDD.n4603 6.59444
R13482 VDD.n4605 VDD.n4604 6.59444
R13483 VDD.n4604 VDD.n4418 6.59444
R13484 VDD.n3722 VDD.n3720 6.59444
R13485 VDD.n3723 VDD.n3722 6.59444
R13486 VDD.n3724 VDD.n3723 6.59444
R13487 VDD.n3724 VDD.n3575 6.59444
R13488 VDD.n3732 VDD.n3575 6.59444
R13489 VDD.n3733 VDD.n3732 6.59444
R13490 VDD.n3734 VDD.n3733 6.59444
R13491 VDD.n3734 VDD.n3571 6.59444
R13492 VDD.n3740 VDD.n3571 6.59444
R13493 VDD.n3741 VDD.n3740 6.59444
R13494 VDD.n3742 VDD.n3741 6.59444
R13495 VDD.n3742 VDD.n3567 6.59444
R13496 VDD.n3748 VDD.n3567 6.59444
R13497 VDD.n3749 VDD.n3748 6.59444
R13498 VDD.n3751 VDD.n3749 6.59444
R13499 VDD.n3751 VDD.n3750 6.59444
R13500 VDD.n3750 VDD.n3564 6.59444
R13501 VDD.n2936 VDD.n2934 6.59444
R13502 VDD.n2937 VDD.n2936 6.59444
R13503 VDD.n2938 VDD.n2937 6.59444
R13504 VDD.n2938 VDD.n2789 6.59444
R13505 VDD.n2946 VDD.n2789 6.59444
R13506 VDD.n2947 VDD.n2946 6.59444
R13507 VDD.n2948 VDD.n2947 6.59444
R13508 VDD.n2948 VDD.n2785 6.59444
R13509 VDD.n2954 VDD.n2785 6.59444
R13510 VDD.n2955 VDD.n2954 6.59444
R13511 VDD.n2956 VDD.n2955 6.59444
R13512 VDD.n2956 VDD.n2781 6.59444
R13513 VDD.n2962 VDD.n2781 6.59444
R13514 VDD.n2963 VDD.n2962 6.59444
R13515 VDD.n2965 VDD.n2963 6.59444
R13516 VDD.n2965 VDD.n2964 6.59444
R13517 VDD.n2964 VDD.n2778 6.59444
R13518 VDD.n2081 VDD.n2079 6.59444
R13519 VDD.n2082 VDD.n2081 6.59444
R13520 VDD.n2083 VDD.n2082 6.59444
R13521 VDD.n2083 VDD.n1934 6.59444
R13522 VDD.n2091 VDD.n1934 6.59444
R13523 VDD.n2092 VDD.n2091 6.59444
R13524 VDD.n2093 VDD.n2092 6.59444
R13525 VDD.n2093 VDD.n1930 6.59444
R13526 VDD.n2099 VDD.n1930 6.59444
R13527 VDD.n2100 VDD.n2099 6.59444
R13528 VDD.n2101 VDD.n2100 6.59444
R13529 VDD.n2101 VDD.n1926 6.59444
R13530 VDD.n2107 VDD.n1926 6.59444
R13531 VDD.n2108 VDD.n2107 6.59444
R13532 VDD.n2110 VDD.n2108 6.59444
R13533 VDD.n2110 VDD.n2109 6.59444
R13534 VDD.n2109 VDD.n1923 6.59444
R13535 VDD.n929 VDD.n926 6.59444
R13536 VDD.n931 VDD.n929 6.59444
R13537 VDD.n935 VDD.n931 6.59444
R13538 VDD.n938 VDD.n935 6.59444
R13539 VDD.n941 VDD.n938 6.59444
R13540 VDD.n944 VDD.n941 6.59444
R13541 VDD.n947 VDD.n944 6.59444
R13542 VDD.n950 VDD.n947 6.59444
R13543 VDD.n953 VDD.n950 6.59444
R13544 VDD.n956 VDD.n953 6.59444
R13545 VDD.n959 VDD.n956 6.59444
R13546 VDD.n962 VDD.n959 6.59444
R13547 VDD.n965 VDD.n962 6.59444
R13548 VDD.n968 VDD.n965 6.59444
R13549 VDD.n971 VDD.n968 6.59444
R13550 VDD.n974 VDD.n971 6.59444
R13551 VDD.n977 VDD.n974 6.59444
R13552 VDD.n483 VDD.n480 6.59444
R13553 VDD.n485 VDD.n483 6.59444
R13554 VDD.n489 VDD.n485 6.59444
R13555 VDD.n492 VDD.n489 6.59444
R13556 VDD.n495 VDD.n492 6.59444
R13557 VDD.n498 VDD.n495 6.59444
R13558 VDD.n501 VDD.n498 6.59444
R13559 VDD.n504 VDD.n501 6.59444
R13560 VDD.n507 VDD.n504 6.59444
R13561 VDD.n510 VDD.n507 6.59444
R13562 VDD.n513 VDD.n510 6.59444
R13563 VDD.n516 VDD.n513 6.59444
R13564 VDD.n519 VDD.n516 6.59444
R13565 VDD.n522 VDD.n519 6.59444
R13566 VDD.n525 VDD.n522 6.59444
R13567 VDD.n528 VDD.n525 6.59444
R13568 VDD.n531 VDD.n528 6.59444
R13569 VDD.t5 VDD.n11232 6.48108
R13570 VDD.n11290 VDD.t43 6.34882
R13571 VDD.n9787 VDD.n9785 6.31678
R13572 VDD.n9812 VDD.n9811 6.31678
R13573 VDD.n9859 VDD.n9857 6.31678
R13574 VDD.n10887 VDD.n10884 6.31678
R13575 VDD.n9765 VDD.n9764 6.31678
R13576 VDD.n9533 VDD.n9531 6.31678
R13577 VDD.n9490 VDD.n9488 6.31678
R13578 VDD.n9120 VDD.n9089 6.31321
R13579 VDD.n9181 VDD.n9180 6.30775
R13580 VDD.n11024 VDD.n8734 6.30775
R13581 VDD.n12690 VDD.n6702 6.29586
R13582 VDD.n10335 VDD.t27 6.29586
R13583 VDD.n6395 VDD.n6394 6.17355
R13584 VDD.n6396 VDD.n6395 6.17355
R13585 VDD.n6396 VDD.n5873 6.17355
R13586 VDD.n6402 VDD.n5873 6.17355
R13587 VDD.n6403 VDD.n6402 6.17355
R13588 VDD.n6404 VDD.n6403 6.17355
R13589 VDD.n6404 VDD.n5869 6.17355
R13590 VDD.n6410 VDD.n5869 6.17355
R13591 VDD.n6411 VDD.n6410 6.17355
R13592 VDD.n6412 VDD.n6411 6.17355
R13593 VDD.n6412 VDD.n5865 6.17355
R13594 VDD.n6418 VDD.n5865 6.17355
R13595 VDD.n5541 VDD.n5540 6.17355
R13596 VDD.n5542 VDD.n5541 6.17355
R13597 VDD.n5542 VDD.n5019 6.17355
R13598 VDD.n5548 VDD.n5019 6.17355
R13599 VDD.n5549 VDD.n5548 6.17355
R13600 VDD.n5550 VDD.n5549 6.17355
R13601 VDD.n5550 VDD.n5015 6.17355
R13602 VDD.n5556 VDD.n5015 6.17355
R13603 VDD.n5557 VDD.n5556 6.17355
R13604 VDD.n5558 VDD.n5557 6.17355
R13605 VDD.n5558 VDD.n5011 6.17355
R13606 VDD.n5564 VDD.n5011 6.17355
R13607 VDD.n4755 VDD.n4754 6.17355
R13608 VDD.n4756 VDD.n4755 6.17355
R13609 VDD.n4756 VDD.n4233 6.17355
R13610 VDD.n4762 VDD.n4233 6.17355
R13611 VDD.n4763 VDD.n4762 6.17355
R13612 VDD.n4764 VDD.n4763 6.17355
R13613 VDD.n4764 VDD.n4229 6.17355
R13614 VDD.n4770 VDD.n4229 6.17355
R13615 VDD.n4771 VDD.n4770 6.17355
R13616 VDD.n4772 VDD.n4771 6.17355
R13617 VDD.n4772 VDD.n4225 6.17355
R13618 VDD.n4778 VDD.n4225 6.17355
R13619 VDD.n3901 VDD.n3900 6.17355
R13620 VDD.n3902 VDD.n3901 6.17355
R13621 VDD.n3902 VDD.n3379 6.17355
R13622 VDD.n3908 VDD.n3379 6.17355
R13623 VDD.n3909 VDD.n3908 6.17355
R13624 VDD.n3910 VDD.n3909 6.17355
R13625 VDD.n3910 VDD.n3375 6.17355
R13626 VDD.n3916 VDD.n3375 6.17355
R13627 VDD.n3917 VDD.n3916 6.17355
R13628 VDD.n3918 VDD.n3917 6.17355
R13629 VDD.n3918 VDD.n3371 6.17355
R13630 VDD.n3924 VDD.n3371 6.17355
R13631 VDD.n3115 VDD.n3114 6.17355
R13632 VDD.n3116 VDD.n3115 6.17355
R13633 VDD.n3116 VDD.n2593 6.17355
R13634 VDD.n3122 VDD.n2593 6.17355
R13635 VDD.n3123 VDD.n3122 6.17355
R13636 VDD.n3124 VDD.n3123 6.17355
R13637 VDD.n3124 VDD.n2589 6.17355
R13638 VDD.n3130 VDD.n2589 6.17355
R13639 VDD.n3131 VDD.n3130 6.17355
R13640 VDD.n3132 VDD.n3131 6.17355
R13641 VDD.n3132 VDD.n2585 6.17355
R13642 VDD.n3138 VDD.n2585 6.17355
R13643 VDD.n2260 VDD.n2259 6.17355
R13644 VDD.n2261 VDD.n2260 6.17355
R13645 VDD.n2261 VDD.n1738 6.17355
R13646 VDD.n2267 VDD.n1738 6.17355
R13647 VDD.n2268 VDD.n2267 6.17355
R13648 VDD.n2269 VDD.n2268 6.17355
R13649 VDD.n2269 VDD.n1734 6.17355
R13650 VDD.n2275 VDD.n1734 6.17355
R13651 VDD.n2276 VDD.n2275 6.17355
R13652 VDD.n2277 VDD.n2276 6.17355
R13653 VDD.n2277 VDD.n1730 6.17355
R13654 VDD.n2283 VDD.n1730 6.17355
R13655 VDD.n1510 VDD.n1507 6.17355
R13656 VDD.n1507 VDD.n1504 6.17355
R13657 VDD.n1504 VDD.n1501 6.17355
R13658 VDD.n1501 VDD.n1498 6.17355
R13659 VDD.n1498 VDD.n1495 6.17355
R13660 VDD.n1495 VDD.n1492 6.17355
R13661 VDD.n1492 VDD.n1489 6.17355
R13662 VDD.n1489 VDD.n1486 6.17355
R13663 VDD.n1486 VDD.n1483 6.17355
R13664 VDD.n1483 VDD.n1480 6.17355
R13665 VDD.n1480 VDD.n1477 6.17355
R13666 VDD.n1477 VDD.n1474 6.17355
R13667 VDD.n282 VDD.n279 6.17355
R13668 VDD.n279 VDD.n276 6.17355
R13669 VDD.n276 VDD.n273 6.17355
R13670 VDD.n273 VDD.n270 6.17355
R13671 VDD.n270 VDD.n267 6.17355
R13672 VDD.n267 VDD.n264 6.17355
R13673 VDD.n264 VDD.n261 6.17355
R13674 VDD.n261 VDD.n258 6.17355
R13675 VDD.n258 VDD.n255 6.17355
R13676 VDD.n255 VDD.n252 6.17355
R13677 VDD.n252 VDD.n249 6.17355
R13678 VDD.n249 VDD.n246 6.17355
R13679 VDD.n11448 VDD.n11447 6.08431
R13680 VDD.n11645 VDD.n7613 6.06366
R13681 VDD.n10049 VDD.n10048 6.02403
R13682 VDD.n10043 VDD.n10039 6.02403
R13683 VDD.n10608 VDD.n10607 6.02403
R13684 VDD.n10602 VDD.n10598 6.02403
R13685 VDD.n10549 VDD.n10539 6.02403
R13686 VDD.n10544 VDD.n10541 6.02403
R13687 VDD.n9628 VDD.n9566 6.02403
R13688 VDD.n9634 VDD.n9633 6.02403
R13689 VDD.n9696 VDD.n9695 6.02403
R13690 VDD.n9702 VDD.n9701 6.02403
R13691 VDD.n10852 VDD.n10851 6.02403
R13692 VDD.n10846 VDD.n10845 6.02403
R13693 VDD.n10728 VDD.n10727 6.02403
R13694 VDD.n10731 VDD.n10729 6.02403
R13695 VDD.n8914 VDD.n8913 6.02403
R13696 VDD.n8896 VDD.n8889 6.02403
R13697 VDD.n9367 VDD.n9365 6.02403
R13698 VDD.n9366 VDD.n9363 6.02403
R13699 VDD.n12476 VDD.n12475 6.02403
R13700 VDD.n12471 VDD.n12432 6.02403
R13701 VDD.n12130 VDD.n12129 6.00276
R13702 VDD.n12596 VDD.t16 5.99608
R13703 VDD.n7983 VDD.n7982 5.96815
R13704 VDD.n11407 VDD.t75 5.95205
R13705 VDD.n11096 VDD.t34 5.95205
R13706 VDD.n11583 VDD.n11582 5.92892
R13707 VDD.n12465 VDD.n12464 5.89705
R13708 VDD.n12486 VDD.n12484 5.80397
R13709 VDD.n5927 VDD.n5900 5.80317
R13710 VDD.n6354 VDD.n5927 5.80317
R13711 VDD.n6354 VDD.n6353 5.80317
R13712 VDD.n6353 VDD.n6352 5.80317
R13713 VDD.n6352 VDD.n5928 5.80317
R13714 VDD.n6329 VDD.n6042 5.80317
R13715 VDD.n6329 VDD.n6328 5.80317
R13716 VDD.n6328 VDD.n6327 5.80317
R13717 VDD.n6327 VDD.n6043 5.80317
R13718 VDD.n6257 VDD.n6043 5.80317
R13719 VDD.n5073 VDD.n5046 5.80317
R13720 VDD.n5500 VDD.n5073 5.80317
R13721 VDD.n5500 VDD.n5499 5.80317
R13722 VDD.n5499 VDD.n5498 5.80317
R13723 VDD.n5498 VDD.n5074 5.80317
R13724 VDD.n5475 VDD.n5188 5.80317
R13725 VDD.n5475 VDD.n5474 5.80317
R13726 VDD.n5474 VDD.n5473 5.80317
R13727 VDD.n5473 VDD.n5189 5.80317
R13728 VDD.n5403 VDD.n5189 5.80317
R13729 VDD.n4287 VDD.n4260 5.80317
R13730 VDD.n4714 VDD.n4287 5.80317
R13731 VDD.n4714 VDD.n4713 5.80317
R13732 VDD.n4713 VDD.n4712 5.80317
R13733 VDD.n4712 VDD.n4288 5.80317
R13734 VDD.n4689 VDD.n4402 5.80317
R13735 VDD.n4689 VDD.n4688 5.80317
R13736 VDD.n4688 VDD.n4687 5.80317
R13737 VDD.n4687 VDD.n4403 5.80317
R13738 VDD.n4617 VDD.n4403 5.80317
R13739 VDD.n3433 VDD.n3406 5.80317
R13740 VDD.n3860 VDD.n3433 5.80317
R13741 VDD.n3860 VDD.n3859 5.80317
R13742 VDD.n3859 VDD.n3858 5.80317
R13743 VDD.n3858 VDD.n3434 5.80317
R13744 VDD.n3835 VDD.n3548 5.80317
R13745 VDD.n3835 VDD.n3834 5.80317
R13746 VDD.n3834 VDD.n3833 5.80317
R13747 VDD.n3833 VDD.n3549 5.80317
R13748 VDD.n3763 VDD.n3549 5.80317
R13749 VDD.n2647 VDD.n2620 5.80317
R13750 VDD.n3074 VDD.n2647 5.80317
R13751 VDD.n3074 VDD.n3073 5.80317
R13752 VDD.n3073 VDD.n3072 5.80317
R13753 VDD.n3072 VDD.n2648 5.80317
R13754 VDD.n3049 VDD.n2762 5.80317
R13755 VDD.n3049 VDD.n3048 5.80317
R13756 VDD.n3048 VDD.n3047 5.80317
R13757 VDD.n3047 VDD.n2763 5.80317
R13758 VDD.n2977 VDD.n2763 5.80317
R13759 VDD.n1792 VDD.n1765 5.80317
R13760 VDD.n2219 VDD.n1792 5.80317
R13761 VDD.n2219 VDD.n2218 5.80317
R13762 VDD.n2218 VDD.n2217 5.80317
R13763 VDD.n2217 VDD.n1793 5.80317
R13764 VDD.n2194 VDD.n1907 5.80317
R13765 VDD.n2194 VDD.n2193 5.80317
R13766 VDD.n2193 VDD.n2192 5.80317
R13767 VDD.n2192 VDD.n1908 5.80317
R13768 VDD.n2122 VDD.n1908 5.80317
R13769 VDD.n1268 VDD.n1266 5.80317
R13770 VDD.n1266 VDD.n1264 5.80317
R13771 VDD.n1264 VDD.n1262 5.80317
R13772 VDD.n865 VDD.n863 5.80317
R13773 VDD.n870 VDD.n868 5.80317
R13774 VDD.n872 VDD.n870 5.80317
R13775 VDD.n874 VDD.n872 5.80317
R13776 VDD.n876 VDD.n874 5.80317
R13777 VDD.n878 VDD.n876 5.80317
R13778 VDD.n40 VDD.n38 5.80317
R13779 VDD.n38 VDD.n36 5.80317
R13780 VDD.n36 VDD.n34 5.80317
R13781 VDD.n419 VDD.n417 5.80317
R13782 VDD.n424 VDD.n422 5.80317
R13783 VDD.n426 VDD.n424 5.80317
R13784 VDD.n428 VDD.n426 5.80317
R13785 VDD.n430 VDD.n428 5.80317
R13786 VDD.n432 VDD.n430 5.80317
R13787 VDD.n12463 VDD.n12426 5.76535
R13788 VDD.n12479 VDD.n12426 5.76535
R13789 VDD.n9422 VDD.n9419 5.73742
R13790 VDD.n10078 VDD.n10077 5.64756
R13791 VDD.n10111 VDD.n10089 5.64756
R13792 VDD.n10637 VDD.n10139 5.64756
R13793 VDD.n10527 VDD.n10516 5.64756
R13794 VDD.n9648 VDD.n9647 5.64756
R13795 VDD.n9656 VDD.n9655 5.64756
R13796 VDD.n9671 VDD.n9670 5.64756
R13797 VDD.n9665 VDD.n9661 5.64756
R13798 VDD.n10791 VDD.n10790 5.64756
R13799 VDD.n10799 VDD.n10798 5.64756
R13800 VDD.n10814 VDD.n10813 5.64756
R13801 VDD.n10808 VDD.n10804 5.64756
R13802 VDD.n8867 VDD.n8866 5.64756
R13803 VDD.n8875 VDD.n8874 5.64756
R13804 VDD.n8958 VDD.n8862 5.64756
R13805 VDD.n8960 VDD.n8860 5.64756
R13806 VDD.n8967 VDD.n8964 5.64756
R13807 VDD.n8973 VDD.n8972 5.64756
R13808 VDD.n9010 VDD.n9009 5.64756
R13809 VDD.n9004 VDD.n9000 5.64756
R13810 VDD.n8981 VDD.n8835 5.64756
R13811 VDD.n8983 VDD.n8832 5.64756
R13812 VDD.n8986 VDD.n8833 5.64756
R13813 VDD.n8995 VDD.n8994 5.64756
R13814 VDD.n9281 VDD.n9278 5.64756
R13815 VDD.n9286 VDD.n9285 5.64756
R13816 VDD.n9411 VDD.n9408 5.64756
R13817 VDD.n9416 VDD.n9415 5.64756
R13818 VDD.n9117 VDD.n9116 5.64756
R13819 VDD.n9121 VDD.n9120 5.64756
R13820 VDD.n9732 VDD.n9730 5.63005
R13821 VDD.n9549 VDD.n9548 5.63005
R13822 VDD.n9775 VDD.n9774 5.63005
R13823 VDD.n9781 VDD.n9518 5.63005
R13824 VDD.n9505 VDD.n9504 5.63005
R13825 VDD.n9822 VDD.n9821 5.63005
R13826 VDD.n10693 VDD.n10692 5.63005
R13827 VDD.n6518 VDD.n6516 5.61598
R13828 VDD.n6516 VDD.n6515 5.61598
R13829 VDD.n6515 VDD.n5811 5.61598
R13830 VDD.n6509 VDD.n5811 5.61598
R13831 VDD.n6509 VDD.n6508 5.61598
R13832 VDD.n6508 VDD.n6507 5.61598
R13833 VDD.n6507 VDD.n5816 5.61598
R13834 VDD.n6501 VDD.n5816 5.61598
R13835 VDD.n6501 VDD.n6500 5.61598
R13836 VDD.n6500 VDD.n6499 5.61598
R13837 VDD.n6499 VDD.n5820 5.61598
R13838 VDD.n6493 VDD.n5820 5.61598
R13839 VDD.n5664 VDD.n5662 5.61598
R13840 VDD.n5662 VDD.n5661 5.61598
R13841 VDD.n5661 VDD.n4957 5.61598
R13842 VDD.n5655 VDD.n4957 5.61598
R13843 VDD.n5655 VDD.n5654 5.61598
R13844 VDD.n5654 VDD.n5653 5.61598
R13845 VDD.n5653 VDD.n4962 5.61598
R13846 VDD.n5647 VDD.n4962 5.61598
R13847 VDD.n5647 VDD.n5646 5.61598
R13848 VDD.n5646 VDD.n5645 5.61598
R13849 VDD.n5645 VDD.n4966 5.61598
R13850 VDD.n5639 VDD.n4966 5.61598
R13851 VDD.n4878 VDD.n4876 5.61598
R13852 VDD.n4876 VDD.n4875 5.61598
R13853 VDD.n4875 VDD.n4171 5.61598
R13854 VDD.n4869 VDD.n4171 5.61598
R13855 VDD.n4869 VDD.n4868 5.61598
R13856 VDD.n4868 VDD.n4867 5.61598
R13857 VDD.n4867 VDD.n4176 5.61598
R13858 VDD.n4861 VDD.n4176 5.61598
R13859 VDD.n4861 VDD.n4860 5.61598
R13860 VDD.n4860 VDD.n4859 5.61598
R13861 VDD.n4859 VDD.n4180 5.61598
R13862 VDD.n4853 VDD.n4180 5.61598
R13863 VDD.n4024 VDD.n4022 5.61598
R13864 VDD.n4022 VDD.n4021 5.61598
R13865 VDD.n4021 VDD.n3317 5.61598
R13866 VDD.n4015 VDD.n3317 5.61598
R13867 VDD.n4015 VDD.n4014 5.61598
R13868 VDD.n4014 VDD.n4013 5.61598
R13869 VDD.n4013 VDD.n3322 5.61598
R13870 VDD.n4007 VDD.n3322 5.61598
R13871 VDD.n4007 VDD.n4006 5.61598
R13872 VDD.n4006 VDD.n4005 5.61598
R13873 VDD.n4005 VDD.n3326 5.61598
R13874 VDD.n3999 VDD.n3326 5.61598
R13875 VDD.n3238 VDD.n3236 5.61598
R13876 VDD.n3236 VDD.n3235 5.61598
R13877 VDD.n3235 VDD.n2531 5.61598
R13878 VDD.n3229 VDD.n2531 5.61598
R13879 VDD.n3229 VDD.n3228 5.61598
R13880 VDD.n3228 VDD.n3227 5.61598
R13881 VDD.n3227 VDD.n2536 5.61598
R13882 VDD.n3221 VDD.n2536 5.61598
R13883 VDD.n3221 VDD.n3220 5.61598
R13884 VDD.n3220 VDD.n3219 5.61598
R13885 VDD.n3219 VDD.n2540 5.61598
R13886 VDD.n3213 VDD.n2540 5.61598
R13887 VDD.n2383 VDD.n2381 5.61598
R13888 VDD.n2381 VDD.n2380 5.61598
R13889 VDD.n2380 VDD.n1676 5.61598
R13890 VDD.n2374 VDD.n1676 5.61598
R13891 VDD.n2374 VDD.n2373 5.61598
R13892 VDD.n2373 VDD.n2372 5.61598
R13893 VDD.n2372 VDD.n1681 5.61598
R13894 VDD.n2366 VDD.n1681 5.61598
R13895 VDD.n2366 VDD.n2365 5.61598
R13896 VDD.n2365 VDD.n2364 5.61598
R13897 VDD.n2364 VDD.n1685 5.61598
R13898 VDD.n2358 VDD.n1685 5.61598
R13899 VDD.n1124 VDD.n1122 5.61598
R13900 VDD.n1122 VDD.n1119 5.61598
R13901 VDD.n1119 VDD.n1116 5.61598
R13902 VDD.n1116 VDD.n1113 5.61598
R13903 VDD.n1113 VDD.n1110 5.61598
R13904 VDD.n1110 VDD.n1107 5.61598
R13905 VDD.n1107 VDD.n1104 5.61598
R13906 VDD.n1104 VDD.n1101 5.61598
R13907 VDD.n1101 VDD.n1098 5.61598
R13908 VDD.n1098 VDD.n1095 5.61598
R13909 VDD.n1095 VDD.n1092 5.61598
R13910 VDD.n1092 VDD.n1089 5.61598
R13911 VDD.n678 VDD.n676 5.61598
R13912 VDD.n676 VDD.n673 5.61598
R13913 VDD.n673 VDD.n670 5.61598
R13914 VDD.n670 VDD.n667 5.61598
R13915 VDD.n667 VDD.n664 5.61598
R13916 VDD.n664 VDD.n661 5.61598
R13917 VDD.n661 VDD.n658 5.61598
R13918 VDD.n658 VDD.n655 5.61598
R13919 VDD.n655 VDD.n652 5.61598
R13920 VDD.n652 VDD.n649 5.61598
R13921 VDD.n649 VDD.n646 5.61598
R13922 VDD.n646 VDD.n643 5.61598
R13923 VDD.n10768 VDD.n10699 5.57349
R13924 VDD.n9597 VDD.n9589 5.57349
R13925 VDD.n10110 VDD.t155 5.5395
R13926 VDD.n10110 VDD.t153 5.5395
R13927 VDD.n9739 VDD.t35 5.5395
R13928 VDD.n9739 VDD.t56 5.5395
R13929 VDD.n9763 VDD.t56 5.5395
R13930 VDD.n9763 VDD.t199 5.5395
R13931 VDD.n9523 VDD.t198 5.5395
R13932 VDD.n9523 VDD.t192 5.5395
R13933 VDD.n9784 VDD.t166 5.5395
R13934 VDD.n9784 VDD.t169 5.5395
R13935 VDD.n9810 VDD.t124 5.5395
R13936 VDD.n9810 VDD.t161 5.5395
R13937 VDD.n9480 VDD.t116 5.5395
R13938 VDD.n9480 VDD.t114 5.5395
R13939 VDD.n9856 VDD.t135 5.5395
R13940 VDD.n9856 VDD.t2 5.5395
R13941 VDD.n10883 VDD.t141 5.5395
R13942 VDD.n10883 VDD.t53 5.5395
R13943 VDD.t53 VDD.n10878 5.5395
R13944 VDD.n10878 VDD.t38 5.5395
R13945 VDD.n8933 VDD.t41 5.5395
R13946 VDD.n8933 VDD.t60 5.5395
R13947 VDD.n9049 VDD.t60 5.5395
R13948 VDD.n9049 VDD.t44 5.5395
R13949 VDD.t44 VDD.n9033 5.5395
R13950 VDD.n9033 VDD.t50 5.5395
R13951 VDD.n9311 VDD.t58 5.5395
R13952 VDD.n9311 VDD.t191 5.5395
R13953 VDD.n10924 VDD.t190 5.5395
R13954 VDD.n10924 VDD.t46 5.5395
R13955 VDD.n12481 VDD.n12429 5.44996
R13956 VDD VDD.n9969 5.43553
R13957 VDD.n8720 VDD.n8719 5.42303
R13958 VDD.n9697 VDD.n9641 5.39401
R13959 VDD.n10850 VDD.n10687 5.39401
R13960 VDD.n9700 VDD.n9641 5.39321
R13961 VDD.n10847 VDD.n10687 5.39321
R13962 VDD.n2471 VDD 5.2805
R13963 VDD.n831 VDD 5.2805
R13964 VDD.n12776 VDD.t176 5.27719
R13965 VDD.n10033 VDD.n10031 5.27109
R13966 VDD.n10038 VDD.n10034 5.27109
R13967 VDD.n10592 VDD.n10590 5.27109
R13968 VDD.n10597 VDD.n10593 5.27109
R13969 VDD.n10556 VDD.n10555 5.27109
R13970 VDD.n10550 VDD.n10535 5.27109
R13971 VDD.n9620 VDD.n9568 5.27109
R13972 VDD.n9629 VDD.n9565 5.27109
R13973 VDD.n9691 VDD.n9690 5.27109
R13974 VDD.n9707 VDD.n9706 5.27109
R13975 VDD.n10857 VDD.n10856 5.27109
R13976 VDD.n10841 VDD.n10840 5.27109
R13977 VDD.n10744 VDD.n10723 5.27109
R13978 VDD.n10739 VDD.n10725 5.27109
R13979 VDD.n12482 VDD.n12428 5.27109
R13980 VDD.n12467 VDD.n12466 5.27109
R13981 VDD.n12442 VDD.n12439 5.27109
R13982 VDD.n10024 VDD.n10018 5.25364
R13983 VDD.n10143 VDD.n10137 5.25364
R13984 VDD.n10530 VDD.n10529 5.25364
R13985 VDD.n5948 VDD.n5947 5.2318
R13986 VDD.n5094 VDD.n5093 5.2318
R13987 VDD.n4308 VDD.n4307 5.2318
R13988 VDD.n3454 VDD.n3453 5.2318
R13989 VDD.n2668 VDD.n2667 5.2318
R13990 VDD.n1813 VDD.n1812 5.2318
R13991 VDD.n1573 VDD.n1570 5.2318
R13992 VDD.n345 VDD.n342 5.2318
R13993 VDD.n9177 VDD.n9176 5.15851
R13994 VDD.n10183 VDD.t150 5.09674
R13995 VDD.n9289 VDD.n9265 4.96787
R13996 VDD.n9729 VDD.n9675 4.95584
R13997 VDD.n10818 VDD.n10690 4.95584
R13998 VDD.n8952 VDD.n8878 4.95584
R13999 VDD.n8855 VDD.n8790 4.95584
R14000 VDD.n9014 VDD.n8797 4.95584
R14001 VDD.n12362 VDD.n6975 4.91801
R14002 VDD.n12312 VDD.n12311 4.91801
R14003 VDD.n7056 VDD.n7053 4.91801
R14004 VDD.n7166 VDD.n7114 4.91801
R14005 VDD.n7221 VDD.n7220 4.91801
R14006 VDD.n7269 VDD.n7266 4.91801
R14007 VDD.n12185 VDD.n7308 4.91801
R14008 VDD.n12135 VDD.n12134 4.91801
R14009 VDD.n12129 VDD.n7351 4.91801
R14010 VDD.n12123 VDD.n7351 4.91801
R14011 VDD.n12123 VDD.n12122 4.91801
R14012 VDD.n12122 VDD.n12121 4.91801
R14013 VDD.n12121 VDD.n7357 4.91801
R14014 VDD.n12115 VDD.n7357 4.91801
R14015 VDD.n12115 VDD.n12114 4.91801
R14016 VDD.n12114 VDD.n12113 4.91801
R14017 VDD.n12113 VDD.n7361 4.91801
R14018 VDD.n12107 VDD.n7361 4.91801
R14019 VDD.n12107 VDD.n12106 4.91801
R14020 VDD.n12106 VDD.n12105 4.91801
R14021 VDD.n12105 VDD.n7365 4.91801
R14022 VDD.n12099 VDD.n7365 4.91801
R14023 VDD.n12099 VDD.n12098 4.91801
R14024 VDD.n12098 VDD.n12097 4.91801
R14025 VDD.n12097 VDD.n7369 4.91801
R14026 VDD.n8909 VDD.n8908 4.89462
R14027 VDD.n9377 VDD.n9376 4.89462
R14028 VDD.n9157 VDD.n9156 4.89462
R14029 VDD.n9130 VDD.n9129 4.89462
R14030 VDD.n9183 VDD.n9172 4.894
R14031 VDD.n12413 VDD.n6930 4.89039
R14032 VDD.n12408 VDD.n6930 4.89039
R14033 VDD.n12363 VDD.n6972 4.8457
R14034 VDD.n7014 VDD.n7013 4.8457
R14035 VDD.n12267 VDD.n12266 4.8457
R14036 VDD.n7160 VDD.n7159 4.8457
R14037 VDD.n7219 VDD.n7092 4.8457
R14038 VDD.n12234 VDD.n12233 4.8457
R14039 VDD.n12186 VDD.n7305 4.8457
R14040 VDD.n7347 VDD.n7346 4.8457
R14041 VDD.n9158 VDD.n9082 4.78705
R14042 VDD.n6346 VDD.n6345 4.78659
R14043 VDD.n5492 VDD.n5491 4.78659
R14044 VDD.n4706 VDD.n4705 4.78659
R14045 VDD.n3852 VDD.n3851 4.78659
R14046 VDD.n3066 VDD.n3065 4.78659
R14047 VDD.n2211 VDD.n2210 4.78659
R14048 VDD.n1604 VDD.n1601 4.78659
R14049 VDD.n376 VDD.n373 4.78659
R14050 VDD.n8201 VDD.n8087 4.7505
R14051 VDD.n8203 VDD.n8202 4.7505
R14052 VDD.n8213 VDD.n8081 4.7505
R14053 VDD.n8214 VDD.n8076 4.7505
R14054 VDD.n8219 VDD.n8217 4.7505
R14055 VDD.n8218 VDD.n8070 4.7505
R14056 VDD.n8230 VDD.n8229 4.7505
R14057 VDD.n8233 VDD.n8065 4.7505
R14058 VDD.n8235 VDD.n8234 4.7505
R14059 VDD.n8245 VDD.n8059 4.7505
R14060 VDD.n8247 VDD.n8246 4.7505
R14061 VDD.n8257 VDD.n8053 4.7505
R14062 VDD.n8258 VDD.n8048 4.7505
R14063 VDD.n8263 VDD.n8261 4.7505
R14064 VDD.n8262 VDD.n8042 4.7505
R14065 VDD.n8274 VDD.n8273 4.7505
R14066 VDD.n8277 VDD.n8037 4.7505
R14067 VDD.n8279 VDD.n8278 4.7505
R14068 VDD.n8288 VDD.n8030 4.7505
R14069 VDD.n8289 VDD.n8025 4.7505
R14070 VDD.n8294 VDD.n8292 4.7505
R14071 VDD.n8293 VDD.n8019 4.7505
R14072 VDD.n8305 VDD.n8304 4.7505
R14073 VDD.n8308 VDD.n8014 4.7505
R14074 VDD.n8310 VDD.n8309 4.7505
R14075 VDD.n8320 VDD.n8008 4.7505
R14076 VDD.n8322 VDD.n8321 4.7505
R14077 VDD.n8332 VDD.n8002 4.7505
R14078 VDD.n8334 VDD.n8333 4.7505
R14079 VDD.n8339 VDD.n7989 4.7505
R14080 VDD.n8488 VDD.n8487 4.7505
R14081 VDD.n8484 VDD.n8340 4.7505
R14082 VDD.n8483 VDD.n8345 4.7505
R14083 VDD.n8355 VDD.n8354 4.7505
R14084 VDD.n8473 VDD.n8472 4.7505
R14085 VDD.n8469 VDD.n8356 4.7505
R14086 VDD.n8468 VDD.n8362 4.7505
R14087 VDD.n8371 VDD.n8370 4.7505
R14088 VDD.n8459 VDD.n8458 4.7505
R14089 VDD.n8455 VDD.n8372 4.7505
R14090 VDD.n8454 VDD.n8378 4.7505
R14091 VDD.n8388 VDD.n8387 4.7505
R14092 VDD.n8444 VDD.n8443 4.7505
R14093 VDD.n8440 VDD.n8389 4.7505
R14094 VDD.n8439 VDD.n8395 4.7505
R14095 VDD.n8405 VDD.n8404 4.7505
R14096 VDD.n8429 VDD.n8428 4.7505
R14097 VDD.n8425 VDD.n8406 4.7505
R14098 VDD.n8424 VDD.n8413 4.7505
R14099 VDD.n8412 VDD.n7764 4.7505
R14100 VDD.n8568 VDD.n8567 4.7505
R14101 VDD.n9658 VDD.n9657 4.73575
R14102 VDD.n9673 VDD.n9659 4.73575
R14103 VDD.n10801 VDD.n10800 4.73575
R14104 VDD.n10816 VDD.n10802 4.73575
R14105 VDD.n8877 VDD.n8876 4.73575
R14106 VDD.n8955 VDD.n8954 4.73575
R14107 VDD.n8975 VDD.n8974 4.73575
R14108 VDD.n9012 VDD.n8998 4.73575
R14109 VDD.n8978 VDD.n8977 4.73575
R14110 VDD.n8997 VDD.n8996 4.73575
R14111 VDD.n9288 VDD.n9287 4.73575
R14112 VDD.n9418 VDD.n9417 4.73575
R14113 VDD.n6155 VDD.n6103 4.73093
R14114 VDD.n6109 VDD.n6103 4.73093
R14115 VDD.n6149 VDD.n6109 4.73093
R14116 VDD.n6149 VDD.n6148 4.73093
R14117 VDD.n6148 VDD.n6147 4.73093
R14118 VDD.n6147 VDD.n6110 4.73093
R14119 VDD.n6141 VDD.n6110 4.73093
R14120 VDD.n6141 VDD.n6140 4.73093
R14121 VDD.n6140 VDD.n6139 4.73093
R14122 VDD.n6139 VDD.n6115 4.73093
R14123 VDD.n6133 VDD.n6115 4.73093
R14124 VDD.n6133 VDD.n6132 4.73093
R14125 VDD.n6132 VDD.n6131 4.73093
R14126 VDD.n6131 VDD.n6119 4.73093
R14127 VDD.n6125 VDD.n6119 4.73093
R14128 VDD.n6125 VDD.n6124 4.73093
R14129 VDD.n6124 VDD.n5899 4.73093
R14130 VDD.n5301 VDD.n5249 4.73093
R14131 VDD.n5255 VDD.n5249 4.73093
R14132 VDD.n5295 VDD.n5255 4.73093
R14133 VDD.n5295 VDD.n5294 4.73093
R14134 VDD.n5294 VDD.n5293 4.73093
R14135 VDD.n5293 VDD.n5256 4.73093
R14136 VDD.n5287 VDD.n5256 4.73093
R14137 VDD.n5287 VDD.n5286 4.73093
R14138 VDD.n5286 VDD.n5285 4.73093
R14139 VDD.n5285 VDD.n5261 4.73093
R14140 VDD.n5279 VDD.n5261 4.73093
R14141 VDD.n5279 VDD.n5278 4.73093
R14142 VDD.n5278 VDD.n5277 4.73093
R14143 VDD.n5277 VDD.n5265 4.73093
R14144 VDD.n5271 VDD.n5265 4.73093
R14145 VDD.n5271 VDD.n5270 4.73093
R14146 VDD.n5270 VDD.n5045 4.73093
R14147 VDD.n4515 VDD.n4463 4.73093
R14148 VDD.n4469 VDD.n4463 4.73093
R14149 VDD.n4509 VDD.n4469 4.73093
R14150 VDD.n4509 VDD.n4508 4.73093
R14151 VDD.n4508 VDD.n4507 4.73093
R14152 VDD.n4507 VDD.n4470 4.73093
R14153 VDD.n4501 VDD.n4470 4.73093
R14154 VDD.n4501 VDD.n4500 4.73093
R14155 VDD.n4500 VDD.n4499 4.73093
R14156 VDD.n4499 VDD.n4475 4.73093
R14157 VDD.n4493 VDD.n4475 4.73093
R14158 VDD.n4493 VDD.n4492 4.73093
R14159 VDD.n4492 VDD.n4491 4.73093
R14160 VDD.n4491 VDD.n4479 4.73093
R14161 VDD.n4485 VDD.n4479 4.73093
R14162 VDD.n4485 VDD.n4484 4.73093
R14163 VDD.n4484 VDD.n4259 4.73093
R14164 VDD.n3661 VDD.n3609 4.73093
R14165 VDD.n3615 VDD.n3609 4.73093
R14166 VDD.n3655 VDD.n3615 4.73093
R14167 VDD.n3655 VDD.n3654 4.73093
R14168 VDD.n3654 VDD.n3653 4.73093
R14169 VDD.n3653 VDD.n3616 4.73093
R14170 VDD.n3647 VDD.n3616 4.73093
R14171 VDD.n3647 VDD.n3646 4.73093
R14172 VDD.n3646 VDD.n3645 4.73093
R14173 VDD.n3645 VDD.n3621 4.73093
R14174 VDD.n3639 VDD.n3621 4.73093
R14175 VDD.n3639 VDD.n3638 4.73093
R14176 VDD.n3638 VDD.n3637 4.73093
R14177 VDD.n3637 VDD.n3625 4.73093
R14178 VDD.n3631 VDD.n3625 4.73093
R14179 VDD.n3631 VDD.n3630 4.73093
R14180 VDD.n3630 VDD.n3405 4.73093
R14181 VDD.n2875 VDD.n2823 4.73093
R14182 VDD.n2829 VDD.n2823 4.73093
R14183 VDD.n2869 VDD.n2829 4.73093
R14184 VDD.n2869 VDD.n2868 4.73093
R14185 VDD.n2868 VDD.n2867 4.73093
R14186 VDD.n2867 VDD.n2830 4.73093
R14187 VDD.n2861 VDD.n2830 4.73093
R14188 VDD.n2861 VDD.n2860 4.73093
R14189 VDD.n2860 VDD.n2859 4.73093
R14190 VDD.n2859 VDD.n2835 4.73093
R14191 VDD.n2853 VDD.n2835 4.73093
R14192 VDD.n2853 VDD.n2852 4.73093
R14193 VDD.n2852 VDD.n2851 4.73093
R14194 VDD.n2851 VDD.n2839 4.73093
R14195 VDD.n2845 VDD.n2839 4.73093
R14196 VDD.n2845 VDD.n2844 4.73093
R14197 VDD.n2844 VDD.n2619 4.73093
R14198 VDD.n2020 VDD.n1968 4.73093
R14199 VDD.n1974 VDD.n1968 4.73093
R14200 VDD.n2014 VDD.n1974 4.73093
R14201 VDD.n2014 VDD.n2013 4.73093
R14202 VDD.n2013 VDD.n2012 4.73093
R14203 VDD.n2012 VDD.n1975 4.73093
R14204 VDD.n2006 VDD.n1975 4.73093
R14205 VDD.n2006 VDD.n2005 4.73093
R14206 VDD.n2005 VDD.n2004 4.73093
R14207 VDD.n2004 VDD.n1980 4.73093
R14208 VDD.n1998 VDD.n1980 4.73093
R14209 VDD.n1998 VDD.n1997 4.73093
R14210 VDD.n1997 VDD.n1996 4.73093
R14211 VDD.n1996 VDD.n1984 4.73093
R14212 VDD.n1990 VDD.n1984 4.73093
R14213 VDD.n1990 VDD.n1989 4.73093
R14214 VDD.n1989 VDD.n1764 4.73093
R14215 VDD.n1316 VDD.n1314 4.73093
R14216 VDD.n1319 VDD.n1316 4.73093
R14217 VDD.n1323 VDD.n1319 4.73093
R14218 VDD.n1326 VDD.n1323 4.73093
R14219 VDD.n1329 VDD.n1326 4.73093
R14220 VDD.n1332 VDD.n1329 4.73093
R14221 VDD.n1335 VDD.n1332 4.73093
R14222 VDD.n1338 VDD.n1335 4.73093
R14223 VDD.n1341 VDD.n1338 4.73093
R14224 VDD.n1344 VDD.n1341 4.73093
R14225 VDD.n1347 VDD.n1344 4.73093
R14226 VDD.n1350 VDD.n1347 4.73093
R14227 VDD.n1353 VDD.n1350 4.73093
R14228 VDD.n1356 VDD.n1353 4.73093
R14229 VDD.n1359 VDD.n1356 4.73093
R14230 VDD.n1362 VDD.n1359 4.73093
R14231 VDD.n1365 VDD.n1362 4.73093
R14232 VDD.n88 VDD.n86 4.73093
R14233 VDD.n91 VDD.n88 4.73093
R14234 VDD.n95 VDD.n91 4.73093
R14235 VDD.n98 VDD.n95 4.73093
R14236 VDD.n101 VDD.n98 4.73093
R14237 VDD.n104 VDD.n101 4.73093
R14238 VDD.n107 VDD.n104 4.73093
R14239 VDD.n110 VDD.n107 4.73093
R14240 VDD.n113 VDD.n110 4.73093
R14241 VDD.n116 VDD.n113 4.73093
R14242 VDD.n119 VDD.n116 4.73093
R14243 VDD.n122 VDD.n119 4.73093
R14244 VDD.n125 VDD.n122 4.73093
R14245 VDD.n128 VDD.n125 4.73093
R14246 VDD.n131 VDD.n128 4.73093
R14247 VDD.n134 VDD.n131 4.73093
R14248 VDD.n137 VDD.n134 4.73093
R14249 VDD.n8553 VDD.n7775 4.70536
R14250 VDD.n12356 VDD.n6979 4.70106
R14251 VDD.n12310 VDD.n7015 4.70106
R14252 VDD.n12263 VDD.n12262 4.70106
R14253 VDD.n7167 VDD.n7112 4.70106
R14254 VDD.n7226 VDD.n7090 4.70106
R14255 VDD.n12230 VDD.n12229 4.70106
R14256 VDD.n12179 VDD.n7312 4.70106
R14257 VDD.n12133 VDD.n7348 4.70106
R14258 VDD.n5726 VDD.n5725 4.6533
R14259 VDD.n4086 VDD.n4085 4.6533
R14260 VDD.n2445 VDD.n2444 4.6533
R14261 VDD.n805 VDD.n804 4.6533
R14262 VDD.n9911 VDD.n9908 4.6505
R14263 VDD.n9967 VDD.n9906 4.6505
R14264 VDD.n9969 VDD.n9968 4.6505
R14265 VDD.n9959 VDD.n9958 4.6505
R14266 VDD.n9949 VDD.n9912 4.6505
R14267 VDD.n9948 VDD.n9913 4.6505
R14268 VDD.n9926 VDD.n9925 4.6505
R14269 VDD.n9936 VDD.n9926 4.6505
R14270 VDD.n9946 VDD.n9945 4.6505
R14271 VDD.n9915 VDD.n9914 4.6505
R14272 VDD.n9924 VDD.n9920 4.6505
R14273 VDD.n9938 VDD.n9937 4.6505
R14274 VDD.n9935 VDD.n9921 4.6505
R14275 VDD.n9934 VDD.n9933 4.6505
R14276 VDD.n9931 VDD.n9930 4.6505
R14277 VDD.n9981 VDD.n9980 4.6505
R14278 VDD.n8991 VDD.n8990 4.6505
R14279 VDD.n8969 VDD.n8968 4.6505
R14280 VDD.n8117 VDD.n8106 4.6505
R14281 VDD.n8193 VDD.n8192 4.6505
R14282 VDD.n8191 VDD.n8190 4.6505
R14283 VDD.n8127 VDD.n8107 4.6505
R14284 VDD.n8182 VDD.n8181 4.6505
R14285 VDD.n8180 VDD.n8179 4.6505
R14286 VDD.n8136 VDD.n8129 4.6505
R14287 VDD.n8172 VDD.n8171 4.6505
R14288 VDD.n8170 VDD.n8169 4.6505
R14289 VDD.n8145 VDD.n8138 4.6505
R14290 VDD.n8161 VDD.n8160 4.6505
R14291 VDD.n8159 VDD.n8158 4.6505
R14292 VDD.n8151 VDD.n7744 4.6505
R14293 VDD.n8604 VDD.n8603 4.6505
R14294 VDD.n8605 VDD.n7722 4.6505
R14295 VDD.n8606 VDD.n7723 4.6505
R14296 VDD.n8608 VDD.n8607 4.6505
R14297 VDD.n8609 VDD.n7740 4.6505
R14298 VDD.n11432 VDD.n11431 4.6505
R14299 VDD.n11430 VDD.n11429 4.6505
R14300 VDD.n8620 VDD.n7741 4.6505
R14301 VDD.n8639 VDD.n8638 4.6505
R14302 VDD.n8640 VDD.n8634 4.6505
R14303 VDD.n11413 VDD.n11412 4.6505
R14304 VDD.n11411 VDD.n11410 4.6505
R14305 VDD.n8651 VDD.n8635 4.6505
R14306 VDD.n8674 VDD.n8673 4.6505
R14307 VDD.n8679 VDD.n8678 4.6505
R14308 VDD.n8680 VDD.n8663 4.6505
R14309 VDD.n11388 VDD.n11387 4.6505
R14310 VDD.n11386 VDD.n11385 4.6505
R14311 VDD.n8689 VDD.n8681 4.6505
R14312 VDD.n8711 VDD.n8710 4.6505
R14313 VDD.n8712 VDD.n8706 4.6505
R14314 VDD.n11369 VDD.n11368 4.6505
R14315 VDD.n11367 VDD.n11366 4.6505
R14316 VDD.n8724 VDD.n8707 4.6505
R14317 VDD.n11044 VDD.n11043 4.6505
R14318 VDD.n11045 VDD.n11039 4.6505
R14319 VDD.n11350 VDD.n11349 4.6505
R14320 VDD.n11348 VDD.n11347 4.6505
R14321 VDD.n11056 VDD.n11040 4.6505
R14322 VDD.n11091 VDD.n11090 4.6505
R14323 VDD.n11092 VDD.n11068 4.6505
R14324 VDD.n11331 VDD.n11330 4.6505
R14325 VDD.n11329 VDD.n11328 4.6505
R14326 VDD.n11084 VDD.n11069 4.6505
R14327 VDD.n11316 VDD.n11315 4.6505
R14328 VDD.n11314 VDD.n11313 4.6505
R14329 VDD.n11109 VDD.n11087 4.6505
R14330 VDD.n11128 VDD.n11127 4.6505
R14331 VDD.n11129 VDD.n11123 4.6505
R14332 VDD.n11297 VDD.n11296 4.6505
R14333 VDD.n11295 VDD.n11294 4.6505
R14334 VDD.n11139 VDD.n11124 4.6505
R14335 VDD.n11159 VDD.n11158 4.6505
R14336 VDD.n11160 VDD.n11154 4.6505
R14337 VDD.n11278 VDD.n11277 4.6505
R14338 VDD.n11276 VDD.n11275 4.6505
R14339 VDD.n11171 VDD.n11155 4.6505
R14340 VDD.n11195 VDD.n11194 4.6505
R14341 VDD.n11200 VDD.n11199 4.6505
R14342 VDD.n11201 VDD.n11184 4.6505
R14343 VDD.n11253 VDD.n11252 4.6505
R14344 VDD.n11251 VDD.n11250 4.6505
R14345 VDD.n11210 VDD.n11202 4.6505
R14346 VDD.n11225 VDD.n11224 4.6505
R14347 VDD.n11227 VDD.n11226 4.6505
R14348 VDD.n11228 VDD.n6605 4.6505
R14349 VDD.n12707 VDD.n12706 4.6505
R14350 VDD.n12705 VDD.n12704 4.6505
R14351 VDD.n12699 VDD.n12698 4.6505
R14352 VDD.n6704 VDD.n6611 4.6505
R14353 VDD.n6708 VDD.n6706 4.6505
R14354 VDD.n12687 VDD.n12686 4.6505
R14355 VDD.n12685 VDD.n12684 4.6505
R14356 VDD.n6710 VDD.n6709 4.6505
R14357 VDD.n10255 VDD.n10254 4.6505
R14358 VDD.n10252 VDD.n10251 4.6505
R14359 VDD.n10261 VDD.n10260 4.6505
R14360 VDD.n10263 VDD.n10262 4.6505
R14361 VDD.n10248 VDD.n10247 4.6505
R14362 VDD.n10269 VDD.n10268 4.6505
R14363 VDD.n10271 VDD.n10270 4.6505
R14364 VDD.n10242 VDD.n10241 4.6505
R14365 VDD.n10277 VDD.n10276 4.6505
R14366 VDD.n10279 VDD.n10278 4.6505
R14367 VDD.n10280 VDD.n10237 4.6505
R14368 VDD.n10287 VDD.n10286 4.6505
R14369 VDD.n10289 VDD.n10288 4.6505
R14370 VDD.n10234 VDD.n10233 4.6505
R14371 VDD.n10295 VDD.n10294 4.6505
R14372 VDD.n10297 VDD.n10296 4.6505
R14373 VDD.n10230 VDD.n10229 4.6505
R14374 VDD.n10303 VDD.n10302 4.6505
R14375 VDD.n10305 VDD.n10304 4.6505
R14376 VDD.n10224 VDD.n10223 4.6505
R14377 VDD.n10311 VDD.n10310 4.6505
R14378 VDD.n10313 VDD.n10312 4.6505
R14379 VDD.n10220 VDD.n10219 4.6505
R14380 VDD.n10319 VDD.n10318 4.6505
R14381 VDD.n10321 VDD.n10320 4.6505
R14382 VDD.n10216 VDD.n10215 4.6505
R14383 VDD.n10328 VDD.n10327 4.6505
R14384 VDD.n10330 VDD.n10329 4.6505
R14385 VDD.n10331 VDD.n10208 4.6505
R14386 VDD.n10340 VDD.n10339 4.6505
R14387 VDD.n10342 VDD.n10341 4.6505
R14388 VDD.n10205 VDD.n10204 4.6505
R14389 VDD.n10348 VDD.n10347 4.6505
R14390 VDD.n10350 VDD.n10349 4.6505
R14391 VDD.n10201 VDD.n10200 4.6505
R14392 VDD.n10356 VDD.n10355 4.6505
R14393 VDD.n10358 VDD.n10357 4.6505
R14394 VDD.n10197 VDD.n10196 4.6505
R14395 VDD.n10364 VDD.n10363 4.6505
R14396 VDD.n10366 VDD.n10365 4.6505
R14397 VDD.n10191 VDD.n10190 4.6505
R14398 VDD.n10372 VDD.n10371 4.6505
R14399 VDD.n10374 VDD.n10373 4.6505
R14400 VDD.n10187 VDD.n10186 4.6505
R14401 VDD.n10381 VDD.n10380 4.6505
R14402 VDD.n10383 VDD.n10382 4.6505
R14403 VDD.n10181 VDD.n10180 4.6505
R14404 VDD.n10390 VDD.n10389 4.6505
R14405 VDD.n10392 VDD.n10391 4.6505
R14406 VDD.n10177 VDD.n10176 4.6505
R14407 VDD.n10398 VDD.n10397 4.6505
R14408 VDD.n10400 VDD.n10399 4.6505
R14409 VDD.n10173 VDD.n10172 4.6505
R14410 VDD.n10406 VDD.n10405 4.6505
R14411 VDD.n10408 VDD.n10407 4.6505
R14412 VDD.n10169 VDD.n10168 4.6505
R14413 VDD.n10414 VDD.n10413 4.6505
R14414 VDD.n10416 VDD.n10415 4.6505
R14415 VDD.n10417 VDD.n6928 4.6505
R14416 VDD.n12417 VDD.n12416 4.6505
R14417 VDD.n12415 VDD.n12414 4.6505
R14418 VDD.n6935 VDD.n6929 4.6505
R14419 VDD.n6945 VDD.n6943 4.6505
R14420 VDD.n12399 VDD.n12398 4.6505
R14421 VDD.n12397 VDD.n12396 4.6505
R14422 VDD.n6947 VDD.n6946 4.6505
R14423 VDD.n6954 VDD.n6952 4.6505
R14424 VDD.n12388 VDD.n12387 4.6505
R14425 VDD.n12386 VDD.n12385 4.6505
R14426 VDD.n6956 VDD.n6955 4.6505
R14427 VDD.n6963 VDD.n6961 4.6505
R14428 VDD.n12377 VDD.n12376 4.6505
R14429 VDD.n12375 VDD.n12374 4.6505
R14430 VDD.n6965 VDD.n6964 4.6505
R14431 VDD.n6973 VDD.n6971 4.6505
R14432 VDD.n12366 VDD.n12365 4.6505
R14433 VDD.n12364 VDD.n12363 4.6505
R14434 VDD.n6979 VDD.n6974 4.6505
R14435 VDD.n12355 VDD.n12354 4.6505
R14436 VDD.n12353 VDD.n12352 4.6505
R14437 VDD.n6982 VDD.n6981 4.6505
R14438 VDD.n6989 VDD.n6987 4.6505
R14439 VDD.n12344 VDD.n12343 4.6505
R14440 VDD.n12342 VDD.n12341 4.6505
R14441 VDD.n6991 VDD.n6990 4.6505
R14442 VDD.n6998 VDD.n6996 4.6505
R14443 VDD.n12333 VDD.n12332 4.6505
R14444 VDD.n12331 VDD.n12330 4.6505
R14445 VDD.n7000 VDD.n6999 4.6505
R14446 VDD.n7007 VDD.n7005 4.6505
R14447 VDD.n12322 VDD.n12321 4.6505
R14448 VDD.n12320 VDD.n12319 4.6505
R14449 VDD.n7009 VDD.n7008 4.6505
R14450 VDD.n7016 VDD.n7014 4.6505
R14451 VDD.n12310 VDD.n12309 4.6505
R14452 VDD.n12308 VDD.n12307 4.6505
R14453 VDD.n7018 VDD.n7017 4.6505
R14454 VDD.n7027 VDD.n7025 4.6505
R14455 VDD.n12299 VDD.n12298 4.6505
R14456 VDD.n12297 VDD.n12296 4.6505
R14457 VDD.n7029 VDD.n7028 4.6505
R14458 VDD.n7036 VDD.n7034 4.6505
R14459 VDD.n12288 VDD.n12287 4.6505
R14460 VDD.n12286 VDD.n12285 4.6505
R14461 VDD.n7038 VDD.n7037 4.6505
R14462 VDD.n7045 VDD.n7043 4.6505
R14463 VDD.n12277 VDD.n12276 4.6505
R14464 VDD.n12275 VDD.n12274 4.6505
R14465 VDD.n7047 VDD.n7046 4.6505
R14466 VDD.n7054 VDD.n7052 4.6505
R14467 VDD.n12266 VDD.n12265 4.6505
R14468 VDD.n12264 VDD.n12263 4.6505
R14469 VDD.n7057 VDD.n7055 4.6505
R14470 VDD.n7066 VDD.n7064 4.6505
R14471 VDD.n12255 VDD.n12254 4.6505
R14472 VDD.n12253 VDD.n12252 4.6505
R14473 VDD.n7068 VDD.n7067 4.6505
R14474 VDD.n7130 VDD.n7129 4.6505
R14475 VDD.n7126 VDD.n7125 4.6505
R14476 VDD.n7137 VDD.n7136 4.6505
R14477 VDD.n7139 VDD.n7138 4.6505
R14478 VDD.n7122 VDD.n7121 4.6505
R14479 VDD.n7147 VDD.n7146 4.6505
R14480 VDD.n7149 VDD.n7148 4.6505
R14481 VDD.n7118 VDD.n7117 4.6505
R14482 VDD.n7156 VDD.n7155 4.6505
R14483 VDD.n7158 VDD.n7157 4.6505
R14484 VDD.n7159 VDD.n7113 4.6505
R14485 VDD.n7168 VDD.n7167 4.6505
R14486 VDD.n7170 VDD.n7169 4.6505
R14487 VDD.n7110 VDD.n7109 4.6505
R14488 VDD.n7178 VDD.n7177 4.6505
R14489 VDD.n7180 VDD.n7179 4.6505
R14490 VDD.n7106 VDD.n7105 4.6505
R14491 VDD.n7187 VDD.n7186 4.6505
R14492 VDD.n7189 VDD.n7188 4.6505
R14493 VDD.n7102 VDD.n7101 4.6505
R14494 VDD.n7197 VDD.n7196 4.6505
R14495 VDD.n7199 VDD.n7198 4.6505
R14496 VDD.n7098 VDD.n7097 4.6505
R14497 VDD.n7206 VDD.n7205 4.6505
R14498 VDD.n7208 VDD.n7207 4.6505
R14499 VDD.n7094 VDD.n7093 4.6505
R14500 VDD.n7217 VDD.n7216 4.6505
R14501 VDD.n7219 VDD.n7218 4.6505
R14502 VDD.n7090 VDD.n7089 4.6505
R14503 VDD.n7228 VDD.n7227 4.6505
R14504 VDD.n7230 VDD.n7229 4.6505
R14505 VDD.n7086 VDD.n7085 4.6505
R14506 VDD.n7237 VDD.n7236 4.6505
R14507 VDD.n7239 VDD.n7238 4.6505
R14508 VDD.n7082 VDD.n7081 4.6505
R14509 VDD.n7247 VDD.n7246 4.6505
R14510 VDD.n7249 VDD.n7248 4.6505
R14511 VDD.n7078 VDD.n7077 4.6505
R14512 VDD.n7257 VDD.n7256 4.6505
R14513 VDD.n7258 VDD.n7075 4.6505
R14514 VDD.n12244 VDD.n12243 4.6505
R14515 VDD.n12242 VDD.n12241 4.6505
R14516 VDD.n7260 VDD.n7259 4.6505
R14517 VDD.n7267 VDD.n7265 4.6505
R14518 VDD.n12233 VDD.n12232 4.6505
R14519 VDD.n12231 VDD.n12230 4.6505
R14520 VDD.n7270 VDD.n7268 4.6505
R14521 VDD.n7279 VDD.n7277 4.6505
R14522 VDD.n12222 VDD.n12221 4.6505
R14523 VDD.n12220 VDD.n12219 4.6505
R14524 VDD.n7281 VDD.n7280 4.6505
R14525 VDD.n7288 VDD.n7286 4.6505
R14526 VDD.n12211 VDD.n12210 4.6505
R14527 VDD.n12209 VDD.n12208 4.6505
R14528 VDD.n7290 VDD.n7289 4.6505
R14529 VDD.n7297 VDD.n7295 4.6505
R14530 VDD.n12200 VDD.n12199 4.6505
R14531 VDD.n12198 VDD.n12197 4.6505
R14532 VDD.n7299 VDD.n7298 4.6505
R14533 VDD.n7306 VDD.n7304 4.6505
R14534 VDD.n12189 VDD.n12188 4.6505
R14535 VDD.n12187 VDD.n12186 4.6505
R14536 VDD.n7312 VDD.n7307 4.6505
R14537 VDD.n12178 VDD.n12177 4.6505
R14538 VDD.n12176 VDD.n12175 4.6505
R14539 VDD.n7315 VDD.n7314 4.6505
R14540 VDD.n7322 VDD.n7320 4.6505
R14541 VDD.n12167 VDD.n12166 4.6505
R14542 VDD.n12165 VDD.n12164 4.6505
R14543 VDD.n7324 VDD.n7323 4.6505
R14544 VDD.n7331 VDD.n7329 4.6505
R14545 VDD.n12156 VDD.n12155 4.6505
R14546 VDD.n12154 VDD.n12153 4.6505
R14547 VDD.n7333 VDD.n7332 4.6505
R14548 VDD.n7340 VDD.n7338 4.6505
R14549 VDD.n12145 VDD.n12144 4.6505
R14550 VDD.n12143 VDD.n12142 4.6505
R14551 VDD.n7342 VDD.n7341 4.6505
R14552 VDD.n12133 VDD.n12132 4.6505
R14553 VDD.n12131 VDD.n12130 4.6505
R14554 VDD.n7373 VDD.n7350 4.6505
R14555 VDD.n7349 VDD.n7347 4.6505
R14556 VDD.n11657 VDD.n11656 4.6505
R14557 VDD.n11658 VDD.n7606 4.6505
R14558 VDD.n11660 VDD.n11659 4.6505
R14559 VDD.n7602 VDD.n7601 4.6505
R14560 VDD.n11669 VDD.n11668 4.6505
R14561 VDD.n11671 VDD.n11670 4.6505
R14562 VDD.n11672 VDD.n7594 4.6505
R14563 VDD.n11681 VDD.n11680 4.6505
R14564 VDD.n11682 VDD.n7592 4.6505
R14565 VDD.n11684 VDD.n11683 4.6505
R14566 VDD.n7588 VDD.n7587 4.6505
R14567 VDD.n11694 VDD.n11693 4.6505
R14568 VDD.n11695 VDD.n7585 4.6505
R14569 VDD.n11697 VDD.n11696 4.6505
R14570 VDD.n7581 VDD.n7580 4.6505
R14571 VDD.n11707 VDD.n11706 4.6505
R14572 VDD.n11708 VDD.n7578 4.6505
R14573 VDD.n11710 VDD.n11709 4.6505
R14574 VDD.n7574 VDD.n7573 4.6505
R14575 VDD.n11720 VDD.n11719 4.6505
R14576 VDD.n11721 VDD.n7571 4.6505
R14577 VDD.n11723 VDD.n11722 4.6505
R14578 VDD.n7567 VDD.n7566 4.6505
R14579 VDD.n11732 VDD.n11731 4.6505
R14580 VDD.n11734 VDD.n11733 4.6505
R14581 VDD.n7561 VDD.n7560 4.6505
R14582 VDD.n11745 VDD.n11744 4.6505
R14583 VDD.n11746 VDD.n7558 4.6505
R14584 VDD.n11748 VDD.n11747 4.6505
R14585 VDD.n7554 VDD.n7553 4.6505
R14586 VDD.n11758 VDD.n11757 4.6505
R14587 VDD.n11759 VDD.n7551 4.6505
R14588 VDD.n11761 VDD.n11760 4.6505
R14589 VDD.n7547 VDD.n7546 4.6505
R14590 VDD.n11771 VDD.n11770 4.6505
R14591 VDD.n11772 VDD.n7544 4.6505
R14592 VDD.n11774 VDD.n11773 4.6505
R14593 VDD.n7540 VDD.n7539 4.6505
R14594 VDD.n11783 VDD.n11782 4.6505
R14595 VDD.n11785 VDD.n11784 4.6505
R14596 VDD.n11786 VDD.n7532 4.6505
R14597 VDD.n11795 VDD.n11794 4.6505
R14598 VDD.n11796 VDD.n7530 4.6505
R14599 VDD.n11798 VDD.n11797 4.6505
R14600 VDD.n7526 VDD.n7525 4.6505
R14601 VDD.n11808 VDD.n11807 4.6505
R14602 VDD.n11809 VDD.n7523 4.6505
R14603 VDD.n11811 VDD.n11810 4.6505
R14604 VDD.n7519 VDD.n7518 4.6505
R14605 VDD.n11821 VDD.n11820 4.6505
R14606 VDD.n11822 VDD.n7516 4.6505
R14607 VDD.n11824 VDD.n11823 4.6505
R14608 VDD.n7512 VDD.n7511 4.6505
R14609 VDD.n11834 VDD.n11833 4.6505
R14610 VDD.n11835 VDD.n7509 4.6505
R14611 VDD.n11837 VDD.n11836 4.6505
R14612 VDD.n7505 VDD.n7504 4.6505
R14613 VDD.n11846 VDD.n11845 4.6505
R14614 VDD.n11848 VDD.n11847 4.6505
R14615 VDD.n7499 VDD.n7498 4.6505
R14616 VDD.n11859 VDD.n11858 4.6505
R14617 VDD.n11860 VDD.n7496 4.6505
R14618 VDD.n11862 VDD.n11861 4.6505
R14619 VDD.n7492 VDD.n7491 4.6505
R14620 VDD.n11872 VDD.n11871 4.6505
R14621 VDD.n11873 VDD.n7489 4.6505
R14622 VDD.n11875 VDD.n11874 4.6505
R14623 VDD.n7485 VDD.n7484 4.6505
R14624 VDD.n11885 VDD.n11884 4.6505
R14625 VDD.n11886 VDD.n7482 4.6505
R14626 VDD.n11888 VDD.n11887 4.6505
R14627 VDD.n7478 VDD.n7477 4.6505
R14628 VDD.n11897 VDD.n11896 4.6505
R14629 VDD.n11899 VDD.n11898 4.6505
R14630 VDD.n11900 VDD.n7470 4.6505
R14631 VDD.n11909 VDD.n11908 4.6505
R14632 VDD.n11910 VDD.n7468 4.6505
R14633 VDD.n11912 VDD.n11911 4.6505
R14634 VDD.n7464 VDD.n7463 4.6505
R14635 VDD.n11922 VDD.n11921 4.6505
R14636 VDD.n11923 VDD.n7461 4.6505
R14637 VDD.n11925 VDD.n11924 4.6505
R14638 VDD.n7457 VDD.n7456 4.6505
R14639 VDD.n11935 VDD.n11934 4.6505
R14640 VDD.n11936 VDD.n7454 4.6505
R14641 VDD.n11938 VDD.n11937 4.6505
R14642 VDD.n7450 VDD.n7449 4.6505
R14643 VDD.n11948 VDD.n11947 4.6505
R14644 VDD.n11949 VDD.n7447 4.6505
R14645 VDD.n11951 VDD.n11950 4.6505
R14646 VDD.n7443 VDD.n7442 4.6505
R14647 VDD.n11960 VDD.n11959 4.6505
R14648 VDD.n11962 VDD.n11961 4.6505
R14649 VDD.n7437 VDD.n7436 4.6505
R14650 VDD.n11973 VDD.n11972 4.6505
R14651 VDD.n11974 VDD.n7434 4.6505
R14652 VDD.n11976 VDD.n11975 4.6505
R14653 VDD.n7430 VDD.n7429 4.6505
R14654 VDD.n11986 VDD.n11985 4.6505
R14655 VDD.n11987 VDD.n7427 4.6505
R14656 VDD.n11989 VDD.n11988 4.6505
R14657 VDD.n7423 VDD.n7422 4.6505
R14658 VDD.n11999 VDD.n11998 4.6505
R14659 VDD.n12000 VDD.n7420 4.6505
R14660 VDD.n12002 VDD.n12001 4.6505
R14661 VDD.n7416 VDD.n7415 4.6505
R14662 VDD.n12011 VDD.n12010 4.6505
R14663 VDD.n12013 VDD.n12012 4.6505
R14664 VDD.n12014 VDD.n7408 4.6505
R14665 VDD.n12023 VDD.n12022 4.6505
R14666 VDD.n12024 VDD.n7406 4.6505
R14667 VDD.n12026 VDD.n12025 4.6505
R14668 VDD.n7402 VDD.n7401 4.6505
R14669 VDD.n12036 VDD.n12035 4.6505
R14670 VDD.n12037 VDD.n7399 4.6505
R14671 VDD.n12039 VDD.n12038 4.6505
R14672 VDD.n7395 VDD.n7394 4.6505
R14673 VDD.n12049 VDD.n12048 4.6505
R14674 VDD.n12050 VDD.n7392 4.6505
R14675 VDD.n12052 VDD.n12051 4.6505
R14676 VDD.n7388 VDD.n7387 4.6505
R14677 VDD.n12062 VDD.n12061 4.6505
R14678 VDD.n12063 VDD.n7385 4.6505
R14679 VDD.n12065 VDD.n12064 4.6505
R14680 VDD.n7381 VDD.n7380 4.6505
R14681 VDD.n12075 VDD.n12074 4.6505
R14682 VDD.n12076 VDD.n7379 4.6505
R14683 VDD.n12079 VDD.n12078 4.6505
R14684 VDD.n12077 VDD.n7374 4.6505
R14685 VDD.n7609 VDD.n7608 4.6505
R14686 VDD.n11634 VDD.n11633 4.6505
R14687 VDD.n11636 VDD.n11635 4.6505
R14688 VDD.n11632 VDD.n7617 4.6505
R14689 VDD.n11631 VDD.n11630 4.6505
R14690 VDD.n7620 VDD.n7619 4.6505
R14691 VDD.n11621 VDD.n11620 4.6505
R14692 VDD.n11619 VDD.n7624 4.6505
R14693 VDD.n11618 VDD.n11617 4.6505
R14694 VDD.n7627 VDD.n7626 4.6505
R14695 VDD.n11608 VDD.n11607 4.6505
R14696 VDD.n11606 VDD.n7631 4.6505
R14697 VDD.n11605 VDD.n11604 4.6505
R14698 VDD.n7634 VDD.n7633 4.6505
R14699 VDD.n11595 VDD.n11594 4.6505
R14700 VDD.n11593 VDD.n7638 4.6505
R14701 VDD.n11592 VDD.n11591 4.6505
R14702 VDD.n11582 VDD.n7640 4.6505
R14703 VDD.n11581 VDD.n11580 4.6505
R14704 VDD.n11579 VDD.n11578 4.6505
R14705 VDD.n7647 VDD.n7646 4.6505
R14706 VDD.n11570 VDD.n11569 4.6505
R14707 VDD.n11568 VDD.n7651 4.6505
R14708 VDD.n11567 VDD.n11566 4.6505
R14709 VDD.n7654 VDD.n7653 4.6505
R14710 VDD.n11557 VDD.n11556 4.6505
R14711 VDD.n11555 VDD.n7658 4.6505
R14712 VDD.n11554 VDD.n11553 4.6505
R14713 VDD.n7661 VDD.n7660 4.6505
R14714 VDD.n11544 VDD.n11543 4.6505
R14715 VDD.n11542 VDD.n7665 4.6505
R14716 VDD.n11541 VDD.n11540 4.6505
R14717 VDD.n7668 VDD.n7667 4.6505
R14718 VDD.n11532 VDD.n11531 4.6505
R14719 VDD.n11530 VDD.n11529 4.6505
R14720 VDD.n7675 VDD.n7674 4.6505
R14721 VDD.n11521 VDD.n11520 4.6505
R14722 VDD.n11519 VDD.n7679 4.6505
R14723 VDD.n11518 VDD.n11517 4.6505
R14724 VDD.n7682 VDD.n7681 4.6505
R14725 VDD.n11508 VDD.n11507 4.6505
R14726 VDD.n11506 VDD.n7686 4.6505
R14727 VDD.n11505 VDD.n11504 4.6505
R14728 VDD.n7689 VDD.n7688 4.6505
R14729 VDD.n11495 VDD.n11494 4.6505
R14730 VDD.n11493 VDD.n7693 4.6505
R14731 VDD.n11492 VDD.n11491 4.6505
R14732 VDD.n7696 VDD.n7695 4.6505
R14733 VDD.n11482 VDD.n11481 4.6505
R14734 VDD.n11480 VDD.n7700 4.6505
R14735 VDD.n11479 VDD.n11478 4.6505
R14736 VDD.n11470 VDD.n7702 4.6505
R14737 VDD.n11469 VDD.n11468 4.6505
R14738 VDD.n11467 VDD.n11466 4.6505
R14739 VDD.n7709 VDD.n7708 4.6505
R14740 VDD.n11458 VDD.n11457 4.6505
R14741 VDD.n11456 VDD.n7713 4.6505
R14742 VDD.n11455 VDD.n11454 4.6505
R14743 VDD.n7716 VDD.n7715 4.6505
R14744 VDD.n7880 VDD.n7878 4.6505
R14745 VDD.n7885 VDD.n7884 4.6505
R14746 VDD.n7887 VDD.n7886 4.6505
R14747 VDD.n7877 VDD.n7875 4.6505
R14748 VDD.n7871 VDD.n7870 4.6505
R14749 VDD.n7895 VDD.n7894 4.6505
R14750 VDD.n7897 VDD.n7896 4.6505
R14751 VDD.n7867 VDD.n7863 4.6505
R14752 VDD.n7904 VDD.n7903 4.6505
R14753 VDD.n7906 VDD.n7905 4.6505
R14754 VDD.n7858 VDD.n7857 4.6505
R14755 VDD.n7913 VDD.n7912 4.6505
R14756 VDD.n7915 VDD.n7914 4.6505
R14757 VDD.n7852 VDD.n7851 4.6505
R14758 VDD.n7922 VDD.n7921 4.6505
R14759 VDD.n7924 VDD.n7923 4.6505
R14760 VDD.n7847 VDD.n7846 4.6505
R14761 VDD.n7931 VDD.n7930 4.6505
R14762 VDD.n7933 VDD.n7932 4.6505
R14763 VDD.n7845 VDD.n7843 4.6505
R14764 VDD.n7839 VDD.n7838 4.6505
R14765 VDD.n7941 VDD.n7940 4.6505
R14766 VDD.n7943 VDD.n7942 4.6505
R14767 VDD.n7834 VDD.n7833 4.6505
R14768 VDD.n7950 VDD.n7949 4.6505
R14769 VDD.n7952 VDD.n7951 4.6505
R14770 VDD.n7827 VDD.n7826 4.6505
R14771 VDD.n7959 VDD.n7958 4.6505
R14772 VDD.n7961 VDD.n7960 4.6505
R14773 VDD.n7821 VDD.n7820 4.6505
R14774 VDD.n7968 VDD.n7967 4.6505
R14775 VDD.n7970 VDD.n7969 4.6505
R14776 VDD.n7814 VDD.n7813 4.6505
R14777 VDD.n7977 VDD.n7976 4.6505
R14778 VDD.n7979 VDD.n7978 4.6505
R14779 VDD.n7981 VDD.n7811 4.6505
R14780 VDD.n7789 VDD.n7787 4.6505
R14781 VDD.n8533 VDD.n8532 4.6505
R14782 VDD.n8531 VDD.n8530 4.6505
R14783 VDD.n7791 VDD.n7790 4.6505
R14784 VDD.n8524 VDD.n8523 4.6505
R14785 VDD.n8522 VDD.n8521 4.6505
R14786 VDD.n7799 VDD.n7795 4.6505
R14787 VDD.n8514 VDD.n8513 4.6505
R14788 VDD.n8512 VDD.n8511 4.6505
R14789 VDD.n7802 VDD.n7801 4.6505
R14790 VDD.n8506 VDD.n8505 4.6505
R14791 VDD.n8504 VDD.n8503 4.6505
R14792 VDD.n7807 VDD.n7806 4.6505
R14793 VDD.n7986 VDD.n7985 4.6505
R14794 VDD.n7984 VDD.n7810 4.6505
R14795 VDD.n7780 VDD.n7779 4.6505
R14796 VDD.n8550 VDD.n8549 4.6505
R14797 VDD.n8552 VDD.n8551 4.6505
R14798 VDD.n7778 VDD.n7777 4.6505
R14799 VDD.n7770 VDD.n7769 4.6505
R14800 VDD.n8420 VDD.n8419 4.6505
R14801 VDD.n8409 VDD.n8400 4.6505
R14802 VDD.n8392 VDD.n8383 4.6505
R14803 VDD.n8450 VDD.n8449 4.6505
R14804 VDD.n8375 VDD.n8365 4.6505
R14805 VDD.n8465 VDD.n8464 4.6505
R14806 VDD.n8479 VDD.n8478 4.6505
R14807 VDD.n8342 VDD.n7995 4.6505
R14808 VDD.n8494 VDD.n8493 4.6505
R14809 VDD.n8006 VDD.n8005 4.6505
R14810 VDD.n8314 VDD.n8313 4.6505
R14811 VDD.n8301 VDD.n8300 4.6505
R14812 VDD.n8028 VDD.n8022 4.6505
R14813 VDD.n8040 VDD.n8033 4.6505
R14814 VDD.n8268 VDD.n8267 4.6505
R14815 VDD.n8254 VDD.n8253 4.6505
R14816 VDD.n8239 VDD.n8238 4.6505
R14817 VDD.n8226 VDD.n8225 4.6505
R14818 VDD.n8078 VDD.n8073 4.6505
R14819 VDD.n8208 VDD.n8207 4.6505
R14820 VDD.n8089 VDD.n8084 4.6505
R14821 VDD.n8210 VDD.n8209 4.6505
R14822 VDD.n8224 VDD.n8223 4.6505
R14823 VDD.n8068 VDD.n8062 4.6505
R14824 VDD.n8241 VDD.n8240 4.6505
R14825 VDD.n8057 VDD.n8056 4.6505
R14826 VDD.n8252 VDD.n8251 4.6505
R14827 VDD.n8050 VDD.n8045 4.6505
R14828 VDD.n8270 VDD.n8269 4.6505
R14829 VDD.n8283 VDD.n8282 4.6505
R14830 VDD.n8285 VDD.n8284 4.6505
R14831 VDD.n8299 VDD.n8298 4.6505
R14832 VDD.n8017 VDD.n8011 4.6505
R14833 VDD.n8316 VDD.n8315 4.6505
R14834 VDD.n8327 VDD.n8326 4.6505
R14835 VDD.n8329 VDD.n8328 4.6505
R14836 VDD.n7999 VDD.n7994 4.6505
R14837 VDD.n8492 VDD.n8491 4.6505
R14838 VDD.n8349 VDD.n8347 4.6505
R14839 VDD.n8477 VDD.n8476 4.6505
R14840 VDD.n8360 VDD.n8350 4.6505
R14841 VDD.n8463 VDD.n8462 4.6505
R14842 VDD.n8382 VDD.n8380 4.6505
R14843 VDD.n8448 VDD.n8447 4.6505
R14844 VDD.n8399 VDD.n8397 4.6505
R14845 VDD.n8435 VDD.n8434 4.6505
R14846 VDD.n8433 VDD.n8432 4.6505
R14847 VDD.n8418 VDD.n8414 4.6505
R14848 VDD.n8415 VDD.n7768 4.6505
R14849 VDD.n8564 VDD.n8563 4.6505
R14850 VDD.n8562 VDD.n8561 4.6505
R14851 VDD.n12702 VDD.n6606 4.6505
R14852 VDD.n5760 VDD.n5746 4.6505
R14853 VDD.n5759 VDD.n5758 4.6505
R14854 VDD.n5757 VDD.n5748 4.6505
R14855 VDD.n5756 VDD.n5755 4.6505
R14856 VDD.n5729 VDD.n5717 4.6505
R14857 VDD.n5736 VDD.n5735 4.6505
R14858 VDD.n5720 VDD.n5713 4.6505
R14859 VDD VDD.n5767 4.6505
R14860 VDD.n5719 VDD.n5712 4.6505
R14861 VDD.n5722 VDD.n5719 4.6505
R14862 VDD.n5728 VDD.n5727 4.6505
R14863 VDD.n4120 VDD.n4106 4.6505
R14864 VDD.n4119 VDD.n4118 4.6505
R14865 VDD.n4117 VDD.n4108 4.6505
R14866 VDD.n4116 VDD.n4115 4.6505
R14867 VDD.n4089 VDD.n4077 4.6505
R14868 VDD.n4096 VDD.n4095 4.6505
R14869 VDD.n4080 VDD.n4073 4.6505
R14870 VDD VDD.n4127 4.6505
R14871 VDD.n4079 VDD.n4072 4.6505
R14872 VDD.n4082 VDD.n4079 4.6505
R14873 VDD.n4088 VDD.n4087 4.6505
R14874 VDD.n2480 VDD.n2465 4.6505
R14875 VDD.n2479 VDD.n2478 4.6505
R14876 VDD.n2477 VDD.n2467 4.6505
R14877 VDD.n2476 VDD.n2475 4.6505
R14878 VDD.n2448 VDD.n2436 4.6505
R14879 VDD.n2455 VDD.n2454 4.6505
R14880 VDD.n2439 VDD.n2432 4.6505
R14881 VDD VDD.n2487 4.6505
R14882 VDD.n2438 VDD.n2431 4.6505
R14883 VDD.n2441 VDD.n2438 4.6505
R14884 VDD.n2447 VDD.n2446 4.6505
R14885 VDD.n840 VDD.n825 4.6505
R14886 VDD.n839 VDD.n838 4.6505
R14887 VDD.n837 VDD.n827 4.6505
R14888 VDD.n836 VDD.n835 4.6505
R14889 VDD.n808 VDD.n796 4.6505
R14890 VDD.n815 VDD.n814 4.6505
R14891 VDD.n799 VDD.n792 4.6505
R14892 VDD VDD.n847 4.6505
R14893 VDD.n798 VDD.n791 4.6505
R14894 VDD.n801 VDD.n798 4.6505
R14895 VDD.n807 VDD.n806 4.6505
R14896 VDD.n7777 VDD.n7772 4.63618
R14897 VDD.n11679 VDD.n7596 4.60579
R14898 VDD.n11736 VDD.n11735 4.60579
R14899 VDD.n11793 VDD.n7534 4.60579
R14900 VDD.n11850 VDD.n11849 4.60579
R14901 VDD.n11907 VDD.n7472 4.60579
R14902 VDD.n11964 VDD.n11963 4.60579
R14903 VDD.n12021 VDD.n7410 4.60579
R14904 VDD.n12081 VDD.n12080 4.60579
R14905 VDD.n7953 VDD.n7952 4.58155
R14906 VDD.n7952 VDD.n7832 4.58155
R14907 VDD.n7903 VDD.n7862 4.58155
R14908 VDD.n7903 VDD.n7902 4.58155
R14909 VDD.n11478 VDD.n7703 4.58155
R14910 VDD.n11478 VDD.n11477 4.58155
R14911 VDD.n11532 VDD.n7672 4.58155
R14912 VDD.n11532 VDD.n7673 4.58155
R14913 VDD.n11589 VDD.n7641 4.58155
R14914 VDD.n12367 VDD.n12366 4.55643
R14915 VDD.n12318 VDD.n7009 4.55643
R14916 VDD.n7052 VDD.n7051 4.55643
R14917 VDD.n7158 VDD.n7116 4.55643
R14918 VDD.n7216 VDD.n7215 4.55643
R14919 VDD.n7265 VDD.n7264 4.55643
R14920 VDD.n12190 VDD.n12189 4.55643
R14921 VDD.n12141 VDD.n7342 4.55643
R14922 VDD.n9069 VDD.n8748 4.53566
R14923 VDD.n11012 VDD.n8740 4.53566
R14924 VDD.n9118 VDD.n9112 4.5337
R14925 VDD.n11016 VDD.n8736 4.53087
R14926 VDD.n11009 VDD.n11008 4.52784
R14927 VDD.n10476 VDD.n10450 4.52055
R14928 VDD.n10072 VDD.n10071 4.51815
R14929 VDD.n10056 VDD.n10055 4.51815
R14930 VDD.n10092 VDD.n10006 4.51815
R14931 VDD.n10632 VDD.n10146 4.51815
R14932 VDD.n10615 VDD.n10614 4.51815
R14933 VDD.n10519 VDD.n10518 4.51815
R14934 VDD.n10534 VDD.n10533 4.51815
R14935 VDD.n9613 VDD.n9572 4.51815
R14936 VDD.n9621 VDD.n9570 4.51815
R14937 VDD.n9686 VDD.n9560 4.51815
R14938 VDD.n9712 VDD.n9711 4.51815
R14939 VDD.n10862 VDD.n10861 4.51815
R14940 VDD.n10836 VDD.n10835 4.51815
R14941 VDD.n10751 VDD.n10750 4.51815
R14942 VDD.n10745 VDD.n10715 4.51815
R14943 VDD.n8922 VDD.n8886 4.51815
R14944 VDD.n9051 VDD.n8781 4.51815
R14945 VDD.n8805 VDD.n8799 4.51815
R14946 VDD.n9059 VDD.n8764 4.51815
R14947 VDD.n9314 VDD.n9313 4.51815
R14948 VDD.n9340 VDD.n9339 4.51815
R14949 VDD.n9443 VDD.n9359 4.51815
R14950 VDD.n9101 VDD.n9100 4.51815
R14951 VDD.n7986 VDD.n7810 4.51815
R14952 VDD.n7982 VDD.n7810 4.51815
R14953 VDD.n12494 VDD.n12493 4.51815
R14954 VDD.n12487 VDD.n6910 4.51815
R14955 VDD.n12461 VDD.n12460 4.51815
R14956 VDD.n12447 VDD.n12440 4.51815
R14957 VDD.n9611 VDD.n9610 4.51417
R14958 VDD.n9747 VDD.n9554 4.51417
R14959 VDD.n9758 VDD.n9546 4.51417
R14960 VDD.n9538 VDD.n9527 4.51417
R14961 VDD.n9792 VDD.n9513 4.51417
R14962 VDD.n9805 VDD.n9502 4.51417
R14963 VDD.n9495 VDD.n9484 4.51417
R14964 VDD.n10864 VDD.n10774 4.51417
R14965 VDD.n10753 VDD.n10708 4.51417
R14966 VDD.n10497 VDD.n10158 4.50958
R14967 VDD.n10079 VDD.n10078 4.5005
R14968 VDD.n10113 VDD.n10089 4.5005
R14969 VDD.n10639 VDD.n10139 4.5005
R14970 VDD.n10454 VDD.n10452 4.5005
R14971 VDD.n10462 VDD.n10461 4.5005
R14972 VDD.n10467 VDD.n10466 4.5005
R14973 VDD.n10488 VDD.n10440 4.5005
R14974 VDD.n10445 VDD.n10441 4.5005
R14975 VDD.n10468 VDD.n10460 4.5005
R14976 VDD.n10463 VDD.n10459 4.5005
R14977 VDD.n10465 VDD.n10464 4.5005
R14978 VDD.n10490 VDD.n10437 4.5005
R14979 VDD.n10426 VDD.n10425 4.5005
R14980 VDD.n10516 VDD.n10510 4.5005
R14981 VDD.n10499 VDD.n10152 4.5005
R14982 VDD.n10568 VDD.n10152 4.5005
R14983 VDD.n10568 VDD.n10150 4.5005
R14984 VDD.n10567 VDD.n10499 4.5005
R14985 VDD.n10568 VDD.n10567 4.5005
R14986 VDD.n10568 VDD.n10149 4.5005
R14987 VDD.n10559 VDD.n10499 4.5005
R14988 VDD.n10498 VDD.n10155 4.5005
R14989 VDD.n10498 VDD.n10497 4.5005
R14990 VDD.n10616 VDD.n10583 4.5005
R14991 VDD.n10630 VDD.n10583 4.5005
R14992 VDD.n10148 VDD.n10131 4.5005
R14993 VDD.n10617 VDD.n10148 4.5005
R14994 VDD.n10629 VDD.n10131 4.5005
R14995 VDD.n10631 VDD.n10131 4.5005
R14996 VDD.n10628 VDD.n10627 4.5005
R14997 VDD.n10630 VDD.n10148 4.5005
R14998 VDD.n10117 VDD.n10116 4.5005
R14999 VDD.n10116 VDD.n10084 4.5005
R15000 VDD.n10116 VDD.n10002 4.5005
R15001 VDD.n10118 VDD.n10003 4.5005
R15002 VDD.n10059 VDD.n10015 4.5005
R15003 VDD.n10059 VDD.n10057 4.5005
R15004 VDD.n10082 VDD.n10013 4.5005
R15005 VDD.n10015 VDD.n10011 4.5005
R15006 VDD.n10015 VDD.n10010 4.5005
R15007 VDD.n10027 VDD.n10009 4.5005
R15008 VDD.n10083 VDD.n10010 4.5005
R15009 VDD.n10630 VDD.n10628 4.5005
R15010 VDD.n10631 VDD.n10630 4.5005
R15011 VDD.n10630 VDD.n10629 4.5005
R15012 VDD.n10629 VDD.n10145 4.5005
R15013 VDD.n10118 VDD.n10004 4.5005
R15014 VDD.n10116 VDD.n10004 4.5005
R15015 VDD.n10098 VDD.n10004 4.5005
R15016 VDD.n10026 VDD.n10011 4.5005
R15017 VDD.n10083 VDD.n10011 4.5005
R15018 VDD.n10083 VDD.n10009 4.5005
R15019 VDD.n10083 VDD.n10082 4.5005
R15020 VDD.n10015 VDD.n10009 4.5005
R15021 VDD.n10100 VDD.n10003 4.5005
R15022 VDD.n10108 VDD.n10002 4.5005
R15023 VDD.n10118 VDD.n10002 4.5005
R15024 VDD.n10102 VDD.n10084 4.5005
R15025 VDD.n10118 VDD.n10117 4.5005
R15026 VDD.n10628 VDD.n10131 4.5005
R15027 VDD.n10559 VDD.n10505 4.5005
R15028 VDD.n10506 VDD.n10149 4.5005
R15029 VDD.n10499 VDD.n10149 4.5005
R15030 VDD.n10567 VDD.n10566 4.5005
R15031 VDD.n10523 VDD.n10152 4.5005
R15032 VDD.n8839 VDD.n8782 4.5005
R15033 VDD.n9031 VDD.n9030 4.5005
R15034 VDD.n8936 VDD.n8935 4.5005
R15035 VDD.n9065 VDD.n8757 4.5005
R15036 VDD.n9058 VDD.n9057 4.5005
R15037 VDD.n8821 VDD.n8812 4.5005
R15038 VDD.n8812 VDD.n8809 4.5005
R15039 VDD.n8821 VDD.n8811 4.5005
R15040 VDD.n8821 VDD.n8820 4.5005
R15041 VDD.n8820 VDD.n8809 4.5005
R15042 VDD.n8809 VDD.n8808 4.5005
R15043 VDD.n9052 VDD.n8779 4.5005
R15044 VDD.n9053 VDD.n8777 4.5005
R15045 VDD.n8787 VDD.n8777 4.5005
R15046 VDD.n8819 VDD.n8813 4.5005
R15047 VDD.n8820 VDD.n8819 4.5005
R15048 VDD.n9056 VDD.n8768 4.5005
R15049 VDD.n9054 VDD.n8769 4.5005
R15050 VDD.n9056 VDD.n8769 4.5005
R15051 VDD.n9056 VDD.n9055 4.5005
R15052 VDD.n9055 VDD.n8771 4.5005
R15053 VDD.n9055 VDD.n9054 4.5005
R15054 VDD.n9054 VDD.n8774 4.5005
R15055 VDD.n9057 VDD.n8756 4.5005
R15056 VDD.n8902 VDD.n8756 4.5005
R15057 VDD.n9065 VDD.n8756 4.5005
R15058 VDD.n9065 VDD.n9064 4.5005
R15059 VDD.n9064 VDD.n8760 4.5005
R15060 VDD.n8927 VDD.n8774 4.5005
R15061 VDD.n8931 VDD.n8768 4.5005
R15062 VDD.n8779 VDD.n8777 4.5005
R15063 VDD.n8779 VDD.n8775 4.5005
R15064 VDD.n9040 VDD.n8775 4.5005
R15065 VDD.n9053 VDD.n8775 4.5005
R15066 VDD.n9053 VDD.n9052 4.5005
R15067 VDD.n9047 VDD.n9046 4.5005
R15068 VDD.n9046 VDD.n8779 4.5005
R15069 VDD.n8812 VDD.n8800 4.5005
R15070 VDD.n8908 VDD.n8757 4.5005
R15071 VDD.n9057 VDD.n8757 4.5005
R15072 VDD.n9069 VDD.n8754 4.5005
R15073 VDD.n8754 VDD.n8747 4.5005
R15074 VDD.n11002 VDD.n8747 4.5005
R15075 VDD.n11002 VDD.n11001 4.5005
R15076 VDD.n11001 VDD.n8754 4.5005
R15077 VDD.n9269 VDD.n9258 4.5005
R15078 VDD.n9394 VDD.n9360 4.5005
R15079 VDD.n9444 VDD.n9356 4.5005
R15080 VDD.n9445 VDD.n9444 4.5005
R15081 VDD.n10928 VDD.n9322 4.5005
R15082 VDD.n9326 VDD.n9322 4.5005
R15083 VDD.n9445 VDD.n9357 4.5005
R15084 VDD.n9377 VDD.n9357 4.5005
R15085 VDD.n10955 VDD.n10946 4.5005
R15086 VDD.n10956 VDD.n9226 4.5005
R15087 VDD.n10956 VDD.n10955 4.5005
R15088 VDD.n10946 VDD.n9226 4.5005
R15089 VDD.n10928 VDD.n9324 4.5005
R15090 VDD.n10928 VDD.n9321 4.5005
R15091 VDD.n10928 VDD.n10927 4.5005
R15092 VDD.n9331 VDD.n9321 4.5005
R15093 VDD.n9326 VDD.n9321 4.5005
R15094 VDD.n10927 VDD.n9326 4.5005
R15095 VDD.n10927 VDD.n10926 4.5005
R15096 VDD.n9318 VDD.n9250 4.5005
R15097 VDD.n9254 VDD.n9250 4.5005
R15098 VDD.n9318 VDD.n9251 4.5005
R15099 VDD.n9261 VDD.n9249 4.5005
R15100 VDD.n9318 VDD.n9249 4.5005
R15101 VDD.n9254 VDD.n9249 4.5005
R15102 VDD.n9309 VDD.n9251 4.5005
R15103 VDD.n9254 VDD.n9251 4.5005
R15104 VDD.n9317 VDD.n9253 4.5005
R15105 VDD.n9318 VDD.n9317 4.5005
R15106 VDD.n9342 VDD.n9324 4.5005
R15107 VDD.n9357 VDD.n9356 4.5005
R15108 VDD.n9446 VDD.n9356 4.5005
R15109 VDD.n9446 VDD.n9355 4.5005
R15110 VDD.n9446 VDD.n9445 4.5005
R15111 VDD.n9387 VDD.n9353 4.5005
R15112 VDD.n9356 VDD.n9353 4.5005
R15113 VDD.n9162 VDD.n9161 4.5005
R15114 VDD.n9096 VDD.n9085 4.5005
R15115 VDD.n9144 VDD.n9143 4.5005
R15116 VDD.n9122 VDD.n9121 4.5005
R15117 VDD.n9126 VDD.n9125 4.5005
R15118 VDD.n9138 VDD.n9137 4.5005
R15119 VDD.n9124 VDD.n9111 4.5005
R15120 VDD.n9127 VDD.n9110 4.5005
R15121 VDD.n9134 VDD.n9133 4.5005
R15122 VDD.n9135 VDD.n9107 4.5005
R15123 VDD.n9114 VDD.n9112 4.5005
R15124 VDD.n9145 VDD.n9095 4.5005
R15125 VDD.n9148 VDD.n9147 4.5005
R15126 VDD.n9103 VDD.n9100 4.5005
R15127 VDD.n9098 VDD.n9097 4.5005
R15128 VDD.n9153 VDD.n9152 4.5005
R15129 VDD.n9157 VDD.n9083 4.5005
R15130 VDD.n9160 VDD.n9081 4.5005
R15131 VDD.n10769 VDD.n10768 4.5005
R15132 VDD.n10866 VDD.n10674 4.5005
R15133 VDD.n10867 VDD.n10866 4.5005
R15134 VDD.n10897 VDD.n10896 4.5005
R15135 VDD.n10675 VDD.n10667 4.5005
R15136 VDD.n10675 VDD.n10670 4.5005
R15137 VDD.n10888 VDD.n10675 4.5005
R15138 VDD.n10895 VDD.n10675 4.5005
R15139 VDD.n10894 VDD.n10667 4.5005
R15140 VDD.n10894 VDD.n10670 4.5005
R15141 VDD.n10894 VDD.n10893 4.5005
R15142 VDD.n9849 VDD.n9830 4.5005
R15143 VDD.n9817 VDD.n9816 4.5005
R15144 VDD.n9817 VDD.n9481 4.5005
R15145 VDD.n10772 VDD.n10770 4.5005
R15146 VDD.n10874 VDD.n10770 4.5005
R15147 VDD.n10874 VDD.n10674 4.5005
R15148 VDD.n10769 VDD.n10696 4.5005
R15149 VDD.n10705 VDD.n10696 4.5005
R15150 VDD.n10712 VDD.n10696 4.5005
R15151 VDD.n10755 VDD.n10712 4.5005
R15152 VDD.n9215 VDD.n9214 4.5005
R15153 VDD.n10969 VDD.n9214 4.5005
R15154 VDD.n10968 VDD.n9215 4.5005
R15155 VDD.n10969 VDD.n10968 4.5005
R15156 VDD.n10709 VDD.n10708 4.5005
R15157 VDD.n10756 VDD.n10755 4.5005
R15158 VDD.n10874 VDD.n10694 4.5005
R15159 VDD.n10896 VDD.n10669 4.5005
R15160 VDD.n10673 VDD.n10667 4.5005
R15161 VDD.n10879 VDD.n10673 4.5005
R15162 VDD.n10895 VDD.n10673 4.5005
R15163 VDD.n9850 VDD.n9827 4.5005
R15164 VDD.n9850 VDD.n9838 4.5005
R15165 VDD.n9850 VDD.n9849 4.5005
R15166 VDD.n9849 VDD.n9835 4.5005
R15167 VDD.n9836 VDD.n9835 4.5005
R15168 VDD.n9867 VDD.n9830 4.5005
R15169 VDD.n9860 VDD.n9830 4.5005
R15170 VDD.n9830 VDD.n9827 4.5005
R15171 VDD.n9797 VDD.n9796 4.5005
R15172 VDD.n9814 VDD.n9500 4.5005
R15173 VDD.n9816 VDD.n9477 4.5005
R15174 VDD.n9491 VDD.n9477 4.5005
R15175 VDD.n9824 VDD.n9477 4.5005
R15176 VDD.n9778 VDD.n9508 4.5005
R15177 VDD.n9788 VDD.n9508 4.5005
R15178 VDD.n9795 VDD.n9508 4.5005
R15179 VDD.n9794 VDD.n9510 4.5005
R15180 VDD.n9796 VDD.n9498 4.5005
R15181 VDD.n9506 VDD.n9498 4.5005
R15182 VDD.n9815 VDD.n9498 4.5005
R15183 VDD.n9770 VDD.n9769 4.5005
R15184 VDD.n9770 VDD.n9524 4.5005
R15185 VDD.n9779 VDD.n9778 4.5005
R15186 VDD.n9751 VDD.n9750 4.5005
R15187 VDD.n9587 VDD.n9553 4.5005
R15188 VDD.n9743 VDD.n9553 4.5005
R15189 VDD.n9599 VDD.n9598 4.5005
R15190 VDD.n9600 VDD.n9599 4.5005
R15191 VDD.n9599 VDD.n9588 4.5005
R15192 VDD.n9582 VDD.n9581 4.5005
R15193 VDD.n11021 VDD.n8738 4.5005
R15194 VDD.n11022 VDD.n11021 4.5005
R15195 VDD.n11023 VDD.n8738 4.5005
R15196 VDD.n9164 VDD.n9079 4.5005
R15197 VDD.n9187 VDD.n9164 4.5005
R15198 VDD.n9186 VDD.n9079 4.5005
R15199 VDD.n9188 VDD.n9187 4.5005
R15200 VDD.n9187 VDD.n9186 4.5005
R15201 VDD.n9749 VDD.n9552 4.5005
R15202 VDD.n9749 VDD.n9551 4.5005
R15203 VDD.n9587 VDD.n9551 4.5005
R15204 VDD.n9750 VDD.n9541 4.5005
R15205 VDD.n9550 VDD.n9541 4.5005
R15206 VDD.n9768 VDD.n9541 4.5005
R15207 VDD.n9768 VDD.n9767 4.5005
R15208 VDD.n9769 VDD.n9520 4.5005
R15209 VDD.n9534 VDD.n9520 4.5005
R15210 VDD.n9777 VDD.n9520 4.5005
R15211 VDD.n9758 VDD.n9542 4.5005
R15212 VDD.n9767 VDD.n9766 4.5005
R15213 VDD.n9735 VDD.n9551 4.5005
R15214 VDD.n9598 VDD.n9597 4.5005
R15215 VDD.n11022 VDD.n8740 4.5005
R15216 VDD.n8740 VDD.n8738 4.5005
R15217 VDD.n9188 VDD.n9079 4.5005
R15218 VDD.n11023 VDD.n11022 4.5005
R15219 VDD.n9610 VDD.n9609 4.5005
R15220 VDD.n9588 VDD.n9581 4.5005
R15221 VDD.n9747 VDD.n9746 4.5005
R15222 VDD.n9777 VDD.n9776 4.5005
R15223 VDD.n9539 VDD.n9538 4.5005
R15224 VDD.n9793 VDD.n9792 4.5005
R15225 VDD.n9795 VDD.n9794 4.5005
R15226 VDD.n9805 VDD.n9499 4.5005
R15227 VDD.n9815 VDD.n9814 4.5005
R15228 VDD.n9824 VDD.n9823 4.5005
R15229 VDD.n9496 VDD.n9495 4.5005
R15230 VDD.n10896 VDD.n10668 4.5005
R15231 VDD.n10895 VDD.n10894 4.5005
R15232 VDD.n10775 VDD.n10774 4.5005
R15233 VDD.n6574 VDD.n6572 4.5005
R15234 VDD.n5776 VDD.n5775 4.5005
R15235 VDD.n4136 VDD.n4135 4.5005
R15236 VDD.n2496 VDD.n2495 4.5005
R15237 VDD.n8552 VDD.n7776 4.4978
R15238 VDD.n9975 VDD.n9972 4.48249
R15239 VDD.n11680 VDD.n7595 4.47034
R15240 VDD.n11685 VDD.n7592 4.47034
R15241 VDD.n11734 VDD.n7565 4.47034
R15242 VDD.n11742 VDD.n7561 4.47034
R15243 VDD.n11794 VDD.n7533 4.47034
R15244 VDD.n11799 VDD.n7530 4.47034
R15245 VDD.n11848 VDD.n7503 4.47034
R15246 VDD.n11856 VDD.n7499 4.47034
R15247 VDD.n11908 VDD.n7471 4.47034
R15248 VDD.n11913 VDD.n7468 4.47034
R15249 VDD.n11962 VDD.n7441 4.47034
R15250 VDD.n11970 VDD.n7437 4.47034
R15251 VDD.n12022 VDD.n7409 4.47034
R15252 VDD.n12027 VDD.n7406 4.47034
R15253 VDD.n12073 VDD.n7379 4.47034
R15254 VDD.n12079 VDD.n7376 4.47034
R15255 VDD.n11591 VDD.n11590 4.44682
R15256 VDD.n6942 VDD.n6935 4.4118
R15257 VDD.n12355 VDD.n6980 4.4118
R15258 VDD.n12307 VDD.n12306 4.4118
R15259 VDD.n7063 VDD.n7057 4.4118
R15260 VDD.n7171 VDD.n7170 4.4118
R15261 VDD.n7227 VDD.n7088 4.4118
R15262 VDD.n7276 VDD.n7270 4.4118
R15263 VDD.n12178 VDD.n7313 4.4118
R15264 VDD.n12484 VDD.n6567 4.38481
R15265 VDD.n7749 VDD.n7748 4.36497
R15266 VDD.n10110 VDD.n10097 4.35817
R15267 VDD.n8560 VDD.n7770 4.3536
R15268 VDD.n10965 VDD.n9218 4.31361
R15269 VDD.n10967 VDD.n9217 4.31361
R15270 VDD.n10972 VDD.n9209 4.31361
R15271 VDD.n11025 VDD.n11024 4.31361
R15272 VDD.n10993 VDD.n8731 4.31361
R15273 VDD.n8742 VDD.n8728 4.31361
R15274 VDD.n10469 VDD.n10448 4.31361
R15275 VDD.n10482 VDD.n10481 4.31361
R15276 VDD.n10478 VDD.n10477 4.31361
R15277 VDD.n10430 VDD.n10426 4.31327
R15278 VDD.n7957 VDD.n7827 4.31208
R15279 VDD.n7949 VDD.n7948 4.31208
R15280 VDD.n7907 VDD.n7906 4.31208
R15281 VDD.n7898 VDD.n7867 4.31208
R15282 VDD.n11471 VDD.n11470 4.31208
R15283 VDD.n11483 VDD.n7700 4.31208
R15284 VDD.n11529 VDD.n11528 4.31208
R15285 VDD.n11538 VDD.n7668 4.31208
R15286 VDD.n8119 VDD.n8091 4.30941
R15287 VDD.n6971 VDD.n6970 4.26717
R15288 VDD.n12319 VDD.n7006 4.26717
R15289 VDD.n12273 VDD.n7047 4.26717
R15290 VDD.n7155 VDD.n7154 4.26717
R15291 VDD.n7209 VDD.n7094 4.26717
R15292 VDD.n12240 VDD.n7260 4.26717
R15293 VDD.n7304 VDD.n7303 4.26717
R15294 VDD.n12142 VDD.n7339 4.26717
R15295 VDD.n8539 VDD.n7784 4.26717
R15296 VDD.n8520 VDD.n7796 4.26717
R15297 VDD.n11646 VDD.n11645 4.24471
R15298 VDD.n10546 VDD.n10540 4.23768
R15299 VDD.n9635 VDD.n9562 4.23768
R15300 VDD.n10734 VDD.n10733 4.23768
R15301 VDD.n8890 VDD.n8887 4.23768
R15302 VDD.n10042 VDD.n10040 4.23684
R15303 VDD.n10601 VDD.n10599 4.23684
R15304 VDD.n9372 VDD.n9369 4.23684
R15305 VDD.n8549 VDD.n8548 4.22104
R15306 VDD.n11673 VDD.n11672 4.19944
R15307 VDD.n11684 VDD.n7593 4.19944
R15308 VDD.n11731 VDD.n11730 4.19944
R15309 VDD.n11744 VDD.n11743 4.19944
R15310 VDD.n11787 VDD.n11786 4.19944
R15311 VDD.n11798 VDD.n7531 4.19944
R15312 VDD.n11845 VDD.n11844 4.19944
R15313 VDD.n11858 VDD.n11857 4.19944
R15314 VDD.n11901 VDD.n11900 4.19944
R15315 VDD.n11912 VDD.n7469 4.19944
R15316 VDD.n11959 VDD.n11958 4.19944
R15317 VDD.n11972 VDD.n11971 4.19944
R15318 VDD.n12015 VDD.n12014 4.19944
R15319 VDD.n12026 VDD.n7407 4.19944
R15320 VDD.n12074 VDD.n12072 4.19944
R15321 VDD.n12088 VDD.n7374 4.19944
R15322 VDD.n9174 VDD.n9169 4.18565
R15323 VDD.n11026 VDD.n8727 4.18565
R15324 VDD.n11596 VDD.n7638 4.17734
R15325 VDD.n11633 VDD.n7618 4.17734
R15326 VDD.n6555 VDD.n5780 4.17441
R15327 VDD.n5701 VDD.n4926 4.17441
R15328 VDD.n4915 VDD.n4140 4.17441
R15329 VDD.n4061 VDD.n3286 4.17441
R15330 VDD.n3275 VDD.n2500 4.17441
R15331 VDD.n2420 VDD.n1645 4.17441
R15332 VDD.n1224 VDD.n1221 4.17441
R15333 VDD.n778 VDD.n775 4.17441
R15334 VDD.n10061 VDD.n10030 4.14168
R15335 VDD.n10103 VDD.n10095 4.14168
R15336 VDD.n10622 VDD.n10589 4.14168
R15337 VDD.n10561 VDD.n10504 4.14168
R15338 VDD.n9595 VDD.n9594 4.14168
R15339 VDD.n9724 VDD.n9676 4.14168
R15340 VDD.n10822 VDD.n10821 4.14168
R15341 VDD.n10766 VDD.n10765 4.14168
R15342 VDD.n8920 VDD.n8917 4.14168
R15343 VDD.n8928 VDD.n8927 4.14168
R15344 VDD.n8949 VDD.n8948 4.14168
R15345 VDD.n9035 VDD.n9034 4.14168
R15346 VDD.n9048 VDD.n9047 4.14168
R15347 VDD.n8852 VDD.n8851 4.14168
R15348 VDD.n8817 VDD.n8816 4.14168
R15349 VDD.n8808 VDD.n8795 4.14168
R15350 VDD.n9018 VDD.n9017 4.14168
R15351 VDD.n8906 VDD.n8897 4.14168
R15352 VDD.n8903 VDD.n8760 4.14168
R15353 VDD.n9304 VDD.n9303 4.14168
R15354 VDD.n9310 VDD.n9253 4.14168
R15355 VDD.n9293 VDD.n9292 4.14168
R15356 VDD.n9336 VDD.n9330 4.14168
R15357 VDD.n10926 VDD.n9328 4.14168
R15358 VDD.n9383 VDD.n9380 4.14168
R15359 VDD.n9387 VDD.n9386 4.14168
R15360 VDD.n9424 VDD.n9401 4.14168
R15361 VDD.n9424 VDD.n9402 4.14168
R15362 VDD.n8521 VDD.n7794 4.14168
R15363 VDD.n8515 VDD.n7799 4.14168
R15364 VDD.n8149 VDD.n8148 4.13172
R15365 VDD.n8157 VDD.n8156 4.13172
R15366 VDD.n8151 VDD.n7745 4.13172
R15367 VDD.n11395 VDD.n11394 4.13172
R15368 VDD.n8667 VDD.n8666 4.13172
R15369 VDD.n11388 VDD.n8672 4.13172
R15370 VDD.n11071 VDD.n11070 4.13172
R15371 VDD.n11327 VDD.n11072 4.13172
R15372 VDD.n11085 VDD.n11084 4.13172
R15373 VDD.n11260 VDD.n11259 4.13172
R15374 VDD.n11188 VDD.n11187 4.13172
R15375 VDD.n11253 VDD.n11193 4.13172
R15376 VDD.n12400 VDD.n6943 4.12253
R15377 VDD.n12352 VDD.n12351 4.12253
R15378 VDD.n7024 VDD.n7018 4.12253
R15379 VDD.n12256 VDD.n7064 4.12253
R15380 VDD.n7176 VDD.n7110 4.12253
R15381 VDD.n7231 VDD.n7230 4.12253
R15382 VDD.n12223 VDD.n7277 4.12253
R15383 VDD.n12175 VDD.n12174 4.12253
R15384 VDD.n11180 VDD.t49 4.10046
R15385 VDD.n12418 VDD.n6925 4.08166
R15386 VDD.n8163 VDD.n8161 4.06399
R15387 VDD.n8678 VDD.n8677 4.06399
R15388 VDD.n11332 VDD.n11331 4.06399
R15389 VDD.n11199 VDD.n11198 4.06399
R15390 VDD.n12407 VDD.n12406 4.05022
R15391 VDD.n7958 VDD.n7825 4.04261
R15392 VDD.n7944 VDD.n7834 4.04261
R15393 VDD.n7911 VDD.n7858 4.04261
R15394 VDD.n7897 VDD.n7869 4.04261
R15395 VDD.n11469 VDD.n7707 4.04261
R15396 VDD.n11482 VDD.n7701 4.04261
R15397 VDD.n7680 VDD.n7675 4.04261
R15398 VDD.n11540 VDD.n11539 4.04261
R15399 VDD.n11581 VDD.n7645 4.04261
R15400 VDD.n9982 VDD.n9904 4.03708
R15401 VDD.n9982 VDD.n9905 4.03708
R15402 VDD.n12781 VDD 3.99913
R15403 VDD.n12373 VDD.n6965 3.9779
R15404 VDD.n12323 VDD.n12322 3.9779
R15405 VDD.n12274 VDD.n7044 3.9779
R15406 VDD.n7150 VDD.n7118 3.9779
R15407 VDD.n7208 VDD.n7096 3.9779
R15408 VDD.n12241 VDD.n7076 3.9779
R15409 VDD.n12196 VDD.n7299 3.9779
R15410 VDD.n12146 VDD.n12145 3.9779
R15411 VDD.t49 VDD.n11179 3.9682
R15412 VDD.n8540 VDD.n7780 3.94428
R15413 VDD.n8091 VDD.n8090 3.92921
R15414 VDD.n8205 VDD.n8085 3.92921
R15415 VDD.n8206 VDD.n8083 3.92921
R15416 VDD.n8035 VDD.n8032 3.92921
R15417 VDD.n8286 VDD.n8029 3.92921
R15418 VDD.n8027 VDD.n8023 3.92921
R15419 VDD.n8359 VDD.n8352 3.92921
R15420 VDD.n8466 VDD.n8361 3.92921
R15421 VDD.n8366 VDD.n8364 3.92921
R15422 VDD.n11671 VDD.n7600 3.92854
R15423 VDD.n11691 VDD.n7588 3.92854
R15424 VDD.n7572 VDD.n7567 3.92854
R15425 VDD.n11749 VDD.n7558 3.92854
R15426 VDD.n11785 VDD.n7538 3.92854
R15427 VDD.n11805 VDD.n7526 3.92854
R15428 VDD.n7510 VDD.n7505 3.92854
R15429 VDD.n11863 VDD.n7496 3.92854
R15430 VDD.n11899 VDD.n7476 3.92854
R15431 VDD.n11919 VDD.n7464 3.92854
R15432 VDD.n7448 VDD.n7443 3.92854
R15433 VDD.n11977 VDD.n7434 3.92854
R15434 VDD.n12013 VDD.n7414 3.92854
R15435 VDD.n12033 VDD.n7402 3.92854
R15436 VDD.n7386 VDD.n7381 3.92854
R15437 VDD.n11595 VDD.n7639 3.90787
R15438 VDD.n11637 VDD.n11636 3.90787
R15439 VDD.n12681 VDD.n12680 3.89763
R15440 VDD.n6722 VDD.n6713 3.89763
R15441 VDD.n12674 VDD.n6720 3.89763
R15442 VDD.n6747 VDD.n6721 3.89763
R15443 VDD.n12668 VDD.n6748 3.89763
R15444 VDD.n6753 VDD.n6749 3.89763
R15445 VDD.n12662 VDD.n6754 3.89763
R15446 VDD.n10244 VDD.n10243 3.89763
R15447 VDD.n12656 VDD.n6758 3.89763
R15448 VDD.n6763 VDD.n6759 3.89763
R15449 VDD.n12650 VDD.n6764 3.89763
R15450 VDD.n6769 VDD.n6765 3.89763
R15451 VDD.n12644 VDD.n6770 3.89763
R15452 VDD.n6775 VDD.n6771 3.89763
R15453 VDD.n12638 VDD.n6776 3.89763
R15454 VDD.n6781 VDD.n6777 3.89763
R15455 VDD.n12632 VDD.n6782 3.89763
R15456 VDD.n6787 VDD.n6783 3.89763
R15457 VDD.n12626 VDD.n6788 3.89763
R15458 VDD.n10225 VDD.n6789 3.89763
R15459 VDD.n6797 VDD.n6793 3.89763
R15460 VDD.n12614 VDD.n6798 3.89763
R15461 VDD.n6803 VDD.n6799 3.89763
R15462 VDD.n12608 VDD.n6804 3.89763
R15463 VDD.n6809 VDD.n6805 3.89763
R15464 VDD.n12602 VDD.n6810 3.89763
R15465 VDD.n6815 VDD.n6811 3.89763
R15466 VDD.n12596 VDD.n6816 3.89763
R15467 VDD.n10212 VDD.n10211 3.89763
R15468 VDD.n12590 VDD.n6820 3.89763
R15469 VDD.n10335 VDD.n10334 3.89763
R15470 VDD.n12584 VDD.n6824 3.89763
R15471 VDD.n6829 VDD.n6825 3.89763
R15472 VDD.n12578 VDD.n6830 3.89763
R15473 VDD.n6835 VDD.n6831 3.89763
R15474 VDD.n12572 VDD.n6836 3.89763
R15475 VDD.n6841 VDD.n6837 3.89763
R15476 VDD.n12566 VDD.n6842 3.89763
R15477 VDD.n6847 VDD.n6843 3.89763
R15478 VDD.n12560 VDD.n6848 3.89763
R15479 VDD.n10192 VDD.n6849 3.89763
R15480 VDD.n6857 VDD.n6853 3.89763
R15481 VDD.n12548 VDD.n6858 3.89763
R15482 VDD.n6863 VDD.n6859 3.89763
R15483 VDD.n12542 VDD.n6864 3.89763
R15484 VDD.n6869 VDD.n6865 3.89763
R15485 VDD.n12536 VDD.n6870 3.89763
R15486 VDD.n10183 VDD.n10182 3.89763
R15487 VDD.n12530 VDD.n6874 3.89763
R15488 VDD.n6879 VDD.n6875 3.89763
R15489 VDD.n12524 VDD.n6880 3.89763
R15490 VDD.n6885 VDD.n6881 3.89763
R15491 VDD.n12518 VDD.n6886 3.89763
R15492 VDD.n6891 VDD.n6887 3.89763
R15493 VDD.n12512 VDD.n6892 3.89763
R15494 VDD.n6897 VDD.n6893 3.89763
R15495 VDD.n12506 VDD.n6898 3.89763
R15496 VDD.n6903 VDD.n6899 3.89763
R15497 VDD.n12500 VDD.n6904 3.89763
R15498 VDD.n10164 VDD.n6905 3.89763
R15499 VDD.n8525 VDD.n8524 3.8907
R15500 VDD.n8514 VDD.n7800 3.8907
R15501 VDD.n12496 VDD.n6907 3.87632
R15502 VDD.n12451 VDD.n12450 3.87632
R15503 VDD.n8603 VDD.n8602 3.86082
R15504 VDD.n11385 VDD.n11384 3.86082
R15505 VDD.n11316 VDD.n11086 3.86082
R15506 VDD.n11250 VDD.n11249 3.86082
R15507 VDD.n12399 VDD.n6944 3.83327
R15508 VDD.n6986 VDD.n6982 3.83327
R15509 VDD.n12300 VDD.n7025 3.83327
R15510 VDD.n12255 VDD.n7065 3.83327
R15511 VDD.n7177 VDD.n7108 3.83327
R15512 VDD.n7235 VDD.n7086 3.83327
R15513 VDD.n12222 VDD.n7278 3.83327
R15514 VDD.n7319 VDD.n7315 3.83327
R15515 VDD.n8145 VDD.n8142 3.79309
R15516 VDD.n8674 VDD.n8653 3.79309
R15517 VDD.n11093 VDD.n11092 3.79309
R15518 VDD.n11195 VDD.n11173 3.79309
R15519 VDD.n9972 VDD.n9971 3.79052
R15520 VDD.n6348 VDD.n5933 3.78485
R15521 VDD.n6335 VDD.n6009 3.78485
R15522 VDD.n6323 VDD.n6322 3.78485
R15523 VDD.n5494 VDD.n5079 3.78485
R15524 VDD.n5481 VDD.n5155 3.78485
R15525 VDD.n5469 VDD.n5468 3.78485
R15526 VDD.n4708 VDD.n4293 3.78485
R15527 VDD.n4695 VDD.n4369 3.78485
R15528 VDD.n4683 VDD.n4682 3.78485
R15529 VDD.n3854 VDD.n3439 3.78485
R15530 VDD.n3841 VDD.n3515 3.78485
R15531 VDD.n3829 VDD.n3828 3.78485
R15532 VDD.n3068 VDD.n2653 3.78485
R15533 VDD.n3055 VDD.n2729 3.78485
R15534 VDD.n3043 VDD.n3042 3.78485
R15535 VDD.n2213 VDD.n1798 3.78485
R15536 VDD.n2200 VDD.n1874 3.78485
R15537 VDD.n2188 VDD.n2187 3.78485
R15538 VDD.n1597 VDD.n1594 3.78485
R15539 VDD.n369 VDD.n366 3.78485
R15540 VDD.n7962 VDD.n7961 3.77313
R15541 VDD.n7943 VDD.n7837 3.77313
R15542 VDD.n7912 VDD.n7856 3.77313
R15543 VDD.n7894 VDD.n7893 3.77313
R15544 VDD.n11466 VDD.n11465 3.77313
R15545 VDD.n11489 VDD.n7696 3.77313
R15546 VDD.n11522 VDD.n11521 3.77313
R15547 VDD.n11545 VDD.n7665 3.77313
R15548 VDD.n11578 VDD.n11577 3.77313
R15549 VDD.n10065 VDD.n10064 3.76521
R15550 VDD.n10626 VDD.n10586 3.76521
R15551 VDD.n10565 VDD.n10501 3.76521
R15552 VDD.n9975 VDD.n9974 3.76521
R15553 VDD.n9602 VDD.n9600 3.76521
R15554 VDD.n9614 VDD.n9574 3.76521
R15555 VDD.n9744 VDD.n9743 3.76521
R15556 VDD.n9717 VDD.n9716 3.76521
R15557 VDD.n9766 VDD.n9545 3.76521
R15558 VDD.n9535 VDD.n9534 3.76521
R15559 VDD.n9789 VDD.n9788 3.76521
R15560 VDD.n9802 VDD.n9500 3.76521
R15561 VDD.n9492 VDD.n9491 3.76521
R15562 VDD.n9862 VDD.n9860 3.76521
R15563 VDD.n10889 VDD.n10888 3.76521
R15564 VDD.n10868 VDD.n10867 3.76521
R15565 VDD.n10831 VDD.n10830 3.76521
R15566 VDD.n10757 VDD.n10756 3.76521
R15567 VDD.n10719 VDD.n10714 3.76521
R15568 VDD.n12422 VDD.n6909 3.76521
R15569 VDD.n12455 VDD.n12454 3.76521
R15570 VDD.n8120 VDD.n8119 3.73911
R15571 VDD.n8210 VDD.n8080 3.73911
R15572 VDD.n8282 VDD.n8034 3.73911
R15573 VDD.n8298 VDD.n8297 3.73911
R15574 VDD.n8476 VDD.n8351 3.73911
R15575 VDD.n8462 VDD.n8461 3.73911
R15576 VDD.n8598 VDD.n7749 3.70369
R15577 VDD.n9960 VDD.n9910 3.70003
R15578 VDD.n12374 VDD.n6962 3.68864
R15579 VDD.n7005 VDD.n7004 3.68864
R15580 VDD.n12278 VDD.n12277 3.68864
R15581 VDD.n7149 VDD.n7120 3.68864
R15582 VDD.n7205 VDD.n7204 3.68864
R15583 VDD.n12245 VDD.n12244 3.68864
R15584 VDD.n12197 VDD.n7296 3.68864
R15585 VDD.n7338 VDD.n7337 3.68864
R15586 VDD.n5745 VDD.n5744 3.67828
R15587 VDD.n4105 VDD.n4104 3.67828
R15588 VDD.n2464 VDD.n2463 3.67828
R15589 VDD.n824 VDD.n823 3.67828
R15590 VDD.n11668 VDD.n11667 3.65764
R15591 VDD.n11693 VDD.n11692 3.65764
R15592 VDD.n11724 VDD.n11723 3.65764
R15593 VDD.n11748 VDD.n7559 3.65764
R15594 VDD.n11782 VDD.n11781 3.65764
R15595 VDD.n11807 VDD.n11806 3.65764
R15596 VDD.n11838 VDD.n11837 3.65764
R15597 VDD.n11862 VDD.n7497 3.65764
R15598 VDD.n11896 VDD.n11895 3.65764
R15599 VDD.n11921 VDD.n11920 3.65764
R15600 VDD.n11952 VDD.n11951 3.65764
R15601 VDD.n11976 VDD.n7435 3.65764
R15602 VDD.n12010 VDD.n12009 3.65764
R15603 VDD.n12035 VDD.n12034 3.65764
R15604 VDD.n12066 VDD.n12065 3.65764
R15605 VDD.n6156 VDD.n6099 3.64278
R15606 VDD.n5302 VDD.n5245 3.64278
R15607 VDD.n4516 VDD.n4459 3.64278
R15608 VDD.n3662 VDD.n3605 3.64278
R15609 VDD.n2876 VDD.n2819 3.64278
R15610 VDD.n2021 VDD.n1964 3.64278
R15611 VDD.n1311 VDD.n1304 3.64278
R15612 VDD.n83 VDD.n76 3.64278
R15613 VDD.n8529 VDD.n7791 3.63972
R15614 VDD.n8511 VDD.n8510 3.63972
R15615 VDD.n11602 VDD.n7634 3.63839
R15616 VDD.n11629 VDD.n7617 3.63839
R15617 VDD.n12554 VDD.t152 3.59785
R15618 VDD.n11445 VDD.n7722 3.58992
R15619 VDD.n8690 VDD.n8689 3.58992
R15620 VDD.n11313 VDD.n11312 3.58992
R15621 VDD.n11211 VDD.n11210 3.58992
R15622 VDD.n12396 VDD.n12395 3.544
R15623 VDD.n12345 VDD.n6987 3.544
R15624 VDD.n12299 VDD.n7026 3.544
R15625 VDD.n12252 VDD.n12251 3.544
R15626 VDD.n7181 VDD.n7180 3.544
R15627 VDD.n7236 VDD.n7084 3.544
R15628 VDD.n12219 VDD.n12218 3.544
R15629 VDD.n12168 VDD.n7320 3.544
R15630 VDD.n9955 VDD 3.53589
R15631 VDD.n8169 VDD.n8140 3.52219
R15632 VDD.n8651 VDD.n8637 3.52219
R15633 VDD.n11091 VDD.n11058 3.52219
R15634 VDD.n11171 VDD.n11157 3.52219
R15635 VDD.n7966 VDD.n7821 3.50366
R15636 VDD.n7940 VDD.n7939 3.50366
R15637 VDD.n7916 VDD.n7915 3.50366
R15638 VDD.n7873 VDD.n7871 3.50366
R15639 VDD.n7714 VDD.n7709 3.50366
R15640 VDD.n11491 VDD.n11490 3.50366
R15641 VDD.n11516 VDD.n7679 3.50366
R15642 VDD.n11544 VDD.n7666 3.50366
R15643 VDD.n7652 VDD.n7647 3.50366
R15644 VDD.n8078 VDD.n8074 3.48565
R15645 VDD.n8041 VDD.n8040 3.48565
R15646 VDD.n8302 VDD.n8301 3.48565
R15647 VDD.n8480 VDD.n8479 3.48565
R15648 VDD.n8376 VDD.n8375 3.48565
R15649 VDD.n8565 VDD.n8564 3.48565
R15650 VDD.n9950 VDD 3.44516
R15651 VDD.n2476 VDD.n2474 3.43528
R15652 VDD.n836 VDD.n834 3.43528
R15653 VDD.n9283 VDD.n9282 3.42768
R15654 VDD.n9413 VDD.n9412 3.42768
R15655 VDD.n9664 VDD.n9662 3.42765
R15656 VDD.n10807 VDD.n10805 3.42765
R15657 VDD.n9003 VDD.n9001 3.42765
R15658 VDD.n9653 VDD.n9652 3.42683
R15659 VDD.n10796 VDD.n10795 3.42683
R15660 VDD.n8872 VDD.n8871 3.42683
R15661 VDD.n10450 VDD.n10442 3.42673
R15662 VDD.n11010 VDD.n11009 3.42318
R15663 VDD.n11005 VDD.n8748 3.42286
R15664 VDD.n6058 VDD.n6055 3.42221
R15665 VDD.n5204 VDD.n5201 3.42221
R15666 VDD.n4418 VDD.n4415 3.42221
R15667 VDD.n3564 VDD.n3561 3.42221
R15668 VDD.n2778 VDD.n2775 3.42221
R15669 VDD.n1923 VDD.n1920 3.42221
R15670 VDD.n980 VDD.n977 3.42221
R15671 VDD.n534 VDD.n531 3.42221
R15672 VDD.n10487 VDD.n10486 3.41892
R15673 VDD.n11012 VDD.n11011 3.41503
R15674 VDD.n10486 VDD.n10485 3.4105
R15675 VDD.n8746 VDD.n8745 3.4105
R15676 VDD.n11004 VDD.n11003 3.4105
R15677 VDD.n11004 VDD.n9066 3.4105
R15678 VDD.n9067 VDD.n9066 3.4105
R15679 VDD.n11003 VDD.n9067 3.4105
R15680 VDD.n9066 VDD.n8752 3.4105
R15681 VDD.n11003 VDD.n8752 3.4105
R15682 VDD.n11006 VDD.n11005 3.4105
R15683 VDD.n11007 VDD.n8752 3.4105
R15684 VDD.n11008 VDD.n11007 3.4105
R15685 VDD.n11019 VDD.n11015 3.4105
R15686 VDD.n11019 VDD.n11018 3.4105
R15687 VDD.n11019 VDD.n8743 3.4105
R15688 VDD.n11018 VDD.n8741 3.4105
R15689 VDD.n8744 VDD.n8739 3.4105
R15690 VDD.n10898 VDD.n10897 3.4105
R15691 VDD.n9867 VDD.n9866 3.4105
R15692 VDD.n10898 VDD.n10669 3.4105
R15693 VDD.n10898 VDD.n10668 3.4105
R15694 VDD.n9469 VDD.n9463 3.4105
R15695 VDD.n9469 VDD.n9464 3.4105
R15696 VDD.n9469 VDD.n9462 3.4105
R15697 VDD.n9469 VDD.n9465 3.4105
R15698 VDD.n9469 VDD.n9461 3.4105
R15699 VDD.n9469 VDD.n9466 3.4105
R15700 VDD.n9469 VDD.n9460 3.4105
R15701 VDD.n9469 VDD.n9467 3.4105
R15702 VDD.n9887 VDD.n9469 3.4105
R15703 VDD.n9888 VDD.n9463 3.4105
R15704 VDD.n9888 VDD.n9464 3.4105
R15705 VDD.n9888 VDD.n9462 3.4105
R15706 VDD.n9888 VDD.n9465 3.4105
R15707 VDD.n9888 VDD.n9461 3.4105
R15708 VDD.n9888 VDD.n9466 3.4105
R15709 VDD.n9888 VDD.n9460 3.4105
R15710 VDD.n9888 VDD.n9467 3.4105
R15711 VDD.n9888 VDD.n9887 3.4105
R15712 VDD.n9465 VDD.n9458 3.4105
R15713 VDD.n9461 VDD.n9458 3.4105
R15714 VDD.n9466 VDD.n9458 3.4105
R15715 VDD.n9460 VDD.n9458 3.4105
R15716 VDD.n9467 VDD.n9458 3.4105
R15717 VDD.n9885 VDD.n9458 3.4105
R15718 VDD.n9887 VDD.n9458 3.4105
R15719 VDD.n9462 VDD.n9458 3.4105
R15720 VDD.n9464 VDD.n9458 3.4105
R15721 VDD.n9463 VDD.n9458 3.4105
R15722 VDD.n9470 VDD.n9462 3.4105
R15723 VDD.n9470 VDD.n9464 3.4105
R15724 VDD.n9470 VDD.n9463 3.4105
R15725 VDD.n9474 VDD.n9463 3.4105
R15726 VDD.n9474 VDD.n9464 3.4105
R15727 VDD.n9474 VDD.n9462 3.4105
R15728 VDD.n9474 VDD.n9465 3.4105
R15729 VDD.n9474 VDD.n9461 3.4105
R15730 VDD.n9474 VDD.n9466 3.4105
R15731 VDD.n9474 VDD.n9460 3.4105
R15732 VDD.n9474 VDD.n9467 3.4105
R15733 VDD.n9474 VDD.n9471 3.4105
R15734 VDD.n9474 VDD.n9468 3.4105
R15735 VDD.n9887 VDD.n9886 3.4105
R15736 VDD.n9886 VDD.n9885 3.4105
R15737 VDD.n9886 VDD.n9467 3.4105
R15738 VDD.n9886 VDD.n9460 3.4105
R15739 VDD.n9886 VDD.n9466 3.4105
R15740 VDD.n9886 VDD.n9461 3.4105
R15741 VDD.n9886 VDD.n9465 3.4105
R15742 VDD.n9886 VDD.n9462 3.4105
R15743 VDD.n9886 VDD.n9464 3.4105
R15744 VDD.n9886 VDD.n9463 3.4105
R15745 VDD.n9470 VDD.n9468 3.4105
R15746 VDD.n9471 VDD.n9470 3.4105
R15747 VDD.n9470 VDD.n9467 3.4105
R15748 VDD.n9470 VDD.n9460 3.4105
R15749 VDD.n9470 VDD.n9466 3.4105
R15750 VDD.n9470 VDD.n9461 3.4105
R15751 VDD.n9470 VDD.n9465 3.4105
R15752 VDD.n10900 VDD.n10662 3.4105
R15753 VDD.n10662 VDD.n9452 3.4105
R15754 VDD.n10902 VDD.n9903 3.4105
R15755 VDD.n9903 VDD.n9452 3.4105
R15756 VDD.n9347 VDD.n9230 3.4105
R15757 VDD.n10906 VDD.n9347 3.4105
R15758 VDD.n9347 VDD.n9238 3.4105
R15759 VDD.n9347 VDD.n9235 3.4105
R15760 VDD.n9347 VDD.n9239 3.4105
R15761 VDD.n9347 VDD.n9234 3.4105
R15762 VDD.n9347 VDD.n9240 3.4105
R15763 VDD.n9347 VDD.n9241 3.4105
R15764 VDD.n10904 VDD.n9347 3.4105
R15765 VDD.n9247 VDD.n9238 3.4105
R15766 VDD.n9247 VDD.n9235 3.4105
R15767 VDD.n9247 VDD.n9239 3.4105
R15768 VDD.n9247 VDD.n9234 3.4105
R15769 VDD.n9247 VDD.n9240 3.4105
R15770 VDD.n9247 VDD.n9233 3.4105
R15771 VDD.n9247 VDD.n9241 3.4105
R15772 VDD.n10942 VDD.n9247 3.4105
R15773 VDD.n10943 VDD.n9236 3.4105
R15774 VDD.n9236 VDD.n9229 3.4105
R15775 VDD.n10942 VDD.n9229 3.4105
R15776 VDD.n9241 VDD.n9229 3.4105
R15777 VDD.n9240 VDD.n9229 3.4105
R15778 VDD.n9234 VDD.n9229 3.4105
R15779 VDD.n9239 VDD.n9229 3.4105
R15780 VDD.n9235 VDD.n9229 3.4105
R15781 VDD.n9238 VDD.n9229 3.4105
R15782 VDD.n10906 VDD.n9229 3.4105
R15783 VDD.n10944 VDD.n9229 3.4105
R15784 VDD.n9232 VDD.n9229 3.4105
R15785 VDD.n10905 VDD.n10904 3.4105
R15786 VDD.n10905 VDD.n9241 3.4105
R15787 VDD.n10905 VDD.n9233 3.4105
R15788 VDD.n10905 VDD.n9240 3.4105
R15789 VDD.n10905 VDD.n9234 3.4105
R15790 VDD.n10905 VDD.n9239 3.4105
R15791 VDD.n10905 VDD.n9235 3.4105
R15792 VDD.n10905 VDD.n9238 3.4105
R15793 VDD.n10906 VDD.n10905 3.4105
R15794 VDD.n10905 VDD.n9230 3.4105
R15795 VDD.n10944 VDD.n10943 3.4105
R15796 VDD.n10943 VDD.n9238 3.4105
R15797 VDD.n10943 VDD.n9235 3.4105
R15798 VDD.n10943 VDD.n9239 3.4105
R15799 VDD.n10943 VDD.n9234 3.4105
R15800 VDD.n10943 VDD.n9240 3.4105
R15801 VDD.n10943 VDD.n9233 3.4105
R15802 VDD.n10943 VDD.n9241 3.4105
R15803 VDD.n10943 VDD.n9232 3.4105
R15804 VDD.n10906 VDD.n9243 3.4105
R15805 VDD.n9243 VDD.n9238 3.4105
R15806 VDD.n9243 VDD.n9235 3.4105
R15807 VDD.n9243 VDD.n9239 3.4105
R15808 VDD.n9243 VDD.n9234 3.4105
R15809 VDD.n9243 VDD.n9240 3.4105
R15810 VDD.n9243 VDD.n9233 3.4105
R15811 VDD.n9243 VDD.n9241 3.4105
R15812 VDD.n10942 VDD.n9243 3.4105
R15813 VDD.n10943 VDD.n10942 3.4105
R15814 VDD.n10902 VDD.n9899 3.4105
R15815 VDD.n10903 VDD.n9452 3.4105
R15816 VDD.n10903 VDD.n9451 3.4105
R15817 VDD.n9899 VDD.n9452 3.4105
R15818 VDD.n10903 VDD.n10902 3.4105
R15819 VDD.n10663 VDD.n10661 3.4105
R15820 VDD.n10663 VDD.n9451 3.4105
R15821 VDD.n10663 VDD.n9452 3.4105
R15822 VDD.n10901 VDD.n9452 3.4105
R15823 VDD.n10902 VDD.n10901 3.4105
R15824 VDD.n10901 VDD.n10900 3.4105
R15825 VDD.n10661 VDD.n9899 3.4105
R15826 VDD.n10904 VDD.n9243 3.4105
R15827 VDD.n10904 VDD.n9247 3.4105
R15828 VDD.n10657 VDD.n9996 3.4105
R15829 VDD.n9996 VDD.n9985 3.4105
R15830 VDD.n9996 VDD.n9993 3.4105
R15831 VDD.n9996 VDD.n9986 3.4105
R15832 VDD.n9996 VDD.n9989 3.4105
R15833 VDD.n9996 VDD.n9988 3.4105
R15834 VDD.n9996 VDD.n9990 3.4105
R15835 VDD.n10650 VDD.n9996 3.4105
R15836 VDD.n9996 VDD.n9991 3.4105
R15837 VDD.n10657 VDD.n10656 3.4105
R15838 VDD.n10656 VDD.n9985 3.4105
R15839 VDD.n10656 VDD.n9993 3.4105
R15840 VDD.n10656 VDD.n9986 3.4105
R15841 VDD.n10656 VDD.n9989 3.4105
R15842 VDD.n10656 VDD.n9988 3.4105
R15843 VDD.n10656 VDD.n9990 3.4105
R15844 VDD.n10656 VDD.n9991 3.4105
R15845 VDD.n10656 VDD.n9992 3.4105
R15846 VDD.n10658 VDD.n9989 3.4105
R15847 VDD.n10658 VDD.n9988 3.4105
R15848 VDD.n10658 VDD.n9990 3.4105
R15849 VDD.n10658 VDD.n9991 3.4105
R15850 VDD.n10658 VDD.n9987 3.4105
R15851 VDD.n10658 VDD.n9992 3.4105
R15852 VDD.n10658 VDD.n9986 3.4105
R15853 VDD.n10658 VDD.n9993 3.4105
R15854 VDD.n10658 VDD.n9985 3.4105
R15855 VDD.n10658 VDD.n10657 3.4105
R15856 VDD.n10652 VDD.n9997 3.4105
R15857 VDD.n10652 VDD.n9994 3.4105
R15858 VDD.n10652 VDD.n9985 3.4105
R15859 VDD.n10652 VDD.n9993 3.4105
R15860 VDD.n10652 VDD.n9986 3.4105
R15861 VDD.n10652 VDD.n9989 3.4105
R15862 VDD.n10652 VDD.n9988 3.4105
R15863 VDD.n10652 VDD.n9990 3.4105
R15864 VDD.n10652 VDD.n10650 3.4105
R15865 VDD.n10652 VDD.n9991 3.4105
R15866 VDD.n10653 VDD.n10652 3.4105
R15867 VDD.n9987 VDD.n6569 3.4105
R15868 VDD.n9991 VDD.n6569 3.4105
R15869 VDD.n10650 VDD.n6569 3.4105
R15870 VDD.n9990 VDD.n6569 3.4105
R15871 VDD.n9988 VDD.n6569 3.4105
R15872 VDD.n9989 VDD.n6569 3.4105
R15873 VDD.n9986 VDD.n6569 3.4105
R15874 VDD.n9993 VDD.n6569 3.4105
R15875 VDD.n9985 VDD.n6569 3.4105
R15876 VDD.n10657 VDD.n6569 3.4105
R15877 VDD.n10654 VDD.n9986 3.4105
R15878 VDD.n10654 VDD.n9993 3.4105
R15879 VDD.n10654 VDD.n9985 3.4105
R15880 VDD.n10654 VDD.n9994 3.4105
R15881 VDD.n10654 VDD.n9997 3.4105
R15882 VDD.n10654 VDD.n10653 3.4105
R15883 VDD.n10654 VDD.n9991 3.4105
R15884 VDD.n10654 VDD.n10650 3.4105
R15885 VDD.n10654 VDD.n9990 3.4105
R15886 VDD.n10654 VDD.n9988 3.4105
R15887 VDD.n10654 VDD.n9989 3.4105
R15888 VDD.n10474 VDD.n10455 3.4105
R15889 VDD.n10474 VDD.n10453 3.4105
R15890 VDD.n10471 VDD.n10453 3.4105
R15891 VDD.n10453 VDD.n10443 3.4105
R15892 VDD.n10455 VDD.n10443 3.4105
R15893 VDD.n10473 VDD.n10443 3.4105
R15894 VDD.n10444 VDD.n10443 3.4105
R15895 VDD.n10473 VDD.n10458 3.4105
R15896 VDD.n10473 VDD.n10457 3.4105
R15897 VDD.n10473 VDD.n10456 3.4105
R15898 VDD.n10474 VDD.n10473 3.4105
R15899 VDD.n10475 VDD.n10474 3.4105
R15900 VDD.n12378 VDD.n12377 3.39937
R15901 VDD.n12329 VDD.n7000 3.39937
R15902 VDD.n7043 VDD.n7042 3.39937
R15903 VDD.n7146 VDD.n7145 3.39937
R15904 VDD.n7200 VDD.n7098 3.39937
R15905 VDD.n7255 VDD.n7075 3.39937
R15906 VDD.n12201 VDD.n12200 3.39937
R15907 VDD.n12152 VDD.n7333 3.39937
R15908 VDD.n6388 VDD.n5899 3.39504
R15909 VDD.n5534 VDD.n5045 3.39504
R15910 VDD.n4748 VDD.n4259 3.39504
R15911 VDD.n3894 VDD.n3405 3.39504
R15912 VDD.n3108 VDD.n2619 3.39504
R15913 VDD.n2253 VDD.n1764 3.39504
R15914 VDD.n1368 VDD.n1365 3.39504
R15915 VDD.n140 VDD.n137 3.39504
R15916 VDD.n9607 VDD.n9582 3.38874
R15917 VDD.n9607 VDD.n9583 3.38874
R15918 VDD.n9735 VDD.n9734 3.38874
R15919 VDD.n9721 VDD.n9720 3.38874
R15920 VDD.n9755 VDD.n9550 3.38874
R15921 VDD.n9529 VDD.n9524 3.38874
R15922 VDD.n9516 VDD.n9510 3.38874
R15923 VDD.n9800 VDD.n9506 3.38874
R15924 VDD.n9486 VDD.n9481 3.38874
R15925 VDD.n9864 VDD.n9836 3.38874
R15926 VDD.n10893 VDD.n10892 3.38874
R15927 VDD.n10871 VDD.n10694 3.38874
R15928 VDD.n10827 VDD.n10826 3.38874
R15929 VDD.n10761 VDD.n10705 3.38874
R15930 VDD.n10761 VDD.n10706 3.38874
R15931 VDD.n8935 VDD.n8934 3.38874
R15932 VDD.n8939 VDD.n8938 3.38874
R15933 VDD.n8944 VDD.n8943 3.38874
R15934 VDD.n9050 VDD.n8782 3.38874
R15935 VDD.n8842 VDD.n8841 3.38874
R15936 VDD.n8847 VDD.n8846 3.38874
R15937 VDD.n9032 VDD.n9031 3.38874
R15938 VDD.n9028 VDD.n9027 3.38874
R15939 VDD.n9023 VDD.n9022 3.38874
R15940 VDD.n9312 VDD.n9258 3.38874
R15941 VDD.n9270 VDD.n9267 3.38874
R15942 VDD.n9297 VDD.n9266 3.38874
R15943 VDD.n9442 VDD.n9360 3.38874
R15944 VDD.n9438 VDD.n9393 3.38874
R15945 VDD.n9429 VDD.n9396 3.38874
R15946 VDD.n9429 VDD.n9428 3.38874
R15947 VDD.n9140 VDD.n9139 3.38874
R15948 VDD.n8530 VDD.n7788 3.38874
R15949 VDD.n8507 VDD.n7802 3.38874
R15950 VDD.n7607 VDD.n7602 3.38674
R15951 VDD.n11698 VDD.n7585 3.38674
R15952 VDD.n11718 VDD.n7571 3.38674
R15953 VDD.n11755 VDD.n7554 3.38674
R15954 VDD.n7545 VDD.n7540 3.38674
R15955 VDD.n11812 VDD.n7523 3.38674
R15956 VDD.n11832 VDD.n7509 3.38674
R15957 VDD.n11869 VDD.n7492 3.38674
R15958 VDD.n7483 VDD.n7478 3.38674
R15959 VDD.n11926 VDD.n7461 3.38674
R15960 VDD.n11946 VDD.n7447 3.38674
R15961 VDD.n11983 VDD.n7430 3.38674
R15962 VDD.n7421 VDD.n7416 3.38674
R15963 VDD.n12040 VDD.n7399 3.38674
R15964 VDD.n12060 VDD.n7385 3.38674
R15965 VDD.n11604 VDD.n11603 3.36892
R15966 VDD.n11630 VDD.n11628 3.36892
R15967 VDD.n10477 VDD.n10449 3.33963
R15968 VDD.n10469 VDD.n10449 3.33963
R15969 VDD.n10469 VDD.n10446 3.33963
R15970 VDD.n10482 VDD.n10446 3.33963
R15971 VDD.n10436 VDD.n10435 3.33963
R15972 VDD.n10435 VDD.n10160 3.33963
R15973 VDD.n10496 VDD.n10160 3.33963
R15974 VDD.n10496 VDD.n10161 3.33963
R15975 VDD.n10972 VDD.n9210 3.33963
R15976 VDD.n10967 VDD.n9210 3.33963
R15977 VDD.n10967 VDD.n10966 3.33963
R15978 VDD.n10966 VDD.n10965 3.33963
R15979 VDD.n10951 VDD.n9219 3.33963
R15980 VDD.n10952 VDD.n10951 3.33963
R15981 VDD.n10952 VDD.n9224 3.33963
R15982 VDD.n10957 VDD.n9224 3.33963
R15983 VDD.n9181 VDD.n9166 3.33963
R15984 VDD.n9185 VDD.n9166 3.33963
R15985 VDD.n9185 VDD.n9077 3.33963
R15986 VDD.n9189 VDD.n9077 3.33963
R15987 VDD.n11024 VDD.n8735 3.33963
R15988 VDD.n8742 VDD.n8735 3.33963
R15989 VDD.n10994 VDD.n8742 3.33963
R15990 VDD.n10994 VDD.n10993 3.33963
R15991 VDD.n10987 VDD.n9068 3.33963
R15992 VDD.n11000 VDD.n9068 3.33963
R15993 VDD.n11000 VDD.n10999 3.33963
R15994 VDD.n10999 VDD.n9070 3.33963
R15995 VDD.n7726 VDD.n7723 3.31902
R15996 VDD.n8714 VDD.n8711 3.31902
R15997 VDD.n11110 VDD.n11109 3.31902
R15998 VDD.n11224 VDD.n11223 3.31902
R15999 VDD.n4116 VDD.n4114 3.29941
R16000 VDD.n7767 VDD.n7761 3.29555
R16001 VDD.n10046 VDD.n10045 3.2936
R16002 VDD.n10605 VDD.n10604 3.2936
R16003 VDD.n10543 VDD.n10538 3.2936
R16004 VDD.n9632 VDD.n9631 3.2936
R16005 VDD.n10736 VDD.n10726 3.2936
R16006 VDD.n8911 VDD.n8888 3.2936
R16007 VDD.n9374 VDD.n9364 3.2936
R16008 VDD.n6951 VDD.n6947 3.25474
R16009 VDD.n12344 VDD.n6988 3.25474
R16010 VDD.n12296 VDD.n12295 3.25474
R16011 VDD.n7128 VDD.n7068 3.25474
R16012 VDD.n7185 VDD.n7106 3.25474
R16013 VDD.n7240 VDD.n7239 3.25474
R16014 VDD.n7285 VDD.n7281 3.25474
R16015 VDD.n12167 VDD.n7321 3.25474
R16016 VDD.n12414 VDD.n6927 3.25377
R16017 VDD.n8174 VDD.n8172 3.25129
R16018 VDD.n11410 VDD.n8636 3.25129
R16019 VDD.n11056 VDD.n11042 3.25129
R16020 VDD.n11275 VDD.n11156 3.25129
R16021 VDD.n12479 VDD.n12478 3.24687
R16022 VDD.n12464 VDD.n12463 3.24687
R16023 VDD.n7967 VDD.n7819 3.23418
R16024 VDD.n7841 VDD.n7839 3.23418
R16025 VDD.n7920 VDD.n7852 3.23418
R16026 VDD.n7888 VDD.n7875 3.23418
R16027 VDD.n11459 VDD.n11458 3.23418
R16028 VDD.n11496 VDD.n7693 3.23418
R16029 VDD.n11517 VDD.n11515 3.23418
R16030 VDD.n11551 VDD.n7661 3.23418
R16031 VDD.n11571 VDD.n11570 3.23418
R16032 VDD.n8223 VDD.n8222 3.23218
R16033 VDD.n8270 VDD.n8044 3.23218
R16034 VDD.n8017 VDD.n8016 3.23218
R16035 VDD.n8347 VDD.n8344 3.23218
R16036 VDD.n8452 VDD.n8380 3.23218
R16037 VDD.n8416 VDD.n8415 3.23218
R16038 VDD.n5756 VDD.n5754 3.20702
R16039 VDD.n9183 VDD.n7735 3.17466
R16040 VDD.n9169 VDD.n9168 3.17466
R16041 VDD.n6361 VDD.n5916 3.17267
R16042 VDD.n6360 VDD.n6359 3.17267
R16043 VDD.n6358 VDD.n5921 3.17267
R16044 VDD.n5507 VDD.n5062 3.17267
R16045 VDD.n5506 VDD.n5505 3.17267
R16046 VDD.n5504 VDD.n5067 3.17267
R16047 VDD.n4721 VDD.n4276 3.17267
R16048 VDD.n4720 VDD.n4719 3.17267
R16049 VDD.n4718 VDD.n4281 3.17267
R16050 VDD.n3867 VDD.n3422 3.17267
R16051 VDD.n3866 VDD.n3865 3.17267
R16052 VDD.n3864 VDD.n3427 3.17267
R16053 VDD.n3081 VDD.n2636 3.17267
R16054 VDD.n3080 VDD.n3079 3.17267
R16055 VDD.n3078 VDD.n2641 3.17267
R16056 VDD.n2226 VDD.n1781 3.17267
R16057 VDD.n2225 VDD.n2224 3.17267
R16058 VDD.n2223 VDD.n1786 3.17267
R16059 VDD.n1579 VDD.n1576 3.17267
R16060 VDD.n1585 VDD.n1582 3.17267
R16061 VDD.n1591 VDD.n1588 3.17267
R16062 VDD.n351 VDD.n348 3.17267
R16063 VDD.n357 VDD.n354 3.17267
R16064 VDD.n363 VDD.n360 3.17267
R16065 VDD.n8498 VDD.n7988 3.16717
R16066 VDD.n10437 VDD.n10436 3.15412
R16067 VDD.n8534 VDD.n8533 3.13775
R16068 VDD.n8506 VDD.n7805 3.13775
R16069 VDD.n11661 VDD.n11660 3.11584
R16070 VDD.n11697 VDD.n7586 3.11584
R16071 VDD.n11719 VDD.n11717 3.11584
R16072 VDD.n11757 VDD.n11756 3.11584
R16073 VDD.n11775 VDD.n11774 3.11584
R16074 VDD.n11811 VDD.n7524 3.11584
R16075 VDD.n11833 VDD.n11831 3.11584
R16076 VDD.n11871 VDD.n11870 3.11584
R16077 VDD.n11889 VDD.n11888 3.11584
R16078 VDD.n11925 VDD.n7462 3.11584
R16079 VDD.n11947 VDD.n11945 3.11584
R16080 VDD.n11985 VDD.n11984 3.11584
R16081 VDD.n12003 VDD.n12002 3.11584
R16082 VDD.n12039 VDD.n7400 3.11584
R16083 VDD.n12061 VDD.n12059 3.11584
R16084 VDD.n6961 VDD.n6960 3.1101
R16085 VDD.n12330 VDD.n6997 3.1101
R16086 VDD.n12284 VDD.n7038 3.1101
R16087 VDD.n7140 VDD.n7122 3.1101
R16088 VDD.n7199 VDD.n7100 3.1101
R16089 VDD.n7256 VDD.n7254 3.1101
R16090 VDD.n7295 VDD.n7294 3.1101
R16091 VDD.n12153 VDD.n7330 3.1101
R16092 VDD.n12764 VDD.n6578 3.10907
R16093 VDD.n12764 VDD.n12763 3.10907
R16094 VDD.n12763 VDD.n6582 3.10907
R16095 VDD.n12757 VDD.n6582 3.10907
R16096 VDD.n12757 VDD.n12756 3.10907
R16097 VDD.n12756 VDD.n6584 3.10907
R16098 VDD.n12750 VDD.n6584 3.10907
R16099 VDD.n12750 VDD.n12749 3.10907
R16100 VDD.n12749 VDD.n6586 3.10907
R16101 VDD.n12743 VDD.n6586 3.10907
R16102 VDD.n12743 VDD.n12742 3.10907
R16103 VDD.n12742 VDD.n6588 3.10907
R16104 VDD.n12736 VDD.n6588 3.10907
R16105 VDD.n12736 VDD.n12735 3.10907
R16106 VDD.n12735 VDD.n6590 3.10907
R16107 VDD.n12729 VDD.n6590 3.10907
R16108 VDD.n12729 VDD.n12728 3.10907
R16109 VDD.n12728 VDD.n6592 3.10907
R16110 VDD.n12722 VDD.n6592 3.10907
R16111 VDD.n12722 VDD.n12721 3.10907
R16112 VDD.n12721 VDD.n6594 3.10907
R16113 VDD.n12715 VDD.n6594 3.10907
R16114 VDD.n12715 VDD.n12714 3.10907
R16115 VDD.n12714 VDD.n6596 3.10907
R16116 VDD.n5727 VDD.n5726 3.10102
R16117 VDD.n4087 VDD.n4086 3.10102
R16118 VDD.n2446 VDD.n2445 3.10102
R16119 VDD.n806 VDD.n805 3.10102
R16120 VDD.n11609 VDD.n7631 3.09945
R16121 VDD.n7625 VDD.n7620 3.09945
R16122 VDD.n9947 VDD.n9912 3.09792
R16123 VDD.n9926 VDD.n9922 3.09792
R16124 VDD.n5719 VDD.n5711 3.09792
R16125 VDD.n4079 VDD.n4071 3.09792
R16126 VDD.n2438 VDD.n2430 3.09792
R16127 VDD.n798 VDD.n790 3.09792
R16128 VDD.n8611 VDD.n8608 3.04812
R16129 VDD.n8712 VDD.n8704 3.04812
R16130 VDD.n11131 VDD.n11128 3.04812
R16131 VDD.n11230 VDD.n11227 3.04812
R16132 VDD.n10072 VDD.n10010 3.03311
R16133 VDD.n10632 VDD.n10631 3.03311
R16134 VDD.n10117 VDD.n10006 3.03311
R16135 VDD.n10519 VDD.n10150 3.03311
R16136 VDD.n9059 VDD.n9058 3.03311
R16137 VDD.n8886 VDD.n8769 3.03311
R16138 VDD.n9052 VDD.n9051 3.03311
R16139 VDD.n8800 VDD.n8799 3.03311
R16140 VDD.n9340 VDD.n9322 3.03311
R16141 VDD.n9313 VDD.n9250 3.03311
R16142 VDD.n9444 VDD.n9443 3.03311
R16143 VDD.n9189 VDD.n9188 3.03311
R16144 VDD.n10957 VDD.n10956 3.03311
R16145 VDD.n10953 VDD.n10952 3.03311
R16146 VDD.n10965 VDD.n9214 3.03311
R16147 VDD.n10946 VDD.n9219 3.03311
R16148 VDD.n11001 VDD.n11000 3.03311
R16149 VDD.n10987 VDD.n8747 3.03311
R16150 VDD.n9070 VDD.n9069 3.03311
R16151 VDD.n11024 VDD.n11023 3.03311
R16152 VDD.n9142 VDD.n9092 3.03311
R16153 VDD.n10968 VDD.n10967 3.03311
R16154 VDD.n11021 VDD.n8742 3.03311
R16155 VDD.n9181 VDD.n9164 3.03311
R16156 VDD.n9186 VDD.n9185 3.03311
R16157 VDD.n10993 VDD.n8740 3.03311
R16158 VDD.n10972 VDD.n10971 3.03311
R16159 VDD.n10470 VDD.n10469 3.03311
R16160 VDD.n10483 VDD.n10482 3.03311
R16161 VDD.n10435 VDD.n10155 3.03311
R16162 VDD.n10497 VDD.n10496 3.03311
R16163 VDD.n10477 VDD.n10476 3.03311
R16164 VDD.n10074 VDD.n10073 3.01226
R16165 VDD.n10634 VDD.n10633 3.01226
R16166 VDD.n10522 VDD.n10521 3.01226
R16167 VDD.n9591 VDD.n9582 3.01226
R16168 VDD.n9603 VDD.n9583 3.01226
R16169 VDD.n9737 VDD.n9735 3.01226
R16170 VDD.n9722 VDD.n9721 3.01226
R16171 VDD.n9761 VDD.n9550 3.01226
R16172 VDD.n9772 VDD.n9524 3.01226
R16173 VDD.n9782 VDD.n9510 3.01226
R16174 VDD.n9808 VDD.n9506 3.01226
R16175 VDD.n9819 VDD.n9481 3.01226
R16176 VDD.n9852 VDD.n9838 3.01226
R16177 VDD.n9854 VDD.n9836 3.01226
R16178 VDD.n10881 VDD.n10879 3.01226
R16179 VDD.n10893 VDD.n10678 3.01226
R16180 VDD.n10876 VDD.n10694 3.01226
R16181 VDD.n10826 VDD.n10825 3.01226
R16182 VDD.n10705 VDD.n10704 3.01226
R16183 VDD.n10710 VDD.n10706 3.01226
R16184 VDD.n8940 VDD.n8939 3.01226
R16185 VDD.n8945 VDD.n8944 3.01226
R16186 VDD.n8843 VDD.n8842 3.01226
R16187 VDD.n8848 VDD.n8847 3.01226
R16188 VDD.n9027 VDD.n9026 3.01226
R16189 VDD.n9022 VDD.n9021 3.01226
R16190 VDD.n9301 VDD.n9267 3.01226
R16191 VDD.n9297 VDD.n9296 3.01226
R16192 VDD.n9434 VDD.n9393 3.01226
R16193 VDD.n9433 VDD.n9396 3.01226
R16194 VDD.n9428 VDD.n9398 3.01226
R16195 VDD.n9148 VDD.n9093 3.01226
R16196 VDD.n9140 VDD.n9092 3.01226
R16197 VDD.t185 VDD.n6775 2.99829
R16198 VDD.n8136 VDD.n8133 2.98039
R16199 VDD.n11414 VDD.n11413 2.98039
R16200 VDD.n11347 VDD.n11041 2.98039
R16201 VDD.n11279 VDD.n11278 2.98039
R16202 VDD.n8227 VDD.n8226 2.97872
R16203 VDD.n8267 VDD.n8265 2.97872
R16204 VDD.n8313 VDD.n8312 2.97872
R16205 VDD.n8342 VDD.n7997 2.97872
R16206 VDD.n8450 VDD.n8381 2.97872
R16207 VDD.n8421 VDD.n8420 2.97872
R16208 VDD.n12389 VDD.n6952 2.96547
R16209 VDD.n12341 VDD.n12340 2.96547
R16210 VDD.n7033 VDD.n7029 2.96547
R16211 VDD.n7131 VDD.n7130 2.96547
R16212 VDD.n7186 VDD.n7104 2.96547
R16213 VDD.n7245 VDD.n7082 2.96547
R16214 VDD.n12212 VDD.n7286 2.96547
R16215 VDD.n12164 VDD.n12163 2.96547
R16216 VDD.n7971 VDD.n7970 2.96471
R16217 VDD.n7934 VDD.n7843 2.96471
R16218 VDD.n7921 VDD.n7850 2.96471
R16219 VDD.n7887 VDD.n7876 2.96471
R16220 VDD.n11453 VDD.n7713 2.96471
R16221 VDD.n11495 VDD.n7694 2.96471
R16222 VDD.n7687 VDD.n7682 2.96471
R16223 VDD.n11553 VDD.n11552 2.96471
R16224 VDD.n11565 VDD.n7651 2.96471
R16225 VDD.n8935 VDD.n8884 2.96007
R16226 VDD.n8783 VDD.n8782 2.96007
R16227 VDD.n9031 VDD.n8791 2.96007
R16228 VDD.n9260 VDD.n9258 2.96007
R16229 VDD.n12697 VDD.n6612 2.91154
R16230 VDD.n10285 VDD.n10236 2.91154
R16231 VDD.n10338 VDD.n10209 2.91154
R16232 VDD.n10385 VDD.n10384 2.91154
R16233 VDD.n9177 VDD.n8659 2.91015
R16234 VDD.n7787 VDD.n7784 2.88677
R16235 VDD.n8503 VDD.n8502 2.88677
R16236 VDD.n10286 VDD.n10238 2.86873
R16237 VDD.n10332 VDD.n10331 2.86873
R16238 VDD.n10383 VDD.n10185 2.86873
R16239 VDD.n10924 VDD.n9341 2.85341
R16240 VDD.n11655 VDD.n7606 2.84494
R16241 VDD.n11704 VDD.n7581 2.84494
R16242 VDD.n7579 VDD.n7574 2.84494
R16243 VDD.n11762 VDD.n7551 2.84494
R16244 VDD.n11769 VDD.n7544 2.84494
R16245 VDD.n11818 VDD.n7519 2.84494
R16246 VDD.n7517 VDD.n7512 2.84494
R16247 VDD.n11876 VDD.n7489 2.84494
R16248 VDD.n11883 VDD.n7482 2.84494
R16249 VDD.n11932 VDD.n7457 2.84494
R16250 VDD.n7455 VDD.n7450 2.84494
R16251 VDD.n11990 VDD.n7427 2.84494
R16252 VDD.n11997 VDD.n7420 2.84494
R16253 VDD.n12046 VDD.n7395 2.84494
R16254 VDD.n7393 VDD.n7388 2.84494
R16255 VDD.n11608 VDD.n7632 2.82997
R16256 VDD.n11622 VDD.n11621 2.82997
R16257 VDD.n12384 VDD.n6956 2.82084
R16258 VDD.n12334 VDD.n12333 2.82084
R16259 VDD.n12285 VDD.n7035 2.82084
R16260 VDD.n7139 VDD.n7124 2.82084
R16261 VDD.n7196 VDD.n7195 2.82084
R16262 VDD.n7250 VDD.n7078 2.82084
R16263 VDD.n12207 VDD.n7290 2.82084
R16264 VDD.n12157 VDD.n12156 2.82084
R16265 VDD.n6705 VDD.n6704 2.78311
R16266 VDD.n10290 VDD.n10289 2.78311
R16267 VDD.n10339 VDD.n10207 2.78311
R16268 VDD.n10388 VDD.n10181 2.78311
R16269 VDD.n8117 VDD.n8104 2.77722
R16270 VDD.n8609 VDD.n7738 2.77722
R16271 VDD.n11369 VDD.n8705 2.77722
R16272 VDD.n11129 VDD.n11121 2.77722
R16273 VDD.n11228 VDD.n6603 2.77722
R16274 VDD.n9150 VDD.t76 2.77
R16275 VDD.n9150 VDD.t68 2.77
R16276 VDD.n8068 VDD.n8067 2.72525
R16277 VDD.n8051 VDD.n8050 2.72525
R16278 VDD.n8317 VDD.n8316 2.72525
R16279 VDD.n8491 VDD.n7996 2.72525
R16280 VDD.n8447 VDD.n8446 2.72525
R16281 VDD.n8414 VDD.n8411 2.72525
R16282 VDD.n8179 VDD.n8131 2.70949
R16283 VDD.n8641 VDD.n8640 2.70949
R16284 VDD.n11351 VDD.n11350 2.70949
R16285 VDD.n11161 VDD.n11160 2.70949
R16286 VDD.n12681 VDD.t183 2.69851
R16287 VDD.n10281 VDD.n10280 2.69749
R16288 VDD.n10330 VDD.n10214 2.69749
R16289 VDD.n10380 VDD.n10379 2.69749
R16290 VDD.n7981 VDD.n7980 2.69524
R16291 VDD.n7975 VDD.n7814 2.69524
R16292 VDD.n7933 VDD.n7844 2.69524
R16293 VDD.n7925 VDD.n7924 2.69524
R16294 VDD.n7884 VDD.n7883 2.69524
R16295 VDD.n11454 VDD.n11452 2.69524
R16296 VDD.n11502 VDD.n7689 2.69524
R16297 VDD.n11509 VDD.n11508 2.69524
R16298 VDD.n11558 VDD.n7658 2.69524
R16299 VDD.n11566 VDD.n11564 2.69524
R16300 VDD.n10477 VDD.n6925 2.69036
R16301 VDD.n12388 VDD.n6953 2.67621
R16302 VDD.n6995 VDD.n6991 2.67621
R16303 VDD.n12289 VDD.n7034 2.67621
R16304 VDD.n7135 VDD.n7126 2.67621
R16305 VDD.n7190 VDD.n7189 2.67621
R16306 VDD.n7246 VDD.n7080 2.67621
R16307 VDD.n12211 VDD.n7287 2.67621
R16308 VDD.n7328 VDD.n7324 2.67621
R16309 VDD.n6523 VDD.n5808 2.64609
R16310 VDD.n5669 VDD.n4954 2.64609
R16311 VDD.n4883 VDD.n4168 2.64609
R16312 VDD.n4029 VDD.n3314 2.64609
R16313 VDD.n3243 VDD.n2528 2.64609
R16314 VDD.n2388 VDD.n1673 2.64609
R16315 VDD.n1155 VDD.n1153 2.64609
R16316 VDD.n709 VDD.n707 2.64609
R16317 VDD.n11363 VDD.n8720 2.64563
R16318 VDD.n11027 VDD.n11026 2.64563
R16319 VDD.n10026 VDD.n10023 2.63579
R16320 VDD.n10098 VDD.n10091 2.63579
R16321 VDD.n10145 VDD.n10141 2.63579
R16322 VDD.n10524 VDD.n10523 2.63579
R16323 VDD.n9979 VDD.n9974 2.63579
R16324 VDD.n9600 VDD.n9586 2.63579
R16325 VDD.n9586 VDD.n9574 2.63579
R16326 VDD.n9743 VDD.n9742 2.63579
R16327 VDD.n9716 VDD.n9715 2.63579
R16328 VDD.n9766 VDD.n9765 2.63579
R16329 VDD.n9534 VDD.n9533 2.63579
R16330 VDD.n9788 VDD.n9787 2.63579
R16331 VDD.n9812 VDD.n9500 2.63579
R16332 VDD.n9491 VDD.n9490 2.63579
R16333 VDD.n9860 VDD.n9859 2.63579
R16334 VDD.n10888 VDD.n10887 2.63579
R16335 VDD.n10867 VDD.n10776 2.63579
R16336 VDD.n10832 VDD.n10831 2.63579
R16337 VDD.n10756 VDD.n10711 2.63579
R16338 VDD.n10719 VDD.n10711 2.63579
R16339 VDD.n9439 VDD.n9438 2.63579
R16340 VDD.n9152 VDD.n9084 2.63579
R16341 VDD.n7987 VDD.n7807 2.63579
R16342 VDD.n12422 VDD.n6907 2.63579
R16343 VDD.n12454 VDD.n12451 2.63579
R16344 VDD.n12688 VDD.n6706 2.61187
R16345 VDD.n10293 VDD.n10234 2.61187
R16346 VDD.n10343 VDD.n10342 2.61187
R16347 VDD.n10389 VDD.n10179 2.61187
R16348 VDD.n11656 VDD.n11654 2.57404
R16349 VDD.n11706 VDD.n11705 2.57404
R16350 VDD.n11711 VDD.n11710 2.57404
R16351 VDD.n11761 VDD.n7552 2.57404
R16352 VDD.n11770 VDD.n11768 2.57404
R16353 VDD.n11820 VDD.n11819 2.57404
R16354 VDD.n11825 VDD.n11824 2.57404
R16355 VDD.n11875 VDD.n7490 2.57404
R16356 VDD.n11884 VDD.n11882 2.57404
R16357 VDD.n11934 VDD.n11933 2.57404
R16358 VDD.n11939 VDD.n11938 2.57404
R16359 VDD.n11989 VDD.n7428 2.57404
R16360 VDD.n11998 VDD.n11996 2.57404
R16361 VDD.n12048 VDD.n12047 2.57404
R16362 VDD.n12053 VDD.n12052 2.57404
R16363 VDD.n6386 VDD.n6385 2.56805
R16364 VDD.n5950 VDD.n5914 2.56805
R16365 VDD.n5951 VDD.n5950 2.56805
R16366 VDD.n5956 VDD.n5954 2.56805
R16367 VDD.n5958 VDD.n5956 2.56805
R16368 VDD.n5977 VDD.n5975 2.56805
R16369 VDD.n5532 VDD.n5531 2.56805
R16370 VDD.n5096 VDD.n5060 2.56805
R16371 VDD.n5097 VDD.n5096 2.56805
R16372 VDD.n5102 VDD.n5100 2.56805
R16373 VDD.n5104 VDD.n5102 2.56805
R16374 VDD.n5123 VDD.n5121 2.56805
R16375 VDD.n4746 VDD.n4745 2.56805
R16376 VDD.n4310 VDD.n4274 2.56805
R16377 VDD.n4311 VDD.n4310 2.56805
R16378 VDD.n4316 VDD.n4314 2.56805
R16379 VDD.n4318 VDD.n4316 2.56805
R16380 VDD.n4337 VDD.n4335 2.56805
R16381 VDD.n3892 VDD.n3891 2.56805
R16382 VDD.n3456 VDD.n3420 2.56805
R16383 VDD.n3457 VDD.n3456 2.56805
R16384 VDD.n3462 VDD.n3460 2.56805
R16385 VDD.n3464 VDD.n3462 2.56805
R16386 VDD.n3483 VDD.n3481 2.56805
R16387 VDD.n3106 VDD.n3105 2.56805
R16388 VDD.n2670 VDD.n2634 2.56805
R16389 VDD.n2671 VDD.n2670 2.56805
R16390 VDD.n2676 VDD.n2674 2.56805
R16391 VDD.n2678 VDD.n2676 2.56805
R16392 VDD.n2697 VDD.n2695 2.56805
R16393 VDD.n2251 VDD.n2250 2.56805
R16394 VDD.n1815 VDD.n1779 2.56805
R16395 VDD.n1816 VDD.n1815 2.56805
R16396 VDD.n1821 VDD.n1819 2.56805
R16397 VDD.n1823 VDD.n1821 2.56805
R16398 VDD.n1842 VDD.n1840 2.56805
R16399 VDD.n1374 VDD.n1371 2.56805
R16400 VDD.n1409 VDD.n1407 2.56805
R16401 VDD.n1414 VDD.n1409 2.56805
R16402 VDD.n1569 VDD.n1566 2.56805
R16403 VDD.n1566 VDD.n1563 2.56805
R16404 VDD.n1530 VDD.n1527 2.56805
R16405 VDD.n146 VDD.n143 2.56805
R16406 VDD.n181 VDD.n179 2.56805
R16407 VDD.n186 VDD.n181 2.56805
R16408 VDD.n341 VDD.n338 2.56805
R16409 VDD.n338 VDD.n335 2.56805
R16410 VDD.n302 VDD.n299 2.56805
R16411 VDD.n10097 VDD.n10087 2.56676
R16412 VDD.n11615 VDD.n7627 2.5605
R16413 VDD.n11616 VDD.n7624 2.5605
R16414 VDD.n6292 VDD.n6021 2.5605
R16415 VDD.n6301 VDD.n6291 2.5605
R16416 VDD.n5438 VDD.n5167 2.5605
R16417 VDD.n5447 VDD.n5437 2.5605
R16418 VDD.n4652 VDD.n4381 2.5605
R16419 VDD.n4661 VDD.n4651 2.5605
R16420 VDD.n3798 VDD.n3527 2.5605
R16421 VDD.n3807 VDD.n3797 2.5605
R16422 VDD.n3012 VDD.n2741 2.5605
R16423 VDD.n3021 VDD.n3011 2.5605
R16424 VDD.n2157 VDD.n1886 2.5605
R16425 VDD.n2166 VDD.n2156 2.5605
R16426 VDD.n1631 VDD.n1628 2.5605
R16427 VDD.n1625 VDD.n1622 2.5605
R16428 VDD.n403 VDD.n400 2.5605
R16429 VDD.n397 VDD.n394 2.5605
R16430 VDD.n12385 VDD.n6953 2.53157
R16431 VDD.n6996 VDD.n6995 2.53157
R16432 VDD.n12289 VDD.n12288 2.53157
R16433 VDD.n7136 VDD.n7135 2.53157
R16434 VDD.n7190 VDD.n7102 2.53157
R16435 VDD.n7249 VDD.n7080 2.53157
R16436 VDD.n12208 VDD.n7287 2.53157
R16437 VDD.n7329 VDD.n7328 2.53157
R16438 VDD.n10279 VDD.n10240 2.52625
R16439 VDD.n10375 VDD.n10187 2.52625
R16440 VDD.n8193 VDD.n8105 2.50632
R16441 VDD.n11432 VDD.n7739 2.50632
R16442 VDD.n11366 VDD.n11365 2.50632
R16443 VDD.n11297 VDD.n11122 2.50632
R16444 VDD.n12707 VDD.n6604 2.50632
R16445 VDD.n8238 VDD.n8237 2.47179
R16446 VDD.n8255 VDD.n8254 2.47179
R16447 VDD.n8324 VDD.n8006 2.47179
R16448 VDD.n8495 VDD.n8494 2.47179
R16449 VDD.n8393 VDD.n8392 2.47179
R16450 VDD.n8409 VDD.n8402 2.47179
R16451 VDD.n12687 VDD.n6707 2.44063
R16452 VDD.n10294 VDD.n10232 2.44063
R16453 VDD.n10346 VDD.n10205 2.44063
R16454 VDD.n10393 VDD.n10392 2.44063
R16455 VDD.n8184 VDD.n8182 2.4386
R16456 VDD.n8639 VDD.n8622 2.4386
R16457 VDD.n11046 VDD.n11045 2.4386
R16458 VDD.n11159 VDD.n11141 2.4386
R16459 VDD.n6543 VDD.n5794 2.43651
R16460 VDD.n5689 VDD.n4940 2.43651
R16461 VDD.n4903 VDD.n4154 2.43651
R16462 VDD.n4049 VDD.n3300 2.43651
R16463 VDD.n3263 VDD.n2514 2.43651
R16464 VDD.n2408 VDD.n1659 2.43651
R16465 VDD.n1189 VDD.n1187 2.43651
R16466 VDD.n743 VDD.n741 2.43651
R16467 VDD.n7979 VDD.n7812 2.42576
R16468 VDD.n7976 VDD.n7812 2.42576
R16469 VDD.n7930 VDD.n7929 2.42576
R16470 VDD.n7929 VDD.n7847 2.42576
R16471 VDD.n7880 VDD.n7879 2.42576
R16472 VDD.n7879 VDD.n7716 2.42576
R16473 VDD.n11504 VDD.n11503 2.42576
R16474 VDD.n11503 VDD.n7686 2.42576
R16475 VDD.n11557 VDD.n7659 2.42576
R16476 VDD.n7659 VDD.n7654 2.42576
R16477 VDD.n2470 VDD.n2469 2.42534
R16478 VDD.n830 VDD.n829 2.42534
R16479 VDD.n12620 VDD.t182 2.39873
R16480 VDD.n12385 VDD.n12384 2.38694
R16481 VDD.n12334 VDD.n6996 2.38694
R16482 VDD.n12288 VDD.n7035 2.38694
R16483 VDD.n7136 VDD.n7124 2.38694
R16484 VDD.n7195 VDD.n7102 2.38694
R16485 VDD.n7250 VDD.n7249 2.38694
R16486 VDD.n12208 VDD.n12207 2.38694
R16487 VDD.n12157 VDD.n7329 2.38694
R16488 VDD.n7373 VDD.n7369 2.38694
R16489 VDD.n12089 VDD.n7373 2.38694
R16490 VDD.n9150 VDD.n9082 2.37942
R16491 VDD.n9982 VDD.n9981 2.3755
R16492 VDD.n12704 VDD.n6604 2.37087
R16493 VDD.n7982 VDD.n7981 2.35839
R16494 VDD.n10276 VDD.n10275 2.35502
R16495 VDD.n10322 VDD.n10216 2.35502
R16496 VDD.n10374 VDD.n10189 2.35502
R16497 VDD.n9928 VDD.n9927 2.31116
R16498 VDD.n5731 VDD.n5723 2.30684
R16499 VDD.n4091 VDD.n4083 2.30684
R16500 VDD.n2450 VDD.n2442 2.30684
R16501 VDD.n810 VDD.n802 2.30684
R16502 VDD.n11654 VDD.n7609 2.30315
R16503 VDD.n11705 VDD.n7578 2.30315
R16504 VDD.n11711 VDD.n7578 2.30315
R16505 VDD.n7552 VDD.n7547 2.30315
R16506 VDD.n11768 VDD.n7547 2.30315
R16507 VDD.n11819 VDD.n7516 2.30315
R16508 VDD.n11825 VDD.n7516 2.30315
R16509 VDD.n7490 VDD.n7485 2.30315
R16510 VDD.n11882 VDD.n7485 2.30315
R16511 VDD.n11933 VDD.n7454 2.30315
R16512 VDD.n11939 VDD.n7454 2.30315
R16513 VDD.n7428 VDD.n7423 2.30315
R16514 VDD.n11996 VDD.n7423 2.30315
R16515 VDD.n12047 VDD.n7392 2.30315
R16516 VDD.n12053 VDD.n7392 2.30315
R16517 VDD.n11617 VDD.n11615 2.29103
R16518 VDD.n11617 VDD.n11616 2.29103
R16519 VDD.n10080 VDD.n10016 2.28225
R16520 VDD.n10114 VDD.n10086 2.28225
R16521 VDD.n10640 VDD.n10132 2.28225
R16522 VDD.n10558 VDD.n10531 2.28225
R16523 VDD.n12684 VDD.n12683 2.2694
R16524 VDD.n10298 VDD.n10297 2.2694
R16525 VDD.n10347 VDD.n10203 2.2694
R16526 VDD.n10396 VDD.n10177 2.2694
R16527 VDD.n10971 VDD.n9211 2.25953
R16528 VDD.n10068 VDD.n10027 2.25932
R16529 VDD.n10030 VDD.n10029 2.25932
R16530 VDD.n10102 VDD.n10094 2.25932
R16531 VDD.n10107 VDD.n10103 2.25932
R16532 VDD.n10627 VDD.n10585 2.25932
R16533 VDD.n10618 VDD.n10589 2.25932
R16534 VDD.n10566 VDD.n10500 2.25932
R16535 VDD.n10507 VDD.n10504 2.25932
R16536 VDD.n9594 VDD.n9592 2.25932
R16537 VDD.n9728 VDD.n9676 2.25932
R16538 VDD.n10821 VDD.n10820 2.25932
R16539 VDD.n10765 VDD.n10701 2.25932
R16540 VDD.n8917 VDD.n8916 2.25932
R16541 VDD.n8950 VDD.n8949 2.25932
R16542 VDD.n9039 VDD.n9034 2.25932
R16543 VDD.n8853 VDD.n8852 2.25932
R16544 VDD.n8816 VDD.n8815 2.25932
R16545 VDD.n9017 VDD.n9016 2.25932
R16546 VDD.n8901 VDD.n8897 2.25932
R16547 VDD.n9308 VDD.n9303 2.25932
R16548 VDD.n9292 VDD.n9291 2.25932
R16549 VDD.n9332 VDD.n9330 2.25932
R16550 VDD.n9380 VDD.n9379 2.25932
R16551 VDD.n9401 VDD.n9400 2.25932
R16552 VDD.n9421 VDD.n9402 2.25932
R16553 VDD.n9139 VDD.n9138 2.25932
R16554 VDD.n10109 VDD.n10102 2.25379
R16555 VDD.n9867 VDD.n9828 2.25051
R16556 VDD.n10885 VDD.n10670 2.25051
R16557 VDD.n5731 VDD.n5730 2.2505
R16558 VDD.n5732 VDD.n5718 2.2505
R16559 VDD.n5734 VDD.n5733 2.2505
R16560 VDD.n5721 VDD.n5710 2.2505
R16561 VDD.n5769 VDD.n5768 2.2505
R16562 VDD.n4091 VDD.n4090 2.2505
R16563 VDD.n4092 VDD.n4078 2.2505
R16564 VDD.n4094 VDD.n4093 2.2505
R16565 VDD.n4081 VDD.n4070 2.2505
R16566 VDD.n4129 VDD.n4128 2.2505
R16567 VDD.n2450 VDD.n2449 2.2505
R16568 VDD.n2451 VDD.n2437 2.2505
R16569 VDD.n2453 VDD.n2452 2.2505
R16570 VDD.n2440 VDD.n2429 2.2505
R16571 VDD.n2489 VDD.n2488 2.2505
R16572 VDD.n810 VDD.n809 2.2505
R16573 VDD.n811 VDD.n797 2.2505
R16574 VDD.n813 VDD.n812 2.2505
R16575 VDD.n800 VDD.n789 2.2505
R16576 VDD.n849 VDD.n848 2.2505
R16577 VDD.n9495 VDD.n9494 2.25002
R16578 VDD.n9792 VDD.n9515 2.25002
R16579 VDD.n9610 VDD.n9578 2.25002
R16580 VDD.n9538 VDD.n9537 2.25002
R16581 VDD.n9867 VDD.n9833 2.24905
R16582 VDD.n10679 VDD.n10670 2.24905
R16583 VDD.n10708 VDD.n10707 2.24807
R16584 VDD.n10873 VDD.n10774 2.24807
R16585 VDD.n9805 VDD.n9799 2.24807
R16586 VDD.n9758 VDD.n9757 2.24807
R16587 VDD.n9747 VDD.n9558 2.24807
R16588 VDD.n10559 VDD.n10151 2.24691
R16589 VDD.n10583 VDD.n10134 2.24691
R16590 VDD.n10115 VDD.n10003 2.24691
R16591 VDD.n10082 VDD.n10081 2.24691
R16592 VDD.n9058 VDD.n8758 2.24691
R16593 VDD.n8819 VDD.n8801 2.24691
R16594 VDD.n8774 VDD.n8767 2.24691
R16595 VDD.n9046 VDD.n8776 2.24691
R16596 VDD.n10954 VDD.n10953 2.24691
R16597 VDD.n9317 VDD.n9255 2.24691
R16598 VDD.n9353 VDD.n9349 2.24691
R16599 VDD.n9069 VDD.n8749 2.24691
R16600 VDD.n10773 VDD.n10772 2.24691
R16601 VDD.n10755 VDD.n10697 2.24691
R16602 VDD.n9835 VDD.n9834 2.24691
R16603 VDD.n9814 VDD.n9501 2.24691
R16604 VDD.n9823 VDD.n9478 2.24691
R16605 VDD.n9794 VDD.n9511 2.24691
R16606 VDD.n9581 VDD.n9576 2.24691
R16607 VDD.n9555 VDD.n9552 2.24691
R16608 VDD.n9767 VDD.n9544 2.24691
R16609 VDD.n9776 VDD.n9521 2.24691
R16610 VDD.n10158 VDD.n10155 2.24671
R16611 VDD.n10084 VDD.n10001 2.24671
R16612 VDD.n10059 VDD.n10008 2.24671
R16613 VDD.n10512 VDD.n10150 2.24671
R16614 VDD.n8802 VDD.n8800 2.24671
R16615 VDD.n9064 VDD.n8761 2.24671
R16616 VDD.n8773 VDD.n8768 2.24671
R16617 VDD.n10953 VDD.n10949 2.24671
R16618 VDD.n9344 VDD.n9324 2.24671
R16619 VDD.n10971 VDD.n10970 2.24671
R16620 VDD.n10768 VDD.n10698 2.24671
R16621 VDD.n10866 VDD.n10777 2.24671
R16622 VDD.n9817 VDD.n9476 2.24671
R16623 VDD.n9797 VDD.n9497 2.24671
R16624 VDD.n9770 VDD.n9519 2.24671
R16625 VDD.n9779 VDD.n9507 2.24671
R16626 VDD.n9751 VDD.n9540 2.24671
R16627 VDD.n9748 VDD.n9553 2.24671
R16628 VDD.n9597 VDD.n9579 2.24671
R16629 VDD.n8823 VDD.n8803 2.24661
R16630 VDD.n8930 VDD.n8929 2.24661
R16631 VDD.n10080 VDD.n10018 2.24613
R16632 VDD.n10114 VDD.n10087 2.24613
R16633 VDD.n10640 VDD.n10137 2.24613
R16634 VDD.n10531 VDD.n10530 2.24613
R16635 VDD.n10439 VDD.n10156 2.24365
R16636 VDD.n12389 VDD.n12388 2.24231
R16637 VDD.n12340 VDD.n6991 2.24231
R16638 VDD.n7034 VDD.n7033 2.24231
R16639 VDD.n7131 VDD.n7126 2.24231
R16640 VDD.n7189 VDD.n7104 2.24231
R16641 VDD.n7246 VDD.n7245 2.24231
R16642 VDD.n12212 VDD.n12211 2.24231
R16643 VDD.n12163 VDD.n7324 2.24231
R16644 VDD.n10870 VDD.n10774 2.23886
R16645 VDD.n10671 VDD.n10670 2.23886
R16646 VDD.n10676 VDD.n10670 2.23886
R16647 VDD.n10759 VDD.n10708 2.23886
R16648 VDD.n9805 VDD.n9804 2.23886
R16649 VDD.n9495 VDD.n9485 2.23886
R16650 VDD.n9792 VDD.n9791 2.23886
R16651 VDD.n9747 VDD.n9557 2.23886
R16652 VDD.n9610 VDD.n9580 2.23886
R16653 VDD.n9758 VDD.n9754 2.23886
R16654 VDD.n9538 VDD.n9528 2.23886
R16655 VDD.n8190 VDD.n8189 2.23542
R16656 VDD.n11429 VDD.n11428 2.23542
R16657 VDD.n8725 VDD.n8724 2.23542
R16658 VDD.n11294 VDD.n11293 2.23542
R16659 VDD.n8927 VDD.n8926 2.22452
R16660 VDD.n9047 VDD.n8785 2.22452
R16661 VDD.n8808 VDD.n8792 2.22452
R16662 VDD.n9257 VDD.n9253 2.22452
R16663 VDD.n10926 VDD.n10925 2.22452
R16664 VDD.n8242 VDD.n8241 2.21832
R16665 VDD.n8251 VDD.n8250 2.21832
R16666 VDD.n8326 VDD.n8004 2.21832
R16667 VDD.n8000 VDD.n7999 2.21832
R16668 VDD.n8437 VDD.n8397 2.21832
R16669 VDD.n8432 VDD.n8401 2.21832
R16670 VDD.n2472 VDD.n2471 2.19693
R16671 VDD.n832 VDD.n831 2.19693
R16672 VDD.n10272 VDD.n10242 2.18378
R16673 VDD.n10321 VDD.n10218 2.18378
R16674 VDD.n10371 VDD.n10370 2.18378
R16675 VDD.n10418 VDD.n10417 2.18378
R16676 VDD.n8127 VDD.n8110 2.1677
R16677 VDD.n8620 VDD.n7743 2.1677
R16678 VDD.n11044 VDD.n8726 2.1677
R16679 VDD.n11139 VDD.n11126 2.1677
R16680 VDD.n7980 VDD.n7979 2.15629
R16681 VDD.n7976 VDD.n7975 2.15629
R16682 VDD.n7930 VDD.n7844 2.15629
R16683 VDD.n7925 VDD.n7847 2.15629
R16684 VDD.n7883 VDD.n7880 2.15629
R16685 VDD.n11452 VDD.n7716 2.15629
R16686 VDD.n11504 VDD.n11502 2.15629
R16687 VDD.n11509 VDD.n7686 2.15629
R16688 VDD.n11558 VDD.n11557 2.15629
R16689 VDD.n11564 VDD.n7654 2.15629
R16690 VDD.n4114 VDD.n4110 2.12973
R16691 VDD.t75 VDD.n8647 2.11661
R16692 VDD.n11340 VDD.t34 2.11661
R16693 VDD.n12431 VDD.n6567 2.11357
R16694 VDD.n12435 VDD.n6567 2.11353
R16695 VDD.n9060 VDD.n8766 2.10401
R16696 VDD.n10253 VDD.n6710 2.09816
R16697 VDD.n10301 VDD.n10230 2.09816
R16698 VDD.n10351 VDD.n10350 2.09816
R16699 VDD.n10397 VDD.n10175 2.09816
R16700 VDD.n6960 VDD.n6956 2.09768
R16701 VDD.n12333 VDD.n6997 2.09768
R16702 VDD.n12285 VDD.n12284 2.09768
R16703 VDD.n7140 VDD.n7139 2.09768
R16704 VDD.n7196 VDD.n7100 2.09768
R16705 VDD.n7254 VDD.n7078 2.09768
R16706 VDD.n7294 VDD.n7290 2.09768
R16707 VDD.n12156 VDD.n7330 2.09768
R16708 VDD.n12770 VDD.n6578 2.07664
R16709 VDD.n5754 VDD.n5750 2.0723
R16710 VDD.n11656 VDD.n11655 2.03225
R16711 VDD.n11706 VDD.n11704 2.03225
R16712 VDD.n11710 VDD.n7579 2.03225
R16713 VDD.n11762 VDD.n11761 2.03225
R16714 VDD.n11770 VDD.n11769 2.03225
R16715 VDD.n11820 VDD.n11818 2.03225
R16716 VDD.n11824 VDD.n7517 2.03225
R16717 VDD.n11876 VDD.n11875 2.03225
R16718 VDD.n11884 VDD.n11883 2.03225
R16719 VDD.n11934 VDD.n11932 2.03225
R16720 VDD.n11938 VDD.n7455 2.03225
R16721 VDD.n11990 VDD.n11989 2.03225
R16722 VDD.n11998 VDD.n11997 2.03225
R16723 VDD.n12048 VDD.n12046 2.03225
R16724 VDD.n12052 VDD.n7393 2.03225
R16725 VDD.n7632 VDD.n7627 2.02155
R16726 VDD.n11622 VDD.n7624 2.02155
R16727 VDD.n10271 VDD.n10246 2.01254
R16728 VDD.n10318 VDD.n10317 2.01254
R16729 VDD.n10367 VDD.n10191 2.01254
R16730 VDD.n10416 VDD.n10167 2.01254
R16731 VDD.n6347 VDD.n6346 2.00398
R16732 VDD.n6345 VDD.n5935 2.00398
R16733 VDD.n6321 VDD.n5780 2.00398
R16734 VDD.n5493 VDD.n5492 2.00398
R16735 VDD.n5491 VDD.n5081 2.00398
R16736 VDD.n5467 VDD.n4926 2.00398
R16737 VDD.n4707 VDD.n4706 2.00398
R16738 VDD.n4705 VDD.n4295 2.00398
R16739 VDD.n4681 VDD.n4140 2.00398
R16740 VDD.n3853 VDD.n3852 2.00398
R16741 VDD.n3851 VDD.n3441 2.00398
R16742 VDD.n3827 VDD.n3286 2.00398
R16743 VDD.n3067 VDD.n3066 2.00398
R16744 VDD.n3065 VDD.n2655 2.00398
R16745 VDD.n3041 VDD.n2500 2.00398
R16746 VDD.n2212 VDD.n2211 2.00398
R16747 VDD.n2210 VDD.n1800 2.00398
R16748 VDD.n2186 VDD.n1645 2.00398
R16749 VDD.n1601 VDD.n1598 2.00398
R16750 VDD.n1605 VDD.n1604 2.00398
R16751 VDD.n1221 VDD.n1218 2.00398
R16752 VDD.n373 VDD.n370 2.00398
R16753 VDD.n377 VDD.n376 2.00398
R16754 VDD.n775 VDD.n772 2.00398
R16755 VDD.n11448 VDD.n7718 1.98435
R16756 VDD.n6076 VDD.n6074 1.97774
R16757 VDD.n5222 VDD.n5220 1.97774
R16758 VDD.n4436 VDD.n4434 1.97774
R16759 VDD.n3582 VDD.n3580 1.97774
R16760 VDD.n2796 VDD.n2794 1.97774
R16761 VDD.n1941 VDD.n1939 1.97774
R16762 VDD.n924 VDD.n923 1.97774
R16763 VDD.n478 VDD.n477 1.97774
R16764 VDD.n12478 VDD.n12430 1.96602
R16765 VDD.n8243 VDD.n8057 1.96486
R16766 VDD.n8249 VDD.n8057 1.96486
R16767 VDD.n8330 VDD.n8329 1.96486
R16768 VDD.n8329 VDD.n8001 1.96486
R16769 VDD.n8436 VDD.n8435 1.96486
R16770 VDD.n8435 VDD.n8398 1.96486
R16771 VDD.n8185 VDD.n8127 1.96452
R16772 VDD.n8621 VDD.n8620 1.96452
R16773 VDD.n11047 VDD.n11044 1.96452
R16774 VDD.n11140 VDD.n11139 1.96452
R16775 VDD.n6385 VDD.n6383 1.96392
R16776 VDD.n5911 VDD.n5902 1.96392
R16777 VDD.n6377 VDD.n5913 1.96392
R16778 VDD.n6376 VDD.n6374 1.96392
R16779 VDD.n6373 VDD.n6371 1.96392
R16780 VDD.n6369 VDD.n6367 1.96392
R16781 VDD.n5531 VDD.n5529 1.96392
R16782 VDD.n5057 VDD.n5048 1.96392
R16783 VDD.n5523 VDD.n5059 1.96392
R16784 VDD.n5522 VDD.n5520 1.96392
R16785 VDD.n5519 VDD.n5517 1.96392
R16786 VDD.n5515 VDD.n5513 1.96392
R16787 VDD.n4745 VDD.n4743 1.96392
R16788 VDD.n4271 VDD.n4262 1.96392
R16789 VDD.n4737 VDD.n4273 1.96392
R16790 VDD.n4736 VDD.n4734 1.96392
R16791 VDD.n4733 VDD.n4731 1.96392
R16792 VDD.n4729 VDD.n4727 1.96392
R16793 VDD.n3891 VDD.n3889 1.96392
R16794 VDD.n3417 VDD.n3408 1.96392
R16795 VDD.n3883 VDD.n3419 1.96392
R16796 VDD.n3882 VDD.n3880 1.96392
R16797 VDD.n3879 VDD.n3877 1.96392
R16798 VDD.n3875 VDD.n3873 1.96392
R16799 VDD.n3105 VDD.n3103 1.96392
R16800 VDD.n2631 VDD.n2622 1.96392
R16801 VDD.n3097 VDD.n2633 1.96392
R16802 VDD.n3096 VDD.n3094 1.96392
R16803 VDD.n3093 VDD.n3091 1.96392
R16804 VDD.n3089 VDD.n3087 1.96392
R16805 VDD.n2250 VDD.n2248 1.96392
R16806 VDD.n1776 VDD.n1767 1.96392
R16807 VDD.n2242 VDD.n1778 1.96392
R16808 VDD.n2241 VDD.n2239 1.96392
R16809 VDD.n2238 VDD.n2236 1.96392
R16810 VDD.n2234 VDD.n2232 1.96392
R16811 VDD.n1376 VDD.n1374 1.96392
R16812 VDD.n1382 VDD.n1379 1.96392
R16813 VDD.n1387 VDD.n1385 1.96392
R16814 VDD.n1393 VDD.n1390 1.96392
R16815 VDD.n1398 VDD.n1396 1.96392
R16816 VDD.n1405 VDD.n1401 1.96392
R16817 VDD.n148 VDD.n146 1.96392
R16818 VDD.n154 VDD.n151 1.96392
R16819 VDD.n159 VDD.n157 1.96392
R16820 VDD.n165 VDD.n162 1.96392
R16821 VDD.n170 VDD.n168 1.96392
R16822 VDD.n177 VDD.n173 1.96392
R16823 VDD.n6952 VDD.n6951 1.95304
R16824 VDD.n12341 VDD.n6988 1.95304
R16825 VDD.n12295 VDD.n7029 1.95304
R16826 VDD.n7130 VDD.n7128 1.95304
R16827 VDD.n7186 VDD.n7185 1.95304
R16828 VDD.n7240 VDD.n7082 1.95304
R16829 VDD.n7286 VDD.n7285 1.95304
R16830 VDD.n12164 VDD.n7321 1.95304
R16831 VDD.n6518 VDD.n6517 1.94579
R16832 VDD.n5664 VDD.n5663 1.94579
R16833 VDD.n4878 VDD.n4877 1.94579
R16834 VDD.n4024 VDD.n4023 1.94579
R16835 VDD.n3238 VDD.n3237 1.94579
R16836 VDD.n2383 VDD.n2382 1.94579
R16837 VDD.n1150 VDD.n1124 1.94579
R16838 VDD.n704 VDD.n678 1.94579
R16839 VDD.n11019 VDD.n8736 1.93951
R16840 VDD.n10256 VDD.n10255 1.92692
R16841 VDD.n10302 VDD.n10228 1.92692
R16842 VDD.n10354 VDD.n10201 1.92692
R16843 VDD.n10401 VDD.n10400 1.92692
R16844 VDD.n12131 VDD.n7350 1.91616
R16845 VDD.n6632 VDD.n6610 1.90031
R16846 VDD.n8120 VDD.n8118 1.8968
R16847 VDD.n8190 VDD.n8108 1.8968
R16848 VDD.n11429 VDD.n7742 1.8968
R16849 VDD.n8724 VDD.n8709 1.8968
R16850 VDD.n11294 VDD.n11125 1.8968
R16851 VDD.n6394 VDD.n5877 1.88841
R16852 VDD.n5540 VDD.n5023 1.88841
R16853 VDD.n4754 VDD.n4237 1.88841
R16854 VDD.n3900 VDD.n3383 1.88841
R16855 VDD.n3114 VDD.n2597 1.88841
R16856 VDD.n2259 VDD.n1742 1.88841
R16857 VDD.n1525 VDD.n1510 1.88841
R16858 VDD.n297 VDD.n282 1.88841
R16859 VDD.n7971 VDD.n7814 1.88682
R16860 VDD.n7934 VDD.n7933 1.88682
R16861 VDD.n7924 VDD.n7850 1.88682
R16862 VDD.n7884 VDD.n7876 1.88682
R16863 VDD.n11454 VDD.n11453 1.88682
R16864 VDD.n7694 VDD.n7689 1.88682
R16865 VDD.n11508 VDD.n7687 1.88682
R16866 VDD.n11552 VDD.n7658 1.88682
R16867 VDD.n11566 VDD.n11565 1.88682
R16868 VDD.n10071 VDD.n10068 1.88285
R16869 VDD.n10094 VDD.n10092 1.88285
R16870 VDD.n10585 VDD.n10146 1.88285
R16871 VDD.n10518 VDD.n10500 1.88285
R16872 VDD.n9617 VDD.n9572 1.88285
R16873 VDD.n9617 VDD.n9570 1.88285
R16874 VDD.n9687 VDD.n9686 1.88285
R16875 VDD.n9711 VDD.n9710 1.88285
R16876 VDD.n10861 VDD.n10860 1.88285
R16877 VDD.n10837 VDD.n10836 1.88285
R16878 VDD.n10750 VDD.n10749 1.88285
R16879 VDD.n10749 VDD.n10715 1.88285
R16880 VDD.n8925 VDD.n8922 1.88285
R16881 VDD.n9044 VDD.n8781 1.88285
R16882 VDD.n8806 VDD.n8805 1.88285
R16883 VDD.n9062 VDD.n8763 1.88285
R16884 VDD.n9062 VDD.n8764 1.88285
R16885 VDD.n9315 VDD.n9314 1.88285
R16886 VDD.n9339 VDD.n9329 1.88285
R16887 VDD.n9390 VDD.n9388 1.88285
R16888 VDD.n9390 VDD.n9359 1.88285
R16889 VDD.n7987 VDD.n7986 1.88285
R16890 VDD.n12493 VDD.n12492 1.88285
R16891 VDD.n12492 VDD.n6910 1.88285
R16892 VDD.n12460 VDD.n12459 1.88285
R16893 VDD.n12459 VDD.n12440 1.88285
R16894 VDD.n10099 VDD.n10098 1.87949
R16895 VDD.n12472 VDD.n12434 1.8537
R16896 VDD.n12703 VDD.n6607 1.85282
R16897 VDD.n10268 VDD.n10267 1.8413
R16898 VDD.n10314 VDD.n10220 1.8413
R16899 VDD.n10366 VDD.n10195 1.8413
R16900 VDD.n10413 VDD.n10412 1.8413
R16901 VDD.n8118 VDD.n8117 1.82907
R16902 VDD.n9739 VDD.n9641 1.81303
R16903 VDD.n10878 VDD.n10687 1.81303
R16904 VDD.n12378 VDD.n6961 1.80841
R16905 VDD.n12330 VDD.n12329 1.80841
R16906 VDD.n7042 VDD.n7038 1.80841
R16907 VDD.n7145 VDD.n7122 1.80841
R16908 VDD.n7200 VDD.n7199 1.80841
R16909 VDD.n7256 VDD.n7255 1.80841
R16910 VDD.n12201 VDD.n7295 1.80841
R16911 VDD.n12153 VDD.n12152 1.80841
R16912 VDD.n12692 VDD.n12691 1.79917
R16913 VDD.t154 VDD.n6835 1.79917
R16914 VDD.n6348 VDD.n6347 1.78137
R16915 VDD.n6322 VDD.n6321 1.78137
R16916 VDD.n5494 VDD.n5493 1.78137
R16917 VDD.n5468 VDD.n5467 1.78137
R16918 VDD.n4708 VDD.n4707 1.78137
R16919 VDD.n4682 VDD.n4681 1.78137
R16920 VDD.n3854 VDD.n3853 1.78137
R16921 VDD.n3828 VDD.n3827 1.78137
R16922 VDD.n3068 VDD.n3067 1.78137
R16923 VDD.n3042 VDD.n3041 1.78137
R16924 VDD.n2213 VDD.n2212 1.78137
R16925 VDD.n2187 VDD.n2186 1.78137
R16926 VDD.n1598 VDD.n1597 1.78137
R16927 VDD.n1218 VDD.n1217 1.78137
R16928 VDD.n370 VDD.n369 1.78137
R16929 VDD.n772 VDD.n771 1.78137
R16930 VDD.n11661 VDD.n7606 1.76135
R16931 VDD.n7586 VDD.n7581 1.76135
R16932 VDD.n11717 VDD.n7574 1.76135
R16933 VDD.n11756 VDD.n7551 1.76135
R16934 VDD.n11775 VDD.n7544 1.76135
R16935 VDD.n7524 VDD.n7519 1.76135
R16936 VDD.n11831 VDD.n7512 1.76135
R16937 VDD.n11870 VDD.n7489 1.76135
R16938 VDD.n11889 VDD.n7482 1.76135
R16939 VDD.n7462 VDD.n7457 1.76135
R16940 VDD.n11945 VDD.n7450 1.76135
R16941 VDD.n11984 VDD.n7427 1.76135
R16942 VDD.n12003 VDD.n7420 1.76135
R16943 VDD.n7400 VDD.n7395 1.76135
R16944 VDD.n12059 VDD.n7388 1.76135
R16945 VDD.n10259 VDD.n10252 1.75568
R16946 VDD.n10306 VDD.n10305 1.75568
R16947 VDD.n10355 VDD.n10199 1.75568
R16948 VDD.n10404 VDD.n10173 1.75568
R16949 VDD.n11609 VDD.n11608 1.75208
R16950 VDD.n11621 VDD.n7625 1.75208
R16951 VDD.n6214 VDD.n6074 1.74595
R16952 VDD.n5360 VDD.n5220 1.74595
R16953 VDD.n4574 VDD.n4434 1.74595
R16954 VDD.n3720 VDD.n3580 1.74595
R16955 VDD.n2934 VDD.n2794 1.74595
R16956 VDD.n2079 VDD.n1939 1.74595
R16957 VDD.n926 VDD.n924 1.74595
R16958 VDD.n480 VDD.n478 1.74595
R16959 VDD.n11142 VDD.t43 1.71984
R16960 VDD.n11018 VDD.n11016 1.71462
R16961 VDD.n6538 VDD.n5798 1.71235
R16962 VDD.n6537 VDD.n5799 1.71235
R16963 VDD.n6534 VDD.n6533 1.71235
R16964 VDD.n6529 VDD.n5802 1.71235
R16965 VDD.n6528 VDD.n5805 1.71235
R16966 VDD.n6524 VDD.n6523 1.71235
R16967 VDD.n5684 VDD.n4944 1.71235
R16968 VDD.n5683 VDD.n4945 1.71235
R16969 VDD.n5680 VDD.n5679 1.71235
R16970 VDD.n5675 VDD.n4948 1.71235
R16971 VDD.n5674 VDD.n4951 1.71235
R16972 VDD.n5670 VDD.n5669 1.71235
R16973 VDD.n4898 VDD.n4158 1.71235
R16974 VDD.n4897 VDD.n4159 1.71235
R16975 VDD.n4894 VDD.n4893 1.71235
R16976 VDD.n4889 VDD.n4162 1.71235
R16977 VDD.n4888 VDD.n4165 1.71235
R16978 VDD.n4884 VDD.n4883 1.71235
R16979 VDD.n4044 VDD.n3304 1.71235
R16980 VDD.n4043 VDD.n3305 1.71235
R16981 VDD.n4040 VDD.n4039 1.71235
R16982 VDD.n4035 VDD.n3308 1.71235
R16983 VDD.n4034 VDD.n3311 1.71235
R16984 VDD.n4030 VDD.n4029 1.71235
R16985 VDD.n3258 VDD.n2518 1.71235
R16986 VDD.n3257 VDD.n2519 1.71235
R16987 VDD.n3254 VDD.n3253 1.71235
R16988 VDD.n3249 VDD.n2522 1.71235
R16989 VDD.n3248 VDD.n2525 1.71235
R16990 VDD.n3244 VDD.n3243 1.71235
R16991 VDD.n2403 VDD.n1663 1.71235
R16992 VDD.n2402 VDD.n1664 1.71235
R16993 VDD.n2399 VDD.n2398 1.71235
R16994 VDD.n2394 VDD.n1667 1.71235
R16995 VDD.n2393 VDD.n1670 1.71235
R16996 VDD.n2389 VDD.n2388 1.71235
R16997 VDD.n1184 VDD.n1180 1.71235
R16998 VDD.n1177 VDD.n1175 1.71235
R16999 VDD.n1173 VDD.n1170 1.71235
R17000 VDD.n1167 VDD.n1165 1.71235
R17001 VDD.n1163 VDD.n1160 1.71235
R17002 VDD.n1157 VDD.n1155 1.71235
R17003 VDD.n738 VDD.n734 1.71235
R17004 VDD.n731 VDD.n729 1.71235
R17005 VDD.n727 VDD.n724 1.71235
R17006 VDD.n721 VDD.n719 1.71235
R17007 VDD.n717 VDD.n714 1.71235
R17008 VDD.n711 VDD.n709 1.71235
R17009 VDD.n8241 VDD.n8061 1.71139
R17010 VDD.n8251 VDD.n8055 1.71139
R17011 VDD.n8326 VDD.n8325 1.71139
R17012 VDD.n7999 VDD.n7992 1.71139
R17013 VDD.n8397 VDD.n8394 1.71139
R17014 VDD.n8432 VDD.n8431 1.71139
R17015 VDD.n10899 VDD.n10664 1.71033
R17016 VDD.n10904 VDD.n9231 1.70907
R17017 VDD.n10906 VDD.n9237 1.70593
R17018 VDD.n9902 VDD.n9451 1.70593
R17019 VDD.n10902 VDD.n9900 1.70592
R17020 VDD.n9346 VDD.n9233 1.70592
R17021 VDD.n9885 VDD.n9459 1.70592
R17022 VDD.n10655 VDD.n9987 1.70591
R17023 VDD.n9885 VDD.n9475 1.70591
R17024 VDD.n10651 VDD.n9987 1.7059
R17025 VDD.n10660 VDD.n9451 1.70583
R17026 VDD.n10942 VDD.n9244 1.70583
R17027 VDD.n9246 VDD.n9230 1.70582
R17028 VDD.n10900 VDD.n9450 1.70582
R17029 VDD.n9890 VDD.n9456 1.7058
R17030 VDD.n9890 VDD.n9889 1.70579
R17031 VDD.n9995 VDD.n9992 1.70578
R17032 VDD.n10650 VDD.n9984 1.70577
R17033 VDD.n9320 VDD.n9242 1.7055
R17034 VDD.n9351 VDD.n9348 1.7055
R17035 VDD.n10908 VDD.n10907 1.7055
R17036 VDD.n10911 VDD.n10910 1.7055
R17037 VDD.n10916 VDD.n10915 1.7055
R17038 VDD.n10919 VDD.n10918 1.7055
R17039 VDD.n10930 VDD.n10929 1.7055
R17040 VDD.n10933 VDD.n10932 1.7055
R17041 VDD.n10936 VDD.n10935 1.7055
R17042 VDD.n10940 VDD.n9245 1.7055
R17043 VDD.n9897 VDD.n9453 1.7055
R17044 VDD.n9895 VDD.n9894 1.7055
R17045 VDD.n9892 VDD.n9891 1.7055
R17046 VDD.n9839 VDD.n9455 1.7055
R17047 VDD.n9842 VDD.n9841 1.7055
R17048 VDD.n9845 VDD.n9844 1.7055
R17049 VDD.n9848 VDD.n9847 1.7055
R17050 VDD.n9826 VDD.n9472 1.7055
R17051 VDD.n9883 VDD.n9473 1.7055
R17052 VDD.n9881 VDD.n9880 1.7055
R17053 VDD.n9876 VDD.n9875 1.7055
R17054 VDD.n9873 VDD.n9872 1.7055
R17055 VDD.n9870 VDD.n9869 1.7055
R17056 VDD.n10665 VDD.n9901 1.7055
R17057 VDD.n9840 VDD.n9463 1.7055
R17058 VDD.n9843 VDD.n9464 1.7055
R17059 VDD.n9825 VDD.n9471 1.7055
R17060 VDD.n9885 VDD.n9884 1.7055
R17061 VDD.n9882 VDD.n9467 1.7055
R17062 VDD.n9877 VDD.n9460 1.7055
R17063 VDD.n9874 VDD.n9466 1.7055
R17064 VDD.n9871 VDD.n9461 1.7055
R17065 VDD.n9832 VDD.n9465 1.7055
R17066 VDD.n9319 VDD.n9236 1.7055
R17067 VDD.n10945 VDD.n10944 1.7055
R17068 VDD.n10906 VDD.n9345 1.7055
R17069 VDD.n10909 VDD.n9238 1.7055
R17070 VDD.n10914 VDD.n9235 1.7055
R17071 VDD.n10917 VDD.n9239 1.7055
R17072 VDD.n10931 VDD.n9240 1.7055
R17073 VDD.n10934 VDD.n9233 1.7055
R17074 VDD.n10939 VDD.n9241 1.7055
R17075 VDD.n10942 VDD.n10941 1.7055
R17076 VDD.n10902 VDD.n9898 1.7055
R17077 VDD.n9896 VDD.n9451 1.7055
R17078 VDD.n9893 VDD.n9452 1.7055
R17079 VDD.n10666 VDD.n10661 1.7055
R17080 VDD.n10582 VDD.n10581 1.7055
R17081 VDD.n10576 VDD.n10575 1.7055
R17082 VDD.n10641 VDD.n10640 1.7055
R17083 VDD.n10130 VDD.n9999 1.7055
R17084 VDD.n10580 VDD.n9986 1.7055
R17085 VDD.n10579 VDD.n10578 1.7055
R17086 VDD.n10577 VDD.n9993 1.7055
R17087 VDD.n10574 VDD.n10573 1.7055
R17088 VDD.n10572 VDD.n9985 1.7055
R17089 VDD.n10571 VDD.n10570 1.7055
R17090 VDD.n10569 VDD.n9994 1.7055
R17091 VDD.n10120 VDD.n10119 1.7055
R17092 VDD.n10122 VDD.n10121 1.7055
R17093 VDD.n10123 VDD.n9987 1.7055
R17094 VDD.n10126 VDD.n10125 1.7055
R17095 VDD.n10127 VDD.n9991 1.7055
R17096 VDD.n10129 VDD.n10128 1.7055
R17097 VDD.n10650 VDD.n10649 1.7055
R17098 VDD.n10648 VDD.n10000 1.7055
R17099 VDD.n10647 VDD.n9990 1.7055
R17100 VDD.n10646 VDD.n10645 1.7055
R17101 VDD.n10643 VDD.n10642 1.7055
R17102 VDD.n10135 VDD.n9989 1.7055
R17103 VDD.n5771 VDD.n5709 1.7055
R17104 VDD.n5771 VDD.n5770 1.7055
R17105 VDD.n4131 VDD.n4069 1.7055
R17106 VDD.n4131 VDD.n4130 1.7055
R17107 VDD.n2491 VDD.n2428 1.7055
R17108 VDD.n2491 VDD.n2490 1.7055
R17109 VDD.n851 VDD.n788 1.7055
R17110 VDD.n851 VDD.n850 1.7055
R17111 VDD.n9890 VDD.n9457 1.70519
R17112 VDD.n10120 VDD.n9998 1.70511
R17113 VDD.n11017 VDD.n8739 1.70413
R17114 VDD.n11006 VDD.n8755 1.70404
R17115 VDD.n11007 VDD.n8751 1.70006
R17116 VDD.n11014 VDD.n8741 1.70006
R17117 VDD.n8182 VDD.n8128 1.69362
R17118 VDD.n8642 VDD.n8639 1.69362
R17119 VDD.n11045 VDD.n11037 1.69362
R17120 VDD.n11162 VDD.n11159 1.69362
R17121 VDD.n10424 VDD.n10161 1.67007
R17122 VDD.n10264 VDD.n10248 1.67007
R17123 VDD.n10313 VDD.n10222 1.67007
R17124 VDD.n10363 VDD.n10362 1.67007
R17125 VDD.n10409 VDD.n10169 1.67007
R17126 VDD.n6556 VDD.n6555 1.67007
R17127 VDD.n5702 VDD.n5701 1.67007
R17128 VDD.n4916 VDD.n4915 1.67007
R17129 VDD.n4062 VDD.n4061 1.67007
R17130 VDD.n3276 VDD.n3275 1.67007
R17131 VDD.n2421 VDD.n2420 1.67007
R17132 VDD.n1225 VDD.n1224 1.67007
R17133 VDD.n779 VDD.n778 1.67007
R17134 VDD.n12395 VDD.n6947 1.66378
R17135 VDD.n12345 VDD.n12344 1.66378
R17136 VDD.n12296 VDD.n7026 1.66378
R17137 VDD.n12251 VDD.n7068 1.66378
R17138 VDD.n7181 VDD.n7106 1.66378
R17139 VDD.n7239 VDD.n7084 1.66378
R17140 VDD.n12218 VDD.n7281 1.66378
R17141 VDD.n12168 VDD.n12167 1.66378
R17142 VDD.n5962 VDD.n5960 1.66186
R17143 VDD.n5963 VDD.n5946 1.66186
R17144 VDD.n5968 VDD.n5966 1.66186
R17145 VDD.n5969 VDD.n5944 1.66186
R17146 VDD.n5974 VDD.n5972 1.66186
R17147 VDD.n5978 VDD.n5977 1.66186
R17148 VDD.n5108 VDD.n5106 1.66186
R17149 VDD.n5109 VDD.n5092 1.66186
R17150 VDD.n5114 VDD.n5112 1.66186
R17151 VDD.n5115 VDD.n5090 1.66186
R17152 VDD.n5120 VDD.n5118 1.66186
R17153 VDD.n5124 VDD.n5123 1.66186
R17154 VDD.n4322 VDD.n4320 1.66186
R17155 VDD.n4323 VDD.n4306 1.66186
R17156 VDD.n4328 VDD.n4326 1.66186
R17157 VDD.n4329 VDD.n4304 1.66186
R17158 VDD.n4334 VDD.n4332 1.66186
R17159 VDD.n4338 VDD.n4337 1.66186
R17160 VDD.n3468 VDD.n3466 1.66186
R17161 VDD.n3469 VDD.n3452 1.66186
R17162 VDD.n3474 VDD.n3472 1.66186
R17163 VDD.n3475 VDD.n3450 1.66186
R17164 VDD.n3480 VDD.n3478 1.66186
R17165 VDD.n3484 VDD.n3483 1.66186
R17166 VDD.n2682 VDD.n2680 1.66186
R17167 VDD.n2683 VDD.n2666 1.66186
R17168 VDD.n2688 VDD.n2686 1.66186
R17169 VDD.n2689 VDD.n2664 1.66186
R17170 VDD.n2694 VDD.n2692 1.66186
R17171 VDD.n2698 VDD.n2697 1.66186
R17172 VDD.n1827 VDD.n1825 1.66186
R17173 VDD.n1828 VDD.n1811 1.66186
R17174 VDD.n1833 VDD.n1831 1.66186
R17175 VDD.n1834 VDD.n1809 1.66186
R17176 VDD.n1839 VDD.n1837 1.66186
R17177 VDD.n1843 VDD.n1842 1.66186
R17178 VDD.n1560 VDD.n1557 1.66186
R17179 VDD.n1554 VDD.n1552 1.66186
R17180 VDD.n1549 VDD.n1546 1.66186
R17181 VDD.n1543 VDD.n1541 1.66186
R17182 VDD.n1538 VDD.n1535 1.66186
R17183 VDD.n1532 VDD.n1530 1.66186
R17184 VDD.n332 VDD.n329 1.66186
R17185 VDD.n326 VDD.n324 1.66186
R17186 VDD.n321 VDD.n318 1.66186
R17187 VDD.n315 VDD.n313 1.66186
R17188 VDD.n310 VDD.n307 1.66186
R17189 VDD.n304 VDD.n302 1.66186
R17190 VDD.n9049 VDD.n8788 1.64452
R17191 VDD.n9033 VDD.n8794 1.64452
R17192 VDD.n8933 VDD.n8932 1.64447
R17193 VDD.n9311 VDD.n9263 1.64446
R17194 VDD.n10924 VDD.n10923 1.64446
R17195 VDD.n8502 VDD.n7807 1.63187
R17196 VDD.n8194 VDD.n8193 1.6259
R17197 VDD.n11433 VDD.n11432 1.6259
R17198 VDD.n11366 VDD.n8708 1.6259
R17199 VDD.n11298 VDD.n11297 1.6259
R17200 VDD.n12708 VDD.n12707 1.6259
R17201 VDD.n9983 VDD.n9982 1.62066
R17202 VDD.n7970 VDD.n7819 1.61734
R17203 VDD.n7843 VDD.n7841 1.61734
R17204 VDD.n7921 VDD.n7920 1.61734
R17205 VDD.n7888 VDD.n7887 1.61734
R17206 VDD.n11459 VDD.n7713 1.61734
R17207 VDD.n11496 VDD.n11495 1.61734
R17208 VDD.n11515 VDD.n7682 1.61734
R17209 VDD.n11553 VDD.n11551 1.61734
R17210 VDD.n11571 VDD.n7651 1.61734
R17211 VDD.n6636 VDD.n6633 1.61534
R17212 VDD.n6637 VDD.n6636 1.61534
R17213 VDD.n6637 VDD.n6630 1.61534
R17214 VDD.n6643 VDD.n6630 1.61534
R17215 VDD.n6644 VDD.n6643 1.61534
R17216 VDD.n6644 VDD.n6628 1.61534
R17217 VDD.n6650 VDD.n6628 1.61534
R17218 VDD.n6651 VDD.n6650 1.61534
R17219 VDD.n6651 VDD.n6626 1.61534
R17220 VDD.n6657 VDD.n6626 1.61534
R17221 VDD.n6658 VDD.n6657 1.61534
R17222 VDD.n6658 VDD.n6623 1.61534
R17223 VDD.n6698 VDD.n6624 1.61534
R17224 VDD.n6692 VDD.n6624 1.61534
R17225 VDD.n6692 VDD.n6691 1.61534
R17226 VDD.n6691 VDD.n6664 1.61534
R17227 VDD.n6685 VDD.n6664 1.61534
R17228 VDD.n6685 VDD.n6684 1.61534
R17229 VDD.n6684 VDD.n6666 1.61534
R17230 VDD.n6678 VDD.n6666 1.61534
R17231 VDD.n6678 VDD.n6677 1.61534
R17232 VDD.n6677 VDD.n6668 1.61534
R17233 VDD.n6671 VDD.n6668 1.61534
R17234 VDD.n6671 VDD.n6575 1.61534
R17235 VDD.n6012 VDD.n6009 1.61441
R17236 VDD.n5158 VDD.n5155 1.61441
R17237 VDD.n4372 VDD.n4369 1.61441
R17238 VDD.n3518 VDD.n3515 1.61441
R17239 VDD.n2732 VDD.n2729 1.61441
R17240 VDD.n1877 VDD.n1874 1.61441
R17241 VDD.n1609 VDD.n1608 1.61441
R17242 VDD.n381 VDD.n380 1.61441
R17243 VDD.n12470 VDD.n12435 1.59629
R17244 VDD.n12477 VDD.n12431 1.59579
R17245 VDD.n11233 VDD.t5 1.58758
R17246 VDD.n10260 VDD.n10250 1.58445
R17247 VDD.n10309 VDD.n10224 1.58445
R17248 VDD.n10326 VDD.n10325 1.58445
R17249 VDD.n10359 VDD.n10358 1.58445
R17250 VDD.n10405 VDD.n10171 1.58445
R17251 VDD.n8498 VDD.n8497 1.58383
R17252 VDD.n10425 VDD.n10424 1.57731
R17253 VDD.n11646 VDD.n7609 1.55817
R17254 VDD.n12702 VDD.n6609 1.5505
R17255 VDD.n12377 VDD.n6962 1.51914
R17256 VDD.n7004 VDD.n7000 1.51914
R17257 VDD.n12278 VDD.n7043 1.51914
R17258 VDD.n7146 VDD.n7120 1.51914
R17259 VDD.n7204 VDD.n7098 1.51914
R17260 VDD.n12245 VDD.n7075 1.51914
R17261 VDD.n12200 VDD.n7296 1.51914
R17262 VDD.n7337 VDD.n7333 1.51914
R17263 VDD.n10531 VDD.n10510 1.51434
R17264 VDD.n10080 VDD.n10079 1.51334
R17265 VDD.n10114 VDD.n10113 1.51334
R17266 VDD.n10640 VDD.n10639 1.51334
R17267 VDD.n10061 VDD.n10057 1.50638
R17268 VDD.n10100 VDD.n10095 1.50638
R17269 VDD.n10622 VDD.n10616 1.50638
R17270 VDD.n10561 VDD.n10505 1.50638
R17271 VDD.n9158 VDD.n9157 1.50638
R17272 VDD.n9131 VDD.n9130 1.50638
R17273 VDD.n9129 VDD.n9110 1.50638
R17274 VDD.n12702 VDD.n12701 1.5044
R17275 VDD.n10110 VDD.n10101 1.50148
R17276 VDD.n10484 VDD.n10483 1.5005
R17277 VDD.n10490 VDD.n10489 1.5005
R17278 VDD.n10476 VDD.n10451 1.5005
R17279 VDD.n9137 VDD.n9136 1.5005
R17280 VDD.n9127 VDD.n9108 1.5005
R17281 VDD.n9123 VDD.n9122 1.5005
R17282 VDD.n9142 VDD.n9105 1.5005
R17283 VDD.n9147 VDD.n9146 1.5005
R17284 VDD.n9104 VDD.n9103 1.5005
R17285 VDD.n9153 VDD.n9087 1.5005
R17286 VDD.n9086 VDD.n9083 1.5005
R17287 VDD.n10226 VDD.t182 1.4994
R17288 VDD.n12426 VDD.n6913 1.4994
R17289 VDD.n10263 VDD.n10250 1.49883
R17290 VDD.n10310 VDD.n10309 1.49883
R17291 VDD.n10359 VDD.n10197 1.49883
R17292 VDD.n10408 VDD.n10171 1.49883
R17293 VDD.n10080 VDD.n10012 1.49119
R17294 VDD.n10114 VDD.n10085 1.49076
R17295 VDD.n8893 VDD.n8759 1.49076
R17296 VDD.n8929 VDD.n8772 1.49076
R17297 VDD.n9043 VDD.n9042 1.49076
R17298 VDD.n9252 VDD.n9248 1.49076
R17299 VDD.n11660 VDD.n7607 1.49045
R17300 VDD.n11698 VDD.n11697 1.49045
R17301 VDD.n11719 VDD.n11718 1.49045
R17302 VDD.n11757 VDD.n11755 1.49045
R17303 VDD.n11774 VDD.n7545 1.49045
R17304 VDD.n11812 VDD.n11811 1.49045
R17305 VDD.n11833 VDD.n11832 1.49045
R17306 VDD.n11871 VDD.n11869 1.49045
R17307 VDD.n11888 VDD.n7483 1.49045
R17308 VDD.n11926 VDD.n11925 1.49045
R17309 VDD.n11947 VDD.n11946 1.49045
R17310 VDD.n11985 VDD.n11983 1.49045
R17311 VDD.n12002 VDD.n7421 1.49045
R17312 VDD.n12040 VDD.n12039 1.49045
R17313 VDD.n12061 VDD.n12060 1.49045
R17314 VDD.n10531 VDD.n10511 1.49033
R17315 VDD.n9042 VDD.n9041 1.4899
R17316 VDD.n8894 VDD.n8893 1.4899
R17317 VDD.n9262 VDD.n9248 1.4899
R17318 VDD.n8931 VDD.n8921 1.4871
R17319 VDD.n8787 VDD.n8786 1.4871
R17320 VDD.n8813 VDD.n8793 1.4871
R17321 VDD.n9261 VDD.n9259 1.4871
R17322 VDD.n9342 VDD.n9337 1.4871
R17323 VDD.n10708 VDD.n10700 1.48392
R17324 VDD.n10774 VDD.n10695 1.48392
R17325 VDD.n9806 VDD.n9805 1.48392
R17326 VDD.n9792 VDD.n9514 1.48392
R17327 VDD.n9759 VDD.n9758 1.48392
R17328 VDD.n9747 VDD.n9556 1.48392
R17329 VDD.n9610 VDD.n9577 1.48392
R17330 VDD.n9538 VDD.n9525 1.48392
R17331 VDD.n9495 VDD.n9482 1.48392
R17332 VDD.n9213 VDD.n9212 1.48264
R17333 VDD.n11603 VDD.n7631 1.48261
R17334 VDD.n11628 VDD.n7620 1.48261
R17335 VDD.n9857 VDD.n9828 1.47597
R17336 VDD.n10885 VDD.n10884 1.47597
R17337 VDD.n9764 VDD.n9546 1.46766
R17338 VDD.n9531 VDD.n9527 1.46766
R17339 VDD.n9488 VDD.n9484 1.46766
R17340 VDD.n9785 VDD.n9513 1.46766
R17341 VDD.n9811 VDD.n9502 1.46766
R17342 VDD.n6255 VDD.n6054 1.45846
R17343 VDD.n6286 VDD.n6048 1.45846
R17344 VDD.n6048 VDD.n5778 1.45846
R17345 VDD.n5401 VDD.n5200 1.45846
R17346 VDD.n5432 VDD.n5194 1.45846
R17347 VDD.n5194 VDD.n4924 1.45846
R17348 VDD.n4615 VDD.n4414 1.45846
R17349 VDD.n4646 VDD.n4408 1.45846
R17350 VDD.n4408 VDD.n4138 1.45846
R17351 VDD.n3761 VDD.n3560 1.45846
R17352 VDD.n3792 VDD.n3554 1.45846
R17353 VDD.n3554 VDD.n3284 1.45846
R17354 VDD.n2975 VDD.n2774 1.45846
R17355 VDD.n3006 VDD.n2768 1.45846
R17356 VDD.n2768 VDD.n2498 1.45846
R17357 VDD.n2120 VDD.n1919 1.45846
R17358 VDD.n2151 VDD.n1913 1.45846
R17359 VDD.n1913 VDD.n1643 1.45846
R17360 VDD.n986 VDD.n983 1.45846
R17361 VDD.n1023 VDD.n1020 1.45846
R17362 VDD.n1026 VDD.n1023 1.45846
R17363 VDD.n540 VDD.n537 1.45846
R17364 VDD.n577 VDD.n574 1.45846
R17365 VDD.n580 VDD.n577 1.45846
R17366 VDD.n8238 VDD.n8063 1.45793
R17367 VDD.n8254 VDD.n8052 1.45793
R17368 VDD.n8318 VDD.n8006 1.45793
R17369 VDD.n8494 VDD.n7993 1.45793
R17370 VDD.n8392 VDD.n8385 1.45793
R17371 VDD.n8410 VDD.n8409 1.45793
R17372 VDD.n12692 VDD.n6622 1.45532
R17373 VDD.n4130 VDD.n4129 1.42802
R17374 VDD.n2490 VDD.n2489 1.42802
R17375 VDD.n850 VDD.n849 1.42802
R17376 VDD.n8179 VDD.n8178 1.42272
R17377 VDD.n8640 VDD.n8632 1.42272
R17378 VDD.n11350 VDD.n11038 1.42272
R17379 VDD.n11160 VDD.n11152 1.42272
R17380 VDD.n5770 VDD.n5769 1.42272
R17381 VDD.n10264 VDD.n10263 1.41321
R17382 VDD.n10310 VDD.n10222 1.41321
R17383 VDD.n10362 VDD.n10197 1.41321
R17384 VDD.n10409 VDD.n10408 1.41321
R17385 VDD.n12418 VDD.n6926 1.41321
R17386 VDD.n10492 VDD.n10434 1.3918
R17387 VDD.n8534 VDD.n7787 1.38089
R17388 VDD.n8503 VDD.n7805 1.38089
R17389 VDD.n12396 VDD.n6944 1.37451
R17390 VDD.n6987 VDD.n6986 1.37451
R17391 VDD.n12300 VDD.n12299 1.37451
R17392 VDD.n12252 VDD.n7065 1.37451
R17393 VDD.n7180 VDD.n7108 1.37451
R17394 VDD.n7236 VDD.n7235 1.37451
R17395 VDD.n12219 VDD.n7278 1.37451
R17396 VDD.n7320 VDD.n7319 1.37451
R17397 VDD.n8610 VDD.n8609 1.355
R17398 VDD.n11370 VDD.n11369 1.355
R17399 VDD.n11130 VDD.n11129 1.355
R17400 VDD.n11229 VDD.n11228 1.355
R17401 VDD.n6544 VDD.n5779 1.35125
R17402 VDD.n5690 VDD.n4925 1.35125
R17403 VDD.n4904 VDD.n4139 1.35125
R17404 VDD.n4050 VDD.n3285 1.35125
R17405 VDD.n3264 VDD.n2499 1.35125
R17406 VDD.n2409 VDD.n1644 1.35125
R17407 VDD.n1200 VDD.n1197 1.35125
R17408 VDD.n754 VDD.n751 1.35125
R17409 VDD.n7967 VDD.n7966 1.34787
R17410 VDD.n7939 VDD.n7839 1.34787
R17411 VDD.n7916 VDD.n7852 1.34787
R17412 VDD.n7875 VDD.n7873 1.34787
R17413 VDD.n11458 VDD.n7714 1.34787
R17414 VDD.n11490 VDD.n7693 1.34787
R17415 VDD.n11517 VDD.n11516 1.34787
R17416 VDD.n7666 VDD.n7661 1.34787
R17417 VDD.n11570 VDD.n7652 1.34787
R17418 VDD.n9448 VDD.n9447 1.3466
R17419 VDD.n10922 VDD.n10921 1.3449
R17420 VDD.n9867 VDD.n9829 1.34458
R17421 VDD.n9867 VDD.n9831 1.34227
R17422 VDD.n6020 VDD.n6017 1.33615
R17423 VDD.n5166 VDD.n5163 1.33615
R17424 VDD.n4380 VDD.n4377 1.33615
R17425 VDD.n3526 VDD.n3523 1.33615
R17426 VDD.n2740 VDD.n2737 1.33615
R17427 VDD.n1885 VDD.n1882 1.33615
R17428 VDD.n1635 VDD.n1634 1.33615
R17429 VDD.n407 VDD.n406 1.33615
R17430 VDD.n10260 VDD.n10259 1.32759
R17431 VDD.n10306 VDD.n10224 1.32759
R17432 VDD.n10358 VDD.n10199 1.32759
R17433 VDD.n10405 VDD.n10404 1.32759
R17434 VDD.n6387 VDD.n6386 1.32203
R17435 VDD.n5954 VDD.n5948 1.32203
R17436 VDD.n5533 VDD.n5532 1.32203
R17437 VDD.n5100 VDD.n5094 1.32203
R17438 VDD.n4747 VDD.n4746 1.32203
R17439 VDD.n4314 VDD.n4308 1.32203
R17440 VDD.n3893 VDD.n3892 1.32203
R17441 VDD.n3460 VDD.n3454 1.32203
R17442 VDD.n3107 VDD.n3106 1.32203
R17443 VDD.n2674 VDD.n2668 1.32203
R17444 VDD.n2252 VDD.n2251 1.32203
R17445 VDD.n1819 VDD.n1813 1.32203
R17446 VDD.n1371 VDD.n1369 1.32203
R17447 VDD.n1570 VDD.n1569 1.32203
R17448 VDD.n143 VDD.n141 1.32203
R17449 VDD.n342 VDD.n341 1.32203
R17450 VDD.n6633 VDD.n6632 1.28287
R17451 VDD.n9118 VDD.n9089 1.26837
R17452 VDD.n6156 VDD.n6155 1.25267
R17453 VDD.n5302 VDD.n5301 1.25267
R17454 VDD.n4516 VDD.n4515 1.25267
R17455 VDD.n3662 VDD.n3661 1.25267
R17456 VDD.n2876 VDD.n2875 1.25267
R17457 VDD.n2021 VDD.n2020 1.25267
R17458 VDD.n1314 VDD.n1311 1.25267
R17459 VDD.n86 VDD.n83 1.25267
R17460 VDD.n6388 VDD.n6387 1.24652
R17461 VDD.n5951 VDD.n5948 1.24652
R17462 VDD.n5534 VDD.n5533 1.24652
R17463 VDD.n5097 VDD.n5094 1.24652
R17464 VDD.n4748 VDD.n4747 1.24652
R17465 VDD.n4311 VDD.n4308 1.24652
R17466 VDD.n3894 VDD.n3893 1.24652
R17467 VDD.n3457 VDD.n3454 1.24652
R17468 VDD.n3108 VDD.n3107 1.24652
R17469 VDD.n2671 VDD.n2668 1.24652
R17470 VDD.n2253 VDD.n2252 1.24652
R17471 VDD.n1816 VDD.n1813 1.24652
R17472 VDD.n1369 VDD.n1368 1.24652
R17473 VDD.n1570 VDD.n1414 1.24652
R17474 VDD.n141 VDD.n140 1.24652
R17475 VDD.n342 VDD.n186 1.24652
R17476 VDD.n10267 VDD.n10248 1.24197
R17477 VDD.n10314 VDD.n10313 1.24197
R17478 VDD.n10363 VDD.n10195 1.24197
R17479 VDD.n10412 VDD.n10169 1.24197
R17480 VDD.n12374 VDD.n12373 1.22988
R17481 VDD.n12323 VDD.n7005 1.22988
R17482 VDD.n12277 VDD.n7044 1.22988
R17483 VDD.n7150 VDD.n7149 1.22988
R17484 VDD.n7205 VDD.n7096 1.22988
R17485 VDD.n12244 VDD.n7076 1.22988
R17486 VDD.n12197 VDD.n12196 1.22988
R17487 VDD.n12146 VDD.n7338 1.22988
R17488 VDD.n6335 VDD.n6334 1.22485
R17489 VDD.n6334 VDD.n6017 1.22485
R17490 VDD.n6021 VDD.n6020 1.22485
R17491 VDD.n6292 VDD.n6291 1.22485
R17492 VDD.n6323 VDD.n6301 1.22485
R17493 VDD.n5481 VDD.n5480 1.22485
R17494 VDD.n5480 VDD.n5163 1.22485
R17495 VDD.n5167 VDD.n5166 1.22485
R17496 VDD.n5438 VDD.n5437 1.22485
R17497 VDD.n5469 VDD.n5447 1.22485
R17498 VDD.n4695 VDD.n4694 1.22485
R17499 VDD.n4694 VDD.n4377 1.22485
R17500 VDD.n4381 VDD.n4380 1.22485
R17501 VDD.n4652 VDD.n4651 1.22485
R17502 VDD.n4683 VDD.n4661 1.22485
R17503 VDD.n3841 VDD.n3840 1.22485
R17504 VDD.n3840 VDD.n3523 1.22485
R17505 VDD.n3527 VDD.n3526 1.22485
R17506 VDD.n3798 VDD.n3797 1.22485
R17507 VDD.n3829 VDD.n3807 1.22485
R17508 VDD.n3055 VDD.n3054 1.22485
R17509 VDD.n3054 VDD.n2737 1.22485
R17510 VDD.n2741 VDD.n2740 1.22485
R17511 VDD.n3012 VDD.n3011 1.22485
R17512 VDD.n3043 VDD.n3021 1.22485
R17513 VDD.n2200 VDD.n2199 1.22485
R17514 VDD.n2199 VDD.n1882 1.22485
R17515 VDD.n1886 VDD.n1885 1.22485
R17516 VDD.n2157 VDD.n2156 1.22485
R17517 VDD.n2188 VDD.n2166 1.22485
R17518 VDD.n1616 VDD.n1613 1.22485
R17519 VDD.n1635 VDD.n1616 1.22485
R17520 VDD.n1634 VDD.n1631 1.22485
R17521 VDD.n1628 VDD.n1625 1.22485
R17522 VDD.n1622 VDD.n1619 1.22485
R17523 VDD.n388 VDD.n385 1.22485
R17524 VDD.n407 VDD.n388 1.22485
R17525 VDD.n406 VDD.n403 1.22485
R17526 VDD.n400 VDD.n397 1.22485
R17527 VDD.n394 VDD.n391 1.22485
R17528 VDD.n11667 VDD.n7602 1.21955
R17529 VDD.n11692 VDD.n7585 1.21955
R17530 VDD.n11724 VDD.n7571 1.21955
R17531 VDD.n7559 VDD.n7554 1.21955
R17532 VDD.n11781 VDD.n7540 1.21955
R17533 VDD.n11806 VDD.n7523 1.21955
R17534 VDD.n11838 VDD.n7509 1.21955
R17535 VDD.n7497 VDD.n7492 1.21955
R17536 VDD.n11895 VDD.n7478 1.21955
R17537 VDD.n11920 VDD.n7461 1.21955
R17538 VDD.n11952 VDD.n7447 1.21955
R17539 VDD.n7435 VDD.n7430 1.21955
R17540 VDD.n12009 VDD.n7416 1.21955
R17541 VDD.n12034 VDD.n7399 1.21955
R17542 VDD.n12066 VDD.n7385 1.21955
R17543 VDD.n11604 VDD.n11602 1.21313
R17544 VDD.n11630 VDD.n11629 1.21313
R17545 VDD.n8069 VDD.n8068 1.20446
R17546 VDD.n8050 VDD.n8046 1.20446
R17547 VDD.n8316 VDD.n8010 1.20446
R17548 VDD.n8491 VDD.n8490 1.20446
R17549 VDD.n8447 VDD.n8384 1.20446
R17550 VDD.n8422 VDD.n8414 1.20446
R17551 VDD.t148 VDD.t16 1.19962
R17552 VDD.n10256 VDD.n10252 1.15635
R17553 VDD.n10305 VDD.n10228 1.15635
R17554 VDD.n10355 VDD.n10354 1.15635
R17555 VDD.n10401 VDD.n10173 1.15635
R17556 VDD.n9983 VDD.n6573 1.15386
R17557 VDD.n8175 VDD.n8136 1.15182
R17558 VDD.n11413 VDD.n8633 1.15182
R17559 VDD.n11347 VDD.n11346 1.15182
R17560 VDD.n11278 VDD.n11153 1.15182
R17561 VDD.n10938 VDD.n10937 1.13717
R17562 VDD.n10921 VDD.n10920 1.13717
R17563 VDD.n10913 VDD.n10912 1.13717
R17564 VDD.n9449 VDD.n9448 1.13717
R17565 VDD.n9228 VDD.n9227 1.13717
R17566 VDD.n10899 VDD.n10898 1.13717
R17567 VDD.n9879 VDD.n9878 1.13717
R17568 VDD.n9868 VDD.n9867 1.13717
R17569 VDD.n10472 VDD.n10471 1.13602
R17570 VDD.n10052 VDD.n10033 1.12991
R17571 VDD.n10052 VDD.n10034 1.12991
R17572 VDD.n10611 VDD.n10592 1.12991
R17573 VDD.n10611 VDD.n10593 1.12991
R17574 VDD.n10555 VDD.n10554 1.12991
R17575 VDD.n10554 VDD.n10535 1.12991
R17576 VDD.n9624 VDD.n9568 1.12991
R17577 VDD.n9624 VDD.n9565 1.12991
R17578 VDD.n9692 VDD.n9691 1.12991
R17579 VDD.n9706 VDD.n9705 1.12991
R17580 VDD.n10856 VDD.n10855 1.12991
R17581 VDD.n10842 VDD.n10841 1.12991
R17582 VDD.n10740 VDD.n10723 1.12991
R17583 VDD.n10740 VDD.n10739 1.12991
R17584 VDD.n8907 VDD.n8906 1.12991
R17585 VDD.n9383 VDD.n9378 1.12991
R17586 VDD.n9156 VDD.n9084 1.12991
R17587 VDD.n9101 VDD.n9093 1.12991
R17588 VDD.n8533 VDD.n7788 1.12991
R17589 VDD.n8507 VDD.n8506 1.12991
R17590 VDD.n12483 VDD.n12482 1.12991
R17591 VDD.n12466 VDD.n12437 1.12991
R17592 VDD.n12442 VDD.n12437 1.12991
R17593 VDD.n6262 VDD.n6054 1.11541
R17594 VDD.n6263 VDD.n6052 1.11541
R17595 VDD.n6269 VDD.n6268 1.11541
R17596 VDD.n6274 VDD.n6050 1.11541
R17597 VDD.n6276 VDD.n6275 1.11541
R17598 VDD.n6287 VDD.n6047 1.11541
R17599 VDD.n5408 VDD.n5200 1.11541
R17600 VDD.n5409 VDD.n5198 1.11541
R17601 VDD.n5415 VDD.n5414 1.11541
R17602 VDD.n5420 VDD.n5196 1.11541
R17603 VDD.n5422 VDD.n5421 1.11541
R17604 VDD.n5433 VDD.n5193 1.11541
R17605 VDD.n4622 VDD.n4414 1.11541
R17606 VDD.n4623 VDD.n4412 1.11541
R17607 VDD.n4629 VDD.n4628 1.11541
R17608 VDD.n4634 VDD.n4410 1.11541
R17609 VDD.n4636 VDD.n4635 1.11541
R17610 VDD.n4647 VDD.n4407 1.11541
R17611 VDD.n3768 VDD.n3560 1.11541
R17612 VDD.n3769 VDD.n3558 1.11541
R17613 VDD.n3775 VDD.n3774 1.11541
R17614 VDD.n3780 VDD.n3556 1.11541
R17615 VDD.n3782 VDD.n3781 1.11541
R17616 VDD.n3793 VDD.n3553 1.11541
R17617 VDD.n2982 VDD.n2774 1.11541
R17618 VDD.n2983 VDD.n2772 1.11541
R17619 VDD.n2989 VDD.n2988 1.11541
R17620 VDD.n2994 VDD.n2770 1.11541
R17621 VDD.n2996 VDD.n2995 1.11541
R17622 VDD.n3007 VDD.n2767 1.11541
R17623 VDD.n2127 VDD.n1919 1.11541
R17624 VDD.n2128 VDD.n1917 1.11541
R17625 VDD.n2134 VDD.n2133 1.11541
R17626 VDD.n2139 VDD.n1915 1.11541
R17627 VDD.n2141 VDD.n2140 1.11541
R17628 VDD.n2152 VDD.n1912 1.11541
R17629 VDD.n989 VDD.n986 1.11541
R17630 VDD.n993 VDD.n991 1.11541
R17631 VDD.n999 VDD.n996 1.11541
R17632 VDD.n1004 VDD.n1001 1.11541
R17633 VDD.n1011 VDD.n1007 1.11541
R17634 VDD.n1015 VDD.n1013 1.11541
R17635 VDD.n543 VDD.n540 1.11541
R17636 VDD.n547 VDD.n545 1.11541
R17637 VDD.n553 VDD.n550 1.11541
R17638 VDD.n558 VDD.n555 1.11541
R17639 VDD.n565 VDD.n561 1.11541
R17640 VDD.n569 VDD.n567 1.11541
R17641 VDD.n10157 VDD.n10156 1.11019
R17642 VDD.n10531 VDD.n10154 1.10959
R17643 VDD.n8823 VDD.n8822 1.10923
R17644 VDD.n10114 VDD.n10005 1.10918
R17645 VDD.n10080 VDD.n10017 1.10899
R17646 VDD.n5754 VDD 1.09833
R17647 VDD.n12777 VDD.n12776 1.09663
R17648 VDD.n12400 VDD.n12399 1.08525
R17649 VDD.n12351 VDD.n6982 1.08525
R17650 VDD.n7025 VDD.n7024 1.08525
R17651 VDD.n12256 VDD.n12255 1.08525
R17652 VDD.n7177 VDD.n7176 1.08525
R17653 VDD.n7231 VDD.n7086 1.08525
R17654 VDD.n12223 VDD.n12222 1.08525
R17655 VDD.n12174 VDD.n7315 1.08525
R17656 VDD.n8608 VDD.n7727 1.0841
R17657 VDD.n8713 VDD.n8712 1.0841
R17658 VDD.n11128 VDD.n11111 1.0841
R17659 VDD.n11227 VDD.n11222 1.0841
R17660 VDD.n7962 VDD.n7821 1.07839
R17661 VDD.n7940 VDD.n7837 1.07839
R17662 VDD.n7915 VDD.n7856 1.07839
R17663 VDD.n7893 VDD.n7871 1.07839
R17664 VDD.n11465 VDD.n7709 1.07839
R17665 VDD.n11491 VDD.n11489 1.07839
R17666 VDD.n11522 VDD.n7679 1.07839
R17667 VDD.n11545 VDD.n11544 1.07839
R17668 VDD.n11577 VDD.n7647 1.07839
R17669 VDD.n12698 VDD.n6610 1.07073
R17670 VDD.n10268 VDD.n10246 1.07073
R17671 VDD.n10317 VDD.n10220 1.07073
R17672 VDD.n10367 VDD.n10366 1.07073
R17673 VDD.n10413 VDD.n10167 1.07073
R17674 VDD.n12775 VDD.n6573 1.04401
R17675 VDD.n12774 VDD.n12773 1.04351
R17676 VDD.n10471 VDD.n10470 1.04225
R17677 VDD.n9448 VDD.n9350 1.02922
R17678 VDD.n10640 VDD.n10136 1.0272
R17679 VDD.n10921 VDD.n9325 1.02676
R17680 VDD.n10640 VDD.n10133 1.02649
R17681 VDD.n12772 VDD.n6575 1.02165
R17682 VDD.n12702 VDD.n6610 0.997903
R17683 VDD.n9649 VDD.n9645 0.994314
R17684 VDD.n9668 VDD.n9667 0.994314
R17685 VDD.n10792 VDD.n10788 0.994314
R17686 VDD.n10811 VDD.n10810 0.994314
R17687 VDD.n8868 VDD.n8864 0.994314
R17688 VDD.n8961 VDD.n8861 0.994314
R17689 VDD.n8965 VDD.n8857 0.994314
R17690 VDD.n9007 VDD.n9006 0.994314
R17691 VDD.n8984 VDD.n8834 0.994314
R17692 VDD.n8987 VDD.n8829 0.994314
R17693 VDD.n9279 VDD.n9275 0.994314
R17694 VDD.n9409 VDD.n9405 0.994314
R17695 VDD.n10255 VDD.n10253 0.985115
R17696 VDD.n10302 VDD.n10301 0.985115
R17697 VDD.n10351 VDD.n10201 0.985115
R17698 VDD.n10400 VDD.n10175 0.985115
R17699 VDD.n8226 VDD.n8072 0.950995
R17700 VDD.n8267 VDD.n8266 0.950995
R17701 VDD.n8313 VDD.n8012 0.950995
R17702 VDD.n8343 VDD.n8342 0.950995
R17703 VDD.n8451 VDD.n8450 0.950995
R17704 VDD.n8420 VDD.n8417 0.950995
R17705 VDD.n11668 VDD.n7600 0.948648
R17706 VDD.n11693 VDD.n11691 0.948648
R17707 VDD.n11723 VDD.n7572 0.948648
R17708 VDD.n11749 VDD.n11748 0.948648
R17709 VDD.n11782 VDD.n7538 0.948648
R17710 VDD.n11807 VDD.n11805 0.948648
R17711 VDD.n11837 VDD.n7510 0.948648
R17712 VDD.n11863 VDD.n11862 0.948648
R17713 VDD.n11896 VDD.n7476 0.948648
R17714 VDD.n11921 VDD.n11919 0.948648
R17715 VDD.n11951 VDD.n7448 0.948648
R17716 VDD.n11977 VDD.n11976 0.948648
R17717 VDD.n12010 VDD.n7414 0.948648
R17718 VDD.n12035 VDD.n12033 0.948648
R17719 VDD.n12065 VDD.n7386 0.948648
R17720 VDD.n7639 VDD.n7634 0.943658
R17721 VDD.n11637 VDD.n7617 0.943658
R17722 VDD.n10327 VDD.n10326 0.942306
R17723 VDD.n12418 VDD.n12417 0.942306
R17724 VDD.n6970 VDD.n6965 0.940613
R17725 VDD.n12322 VDD.n7006 0.940613
R17726 VDD.n12274 VDD.n12273 0.940613
R17727 VDD.n7154 VDD.n7118 0.940613
R17728 VDD.n7209 VDD.n7208 0.940613
R17729 VDD.n12241 VDD.n12240 0.940613
R17730 VDD.n7303 VDD.n7299 0.940613
R17731 VDD.n12145 VDD.n7339 0.940613
R17732 VDD.n5798 VDD.n5794 0.934239
R17733 VDD.n6538 VDD.n6537 0.934239
R17734 VDD.n6534 VDD.n5799 0.934239
R17735 VDD.n6533 VDD.n5802 0.934239
R17736 VDD.n6529 VDD.n6528 0.934239
R17737 VDD.n6524 VDD.n5805 0.934239
R17738 VDD.n4944 VDD.n4940 0.934239
R17739 VDD.n5684 VDD.n5683 0.934239
R17740 VDD.n5680 VDD.n4945 0.934239
R17741 VDD.n5679 VDD.n4948 0.934239
R17742 VDD.n5675 VDD.n5674 0.934239
R17743 VDD.n5670 VDD.n4951 0.934239
R17744 VDD.n4158 VDD.n4154 0.934239
R17745 VDD.n4898 VDD.n4897 0.934239
R17746 VDD.n4894 VDD.n4159 0.934239
R17747 VDD.n4893 VDD.n4162 0.934239
R17748 VDD.n4889 VDD.n4888 0.934239
R17749 VDD.n4884 VDD.n4165 0.934239
R17750 VDD.n3304 VDD.n3300 0.934239
R17751 VDD.n4044 VDD.n4043 0.934239
R17752 VDD.n4040 VDD.n3305 0.934239
R17753 VDD.n4039 VDD.n3308 0.934239
R17754 VDD.n4035 VDD.n4034 0.934239
R17755 VDD.n4030 VDD.n3311 0.934239
R17756 VDD.n2518 VDD.n2514 0.934239
R17757 VDD.n3258 VDD.n3257 0.934239
R17758 VDD.n3254 VDD.n2519 0.934239
R17759 VDD.n3253 VDD.n2522 0.934239
R17760 VDD.n3249 VDD.n3248 0.934239
R17761 VDD.n3244 VDD.n2525 0.934239
R17762 VDD.n1663 VDD.n1659 0.934239
R17763 VDD.n2403 VDD.n2402 0.934239
R17764 VDD.n2399 VDD.n1664 0.934239
R17765 VDD.n2398 VDD.n1667 0.934239
R17766 VDD.n2394 VDD.n2393 0.934239
R17767 VDD.n2389 VDD.n1670 0.934239
R17768 VDD.n1187 VDD.n1184 0.934239
R17769 VDD.n1180 VDD.n1177 0.934239
R17770 VDD.n1175 VDD.n1173 0.934239
R17771 VDD.n1170 VDD.n1167 0.934239
R17772 VDD.n1165 VDD.n1163 0.934239
R17773 VDD.n1160 VDD.n1157 0.934239
R17774 VDD.n741 VDD.n738 0.934239
R17775 VDD.n734 VDD.n731 0.934239
R17776 VDD.n729 VDD.n727 0.934239
R17777 VDD.n724 VDD.n721 0.934239
R17778 VDD.n719 VDD.n717 0.934239
R17779 VDD.n714 VDD.n711 0.934239
R17780 VDD.n8499 VDD.n8498 0.926297
R17781 VDD.n8598 VDD.n7747 0.926297
R17782 VDD.n7748 VDD.n7718 0.926297
R17783 VDD.n11447 VDD.n7719 0.926297
R17784 VDD.n11441 VDD.n7728 0.926297
R17785 VDD.n9172 VDD.n7729 0.926297
R17786 VDD.n11435 VDD.n7735 0.926297
R17787 VDD.n9168 VDD.n8616 0.926297
R17788 VDD.n11426 VDD.n11425 0.926297
R17789 VDD.n11422 VDD.n8617 0.926297
R17790 VDD.n8628 VDD.n8623 0.926297
R17791 VDD.n11416 VDD.n8629 0.926297
R17792 VDD.n8647 VDD.n8630 0.926297
R17793 VDD.n11407 VDD.n11406 0.926297
R17794 VDD.n11403 VDD.n8648 0.926297
R17795 VDD.n9176 VDD.n8654 0.926297
R17796 VDD.n11397 VDD.n8659 0.926297
R17797 VDD.n8668 VDD.n8660 0.926297
R17798 VDD.n11391 VDD.n11390 0.926297
R17799 VDD.n11382 VDD.n11381 0.926297
R17800 VDD.n11378 VDD.n8686 0.926297
R17801 VDD.n8700 VDD.n8692 0.926297
R17802 VDD.n11372 VDD.n8701 0.926297
R17803 VDD.n8719 VDD.n8702 0.926297
R17804 VDD.n11363 VDD.n11362 0.926297
R17805 VDD.n11359 VDD.n11027 0.926297
R17806 VDD.n11033 VDD.n11028 0.926297
R17807 VDD.n11353 VDD.n11034 0.926297
R17808 VDD.n11052 VDD.n11035 0.926297
R17809 VDD.n11344 VDD.n11343 0.926297
R17810 VDD.n11340 VDD.n11053 0.926297
R17811 VDD.n11096 VDD.n11095 0.926297
R17812 VDD.n11334 VDD.n11063 0.926297
R17813 VDD.n11074 VDD.n11064 0.926297
R17814 VDD.n11325 VDD.n11075 0.926297
R17815 VDD.n11080 VDD.n11076 0.926297
R17816 VDD.n11319 VDD.n11081 0.926297
R17817 VDD.n11310 VDD.n11309 0.926297
R17818 VDD.n11306 VDD.n11106 0.926297
R17819 VDD.n11117 VDD.n11112 0.926297
R17820 VDD.n11300 VDD.n11118 0.926297
R17821 VDD.n11136 VDD.n11119 0.926297
R17822 VDD.n11291 VDD.n11290 0.926297
R17823 VDD.n11287 VDD.n11142 0.926297
R17824 VDD.n11148 VDD.n11143 0.926297
R17825 VDD.n11281 VDD.n11149 0.926297
R17826 VDD.n11167 VDD.n11150 0.926297
R17827 VDD.n11272 VDD.n11271 0.926297
R17828 VDD.n11268 VDD.n11168 0.926297
R17829 VDD.n11179 VDD.n11174 0.926297
R17830 VDD.n11262 VDD.n11180 0.926297
R17831 VDD.n11189 VDD.n11181 0.926297
R17832 VDD.n11256 VDD.n11255 0.926297
R17833 VDD.n11206 VDD.n11190 0.926297
R17834 VDD.n11247 VDD.n11246 0.926297
R17835 VDD.n11243 VDD.n11207 0.926297
R17836 VDD.n11233 VDD.n11213 0.926297
R17837 VDD.n11232 VDD.n11214 0.926297
R17838 VDD.n12710 VDD.n6599 0.926297
R17839 VDD.n4113 VDD 0.913543
R17840 VDD.n5960 VDD.n5958 0.906695
R17841 VDD.n5963 VDD.n5962 0.906695
R17842 VDD.n5966 VDD.n5946 0.906695
R17843 VDD.n5969 VDD.n5968 0.906695
R17844 VDD.n5972 VDD.n5944 0.906695
R17845 VDD.n5978 VDD.n5974 0.906695
R17846 VDD.n5106 VDD.n5104 0.906695
R17847 VDD.n5109 VDD.n5108 0.906695
R17848 VDD.n5112 VDD.n5092 0.906695
R17849 VDD.n5115 VDD.n5114 0.906695
R17850 VDD.n5118 VDD.n5090 0.906695
R17851 VDD.n5124 VDD.n5120 0.906695
R17852 VDD.n4320 VDD.n4318 0.906695
R17853 VDD.n4323 VDD.n4322 0.906695
R17854 VDD.n4326 VDD.n4306 0.906695
R17855 VDD.n4329 VDD.n4328 0.906695
R17856 VDD.n4332 VDD.n4304 0.906695
R17857 VDD.n4338 VDD.n4334 0.906695
R17858 VDD.n3466 VDD.n3464 0.906695
R17859 VDD.n3469 VDD.n3468 0.906695
R17860 VDD.n3472 VDD.n3452 0.906695
R17861 VDD.n3475 VDD.n3474 0.906695
R17862 VDD.n3478 VDD.n3450 0.906695
R17863 VDD.n3484 VDD.n3480 0.906695
R17864 VDD.n2680 VDD.n2678 0.906695
R17865 VDD.n2683 VDD.n2682 0.906695
R17866 VDD.n2686 VDD.n2666 0.906695
R17867 VDD.n2689 VDD.n2688 0.906695
R17868 VDD.n2692 VDD.n2664 0.906695
R17869 VDD.n2698 VDD.n2694 0.906695
R17870 VDD.n1825 VDD.n1823 0.906695
R17871 VDD.n1828 VDD.n1827 0.906695
R17872 VDD.n1831 VDD.n1811 0.906695
R17873 VDD.n1834 VDD.n1833 0.906695
R17874 VDD.n1837 VDD.n1809 0.906695
R17875 VDD.n1843 VDD.n1839 0.906695
R17876 VDD.n1563 VDD.n1560 0.906695
R17877 VDD.n1557 VDD.n1554 0.906695
R17878 VDD.n1552 VDD.n1549 0.906695
R17879 VDD.n1546 VDD.n1543 0.906695
R17880 VDD.n1541 VDD.n1538 0.906695
R17881 VDD.n1535 VDD.n1532 0.906695
R17882 VDD.n335 VDD.n332 0.906695
R17883 VDD.n329 VDD.n326 0.906695
R17884 VDD.n324 VDD.n321 0.906695
R17885 VDD.n318 VDD.n315 0.906695
R17886 VDD.n313 VDD.n310 0.906695
R17887 VDD.n307 VDD.n304 0.906695
R17888 VDD.n8824 VDD.n8823 0.903353
R17889 VDD.n8893 VDD.n8766 0.903353
R17890 VDD.n6699 VDD.n6698 0.902912
R17891 VDD.n8541 VDD.n8540 0.899959
R17892 VDD.n10272 VDD.n10271 0.899497
R17893 VDD.n10318 VDD.n10218 0.899497
R17894 VDD.n10370 VDD.n10191 0.899497
R17895 VDD.n10418 VDD.n10416 0.899497
R17896 VDD.n10947 VDD.n9225 0.884222
R17897 VDD.n10948 VDD.n10947 0.883499
R17898 VDD.n8172 VDD.n8137 0.880923
R17899 VDD.n11410 VDD.n11409 0.880923
R17900 VDD.n11057 VDD.n11056 0.880923
R17901 VDD.n11275 VDD.n11274 0.880923
R17902 VDD.n12089 VDD.n12088 0.880923
R17903 VDD.n8530 VDD.n8529 0.878931
R17904 VDD.n8510 VDD.n7802 0.878931
R17905 VDD.n5753 VDD.n5751 0.8405
R17906 VDD.n5751 VDD 0.8405
R17907 VDD.n4113 VDD.n4112 0.8405
R17908 VDD.n4112 VDD 0.8405
R17909 VDD.n11019 VDD.n8737 0.825441
R17910 VDD.n8564 VDD.n7767 0.824262
R17911 VDD.n11007 VDD.n8750 0.82077
R17912 VDD.n12683 VDD.n6710 0.813878
R17913 VDD.n10298 VDD.n10230 0.813878
R17914 VDD.n10350 VDD.n10203 0.813878
R17915 VDD.n10397 VDD.n10396 0.813878
R17916 VDD.n11444 VDD.n7723 0.813198
R17917 VDD.n8711 VDD.n8691 0.813198
R17918 VDD.n11109 VDD.n11089 0.813198
R17919 VDD.n11224 VDD.n11212 0.813198
R17920 VDD.n12704 VDD.n12703 0.813198
R17921 VDD.n7961 VDD.n7825 0.808921
R17922 VDD.n7944 VDD.n7943 0.808921
R17923 VDD.n7912 VDD.n7911 0.808921
R17924 VDD.n7894 VDD.n7869 0.808921
R17925 VDD.n11466 VDD.n7707 0.808921
R17926 VDD.n7701 VDD.n7696 0.808921
R17927 VDD.n11521 VDD.n7680 0.808921
R17928 VDD.n11539 VDD.n7665 0.808921
R17929 VDD.n11578 VDD.n7645 0.808921
R17930 VDD.n6943 VDD.n6942 0.79598
R17931 VDD.n12352 VDD.n6980 0.79598
R17932 VDD.n12306 VDD.n7018 0.79598
R17933 VDD.n7064 VDD.n7063 0.79598
R17934 VDD.n7171 VDD.n7110 0.79598
R17935 VDD.n7230 VDD.n7088 0.79598
R17936 VDD.n7277 VDD.n7276 0.79598
R17937 VDD.n12175 VDD.n7313 0.79598
R17938 VDD.n11362 VDD.n8721 0.79404
R17939 VDD.n9837 VDD.n9833 0.775778
R17940 VDD.n10680 VDD.n10679 0.775778
R17941 VDD.n5746 VDD.n5745 0.761777
R17942 VDD.n4106 VDD.n4105 0.761777
R17943 VDD.n2465 VDD.n2464 0.761777
R17944 VDD.n825 VDD.n824 0.761777
R17945 VDD.n8548 VDD.n7780 0.761581
R17946 VDD.n10078 VDD.n10021 0.753441
R17947 VDD.n10029 VDD.n10013 0.753441
R17948 VDD.n10096 VDD.n10089 0.753441
R17949 VDD.n10108 VDD.n10107 0.753441
R17950 VDD.n10142 VDD.n10139 0.753441
R17951 VDD.n10618 VDD.n10617 0.753441
R17952 VDD.n10516 VDD.n10514 0.753441
R17953 VDD.n10507 VDD.n10506 0.753441
R17954 VDD.n9648 VDD.n9646 0.753441
R17955 VDD.n9655 VDD.n9646 0.753441
R17956 VDD.n9670 VDD.n9669 0.753441
R17957 VDD.n9669 VDD.n9661 0.753441
R17958 VDD.n10791 VDD.n10789 0.753441
R17959 VDD.n10798 VDD.n10789 0.753441
R17960 VDD.n10813 VDD.n10812 0.753441
R17961 VDD.n10812 VDD.n10804 0.753441
R17962 VDD.n8916 VDD.n8771 0.753441
R17963 VDD.n8867 VDD.n8865 0.753441
R17964 VDD.n8874 VDD.n8865 0.753441
R17965 VDD.n8959 VDD.n8958 0.753441
R17966 VDD.n8960 VDD.n8959 0.753441
R17967 VDD.n8964 VDD.n8858 0.753441
R17968 VDD.n8972 VDD.n8858 0.753441
R17969 VDD.n9009 VDD.n9008 0.753441
R17970 VDD.n9008 VDD.n9000 0.753441
R17971 VDD.n8982 VDD.n8981 0.753441
R17972 VDD.n8983 VDD.n8982 0.753441
R17973 VDD.n8986 VDD.n8830 0.753441
R17974 VDD.n8994 VDD.n8830 0.753441
R17975 VDD.n9040 VDD.n9039 0.753441
R17976 VDD.n8815 VDD.n8811 0.753441
R17977 VDD.n8902 VDD.n8901 0.753441
R17978 VDD.n9309 VDD.n9308 0.753441
R17979 VDD.n9278 VDD.n9276 0.753441
R17980 VDD.n9285 VDD.n9276 0.753441
R17981 VDD.n9332 VDD.n9331 0.753441
R17982 VDD.n9379 VDD.n9355 0.753441
R17983 VDD.n9408 VDD.n9406 0.753441
R17984 VDD.n9415 VDD.n9406 0.753441
R17985 VDD.n9100 VDD.n9088 0.753441
R17986 VDD.n9121 VDD.n9117 0.753441
R17987 VDD.n6565 VDD.n6564 0.751569
R17988 VDD.n6256 VDD.n6255 0.750919
R17989 VDD.n6556 VDD.n5779 0.750919
R17990 VDD.n5402 VDD.n5401 0.750919
R17991 VDD.n5702 VDD.n4925 0.750919
R17992 VDD.n4616 VDD.n4615 0.750919
R17993 VDD.n4916 VDD.n4139 0.750919
R17994 VDD.n3762 VDD.n3761 0.750919
R17995 VDD.n4062 VDD.n3285 0.750919
R17996 VDD.n2976 VDD.n2975 0.750919
R17997 VDD.n3276 VDD.n2499 0.750919
R17998 VDD.n2121 VDD.n2120 0.750919
R17999 VDD.n2421 VDD.n1644 0.750919
R18000 VDD.n983 VDD.n981 0.750919
R18001 VDD.n1225 VDD.n1200 0.750919
R18002 VDD.n537 VDD.n535 0.750919
R18003 VDD.n779 VDD.n754 0.750919
R18004 VDD.n9042 VDD.n8780 0.743006
R18005 VDD.n9268 VDD.n9248 0.743006
R18006 VDD.n8929 VDD.n8885 0.742904
R18007 VDD.n10275 VDD.n10242 0.728259
R18008 VDD.n10322 VDD.n10321 0.728259
R18009 VDD.n10371 VDD.n10189 0.728259
R18010 VDD.n10417 VDD.n6926 0.728259
R18011 VDD.n9080 VDD.n9078 0.724685
R18012 VDD.n9165 VDD.n9080 0.724297
R18013 VDD.n6699 VDD.n6623 0.71293
R18014 VDD.n6256 VDD.n6055 0.708038
R18015 VDD.n5402 VDD.n5201 0.708038
R18016 VDD.n4616 VDD.n4415 0.708038
R18017 VDD.n3762 VDD.n3561 0.708038
R18018 VDD.n2976 VDD.n2775 0.708038
R18019 VDD.n2121 VDD.n1920 0.708038
R18020 VDD.n981 VDD.n980 0.708038
R18021 VDD.n535 VDD.n534 0.708038
R18022 VDD.n6517 VDD.n5808 0.700804
R18023 VDD.n5663 VDD.n4954 0.700804
R18024 VDD.n4877 VDD.n4168 0.700804
R18025 VDD.n4023 VDD.n3314 0.700804
R18026 VDD.n3237 VDD.n2528 0.700804
R18027 VDD.n2382 VDD.n1673 0.700804
R18028 VDD.n1153 VDD.n1150 0.700804
R18029 VDD.n707 VDD.n704 0.700804
R18030 VDD.n10659 VDD.n9983 0.699924
R18031 VDD.n8223 VDD.n8221 0.69753
R18032 VDD.n8271 VDD.n8270 0.69753
R18033 VDD.n8018 VDD.n8017 0.69753
R18034 VDD.n8481 VDD.n8347 0.69753
R18035 VDD.n8380 VDD.n8377 0.69753
R18036 VDD.n8415 VDD.n7763 0.69753
R18037 VDD.n11020 VDD.n11019 0.692441
R18038 VDD.n11007 VDD.n8753 0.689368
R18039 VDD.n10431 VDD.n10430 0.687554
R18040 VDD.n5754 VDD 0.682932
R18041 VDD.n5754 VDD 0.682932
R18042 VDD.n10116 VDD.n10083 0.682531
R18043 VDD.n9769 VDD.n9768 0.682531
R18044 VDD.n9778 VDD.n9777 0.682531
R18045 VDD.n9796 VDD.n9795 0.682531
R18046 VDD.n9816 VDD.n9815 0.682531
R18047 VDD.n9890 VDD.n9454 0.6825
R18048 VDD.n9846 VDD.n9462 0.6825
R18049 VDD.n9323 VDD.n9234 0.6825
R18050 VDD.n5975 VDD.n5877 0.680146
R18051 VDD.n5121 VDD.n5023 0.680146
R18052 VDD.n4335 VDD.n4237 0.680146
R18053 VDD.n3481 VDD.n3383 0.680146
R18054 VDD.n2695 VDD.n2597 0.680146
R18055 VDD.n1840 VDD.n1742 0.680146
R18056 VDD.n1527 VDD.n1525 0.680146
R18057 VDD.n299 VDD.n297 0.680146
R18058 VDD.n11673 VDD.n11671 0.677749
R18059 VDD.n7593 VDD.n7588 0.677749
R18060 VDD.n11730 VDD.n7567 0.677749
R18061 VDD.n11743 VDD.n7558 0.677749
R18062 VDD.n11787 VDD.n11785 0.677749
R18063 VDD.n7531 VDD.n7526 0.677749
R18064 VDD.n11844 VDD.n7505 0.677749
R18065 VDD.n11857 VDD.n7496 0.677749
R18066 VDD.n11901 VDD.n11899 0.677749
R18067 VDD.n7469 VDD.n7464 0.677749
R18068 VDD.n11958 VDD.n7443 0.677749
R18069 VDD.n11971 VDD.n7434 0.677749
R18070 VDD.n12015 VDD.n12013 0.677749
R18071 VDD.n7407 VDD.n7402 0.677749
R18072 VDD.n12072 VDD.n7381 0.677749
R18073 VDD.n11596 VDD.n11595 0.674184
R18074 VDD.n11636 VDD.n7618 0.674184
R18075 VDD.t67 VDD.n8669 0.661784
R18076 VDD.t55 VDD.n11082 0.661784
R18077 VDD.n12367 VDD.n6971 0.651347
R18078 VDD.n12319 VDD.n12318 0.651347
R18079 VDD.n7051 VDD.n7047 0.651347
R18080 VDD.n7155 VDD.n7116 0.651347
R18081 VDD.n7215 VDD.n7094 0.651347
R18082 VDD.n7264 VDD.n7260 0.651347
R18083 VDD.n12190 VDD.n7304 0.651347
R18084 VDD.n12142 VDD.n12141 0.651347
R18085 VDD.n12414 VDD.n12413 0.647691
R18086 VDD.n6562 VDD.n6561 0.64299
R18087 VDD.n6564 VDD.n4921 0.64299
R18088 VDD.n6565 VDD.n3281 0.64299
R18089 VDD.n6566 VDD.n1640 0.64299
R18090 VDD.n12684 VDD.n6707 0.64264
R18091 VDD.n10297 VDD.n10232 0.64264
R18092 VDD.n10347 VDD.n10346 0.64264
R18093 VDD.n10393 VDD.n10177 0.64264
R18094 VDD VDD.n5771 0.63923
R18095 VDD VDD.n4131 0.63923
R18096 VDD VDD.n2491 0.63923
R18097 VDD VDD.n851 0.63923
R18098 VDD.n10159 VDD.n10156 0.629672
R18099 VDD.n8525 VDD.n7791 0.627951
R18100 VDD.n8511 VDD.n7800 0.627951
R18101 VDD.n12425 VDD.n12424 0.615996
R18102 VDD.n9216 VDD.n9213 0.614024
R18103 VDD.n5947 VDD.n5916 0.612674
R18104 VDD.n6361 VDD.n6360 0.612674
R18105 VDD.n6359 VDD.n6358 0.612674
R18106 VDD.n5933 VDD.n5921 0.612674
R18107 VDD.n5093 VDD.n5062 0.612674
R18108 VDD.n5507 VDD.n5506 0.612674
R18109 VDD.n5505 VDD.n5504 0.612674
R18110 VDD.n5079 VDD.n5067 0.612674
R18111 VDD.n4307 VDD.n4276 0.612674
R18112 VDD.n4721 VDD.n4720 0.612674
R18113 VDD.n4719 VDD.n4718 0.612674
R18114 VDD.n4293 VDD.n4281 0.612674
R18115 VDD.n3453 VDD.n3422 0.612674
R18116 VDD.n3867 VDD.n3866 0.612674
R18117 VDD.n3865 VDD.n3864 0.612674
R18118 VDD.n3439 VDD.n3427 0.612674
R18119 VDD.n2667 VDD.n2636 0.612674
R18120 VDD.n3081 VDD.n3080 0.612674
R18121 VDD.n3079 VDD.n3078 0.612674
R18122 VDD.n2653 VDD.n2641 0.612674
R18123 VDD.n1812 VDD.n1781 0.612674
R18124 VDD.n2226 VDD.n2225 0.612674
R18125 VDD.n2224 VDD.n2223 0.612674
R18126 VDD.n1798 VDD.n1786 0.612674
R18127 VDD.n1576 VDD.n1573 0.612674
R18128 VDD.n1582 VDD.n1579 0.612674
R18129 VDD.n1588 VDD.n1585 0.612674
R18130 VDD.n1594 VDD.n1591 0.612674
R18131 VDD.n348 VDD.n345 0.612674
R18132 VDD.n354 VDD.n351 0.612674
R18133 VDD.n360 VDD.n357 0.612674
R18134 VDD.n366 VDD.n363 0.612674
R18135 VDD.n8169 VDD.n8168 0.610024
R18136 VDD.n8652 VDD.n8651 0.610024
R18137 VDD.n11094 VDD.n11091 0.610024
R18138 VDD.n11172 VDD.n11171 0.610024
R18139 VDD.n6383 VDD.n5902 0.60463
R18140 VDD.n5913 VDD.n5911 0.60463
R18141 VDD.n6377 VDD.n6376 0.60463
R18142 VDD.n6374 VDD.n6373 0.60463
R18143 VDD.n6371 VDD.n6369 0.60463
R18144 VDD.n6367 VDD.n5914 0.60463
R18145 VDD.n5529 VDD.n5048 0.60463
R18146 VDD.n5059 VDD.n5057 0.60463
R18147 VDD.n5523 VDD.n5522 0.60463
R18148 VDD.n5520 VDD.n5519 0.60463
R18149 VDD.n5517 VDD.n5515 0.60463
R18150 VDD.n5513 VDD.n5060 0.60463
R18151 VDD.n4743 VDD.n4262 0.60463
R18152 VDD.n4273 VDD.n4271 0.60463
R18153 VDD.n4737 VDD.n4736 0.60463
R18154 VDD.n4734 VDD.n4733 0.60463
R18155 VDD.n4731 VDD.n4729 0.60463
R18156 VDD.n4727 VDD.n4274 0.60463
R18157 VDD.n3889 VDD.n3408 0.60463
R18158 VDD.n3419 VDD.n3417 0.60463
R18159 VDD.n3883 VDD.n3882 0.60463
R18160 VDD.n3880 VDD.n3879 0.60463
R18161 VDD.n3877 VDD.n3875 0.60463
R18162 VDD.n3873 VDD.n3420 0.60463
R18163 VDD.n3103 VDD.n2622 0.60463
R18164 VDD.n2633 VDD.n2631 0.60463
R18165 VDD.n3097 VDD.n3096 0.60463
R18166 VDD.n3094 VDD.n3093 0.60463
R18167 VDD.n3091 VDD.n3089 0.60463
R18168 VDD.n3087 VDD.n2634 0.60463
R18169 VDD.n2248 VDD.n1767 0.60463
R18170 VDD.n1778 VDD.n1776 0.60463
R18171 VDD.n2242 VDD.n2241 0.60463
R18172 VDD.n2239 VDD.n2238 0.60463
R18173 VDD.n2236 VDD.n2234 0.60463
R18174 VDD.n2232 VDD.n1779 0.60463
R18175 VDD.n1379 VDD.n1376 0.60463
R18176 VDD.n1385 VDD.n1382 0.60463
R18177 VDD.n1390 VDD.n1387 0.60463
R18178 VDD.n1396 VDD.n1393 0.60463
R18179 VDD.n1401 VDD.n1398 0.60463
R18180 VDD.n1407 VDD.n1405 0.60463
R18181 VDD.n151 VDD.n148 0.60463
R18182 VDD.n157 VDD.n154 0.60463
R18183 VDD.n162 VDD.n159 0.60463
R18184 VDD.n168 VDD.n165 0.60463
R18185 VDD.n173 VDD.n170 0.60463
R18186 VDD.n179 VDD.n177 0.60463
R18187 VDD.n9448 VDD.n9352 0.604026
R18188 VDD.n10921 VDD.n9343 0.603703
R18189 VDD.t28 VDD.n6897 0.600058
R18190 VDD.n9957 VDD 0.592891
R18191 VDD.n9343 VDD.n9341 0.576974
R18192 VDD.n8122 VDD.n8120 0.570797
R18193 VDD.n8561 VDD.n8560 0.570797
R18194 VDD.n10644 VDD.n9988 0.568833
R18195 VDD.n4113 VDD 0.568068
R18196 VDD.n4113 VDD 0.568068
R18197 VDD.n12778 VDD.n12777 0.55916
R18198 VDD.n10276 VDD.n10240 0.557022
R18199 VDD.n10325 VDD.n10216 0.557022
R18200 VDD.n10375 VDD.n10374 0.557022
R18201 VDD.n12417 VDD.n6927 0.557022
R18202 VDD.n8601 VDD.n7722 0.542299
R18203 VDD.n8689 VDD.n8683 0.542299
R18204 VDD.n11313 VDD.n11088 0.542299
R18205 VDD.n11210 VDD.n11204 0.542299
R18206 VDD.n6564 VDD 0.54194
R18207 VDD.n7958 VDD.n7957 0.539447
R18208 VDD.n7948 VDD.n7834 0.539447
R18209 VDD.n7907 VDD.n7858 0.539447
R18210 VDD.n7898 VDD.n7897 0.539447
R18211 VDD.n11471 VDD.n11469 0.539447
R18212 VDD.n11483 VDD.n11482 0.539447
R18213 VDD.n11528 VDD.n7675 0.539447
R18214 VDD.n11540 VDD.n11538 0.539447
R18215 VDD.n11583 VDD.n11581 0.539447
R18216 VDD.n12484 VDD.n12483 0.533379
R18217 VDD.n6566 VDD 0.531324
R18218 VDD.n2473 VDD 0.530391
R18219 VDD.n833 VDD 0.530391
R18220 VDD.n11218 VDD.n6580 0.529527
R18221 VDD.n12771 VDD.n12770 0.522949
R18222 VDD.n6557 VDD.n5778 0.515073
R18223 VDD.n5703 VDD.n4924 0.515073
R18224 VDD.n4917 VDD.n4138 0.515073
R18225 VDD.n4063 VDD.n3284 0.515073
R18226 VDD.n3277 VDD.n2498 0.515073
R18227 VDD.n2422 VDD.n1643 0.515073
R18228 VDD.n1226 VDD.n1026 0.515073
R18229 VDD.n780 VDD.n580 0.515073
R18230 VDD.n12406 VDD.n6935 0.506715
R18231 VDD.n12356 VDD.n12355 0.506715
R18232 VDD.n12307 VDD.n7015 0.506715
R18233 VDD.n12262 VDD.n7057 0.506715
R18234 VDD.n7170 VDD.n7112 0.506715
R18235 VDD.n7227 VDD.n7226 0.506715
R18236 VDD.n12229 VDD.n7270 0.506715
R18237 VDD.n12179 VDD.n12178 0.506715
R18238 VDD.n12130 VDD.n7348 0.506715
R18239 VDD.n8541 VDD.n8539 0.502461
R18240 VDD.n2472 VDD 0.497949
R18241 VDD.n832 VDD 0.497949
R18242 VDD.n9187 VDD.n9163 0.491125
R18243 VDD.n6562 VDD.n5707 0.489126
R18244 VDD.n6564 VDD.n4067 0.489126
R18245 VDD.n11011 VDD.n11010 0.488891
R18246 VDD.n6565 VDD.n2426 0.488186
R18247 VDD.n6566 VDD.n785 0.488186
R18248 VDD.n9163 VDD.n8738 0.488
R18249 VDD.n8549 VDD.n7776 0.484824
R18250 VDD.n9041 VDD.n8788 0.48381
R18251 VDD.n9263 VDD.n9262 0.483797
R18252 VDD.n9957 VDD.n9910 0.477082
R18253 VDD.n10101 VDD.n10086 0.476817
R18254 VDD.n8194 VDD.n8104 0.474574
R18255 VDD.n8108 VDD.n8105 0.474574
R18256 VDD.n8189 VDD.n8110 0.474574
R18257 VDD.n8185 VDD.n8184 0.474574
R18258 VDD.n8131 VDD.n8128 0.474574
R18259 VDD.n8178 VDD.n8133 0.474574
R18260 VDD.n8175 VDD.n8174 0.474574
R18261 VDD.n8140 VDD.n8137 0.474574
R18262 VDD.n8168 VDD.n8142 0.474574
R18263 VDD.n8164 VDD.n8163 0.474574
R18264 VDD.n8148 VDD.n8146 0.474574
R18265 VDD.n8156 VDD.n8151 0.474574
R18266 VDD.n8600 VDD.n7745 0.474574
R18267 VDD.n8602 VDD.n8601 0.474574
R18268 VDD.n11445 VDD.n11444 0.474574
R18269 VDD.n7727 VDD.n7726 0.474574
R18270 VDD.n8611 VDD.n8610 0.474574
R18271 VDD.n11433 VDD.n7738 0.474574
R18272 VDD.n7742 VDD.n7739 0.474574
R18273 VDD.n11428 VDD.n7743 0.474574
R18274 VDD.n8622 VDD.n8621 0.474574
R18275 VDD.n8642 VDD.n8641 0.474574
R18276 VDD.n11414 VDD.n8632 0.474574
R18277 VDD.n8636 VDD.n8633 0.474574
R18278 VDD.n11409 VDD.n8637 0.474574
R18279 VDD.n8653 VDD.n8652 0.474574
R18280 VDD.n8677 VDD.n8676 0.474574
R18281 VDD.n11395 VDD.n8662 0.474574
R18282 VDD.n11388 VDD.n8667 0.474574
R18283 VDD.n8682 VDD.n8672 0.474574
R18284 VDD.n11384 VDD.n8683 0.474574
R18285 VDD.n8691 VDD.n8690 0.474574
R18286 VDD.n8714 VDD.n8713 0.474574
R18287 VDD.n11370 VDD.n8704 0.474574
R18288 VDD.n8708 VDD.n8705 0.474574
R18289 VDD.n11365 VDD.n8709 0.474574
R18290 VDD.n8726 VDD.n8725 0.474574
R18291 VDD.n11047 VDD.n11046 0.474574
R18292 VDD.n11351 VDD.n11037 0.474574
R18293 VDD.n11041 VDD.n11038 0.474574
R18294 VDD.n11346 VDD.n11042 0.474574
R18295 VDD.n11058 VDD.n11057 0.474574
R18296 VDD.n11094 VDD.n11093 0.474574
R18297 VDD.n11332 VDD.n11066 0.474574
R18298 VDD.n11070 VDD.n11067 0.474574
R18299 VDD.n11084 VDD.n11072 0.474574
R18300 VDD.n11317 VDD.n11085 0.474574
R18301 VDD.n11088 VDD.n11086 0.474574
R18302 VDD.n11312 VDD.n11089 0.474574
R18303 VDD.n11111 VDD.n11110 0.474574
R18304 VDD.n11131 VDD.n11130 0.474574
R18305 VDD.n11298 VDD.n11121 0.474574
R18306 VDD.n11125 VDD.n11122 0.474574
R18307 VDD.n11293 VDD.n11126 0.474574
R18308 VDD.n11141 VDD.n11140 0.474574
R18309 VDD.n11162 VDD.n11161 0.474574
R18310 VDD.n11279 VDD.n11152 0.474574
R18311 VDD.n11156 VDD.n11153 0.474574
R18312 VDD.n11274 VDD.n11157 0.474574
R18313 VDD.n11173 VDD.n11172 0.474574
R18314 VDD.n11198 VDD.n11197 0.474574
R18315 VDD.n11260 VDD.n11183 0.474574
R18316 VDD.n11253 VDD.n11188 0.474574
R18317 VDD.n11203 VDD.n11193 0.474574
R18318 VDD.n11249 VDD.n11204 0.474574
R18319 VDD.n11212 VDD.n11211 0.474574
R18320 VDD.n11223 VDD.n11222 0.474574
R18321 VDD.n11230 VDD.n11229 0.474574
R18322 VDD.n12708 VDD.n6603 0.474574
R18323 VDD.n10923 VDD.n10922 0.473002
R18324 VDD.n12688 VDD.n12687 0.471403
R18325 VDD.n10294 VDD.n10293 0.471403
R18326 VDD.n10343 VDD.n10205 0.471403
R18327 VDD.n10392 VDD.n10179 0.471403
R18328 VDD.n8803 VDD.n8794 0.469257
R18329 VDD.n8932 VDD.n8930 0.469245
R18330 VDD.n12496 VDD.n12495 0.466716
R18331 VDD.n12450 VDD.n12449 0.466716
R18332 VDD.n5752 VDD.n5709 0.465811
R18333 VDD.n4111 VDD.n4069 0.465811
R18334 VDD.n2474 VDD.n2428 0.465811
R18335 VDD.n834 VDD.n788 0.465811
R18336 VDD.n10489 VDD.n10487 0.461585
R18337 VDD.n12779 VDD.n6567 0.457934
R18338 VDD.n10445 VDD.n10438 0.452151
R18339 VDD.n12491 VDD.n12490 0.448742
R18340 VDD.n12458 VDD.n12457 0.448742
R18341 VDD.n9419 VDD.n9418 0.444775
R18342 VDD.n8079 VDD.n8078 0.444064
R18343 VDD.n8040 VDD.n8039 0.444064
R18344 VDD.n8301 VDD.n8021 0.444064
R18345 VDD.n8479 VDD.n8348 0.444064
R18346 VDD.n8375 VDD.n8368 0.444064
R18347 VDD.n8561 VDD.n7761 0.444064
R18348 VDD.n12408 VDD.n12407 0.431961
R18349 VDD.n8106 VDD.n8084 0.428211
R18350 VDD.n9952 VDD.n9950 0.424187
R18351 VDD.n11672 VDD.n7595 0.406849
R18352 VDD.n11685 VDD.n11684 0.406849
R18353 VDD.n11731 VDD.n7565 0.406849
R18354 VDD.n11744 VDD.n11742 0.406849
R18355 VDD.n11786 VDD.n7533 0.406849
R18356 VDD.n11799 VDD.n11798 0.406849
R18357 VDD.n11845 VDD.n7503 0.406849
R18358 VDD.n11858 VDD.n11856 0.406849
R18359 VDD.n11900 VDD.n7471 0.406849
R18360 VDD.n11913 VDD.n11912 0.406849
R18361 VDD.n11959 VDD.n7441 0.406849
R18362 VDD.n11972 VDD.n11970 0.406849
R18363 VDD.n12014 VDD.n7409 0.406849
R18364 VDD.n12027 VDD.n12026 0.406849
R18365 VDD.n12074 VDD.n12073 0.406849
R18366 VDD.n7376 VDD.n7374 0.406849
R18367 VDD.n11590 VDD.n7638 0.404711
R18368 VDD.n11633 VDD.n7613 0.404711
R18369 VDD.n9764 VDD.n9763 0.400769
R18370 VDD.n9531 VDD.n9523 0.400769
R18371 VDD.n9488 VDD.n9480 0.400769
R18372 VDD.n9785 VDD.n9784 0.400768
R18373 VDD.n9811 VDD.n9810 0.400768
R18374 VDD.n9857 VDD.n9856 0.400768
R18375 VDD.n10884 VDD.n10883 0.400768
R18376 VDD.n11435 VDD.n7736 0.39727
R18377 VDD.n9956 VDD.n9955 0.395485
R18378 VDD.n10281 VDD.n10279 0.385784
R18379 VDD.n10327 VDD.n10214 0.385784
R18380 VDD.n10379 VDD.n10187 0.385784
R18381 VDD.n8211 VDD.n8083 0.380698
R18382 VDD.n8080 VDD.n8079 0.380698
R18383 VDD.n8221 VDD.n8074 0.380698
R18384 VDD.n8222 VDD.n8072 0.380698
R18385 VDD.n8227 VDD.n8069 0.380698
R18386 VDD.n8067 VDD.n8063 0.380698
R18387 VDD.n8237 VDD.n8061 0.380698
R18388 VDD.n8243 VDD.n8242 0.380698
R18389 VDD.n8250 VDD.n8249 0.380698
R18390 VDD.n8255 VDD.n8055 0.380698
R18391 VDD.n8052 VDD.n8051 0.380698
R18392 VDD.n8265 VDD.n8046 0.380698
R18393 VDD.n8266 VDD.n8044 0.380698
R18394 VDD.n8271 VDD.n8041 0.380698
R18395 VDD.n8039 VDD.n8034 0.380698
R18396 VDD.n8281 VDD.n8035 0.380698
R18397 VDD.n8296 VDD.n8023 0.380698
R18398 VDD.n8297 VDD.n8021 0.380698
R18399 VDD.n8302 VDD.n8018 0.380698
R18400 VDD.n8016 VDD.n8012 0.380698
R18401 VDD.n8312 VDD.n8010 0.380698
R18402 VDD.n8318 VDD.n8317 0.380698
R18403 VDD.n8325 VDD.n8324 0.380698
R18404 VDD.n8330 VDD.n8004 0.380698
R18405 VDD.n8001 VDD.n8000 0.380698
R18406 VDD.n8495 VDD.n7992 0.380698
R18407 VDD.n7996 VDD.n7993 0.380698
R18408 VDD.n8490 VDD.n7997 0.380698
R18409 VDD.n8344 VDD.n8343 0.380698
R18410 VDD.n8481 VDD.n8480 0.380698
R18411 VDD.n8351 VDD.n8348 0.380698
R18412 VDD.n8475 VDD.n8352 0.380698
R18413 VDD.n8367 VDD.n8366 0.380698
R18414 VDD.n8461 VDD.n8368 0.380698
R18415 VDD.n8377 VDD.n8376 0.380698
R18416 VDD.n8452 VDD.n8451 0.380698
R18417 VDD.n8384 VDD.n8381 0.380698
R18418 VDD.n8446 VDD.n8385 0.380698
R18419 VDD.n8394 VDD.n8393 0.380698
R18420 VDD.n8437 VDD.n8436 0.380698
R18421 VDD.n8401 VDD.n8398 0.380698
R18422 VDD.n8431 VDD.n8402 0.380698
R18423 VDD.n8411 VDD.n8410 0.380698
R18424 VDD.n8422 VDD.n8421 0.380698
R18425 VDD.n8417 VDD.n8416 0.380698
R18426 VDD.n8565 VDD.n7763 0.380698
R18427 VDD.n12415 VDD.n6929 0.378512
R18428 VDD.n10077 VDD.n10023 0.376971
R18429 VDD.n10074 VDD.n10026 0.376971
R18430 VDD.n10065 VDD.n10027 0.376971
R18431 VDD.n10057 VDD.n10056 0.376971
R18432 VDD.n10048 VDD.n10047 0.376971
R18433 VDD.n10047 VDD.n10039 0.376971
R18434 VDD.n10111 VDD.n10091 0.376971
R18435 VDD.n10637 VDD.n10141 0.376971
R18436 VDD.n10634 VDD.n10145 0.376971
R18437 VDD.n10627 VDD.n10626 0.376971
R18438 VDD.n10616 VDD.n10615 0.376971
R18439 VDD.n10607 VDD.n10606 0.376971
R18440 VDD.n10606 VDD.n10598 0.376971
R18441 VDD.n10527 VDD.n10524 0.376971
R18442 VDD.n10523 VDD.n10522 0.376971
R18443 VDD.n10566 VDD.n10565 0.376971
R18444 VDD.n10533 VDD.n10505 0.376971
R18445 VDD.n10545 VDD.n10539 0.376971
R18446 VDD.n10545 VDD.n10544 0.376971
R18447 VDD.n9566 VDD.n9563 0.376971
R18448 VDD.n9633 VDD.n9563 0.376971
R18449 VDD.n9697 VDD.n9696 0.376971
R18450 VDD.n9701 VDD.n9700 0.376971
R18451 VDD.n10851 VDD.n10850 0.376971
R18452 VDD.n10847 VDD.n10846 0.376971
R18453 VDD.n10735 VDD.n10728 0.376971
R18454 VDD.n10735 VDD.n10729 0.376971
R18455 VDD.n8913 VDD.n8912 0.376971
R18456 VDD.n8912 VDD.n8889 0.376971
R18457 VDD.n8908 VDD.n8907 0.376971
R18458 VDD.n8763 VDD.n8760 0.376971
R18459 VDD.n9373 VDD.n9365 0.376971
R18460 VDD.n9373 VDD.n9366 0.376971
R18461 VDD.n9378 VDD.n9377 0.376971
R18462 VDD.n9388 VDD.n9387 0.376971
R18463 VDD.n9439 VDD.n9360 0.376971
R18464 VDD.n8524 VDD.n7794 0.376971
R18465 VDD.n8515 VDD.n8514 0.376971
R18466 VDD.n12477 VDD.n12476 0.376971
R18467 VDD.n12471 VDD.n12470 0.376971
R18468 VDD.n9953 VDD 0.368743
R18469 VDD.n9956 VDD 0.368743
R18470 VDD.n12366 VDD.n6972 0.362082
R18471 VDD.n7013 VDD.n7009 0.362082
R18472 VDD.n12267 VDD.n7052 0.362082
R18473 VDD.n7160 VDD.n7158 0.362082
R18474 VDD.n7216 VDD.n7092 0.362082
R18475 VDD.n12234 VDD.n7265 0.362082
R18476 VDD.n12189 VDD.n7305 0.362082
R18477 VDD.n7346 VDD.n7342 0.362082
R18478 VDD.n12781 VDD.n6566 0.361524
R18479 VDD.n9150 VDD.n9089 0.357498
R18480 VDD.n7772 VDD.n7770 0.346446
R18481 VDD.n9954 VDD.n9949 0.344641
R18482 VDD.n6263 VDD.n6262 0.343549
R18483 VDD.n6268 VDD.n6052 0.343549
R18484 VDD.n6269 VDD.n6050 0.343549
R18485 VDD.n6276 VDD.n6274 0.343549
R18486 VDD.n6275 VDD.n6047 0.343549
R18487 VDD.n6287 VDD.n6286 0.343549
R18488 VDD.n5409 VDD.n5408 0.343549
R18489 VDD.n5414 VDD.n5198 0.343549
R18490 VDD.n5415 VDD.n5196 0.343549
R18491 VDD.n5422 VDD.n5420 0.343549
R18492 VDD.n5421 VDD.n5193 0.343549
R18493 VDD.n5433 VDD.n5432 0.343549
R18494 VDD.n4623 VDD.n4622 0.343549
R18495 VDD.n4628 VDD.n4412 0.343549
R18496 VDD.n4629 VDD.n4410 0.343549
R18497 VDD.n4636 VDD.n4634 0.343549
R18498 VDD.n4635 VDD.n4407 0.343549
R18499 VDD.n4647 VDD.n4646 0.343549
R18500 VDD.n3769 VDD.n3768 0.343549
R18501 VDD.n3774 VDD.n3558 0.343549
R18502 VDD.n3775 VDD.n3556 0.343549
R18503 VDD.n3782 VDD.n3780 0.343549
R18504 VDD.n3781 VDD.n3553 0.343549
R18505 VDD.n3793 VDD.n3792 0.343549
R18506 VDD.n2983 VDD.n2982 0.343549
R18507 VDD.n2988 VDD.n2772 0.343549
R18508 VDD.n2989 VDD.n2770 0.343549
R18509 VDD.n2996 VDD.n2994 0.343549
R18510 VDD.n2995 VDD.n2767 0.343549
R18511 VDD.n3007 VDD.n3006 0.343549
R18512 VDD.n2128 VDD.n2127 0.343549
R18513 VDD.n2133 VDD.n1917 0.343549
R18514 VDD.n2134 VDD.n1915 0.343549
R18515 VDD.n2141 VDD.n2139 0.343549
R18516 VDD.n2140 VDD.n1912 0.343549
R18517 VDD.n2152 VDD.n2151 0.343549
R18518 VDD.n991 VDD.n989 0.343549
R18519 VDD.n996 VDD.n993 0.343549
R18520 VDD.n1001 VDD.n999 0.343549
R18521 VDD.n1007 VDD.n1004 0.343549
R18522 VDD.n1013 VDD.n1011 0.343549
R18523 VDD.n1020 VDD.n1015 0.343549
R18524 VDD.n545 VDD.n543 0.343549
R18525 VDD.n550 VDD.n547 0.343549
R18526 VDD.n555 VDD.n553 0.343549
R18527 VDD.n561 VDD.n558 0.343549
R18528 VDD.n567 VDD.n565 0.343549
R18529 VDD.n574 VDD.n569 0.343549
R18530 VDD.n9289 VDD.n9288 0.34084
R18531 VDD.n8164 VDD.n8145 0.339124
R18532 VDD.n8676 VDD.n8674 0.339124
R18533 VDD.n11092 VDD.n11066 0.339124
R18534 VDD.n11197 VDD.n11195 0.339124
R18535 VDD.n11647 VDD.n11646 0.337342
R18536 VDD.n12782 VDD 0.336214
R18537 VDD.n9221 VDD.n9199 0.33059
R18538 VDD.n10978 VDD.n9205 0.33059
R18539 VDD.n10959 VDD.n7070 0.33059
R18540 VDD.n2470 VDD 0.329892
R18541 VDD.n830 VDD 0.329892
R18542 VDD.n9057 VDD.n9056 0.324719
R18543 VDD.n9054 VDD.n9053 0.324719
R18544 VDD.n8812 VDD.n8779 0.324719
R18545 VDD.n9588 VDD.n9587 0.324719
R18546 VDD.n9750 VDD.n9749 0.324719
R18547 VDD.n10895 VDD.n10674 0.324719
R18548 VDD.n10770 VDD.n10769 0.324719
R18549 VDD.n8089 VDD.n8085 0.317332
R18550 VDD.n8207 VDD.n8205 0.317332
R18551 VDD.n8286 VDD.n8285 0.317332
R18552 VDD.n8029 VDD.n8028 0.317332
R18553 VDD.n8361 VDD.n8360 0.317332
R18554 VDD.n8466 VDD.n8465 0.317332
R18555 VDD.n7789 VDD.n7779 0.313753
R18556 VDD.n11634 VDD.n7608 0.309235
R18557 VDD.n12703 VDD.n12702 0.30922
R18558 VDD.n10193 VDD.t152 0.300279
R18559 VDD.n10494 VDD.n6913 0.300279
R18560 VDD.n12421 VDD.n6920 0.300279
R18561 VDD.n10479 VDD.n10162 0.300279
R18562 VDD.n6706 VDD.n6705 0.300166
R18563 VDD.n10290 VDD.n10234 0.300166
R18564 VDD.n10342 VDD.n10207 0.300166
R18565 VDD.n10389 VDD.n10388 0.300166
R18566 VDD.n2474 VDD 0.299413
R18567 VDD.n834 VDD 0.299413
R18568 VDD.n9823 VDD.n9822 0.278729
R18569 VDD.n9776 VDD.n9775 0.278729
R18570 VDD.n9751 VDD.n9548 0.278729
R18571 VDD.n9797 VDD.n9504 0.278729
R18572 VDD.n10772 VDD.n10692 0.278729
R18573 VDD.n9779 VDD.n9518 0.278729
R18574 VDD.n9730 VDD.n9552 0.278729
R18575 VDD.n12429 VDD.n12427 0.27492
R18576 VDD.n8158 VDD.n8157 0.271399
R18577 VDD.n8603 VDD.n8600 0.271399
R18578 VDD.n8666 VDD.n8663 0.271399
R18579 VDD.n11385 VDD.n8682 0.271399
R18580 VDD.n11328 VDD.n11327 0.271399
R18581 VDD.n11317 VDD.n11316 0.271399
R18582 VDD.n11187 VDD.n11184 0.271399
R18583 VDD.n11250 VDD.n11203 0.271399
R18584 VDD.n7953 VDD.n7827 0.269974
R18585 VDD.n7949 VDD.n7832 0.269974
R18586 VDD.n7906 VDD.n7862 0.269974
R18587 VDD.n7902 VDD.n7867 0.269974
R18588 VDD.n11470 VDD.n7703 0.269974
R18589 VDD.n11477 VDD.n7700 0.269974
R18590 VDD.n11529 VDD.n7672 0.269974
R18591 VDD.n7673 VDD.n7668 0.269974
R18592 VDD.n9319 VDD.n9318 0.26925
R18593 VDD.n8685 VDD.t67 0.265013
R18594 VDD.n11105 VDD.t55 0.265013
R18595 VDD.n9969 VDD.n9906 0.26137
R18596 VDD.n9911 VDD.n9906 0.26137
R18597 VDD.n9958 VDD.n9911 0.26137
R18598 VDD.n5758 VDD.n5746 0.26137
R18599 VDD.n5758 VDD.n5757 0.26137
R18600 VDD.n5757 VDD.n5756 0.26137
R18601 VDD.n4118 VDD.n4106 0.26137
R18602 VDD.n4118 VDD.n4117 0.26137
R18603 VDD.n4117 VDD.n4116 0.26137
R18604 VDD.n2478 VDD.n2465 0.26137
R18605 VDD.n2478 VDD.n2477 0.26137
R18606 VDD.n2477 VDD.n2476 0.26137
R18607 VDD.n838 VDD.n825 0.26137
R18608 VDD.n838 VDD.n837 0.26137
R18609 VDD.n837 VDD.n836 0.26137
R18610 VDD.n9971 VDD 0.260619
R18611 VDD.n9981 VDD.n9972 0.25512
R18612 VDD VDD.n6565 0.25301
R18613 VDD.n5161 VDD.n4923 0.247601
R18614 VDD.n3521 VDD.n3283 0.247601
R18615 VDD.n1880 VDD.n1642 0.247601
R18616 VDD.n410 VDD.n409 0.247601
R18617 VDD.n6015 VDD.n5772 0.242094
R18618 VDD.n4375 VDD.n4132 0.242094
R18619 VDD.n2735 VDD.n2492 0.242094
R18620 VDD.n1638 VDD.n1637 0.242094
R18621 VDD.n12077 VDD.n7350 0.236946
R18622 VDD.n6563 VDD.n6562 0.23456
R18623 VDD.n5763 VDD.n5740 0.231925
R18624 VDD.n4123 VDD.n4100 0.231925
R18625 VDD.n2483 VDD.n2459 0.231925
R18626 VDD.n843 VDD.n819 0.231925
R18627 VDD.n9964 VDD.n9963 0.231891
R18628 VDD.n9963 VDD.n9907 0.231891
R18629 VDD.n9963 VDD.n9962 0.231891
R18630 VDD.n9941 VDD.n9916 0.231891
R18631 VDD.n9942 VDD.n9941 0.231891
R18632 VDD.n9941 VDD.n9940 0.231891
R18633 VDD.n9941 VDD.n9918 0.231891
R18634 VDD.n5763 VDD.n5762 0.231891
R18635 VDD.n5763 VDD.n5741 0.231891
R18636 VDD.n4123 VDD.n4122 0.231891
R18637 VDD.n4123 VDD.n4101 0.231891
R18638 VDD.n2483 VDD.n2482 0.231891
R18639 VDD.n2483 VDD.n2460 0.231891
R18640 VDD.n843 VDD.n842 0.231891
R18641 VDD.n843 VDD.n820 0.231891
R18642 VDD.n12782 VDD.n12781 0.230181
R18643 VDD.n9674 VDD.n9658 0.229427
R18644 VDD.n9674 VDD.n9673 0.229427
R18645 VDD.n10817 VDD.n10801 0.229427
R18646 VDD.n10817 VDD.n10816 0.229427
R18647 VDD.n8953 VDD.n8877 0.229427
R18648 VDD.n8955 VDD.n8953 0.229427
R18649 VDD.n8976 VDD.n8975 0.229427
R18650 VDD.n8978 VDD.n8976 0.229427
R18651 VDD.n9013 VDD.n8997 0.229427
R18652 VDD.n9013 VDD.n9012 0.229427
R18653 VDD.n6979 VDD.n6975 0.217449
R18654 VDD.n12311 VDD.n12310 0.217449
R18655 VDD.n12263 VDD.n7056 0.217449
R18656 VDD.n7167 VDD.n7166 0.217449
R18657 VDD.n7221 VDD.n7090 0.217449
R18658 VDD.n12230 VDD.n7269 0.217449
R18659 VDD.n7312 VDD.n7308 0.217449
R18660 VDD.n12134 VDD.n12133 0.217449
R18661 VDD.n12701 VDD.n12699 0.216346
R18662 VDD.n9675 VDD.n9674 0.215848
R18663 VDD.n10818 VDD.n10817 0.215848
R18664 VDD.n8976 VDD.n8855 0.215848
R18665 VDD.n9014 VDD.n9013 0.215848
R18666 VDD.n8953 VDD.n8952 0.215848
R18667 VDD.n6011 VDD 0.215174
R18668 VDD.n5157 VDD 0.215174
R18669 VDD.n4371 VDD 0.215174
R18670 VDD.n3517 VDD 0.215174
R18671 VDD.n2731 VDD 0.215174
R18672 VDD.n1876 VDD 0.215174
R18673 VDD.n1230 VDD 0.215174
R18674 VDD.n2 VDD 0.215174
R18675 VDD.n10280 VDD.n10238 0.214547
R18676 VDD.n10332 VDD.n10330 0.214547
R18677 VDD.n10380 VDD.n10185 0.214547
R18678 VDD.n7984 VDD.n7983 0.214355
R18679 VDD.n12701 VDD.n12700 0.211367
R18680 VDD.n9174 VDD.n7736 0.211364
R18681 VDD.n10996 VDD.n8727 0.211364
R18682 VDD.n10119 VDD.n10118 0.210656
R18683 VDD.n9595 VDD.n9589 0.210461
R18684 VDD.n10766 VDD.n10699 0.210461
R18685 VDD.n8553 VDD.n8552 0.208068
R18686 VDD.n10453 VDD.n6568 0.204334
R18687 VDD.n8158 VDD.n8149 0.203675
R18688 VDD.n11394 VDD.n8663 0.203675
R18689 VDD.n11328 VDD.n11071 0.203675
R18690 VDD.n11259 VDD.n11184 0.203675
R18691 VDD.n9825 VDD.n9824 0.202844
R18692 VDD.n6557 VDD.n6556 0.193465
R18693 VDD.n5703 VDD.n5702 0.193465
R18694 VDD.n4917 VDD.n4916 0.193465
R18695 VDD.n4063 VDD.n4062 0.193465
R18696 VDD.n3277 VDD.n3276 0.193465
R18697 VDD.n2422 VDD.n2421 0.193465
R18698 VDD.n1226 VDD.n1225 0.193465
R18699 VDD.n780 VDD.n779 0.193465
R18700 VDD.n9699 VDD.n9698 0.190717
R18701 VDD.n10849 VDD.n10848 0.190717
R18702 VDD.n8969 VDD.n8859 0.190717
R18703 VDD.n8970 VDD.n8969 0.190717
R18704 VDD.n8991 VDD.n8831 0.190717
R18705 VDD.n8992 VDD.n8991 0.190717
R18706 VDD.n8211 VDD.n8210 0.190599
R18707 VDD.n8282 VDD.n8281 0.190599
R18708 VDD.n8298 VDD.n8296 0.190599
R18709 VDD.n8476 VDD.n8475 0.190599
R18710 VDD.n8462 VDD.n8367 0.190599
R18711 VDD.n9131 VDD.n9090 0.189124
R18712 VDD.n10492 VDD.n10437 0.186007
R18713 VDD.n9149 VDD.n9092 0.178063
R18714 VDD.n5753 VDD 0.167831
R18715 VDD.n6012 VDD.n5935 0.167457
R18716 VDD.n5158 VDD.n5081 0.167457
R18717 VDD.n4372 VDD.n4295 0.167457
R18718 VDD.n3518 VDD.n3441 0.167457
R18719 VDD.n2732 VDD.n2655 0.167457
R18720 VDD.n1877 VDD.n1800 0.167457
R18721 VDD.n1609 VDD.n1605 0.167457
R18722 VDD.n381 VDD.n377 0.167457
R18723 VDD.n9151 VDD.n9088 0.166946
R18724 VDD.n9727 VDD.n9675 0.164777
R18725 VDD.n10819 VDD.n10818 0.164777
R18726 VDD.n8855 VDD.n8854 0.164777
R18727 VDD.n9015 VDD.n9014 0.164777
R18728 VDD.n8952 VDD.n8951 0.164777
R18729 VDD.n9420 VDD.n9419 0.164777
R18730 VDD.n9738 VDD.n9732 0.161367
R18731 VDD.n9724 VDD.n9636 0.161367
R18732 VDD.n9762 VDD.n9549 0.161367
R18733 VDD.n9774 VDD.n9773 0.161367
R18734 VDD.n9783 VDD.n9781 0.161367
R18735 VDD.n9809 VDD.n9505 0.161367
R18736 VDD.n9821 VDD.n9820 0.161367
R18737 VDD.n9855 VDD.n9852 0.161367
R18738 VDD.n10882 VDD.n10881 0.161367
R18739 VDD.n10877 VDD.n10693 0.161367
R18740 VDD.n10822 VDD.n10682 0.161367
R18741 VDD.n8948 VDD.n8880 0.161367
R18742 VDD.n8851 VDD.n8789 0.161367
R18743 VDD.n9018 VDD.n8796 0.161367
R18744 VDD.n9293 VDD.n9264 0.161367
R18745 VDD.n9658 VDD.n9644 0.15935
R18746 VDD.n9673 VDD.n9672 0.15935
R18747 VDD.n10801 VDD.n10787 0.15935
R18748 VDD.n10816 VDD.n10815 0.15935
R18749 VDD.n8877 VDD.n8863 0.15935
R18750 VDD.n8956 VDD.n8955 0.15935
R18751 VDD.n8975 VDD.n8856 0.15935
R18752 VDD.n8979 VDD.n8978 0.15935
R18753 VDD.n8997 VDD.n8828 0.15935
R18754 VDD.n9012 VDD.n9011 0.15935
R18755 VDD.n9288 VDD.n9274 0.15935
R18756 VDD.n9418 VDD.n9404 0.15935
R18757 VDD.n6609 VDD.n6608 0.157987
R18758 VDD.n9734 VDD.n9559 0.150167
R18759 VDD.n9720 VDD.n9637 0.150167
R18760 VDD.n9755 VDD.n9547 0.150167
R18761 VDD.n9530 VDD.n9529 0.150167
R18762 VDD.n9517 VDD.n9516 0.150167
R18763 VDD.n9800 VDD.n9503 0.150167
R18764 VDD.n9487 VDD.n9486 0.150167
R18765 VDD.n9864 VDD.n9863 0.150167
R18766 VDD.n10892 VDD.n10890 0.150167
R18767 VDD.n10871 VDD.n10691 0.150167
R18768 VDD.n10827 VDD.n10683 0.150167
R18769 VDD.n8943 VDD.n8882 0.150167
R18770 VDD.n8846 VDD.n8784 0.150167
R18771 VDD.n9023 VDD.n8798 0.150167
R18772 VDD.n9302 VDD.n9266 0.150167
R18773 VDD.n11580 VDD.n7640 0.145078
R18774 VDD.n12485 VDD.n6911 0.144522
R18775 VDD.n12445 VDD.n12444 0.144522
R18776 VDD.n10051 VDD.n10050 0.144522
R18777 VDD.n10610 VDD.n10609 0.144522
R18778 VDD.n10548 VDD.n10536 0.144522
R18779 VDD.n9619 VDD.n9618 0.144522
R18780 VDD.n9627 VDD.n9625 0.144522
R18781 VDD.n9689 VDD.n9688 0.144522
R18782 VDD.n9694 VDD.n9693 0.144522
R18783 VDD.n9704 VDD.n9703 0.144522
R18784 VDD.n9709 VDD.n9708 0.144522
R18785 VDD.n9714 VDD.n9713 0.144522
R18786 VDD.n9719 VDD.n9718 0.144522
R18787 VDD.n9725 VDD.n9723 0.144522
R18788 VDD.n10859 VDD.n10858 0.144522
R18789 VDD.n10854 VDD.n10853 0.144522
R18790 VDD.n10844 VDD.n10843 0.144522
R18791 VDD.n10839 VDD.n10838 0.144522
R18792 VDD.n10834 VDD.n10833 0.144522
R18793 VDD.n10829 VDD.n10828 0.144522
R18794 VDD.n10824 VDD.n10823 0.144522
R18795 VDD.n10743 VDD.n10716 0.144522
R18796 VDD.n10741 VDD.n10724 0.144522
R18797 VDD.n8845 VDD.n8844 0.144522
R18798 VDD.n8850 VDD.n8849 0.144522
R18799 VDD.n9025 VDD.n9024 0.144522
R18800 VDD.n9020 VDD.n9019 0.144522
R18801 VDD.n8942 VDD.n8941 0.144522
R18802 VDD.n8947 VDD.n8946 0.144522
R18803 VDD.n9300 VDD.n9299 0.144522
R18804 VDD.n9295 VDD.n9294 0.144522
R18805 VDD.n9435 VDD.n9395 0.144522
R18806 VDD.n9426 VDD.n9425 0.144522
R18807 VDD.n12779 VDD.n12778 0.142354
R18808 VDD.n9290 VDD.n9289 0.141804
R18809 VDD.n9742 VDD.n9740 0.138912
R18810 VDD.n9715 VDD.n9638 0.138912
R18811 VDD.n10776 VDD.n10681 0.138912
R18812 VDD.n10832 VDD.n10684 0.138912
R18813 VDD.n11680 VDD.n11679 0.13595
R18814 VDD.n7596 VDD.n7592 0.13595
R18815 VDD.n11736 VDD.n11734 0.13595
R18816 VDD.n11735 VDD.n7561 0.13595
R18817 VDD.n11794 VDD.n11793 0.13595
R18818 VDD.n7534 VDD.n7530 0.13595
R18819 VDD.n11850 VDD.n11848 0.13595
R18820 VDD.n11849 VDD.n7499 0.13595
R18821 VDD.n11908 VDD.n11907 0.13595
R18822 VDD.n7472 VDD.n7468 0.13595
R18823 VDD.n11964 VDD.n11962 0.13595
R18824 VDD.n11963 VDD.n7437 0.13595
R18825 VDD.n12022 VDD.n12021 0.13595
R18826 VDD.n7410 VDD.n7406 0.13595
R18827 VDD.n12081 VDD.n7379 0.13595
R18828 VDD.n12080 VDD.n12079 0.13595
R18829 VDD.n11582 VDD.n7641 0.135237
R18830 VDD.n11591 VDD.n11589 0.135237
R18831 VDD.n6013 VDD.n6011 0.134558
R18832 VDD.n5159 VDD.n5157 0.134558
R18833 VDD.n4373 VDD.n4371 0.134558
R18834 VDD.n3519 VDD.n3517 0.134558
R18835 VDD.n2733 VDD.n2731 0.134558
R18836 VDD.n1878 VDD.n1876 0.134558
R18837 VDD.n1610 VDD.n1230 0.134558
R18838 VDD.n382 VDD.n2 0.134558
R18839 VDD.n10996 VDD.n8721 0.132757
R18840 VDD.n6704 VDD.n6612 0.128928
R18841 VDD.n10289 VDD.n10236 0.128928
R18842 VDD.n10339 VDD.n10338 0.128928
R18843 VDD.n10385 VDD.n10181 0.128928
R18844 VDD.n9687 VDD.n9643 0.127599
R18845 VDD.n9710 VDD.n9639 0.127599
R18846 VDD.n10860 VDD.n10689 0.127599
R18847 VDD.n10837 VDD.n10685 0.127599
R18848 VDD.n10124 VDD.n6570 0.1274
R18849 VDD.n8521 VDD.n8520 0.12599
R18850 VDD.n7799 VDD.n7796 0.12599
R18851 VDD.n6570 VDD.n6568 0.122353
R18852 VDD.n12778 VDD.n6568 0.119879
R18853 VDD.n10659 VDD.n10658 0.117099
R18854 VDD.n9692 VDD.n9642 0.116231
R18855 VDD.n9705 VDD.n9640 0.116231
R18856 VDD.n10855 VDD.n10688 0.116231
R18857 VDD.n10842 VDD.n10686 0.116231
R18858 VDD VDD.n9904 0.116103
R18859 VDD VDD.n9905 0.116103
R18860 VDD.n9458 VDD.n9243 0.110519
R18861 VDD.n10953 VDD.n9225 0.110215
R18862 VDD.n9598 VDD.n8741 0.109875
R18863 VDD.n9066 VDD.n9065 0.109094
R18864 VDD.n8192 VDD.n8106 0.108934
R18865 VDD.n8192 VDD.n8191 0.108934
R18866 VDD.n8191 VDD.n8107 0.108934
R18867 VDD.n8181 VDD.n8107 0.108934
R18868 VDD.n8181 VDD.n8180 0.108934
R18869 VDD.n8180 VDD.n8129 0.108934
R18870 VDD.n8171 VDD.n8129 0.108934
R18871 VDD.n8171 VDD.n8170 0.108934
R18872 VDD.n8170 VDD.n8138 0.108934
R18873 VDD.n8160 VDD.n8138 0.108934
R18874 VDD.n8160 VDD.n8159 0.108934
R18875 VDD.n8159 VDD.n7744 0.108934
R18876 VDD.n8604 VDD.n7744 0.108934
R18877 VDD.n8605 VDD.n8604 0.108934
R18878 VDD.n8606 VDD.n8605 0.108934
R18879 VDD.n8607 VDD.n8606 0.108934
R18880 VDD.n8607 VDD.n7740 0.108934
R18881 VDD.n11431 VDD.n7740 0.108934
R18882 VDD.n11431 VDD.n11430 0.108934
R18883 VDD.n11430 VDD.n7741 0.108934
R18884 VDD.n8638 VDD.n7741 0.108934
R18885 VDD.n8638 VDD.n8634 0.108934
R18886 VDD.n11412 VDD.n8634 0.108934
R18887 VDD.n11412 VDD.n11411 0.108934
R18888 VDD.n11411 VDD.n8635 0.108934
R18889 VDD.n8673 VDD.n8635 0.108934
R18890 VDD.n8679 VDD.n8673 0.108934
R18891 VDD.n8680 VDD.n8679 0.108934
R18892 VDD.n11387 VDD.n8680 0.108934
R18893 VDD.n11387 VDD.n11386 0.108934
R18894 VDD.n11386 VDD.n8681 0.108934
R18895 VDD.n8710 VDD.n8681 0.108934
R18896 VDD.n8710 VDD.n8706 0.108934
R18897 VDD.n11368 VDD.n8706 0.108934
R18898 VDD.n11368 VDD.n11367 0.108934
R18899 VDD.n11367 VDD.n8707 0.108934
R18900 VDD.n11043 VDD.n8707 0.108934
R18901 VDD.n11043 VDD.n11039 0.108934
R18902 VDD.n11349 VDD.n11039 0.108934
R18903 VDD.n11349 VDD.n11348 0.108934
R18904 VDD.n11348 VDD.n11040 0.108934
R18905 VDD.n11090 VDD.n11040 0.108934
R18906 VDD.n11090 VDD.n11068 0.108934
R18907 VDD.n11330 VDD.n11068 0.108934
R18908 VDD.n11330 VDD.n11329 0.108934
R18909 VDD.n11329 VDD.n11069 0.108934
R18910 VDD.n11315 VDD.n11069 0.108934
R18911 VDD.n11315 VDD.n11314 0.108934
R18912 VDD.n11314 VDD.n11087 0.108934
R18913 VDD.n11127 VDD.n11087 0.108934
R18914 VDD.n11127 VDD.n11123 0.108934
R18915 VDD.n11296 VDD.n11123 0.108934
R18916 VDD.n11296 VDD.n11295 0.108934
R18917 VDD.n11295 VDD.n11124 0.108934
R18918 VDD.n11158 VDD.n11124 0.108934
R18919 VDD.n11158 VDD.n11154 0.108934
R18920 VDD.n11277 VDD.n11154 0.108934
R18921 VDD.n11277 VDD.n11276 0.108934
R18922 VDD.n11276 VDD.n11155 0.108934
R18923 VDD.n11194 VDD.n11155 0.108934
R18924 VDD.n11200 VDD.n11194 0.108934
R18925 VDD.n11201 VDD.n11200 0.108934
R18926 VDD.n11252 VDD.n11201 0.108934
R18927 VDD.n11252 VDD.n11251 0.108934
R18928 VDD.n11251 VDD.n11202 0.108934
R18929 VDD.n11225 VDD.n11202 0.108934
R18930 VDD.n11226 VDD.n11225 0.108934
R18931 VDD.n11226 VDD.n6605 0.108934
R18932 VDD.n12706 VDD.n6605 0.108934
R18933 VDD.n12706 VDD.n12705 0.108934
R18934 VDD.n12705 VDD.n6606 0.108934
R18935 VDD.n8208 VDD.n8084 0.108934
R18936 VDD.n8209 VDD.n8208 0.108934
R18937 VDD.n8209 VDD.n8073 0.108934
R18938 VDD.n8224 VDD.n8073 0.108934
R18939 VDD.n8225 VDD.n8224 0.108934
R18940 VDD.n8225 VDD.n8062 0.108934
R18941 VDD.n8239 VDD.n8062 0.108934
R18942 VDD.n8240 VDD.n8239 0.108934
R18943 VDD.n8240 VDD.n8056 0.108934
R18944 VDD.n8252 VDD.n8056 0.108934
R18945 VDD.n8253 VDD.n8252 0.108934
R18946 VDD.n8253 VDD.n8045 0.108934
R18947 VDD.n8268 VDD.n8045 0.108934
R18948 VDD.n8269 VDD.n8268 0.108934
R18949 VDD.n8269 VDD.n8033 0.108934
R18950 VDD.n8283 VDD.n8033 0.108934
R18951 VDD.n8284 VDD.n8283 0.108934
R18952 VDD.n8284 VDD.n8022 0.108934
R18953 VDD.n8299 VDD.n8022 0.108934
R18954 VDD.n8300 VDD.n8299 0.108934
R18955 VDD.n8300 VDD.n8011 0.108934
R18956 VDD.n8314 VDD.n8011 0.108934
R18957 VDD.n8315 VDD.n8314 0.108934
R18958 VDD.n8315 VDD.n8005 0.108934
R18959 VDD.n8327 VDD.n8005 0.108934
R18960 VDD.n8328 VDD.n8327 0.108934
R18961 VDD.n8328 VDD.n7994 0.108934
R18962 VDD.n8493 VDD.n7994 0.108934
R18963 VDD.n8493 VDD.n8492 0.108934
R18964 VDD.n8492 VDD.n7995 0.108934
R18965 VDD.n8349 VDD.n7995 0.108934
R18966 VDD.n8478 VDD.n8349 0.108934
R18967 VDD.n8478 VDD.n8477 0.108934
R18968 VDD.n8477 VDD.n8350 0.108934
R18969 VDD.n8464 VDD.n8350 0.108934
R18970 VDD.n8464 VDD.n8463 0.108934
R18971 VDD.n8463 VDD.n8365 0.108934
R18972 VDD.n8382 VDD.n8365 0.108934
R18973 VDD.n8449 VDD.n8382 0.108934
R18974 VDD.n8449 VDD.n8448 0.108934
R18975 VDD.n8448 VDD.n8383 0.108934
R18976 VDD.n8399 VDD.n8383 0.108934
R18977 VDD.n8434 VDD.n8399 0.108934
R18978 VDD.n8434 VDD.n8433 0.108934
R18979 VDD.n8433 VDD.n8400 0.108934
R18980 VDD.n8418 VDD.n8400 0.108934
R18981 VDD.n8419 VDD.n8418 0.108934
R18982 VDD.n8419 VDD.n7768 0.108934
R18983 VDD.n8563 VDD.n7768 0.108934
R18984 VDD.n8563 VDD.n8562 0.108934
R18985 VDD.n8562 VDD.n7769 0.108934
R18986 VDD.n7778 VDD.n7769 0.108934
R18987 VDD.n8551 VDD.n7778 0.108934
R18988 VDD.n8551 VDD.n8550 0.108934
R18989 VDD.n8550 VDD.n7779 0.108934
R18990 VDD.n8532 VDD.n7789 0.108934
R18991 VDD.n8532 VDD.n8531 0.108934
R18992 VDD.n8531 VDD.n7790 0.108934
R18993 VDD.n8523 VDD.n7790 0.108934
R18994 VDD.n8523 VDD.n8522 0.108934
R18995 VDD.n8522 VDD.n7795 0.108934
R18996 VDD.n8513 VDD.n7795 0.108934
R18997 VDD.n8513 VDD.n8512 0.108934
R18998 VDD.n8512 VDD.n7801 0.108934
R18999 VDD.n8505 VDD.n7801 0.108934
R19000 VDD.n8505 VDD.n8504 0.108934
R19001 VDD.n8504 VDD.n7806 0.108934
R19002 VDD.n7985 VDD.n7806 0.108934
R19003 VDD.n7985 VDD.n7984 0.108934
R19004 VDD.n7983 VDD.n7811 0.108934
R19005 VDD.n7978 VDD.n7811 0.108934
R19006 VDD.n7978 VDD.n7977 0.108934
R19007 VDD.n7977 VDD.n7813 0.108934
R19008 VDD.n7969 VDD.n7813 0.108934
R19009 VDD.n7969 VDD.n7968 0.108934
R19010 VDD.n7968 VDD.n7820 0.108934
R19011 VDD.n7960 VDD.n7820 0.108934
R19012 VDD.n7960 VDD.n7959 0.108934
R19013 VDD.n7959 VDD.n7826 0.108934
R19014 VDD.n7951 VDD.n7826 0.108934
R19015 VDD.n7951 VDD.n7950 0.108934
R19016 VDD.n7950 VDD.n7833 0.108934
R19017 VDD.n7942 VDD.n7833 0.108934
R19018 VDD.n7942 VDD.n7941 0.108934
R19019 VDD.n7941 VDD.n7838 0.108934
R19020 VDD.n7845 VDD.n7838 0.108934
R19021 VDD.n7932 VDD.n7845 0.108934
R19022 VDD.n7932 VDD.n7931 0.108934
R19023 VDD.n7931 VDD.n7846 0.108934
R19024 VDD.n7923 VDD.n7846 0.108934
R19025 VDD.n7923 VDD.n7922 0.108934
R19026 VDD.n7922 VDD.n7851 0.108934
R19027 VDD.n7914 VDD.n7851 0.108934
R19028 VDD.n7914 VDD.n7913 0.108934
R19029 VDD.n7913 VDD.n7857 0.108934
R19030 VDD.n7905 VDD.n7857 0.108934
R19031 VDD.n7905 VDD.n7904 0.108934
R19032 VDD.n7904 VDD.n7863 0.108934
R19033 VDD.n7896 VDD.n7863 0.108934
R19034 VDD.n7896 VDD.n7895 0.108934
R19035 VDD.n7895 VDD.n7870 0.108934
R19036 VDD.n7877 VDD.n7870 0.108934
R19037 VDD.n7886 VDD.n7877 0.108934
R19038 VDD.n7886 VDD.n7885 0.108934
R19039 VDD.n7885 VDD.n7878 0.108934
R19040 VDD.n7878 VDD.n7715 0.108934
R19041 VDD.n11455 VDD.n7715 0.108934
R19042 VDD.n11456 VDD.n11455 0.108934
R19043 VDD.n11457 VDD.n11456 0.108934
R19044 VDD.n11457 VDD.n7708 0.108934
R19045 VDD.n11467 VDD.n7708 0.108934
R19046 VDD.n11468 VDD.n11467 0.108934
R19047 VDD.n11468 VDD.n7702 0.108934
R19048 VDD.n11479 VDD.n7702 0.108934
R19049 VDD.n11480 VDD.n11479 0.108934
R19050 VDD.n11481 VDD.n11480 0.108934
R19051 VDD.n11481 VDD.n7695 0.108934
R19052 VDD.n11492 VDD.n7695 0.108934
R19053 VDD.n11493 VDD.n11492 0.108934
R19054 VDD.n11494 VDD.n11493 0.108934
R19055 VDD.n11494 VDD.n7688 0.108934
R19056 VDD.n11505 VDD.n7688 0.108934
R19057 VDD.n11506 VDD.n11505 0.108934
R19058 VDD.n11507 VDD.n11506 0.108934
R19059 VDD.n11507 VDD.n7681 0.108934
R19060 VDD.n11518 VDD.n7681 0.108934
R19061 VDD.n11519 VDD.n11518 0.108934
R19062 VDD.n11520 VDD.n11519 0.108934
R19063 VDD.n11520 VDD.n7674 0.108934
R19064 VDD.n11530 VDD.n7674 0.108934
R19065 VDD.n11531 VDD.n11530 0.108934
R19066 VDD.n11531 VDD.n7667 0.108934
R19067 VDD.n11541 VDD.n7667 0.108934
R19068 VDD.n11542 VDD.n11541 0.108934
R19069 VDD.n11543 VDD.n11542 0.108934
R19070 VDD.n11543 VDD.n7660 0.108934
R19071 VDD.n11554 VDD.n7660 0.108934
R19072 VDD.n11555 VDD.n11554 0.108934
R19073 VDD.n11556 VDD.n11555 0.108934
R19074 VDD.n11556 VDD.n7653 0.108934
R19075 VDD.n11567 VDD.n7653 0.108934
R19076 VDD.n11568 VDD.n11567 0.108934
R19077 VDD.n11569 VDD.n11568 0.108934
R19078 VDD.n11569 VDD.n7646 0.108934
R19079 VDD.n11579 VDD.n7646 0.108934
R19080 VDD.n11580 VDD.n11579 0.108934
R19081 VDD.n11592 VDD.n7640 0.108934
R19082 VDD.n11593 VDD.n11592 0.108934
R19083 VDD.n11594 VDD.n11593 0.108934
R19084 VDD.n11594 VDD.n7633 0.108934
R19085 VDD.n11605 VDD.n7633 0.108934
R19086 VDD.n11606 VDD.n11605 0.108934
R19087 VDD.n11607 VDD.n11606 0.108934
R19088 VDD.n11607 VDD.n7626 0.108934
R19089 VDD.n11618 VDD.n7626 0.108934
R19090 VDD.n11619 VDD.n11618 0.108934
R19091 VDD.n11620 VDD.n11619 0.108934
R19092 VDD.n11620 VDD.n7619 0.108934
R19093 VDD.n11631 VDD.n7619 0.108934
R19094 VDD.n11632 VDD.n11631 0.108934
R19095 VDD.n11635 VDD.n11632 0.108934
R19096 VDD.n11635 VDD.n11634 0.108934
R19097 VDD.n11657 VDD.n7608 0.108934
R19098 VDD.n11658 VDD.n11657 0.108934
R19099 VDD.n11659 VDD.n11658 0.108934
R19100 VDD.n11659 VDD.n7601 0.108934
R19101 VDD.n11669 VDD.n7601 0.108934
R19102 VDD.n11670 VDD.n11669 0.108934
R19103 VDD.n11670 VDD.n7594 0.108934
R19104 VDD.n11681 VDD.n7594 0.108934
R19105 VDD.n11682 VDD.n11681 0.108934
R19106 VDD.n11683 VDD.n11682 0.108934
R19107 VDD.n11683 VDD.n7587 0.108934
R19108 VDD.n11694 VDD.n7587 0.108934
R19109 VDD.n11695 VDD.n11694 0.108934
R19110 VDD.n11696 VDD.n11695 0.108934
R19111 VDD.n11696 VDD.n7580 0.108934
R19112 VDD.n11707 VDD.n7580 0.108934
R19113 VDD.n11708 VDD.n11707 0.108934
R19114 VDD.n11709 VDD.n11708 0.108934
R19115 VDD.n11709 VDD.n7573 0.108934
R19116 VDD.n11720 VDD.n7573 0.108934
R19117 VDD.n11721 VDD.n11720 0.108934
R19118 VDD.n11722 VDD.n11721 0.108934
R19119 VDD.n11722 VDD.n7566 0.108934
R19120 VDD.n11732 VDD.n7566 0.108934
R19121 VDD.n11733 VDD.n11732 0.108934
R19122 VDD.n11733 VDD.n7560 0.108934
R19123 VDD.n11745 VDD.n7560 0.108934
R19124 VDD.n11746 VDD.n11745 0.108934
R19125 VDD.n11747 VDD.n11746 0.108934
R19126 VDD.n11747 VDD.n7553 0.108934
R19127 VDD.n11758 VDD.n7553 0.108934
R19128 VDD.n11759 VDD.n11758 0.108934
R19129 VDD.n11760 VDD.n11759 0.108934
R19130 VDD.n11760 VDD.n7546 0.108934
R19131 VDD.n11771 VDD.n7546 0.108934
R19132 VDD.n11772 VDD.n11771 0.108934
R19133 VDD.n11773 VDD.n11772 0.108934
R19134 VDD.n11773 VDD.n7539 0.108934
R19135 VDD.n11783 VDD.n7539 0.108934
R19136 VDD.n11784 VDD.n11783 0.108934
R19137 VDD.n11784 VDD.n7532 0.108934
R19138 VDD.n11795 VDD.n7532 0.108934
R19139 VDD.n11796 VDD.n11795 0.108934
R19140 VDD.n11797 VDD.n11796 0.108934
R19141 VDD.n11797 VDD.n7525 0.108934
R19142 VDD.n11808 VDD.n7525 0.108934
R19143 VDD.n11809 VDD.n11808 0.108934
R19144 VDD.n11810 VDD.n11809 0.108934
R19145 VDD.n11810 VDD.n7518 0.108934
R19146 VDD.n11821 VDD.n7518 0.108934
R19147 VDD.n11822 VDD.n11821 0.108934
R19148 VDD.n11823 VDD.n11822 0.108934
R19149 VDD.n11823 VDD.n7511 0.108934
R19150 VDD.n11834 VDD.n7511 0.108934
R19151 VDD.n11835 VDD.n11834 0.108934
R19152 VDD.n11836 VDD.n11835 0.108934
R19153 VDD.n11836 VDD.n7504 0.108934
R19154 VDD.n11846 VDD.n7504 0.108934
R19155 VDD.n11847 VDD.n11846 0.108934
R19156 VDD.n11847 VDD.n7498 0.108934
R19157 VDD.n11859 VDD.n7498 0.108934
R19158 VDD.n11860 VDD.n11859 0.108934
R19159 VDD.n11861 VDD.n11860 0.108934
R19160 VDD.n11861 VDD.n7491 0.108934
R19161 VDD.n11872 VDD.n7491 0.108934
R19162 VDD.n11873 VDD.n11872 0.108934
R19163 VDD.n11874 VDD.n11873 0.108934
R19164 VDD.n11874 VDD.n7484 0.108934
R19165 VDD.n11885 VDD.n7484 0.108934
R19166 VDD.n11886 VDD.n11885 0.108934
R19167 VDD.n11887 VDD.n11886 0.108934
R19168 VDD.n11887 VDD.n7477 0.108934
R19169 VDD.n11897 VDD.n7477 0.108934
R19170 VDD.n11898 VDD.n11897 0.108934
R19171 VDD.n11898 VDD.n7470 0.108934
R19172 VDD.n11909 VDD.n7470 0.108934
R19173 VDD.n11910 VDD.n11909 0.108934
R19174 VDD.n11911 VDD.n11910 0.108934
R19175 VDD.n11911 VDD.n7463 0.108934
R19176 VDD.n11922 VDD.n7463 0.108934
R19177 VDD.n11923 VDD.n11922 0.108934
R19178 VDD.n11924 VDD.n11923 0.108934
R19179 VDD.n11924 VDD.n7456 0.108934
R19180 VDD.n11935 VDD.n7456 0.108934
R19181 VDD.n11936 VDD.n11935 0.108934
R19182 VDD.n11937 VDD.n11936 0.108934
R19183 VDD.n11937 VDD.n7449 0.108934
R19184 VDD.n11948 VDD.n7449 0.108934
R19185 VDD.n11949 VDD.n11948 0.108934
R19186 VDD.n11950 VDD.n11949 0.108934
R19187 VDD.n11950 VDD.n7442 0.108934
R19188 VDD.n11960 VDD.n7442 0.108934
R19189 VDD.n11961 VDD.n11960 0.108934
R19190 VDD.n11961 VDD.n7436 0.108934
R19191 VDD.n11973 VDD.n7436 0.108934
R19192 VDD.n11974 VDD.n11973 0.108934
R19193 VDD.n11975 VDD.n11974 0.108934
R19194 VDD.n11975 VDD.n7429 0.108934
R19195 VDD.n11986 VDD.n7429 0.108934
R19196 VDD.n11987 VDD.n11986 0.108934
R19197 VDD.n11988 VDD.n11987 0.108934
R19198 VDD.n11988 VDD.n7422 0.108934
R19199 VDD.n11999 VDD.n7422 0.108934
R19200 VDD.n12000 VDD.n11999 0.108934
R19201 VDD.n12001 VDD.n12000 0.108934
R19202 VDD.n12001 VDD.n7415 0.108934
R19203 VDD.n12011 VDD.n7415 0.108934
R19204 VDD.n12012 VDD.n12011 0.108934
R19205 VDD.n12012 VDD.n7408 0.108934
R19206 VDD.n12023 VDD.n7408 0.108934
R19207 VDD.n12024 VDD.n12023 0.108934
R19208 VDD.n12025 VDD.n12024 0.108934
R19209 VDD.n12025 VDD.n7401 0.108934
R19210 VDD.n12036 VDD.n7401 0.108934
R19211 VDD.n12037 VDD.n12036 0.108934
R19212 VDD.n12038 VDD.n12037 0.108934
R19213 VDD.n12038 VDD.n7394 0.108934
R19214 VDD.n12049 VDD.n7394 0.108934
R19215 VDD.n12050 VDD.n12049 0.108934
R19216 VDD.n12051 VDD.n12050 0.108934
R19217 VDD.n12051 VDD.n7387 0.108934
R19218 VDD.n12062 VDD.n7387 0.108934
R19219 VDD.n12063 VDD.n12062 0.108934
R19220 VDD.n12064 VDD.n12063 0.108934
R19221 VDD.n12064 VDD.n7380 0.108934
R19222 VDD.n12075 VDD.n7380 0.108934
R19223 VDD.n12076 VDD.n12075 0.108934
R19224 VDD.n12078 VDD.n12076 0.108934
R19225 VDD.n12078 VDD.n12077 0.108934
R19226 VDD.n6945 VDD.n6929 0.108934
R19227 VDD.n12398 VDD.n6945 0.108934
R19228 VDD.n12398 VDD.n12397 0.108934
R19229 VDD.n12397 VDD.n6946 0.108934
R19230 VDD.n6954 VDD.n6946 0.108934
R19231 VDD.n12387 VDD.n6954 0.108934
R19232 VDD.n12387 VDD.n12386 0.108934
R19233 VDD.n12386 VDD.n6955 0.108934
R19234 VDD.n6963 VDD.n6955 0.108934
R19235 VDD.n12376 VDD.n6963 0.108934
R19236 VDD.n12376 VDD.n12375 0.108934
R19237 VDD.n12375 VDD.n6964 0.108934
R19238 VDD.n6973 VDD.n6964 0.108934
R19239 VDD.n12365 VDD.n6973 0.108934
R19240 VDD.n12365 VDD.n12364 0.108934
R19241 VDD.n12364 VDD.n6974 0.108934
R19242 VDD.n12354 VDD.n6974 0.108934
R19243 VDD.n12354 VDD.n12353 0.108934
R19244 VDD.n12353 VDD.n6981 0.108934
R19245 VDD.n6989 VDD.n6981 0.108934
R19246 VDD.n12343 VDD.n6989 0.108934
R19247 VDD.n12343 VDD.n12342 0.108934
R19248 VDD.n12342 VDD.n6990 0.108934
R19249 VDD.n6998 VDD.n6990 0.108934
R19250 VDD.n12332 VDD.n6998 0.108934
R19251 VDD.n12332 VDD.n12331 0.108934
R19252 VDD.n12331 VDD.n6999 0.108934
R19253 VDD.n7007 VDD.n6999 0.108934
R19254 VDD.n12321 VDD.n7007 0.108934
R19255 VDD.n12321 VDD.n12320 0.108934
R19256 VDD.n12320 VDD.n7008 0.108934
R19257 VDD.n7016 VDD.n7008 0.108934
R19258 VDD.n12309 VDD.n7016 0.108934
R19259 VDD.n12309 VDD.n12308 0.108934
R19260 VDD.n12308 VDD.n7017 0.108934
R19261 VDD.n7027 VDD.n7017 0.108934
R19262 VDD.n12298 VDD.n7027 0.108934
R19263 VDD.n12298 VDD.n12297 0.108934
R19264 VDD.n12297 VDD.n7028 0.108934
R19265 VDD.n7036 VDD.n7028 0.108934
R19266 VDD.n12287 VDD.n7036 0.108934
R19267 VDD.n12287 VDD.n12286 0.108934
R19268 VDD.n12286 VDD.n7037 0.108934
R19269 VDD.n7045 VDD.n7037 0.108934
R19270 VDD.n12276 VDD.n7045 0.108934
R19271 VDD.n12276 VDD.n12275 0.108934
R19272 VDD.n12275 VDD.n7046 0.108934
R19273 VDD.n7054 VDD.n7046 0.108934
R19274 VDD.n12265 VDD.n7054 0.108934
R19275 VDD.n12265 VDD.n12264 0.108934
R19276 VDD.n12264 VDD.n7055 0.108934
R19277 VDD.n7066 VDD.n7055 0.108934
R19278 VDD.n12254 VDD.n7066 0.108934
R19279 VDD.n12254 VDD.n12253 0.108934
R19280 VDD.n12253 VDD.n7067 0.108934
R19281 VDD.n7129 VDD.n7067 0.108934
R19282 VDD.n7129 VDD.n7125 0.108934
R19283 VDD.n7137 VDD.n7125 0.108934
R19284 VDD.n7138 VDD.n7137 0.108934
R19285 VDD.n7138 VDD.n7121 0.108934
R19286 VDD.n7147 VDD.n7121 0.108934
R19287 VDD.n7148 VDD.n7147 0.108934
R19288 VDD.n7148 VDD.n7117 0.108934
R19289 VDD.n7156 VDD.n7117 0.108934
R19290 VDD.n7157 VDD.n7156 0.108934
R19291 VDD.n7157 VDD.n7113 0.108934
R19292 VDD.n7168 VDD.n7113 0.108934
R19293 VDD.n7169 VDD.n7168 0.108934
R19294 VDD.n7169 VDD.n7109 0.108934
R19295 VDD.n7178 VDD.n7109 0.108934
R19296 VDD.n7179 VDD.n7178 0.108934
R19297 VDD.n7179 VDD.n7105 0.108934
R19298 VDD.n7187 VDD.n7105 0.108934
R19299 VDD.n7188 VDD.n7187 0.108934
R19300 VDD.n7188 VDD.n7101 0.108934
R19301 VDD.n7197 VDD.n7101 0.108934
R19302 VDD.n7198 VDD.n7197 0.108934
R19303 VDD.n7198 VDD.n7097 0.108934
R19304 VDD.n7206 VDD.n7097 0.108934
R19305 VDD.n7207 VDD.n7206 0.108934
R19306 VDD.n7207 VDD.n7093 0.108934
R19307 VDD.n7217 VDD.n7093 0.108934
R19308 VDD.n7218 VDD.n7217 0.108934
R19309 VDD.n7218 VDD.n7089 0.108934
R19310 VDD.n7228 VDD.n7089 0.108934
R19311 VDD.n7229 VDD.n7228 0.108934
R19312 VDD.n7229 VDD.n7085 0.108934
R19313 VDD.n7237 VDD.n7085 0.108934
R19314 VDD.n7238 VDD.n7237 0.108934
R19315 VDD.n7238 VDD.n7081 0.108934
R19316 VDD.n7247 VDD.n7081 0.108934
R19317 VDD.n7248 VDD.n7247 0.108934
R19318 VDD.n7248 VDD.n7077 0.108934
R19319 VDD.n7257 VDD.n7077 0.108934
R19320 VDD.n7258 VDD.n7257 0.108934
R19321 VDD.n12243 VDD.n7258 0.108934
R19322 VDD.n12243 VDD.n12242 0.108934
R19323 VDD.n12242 VDD.n7259 0.108934
R19324 VDD.n7267 VDD.n7259 0.108934
R19325 VDD.n12232 VDD.n7267 0.108934
R19326 VDD.n12232 VDD.n12231 0.108934
R19327 VDD.n12231 VDD.n7268 0.108934
R19328 VDD.n7279 VDD.n7268 0.108934
R19329 VDD.n12221 VDD.n7279 0.108934
R19330 VDD.n12221 VDD.n12220 0.108934
R19331 VDD.n12220 VDD.n7280 0.108934
R19332 VDD.n7288 VDD.n7280 0.108934
R19333 VDD.n12210 VDD.n7288 0.108934
R19334 VDD.n12210 VDD.n12209 0.108934
R19335 VDD.n12209 VDD.n7289 0.108934
R19336 VDD.n7297 VDD.n7289 0.108934
R19337 VDD.n12199 VDD.n7297 0.108934
R19338 VDD.n12199 VDD.n12198 0.108934
R19339 VDD.n12198 VDD.n7298 0.108934
R19340 VDD.n7306 VDD.n7298 0.108934
R19341 VDD.n12188 VDD.n7306 0.108934
R19342 VDD.n12188 VDD.n12187 0.108934
R19343 VDD.n12187 VDD.n7307 0.108934
R19344 VDD.n12177 VDD.n7307 0.108934
R19345 VDD.n12177 VDD.n12176 0.108934
R19346 VDD.n12176 VDD.n7314 0.108934
R19347 VDD.n7322 VDD.n7314 0.108934
R19348 VDD.n12166 VDD.n7322 0.108934
R19349 VDD.n12166 VDD.n12165 0.108934
R19350 VDD.n12165 VDD.n7323 0.108934
R19351 VDD.n7331 VDD.n7323 0.108934
R19352 VDD.n12155 VDD.n7331 0.108934
R19353 VDD.n12155 VDD.n12154 0.108934
R19354 VDD.n12154 VDD.n7332 0.108934
R19355 VDD.n7340 VDD.n7332 0.108934
R19356 VDD.n12144 VDD.n7340 0.108934
R19357 VDD.n12144 VDD.n12143 0.108934
R19358 VDD.n12143 VDD.n7341 0.108934
R19359 VDD.n7349 VDD.n7341 0.108934
R19360 VDD.n12132 VDD.n7349 0.108934
R19361 VDD.n12132 VDD.n12131 0.108934
R19362 VDD.n12699 VDD.n6611 0.108934
R19363 VDD.n6708 VDD.n6611 0.108934
R19364 VDD.n12686 VDD.n6708 0.108934
R19365 VDD.n12686 VDD.n12685 0.108934
R19366 VDD.n12685 VDD.n6709 0.108934
R19367 VDD.n10254 VDD.n6709 0.108934
R19368 VDD.n10254 VDD.n10251 0.108934
R19369 VDD.n10261 VDD.n10251 0.108934
R19370 VDD.n10262 VDD.n10261 0.108934
R19371 VDD.n10262 VDD.n10247 0.108934
R19372 VDD.n10269 VDD.n10247 0.108934
R19373 VDD.n10270 VDD.n10269 0.108934
R19374 VDD.n10270 VDD.n10241 0.108934
R19375 VDD.n10277 VDD.n10241 0.108934
R19376 VDD.n10278 VDD.n10277 0.108934
R19377 VDD.n10278 VDD.n10237 0.108934
R19378 VDD.n10287 VDD.n10237 0.108934
R19379 VDD.n10288 VDD.n10287 0.108934
R19380 VDD.n10288 VDD.n10233 0.108934
R19381 VDD.n10295 VDD.n10233 0.108934
R19382 VDD.n10296 VDD.n10295 0.108934
R19383 VDD.n10296 VDD.n10229 0.108934
R19384 VDD.n10303 VDD.n10229 0.108934
R19385 VDD.n10304 VDD.n10303 0.108934
R19386 VDD.n10304 VDD.n10223 0.108934
R19387 VDD.n10311 VDD.n10223 0.108934
R19388 VDD.n10312 VDD.n10311 0.108934
R19389 VDD.n10312 VDD.n10219 0.108934
R19390 VDD.n10319 VDD.n10219 0.108934
R19391 VDD.n10320 VDD.n10319 0.108934
R19392 VDD.n10320 VDD.n10215 0.108934
R19393 VDD.n10328 VDD.n10215 0.108934
R19394 VDD.n10329 VDD.n10328 0.108934
R19395 VDD.n10329 VDD.n10208 0.108934
R19396 VDD.n10340 VDD.n10208 0.108934
R19397 VDD.n10341 VDD.n10340 0.108934
R19398 VDD.n10341 VDD.n10204 0.108934
R19399 VDD.n10348 VDD.n10204 0.108934
R19400 VDD.n10349 VDD.n10348 0.108934
R19401 VDD.n10349 VDD.n10200 0.108934
R19402 VDD.n10356 VDD.n10200 0.108934
R19403 VDD.n10357 VDD.n10356 0.108934
R19404 VDD.n10357 VDD.n10196 0.108934
R19405 VDD.n10364 VDD.n10196 0.108934
R19406 VDD.n10365 VDD.n10364 0.108934
R19407 VDD.n10365 VDD.n10190 0.108934
R19408 VDD.n10372 VDD.n10190 0.108934
R19409 VDD.n10373 VDD.n10372 0.108934
R19410 VDD.n10373 VDD.n10186 0.108934
R19411 VDD.n10381 VDD.n10186 0.108934
R19412 VDD.n10382 VDD.n10381 0.108934
R19413 VDD.n10382 VDD.n10180 0.108934
R19414 VDD.n10390 VDD.n10180 0.108934
R19415 VDD.n10391 VDD.n10390 0.108934
R19416 VDD.n10391 VDD.n10176 0.108934
R19417 VDD.n10398 VDD.n10176 0.108934
R19418 VDD.n10399 VDD.n10398 0.108934
R19419 VDD.n10399 VDD.n10172 0.108934
R19420 VDD.n10406 VDD.n10172 0.108934
R19421 VDD.n10407 VDD.n10406 0.108934
R19422 VDD.n10407 VDD.n10168 0.108934
R19423 VDD.n10414 VDD.n10168 0.108934
R19424 VDD.n10415 VDD.n10414 0.108934
R19425 VDD.n10415 VDD.n6928 0.108934
R19426 VDD.n12416 VDD.n6928 0.108934
R19427 VDD.n12416 VDD.n12415 0.108934
R19428 VDD.n10953 VDD.n10948 0.10877
R19429 VDD.n6544 VDD.n6543 0.107703
R19430 VDD.n5690 VDD.n5689 0.107703
R19431 VDD.n4904 VDD.n4903 0.107703
R19432 VDD.n4050 VDD.n4049 0.107703
R19433 VDD.n3264 VDD.n3263 0.107703
R19434 VDD.n2409 VDD.n2408 0.107703
R19435 VDD.n1197 VDD.n1189 0.107703
R19436 VDD.n751 VDD.n743 0.107703
R19437 VDD.n9612 VDD.n9611 0.0995999
R19438 VDD.n9684 VDD.n9554 0.0995999
R19439 VDD.n10864 VDD.n10863 0.0995999
R19440 VDD.n10753 VDD.n10752 0.0995999
R19441 VDD.n11023 VDD.n8737 0.0980399
R19442 VDD.n12469 VDD.n12434 0.0941356
R19443 VDD.n10431 VDD.n10425 0.0932536
R19444 VDD.n5751 VDD 0.0926053
R19445 VDD.n4112 VDD 0.0926053
R19446 VDD.n11021 VDD.n11020 0.0923441
R19447 VDD.n9186 VDD.n9078 0.0905941
R19448 VDD.n9186 VDD.n9165 0.0897616
R19449 VDD.n10569 VDD.n10568 0.0895625
R19450 VDD.n10968 VDD.n9212 0.0861908
R19451 VDD.n10955 VDD.n10945 0.0856562
R19452 VDD.n9134 VDD.n9108 0.0825312
R19453 VDD.n9124 VDD.n9123 0.0825312
R19454 VDD.n9946 VDD.n9914 0.0815811
R19455 VDD.n9935 VDD.n9934 0.0815811
R19456 VDD.n9925 VDD.n9914 0.0790473
R19457 VDD.n10968 VDD.n9216 0.0777426
R19458 VDD.n12780 VDD.n12779 0.0769364
R19459 VDD VDD.n9215 0.0739375
R19460 VDD.n9865 VDD.n9831 0.0736942
R19461 VDD.n9069 VDD.n8753 0.0736373
R19462 VDD.n12363 VDD.n12362 0.0728164
R19463 VDD.n12312 VDD.n7014 0.0728164
R19464 VDD.n12266 VDD.n7053 0.0728164
R19465 VDD.n7159 VDD.n7114 0.0728164
R19466 VDD.n7220 VDD.n7219 0.0728164
R19467 VDD.n12233 VDD.n7266 0.0728164
R19468 VDD.n12186 VDD.n12185 0.0728164
R19469 VDD.n12135 VDD.n7347 0.0728164
R19470 VDD.n11001 VDD.n8750 0.0717614
R19471 VDD.n12772 VDD.n12771 0.071743
R19472 VDD.n8750 VDD.n8747 0.0711193
R19473 VDD.n8824 VDD.n8800 0.0707228
R19474 VDD.n9058 VDD.n8766 0.0707228
R19475 VDD.n11001 VDD.n8753 0.0703248
R19476 VDD.n7777 VDD.n7775 0.0696892
R19477 VDD.n8895 VDD.n8894 0.0692474
R19478 VDD.n6016 VDD.n6015 0.0688877
R19479 VDD.n5162 VDD.n5161 0.0688877
R19480 VDD.n4376 VDD.n4375 0.0688877
R19481 VDD.n3522 VDD.n3521 0.0688877
R19482 VDD.n2736 VDD.n2735 0.0688877
R19483 VDD.n1881 VDD.n1880 0.0688877
R19484 VDD.n1637 VDD.n1636 0.0688877
R19485 VDD.n409 VDD.n408 0.0688877
R19486 VDD.n8161 VDD.n8146 0.0682249
R19487 VDD.n8678 VDD.n8662 0.0682249
R19488 VDD.n11331 VDD.n11067 0.0682249
R19489 VDD.n11199 VDD.n11183 0.0682249
R19490 VDD.n9370 VDD.n9350 0.0679494
R19491 VDD.n10499 VDD 0.0645625
R19492 VDD.n6016 VDD.n6013 0.0643587
R19493 VDD.n5162 VDD.n5159 0.0643587
R19494 VDD.n4376 VDD.n4373 0.0643587
R19495 VDD.n3522 VDD.n3519 0.0643587
R19496 VDD.n2736 VDD.n2733 0.0643587
R19497 VDD.n1881 VDD.n1878 0.0643587
R19498 VDD.n1636 VDD.n1610 0.0643587
R19499 VDD.n408 VDD.n382 0.0643587
R19500 VDD.n8090 VDD.n8089 0.0638663
R19501 VDD.n8207 VDD.n8206 0.0638663
R19502 VDD.n8285 VDD.n8032 0.0638663
R19503 VDD.n8028 VDD.n8027 0.0638663
R19504 VDD.n8360 VDD.n8359 0.0638663
R19505 VDD.n8465 VDD.n8364 0.0638663
R19506 VDD.n9216 VDD.n9214 0.0636644
R19507 VDD.n9760 VDD.n9759 0.0631347
R19508 VDD.n9807 VDD.n9806 0.0631347
R19509 VDD.n10703 VDD.n10700 0.0631347
R19510 VDD.n10875 VDD.n10695 0.0631347
R19511 VDD.n9514 VDD.n9509 0.0631347
R19512 VDD.n9590 VDD.n9577 0.0631347
R19513 VDD.n9736 VDD.n9556 0.0631347
R19514 VDD.n9771 VDD.n9525 0.0627929
R19515 VDD.n9818 VDD.n9482 0.0627929
R19516 VDD.n9924 VDD.n9922 0.0624727
R19517 VDD.n10082 VDD.n10012 0.0608156
R19518 VDD.n5752 VDD 0.060807
R19519 VDD VDD.n4111 0.060807
R19520 VDD.n9046 VDD.n9043 0.0604712
R19521 VDD.n8774 VDD.n8772 0.0604712
R19522 VDD.n9064 VDD.n8759 0.0604712
R19523 VDD.n9317 VDD.n9252 0.0604712
R19524 VDD.n10511 VDD.n10150 0.060461
R19525 VDD VDD.n5709 0.0603214
R19526 VDD VDD.n4069 0.0603214
R19527 VDD VDD.n2428 0.0603214
R19528 VDD VDD.n788 0.0603214
R19529 VDD.n9958 VDD.n9957 0.0602826
R19530 VDD.n8885 VDD.n8769 0.0595872
R19531 VDD.n10497 VDD.n10159 0.0592243
R19532 VDD.n10085 VDD.n10084 0.0591683
R19533 VDD.n9052 VDD.n8780 0.0591603
R19534 VDD.n9268 VDD.n9250 0.0591603
R19535 VDD.n9447 VDD.n9353 0.0586853
R19536 VDD.n9853 VDD.n9829 0.0581563
R19537 VDD.n12441 VDD.n6567 0.0575652
R19538 VDD.n5732 VDD.n5731 0.056838
R19539 VDD.n5733 VDD.n5732 0.056838
R19540 VDD.n5733 VDD.n5710 0.056838
R19541 VDD.n5769 VDD.n5710 0.056838
R19542 VDD.n4092 VDD.n4091 0.056838
R19543 VDD.n4093 VDD.n4092 0.056838
R19544 VDD.n4093 VDD.n4070 0.056838
R19545 VDD.n4129 VDD.n4070 0.056838
R19546 VDD.n2451 VDD.n2450 0.056838
R19547 VDD.n2452 VDD.n2451 0.056838
R19548 VDD.n2452 VDD.n2429 0.056838
R19549 VDD.n2489 VDD.n2429 0.056838
R19550 VDD.n811 VDD.n810 0.056838
R19551 VDD.n812 VDD.n811 0.056838
R19552 VDD.n812 VDD.n789 0.056838
R19553 VDD.n849 VDD.n789 0.056838
R19554 VDD VDD.n10498 0.05675
R19555 VDD.n10971 VDD.n9212 0.0566413
R19556 VDD.n9608 VDD.n9580 0.0565323
R19557 VDD.n9733 VDD.n9557 0.0565323
R19558 VDD.n9756 VDD.n9754 0.0565323
R19559 VDD.n9528 VDD.n9526 0.0565323
R19560 VDD.n9791 VDD.n9512 0.0565323
R19561 VDD.n9804 VDD.n9801 0.0565323
R19562 VDD.n9485 VDD.n9483 0.0565323
R19563 VDD.n10891 VDD.n10671 0.0565323
R19564 VDD.n10872 VDD.n10870 0.0565323
R19565 VDD.n10760 VDD.n10759 0.0565323
R19566 VDD.n9343 VDD.n9322 0.0561943
R19567 VDD.n9444 VDD.n9352 0.0558794
R19568 VDD.n10035 VDD.n10016 0.0547109
R19569 VDD.n10594 VDD.n10132 0.0547109
R19570 VDD.n10558 VDD.n10557 0.0547109
R19571 VDD.n9948 VDD.n9947 0.0531263
R19572 VDD.n11020 VDD.n8740 0.0521995
R19573 VDD.n9165 VDD.n9164 0.0521189
R19574 VDD.n12700 VDD.n6606 0.0517048
R19575 VDD.n9188 VDD.n9078 0.0513458
R19576 VDD.n9934 VDD.n9927 0.0498396
R19577 VDD.n9115 VDD.n9111 0.0493281
R19578 VDD.n9601 VDD.n9580 0.0487198
R19579 VDD.n9745 VDD.n9557 0.0487198
R19580 VDD.n9754 VDD.n9753 0.0487198
R19581 VDD.n9536 VDD.n9528 0.0487198
R19582 VDD.n9791 VDD.n9790 0.0487198
R19583 VDD.n9804 VDD.n9803 0.0487198
R19584 VDD.n9493 VDD.n9485 0.0487198
R19585 VDD.n10870 VDD.n10869 0.0487198
R19586 VDD.n10759 VDD.n10758 0.0487198
R19587 VDD.n9851 VDD.n9829 0.0479088
R19588 VDD.n10905 VDD.n10903 0.0472468
R19589 VDD.n6563 VDD 0.04656
R19590 VDD.n10148 VDD.n10136 0.0462851
R19591 VDD.n10154 VDD.n10149 0.0461165
R19592 VDD.n5728 VDD.n5723 0.0461081
R19593 VDD.n4088 VDD.n4083 0.0461081
R19594 VDD.n2447 VDD.n2442 0.0461081
R19595 VDD.n807 VDD.n802 0.0461081
R19596 VDD.n8822 VDD.n8809 0.0459877
R19597 VDD.n10017 VDD.n10010 0.0459833
R19598 VDD.n10927 VDD.n9325 0.0457021
R19599 VDD.n11021 VDD.n8737 0.0456313
R19600 VDD.n10117 VDD.n10005 0.0456006
R19601 VDD.n10631 VDD.n10133 0.0455549
R19602 VDD.n10629 VDD.n10133 0.0454465
R19603 VDD.n9087 VDD.n9086 0.0454219
R19604 VDD.n9146 VDD.n9104 0.0454219
R19605 VDD.n9136 VDD.n9105 0.0454219
R19606 VDD.n10005 VDD.n10004 0.0454042
R19607 VDD.n9325 VDD.n9321 0.0453096
R19608 VDD.n8822 VDD.n8821 0.045025
R19609 VDD.n10017 VDD.n10011 0.0450203
R19610 VDD.n10567 VDD.n10154 0.0448933
R19611 VDD.n10677 VDD.n10676 0.0448136
R19612 VDD.n10628 VDD.n10136 0.0447244
R19613 VDD.n10157 VDD.n10155 0.0443717
R19614 VDD.n10050 VDD.n10037 0.0439783
R19615 VDD.n10609 VDD.n10596 0.0439783
R19616 VDD.n10548 VDD.n10547 0.0439783
R19617 VDD.n9627 VDD.n9626 0.0439783
R19618 VDD.n9694 VDD.n9682 0.0439783
R19619 VDD.n9703 VDD.n9681 0.0439783
R19620 VDD.n10853 VDD.n10780 0.0439783
R19621 VDD.n10844 VDD.n10781 0.0439783
R19622 VDD.n10730 VDD.n10724 0.0439783
R19623 VDD.n8895 VDD.n8892 0.0439783
R19624 VDD.n9371 VDD.n9370 0.0439783
R19625 VDD.n10497 VDD.n10157 0.0437886
R19626 VDD.n9936 VDD.n9935 0.0435743
R19627 VDD.n5729 VDD.n5718 0.0435743
R19628 VDD.n4089 VDD.n4078 0.0435743
R19629 VDD.n2448 VDD.n2437 0.0435743
R19630 VDD.n808 VDD.n797 0.0435743
R19631 VDD.n10123 VDD.n10122 0.0434688
R19632 VDD.n10126 VDD.n10123 0.0434688
R19633 VDD.n10127 VDD.n10126 0.0434688
R19634 VDD.n10129 VDD.n10127 0.0434688
R19635 VDD.n10649 VDD.n10648 0.0434688
R19636 VDD.n10648 VDD.n10647 0.0434688
R19637 VDD.n10647 VDD.n10646 0.0434688
R19638 VDD.n10646 VDD.n10644 0.0434688
R19639 VDD.n10644 VDD.n10643 0.0434688
R19640 VDD.n10582 VDD.n10580 0.0434688
R19641 VDD.n10580 VDD.n10579 0.0434688
R19642 VDD.n10579 VDD.n10577 0.0434688
R19643 VDD.n10573 VDD.n10572 0.0434688
R19644 VDD.n10572 VDD.n10571 0.0434688
R19645 VDD.n10941 VDD.n9320 0.0434688
R19646 VDD.n10941 VDD.n10940 0.0434688
R19647 VDD.n10940 VDD.n10939 0.0434688
R19648 VDD.n10935 VDD.n10934 0.0434688
R19649 VDD.n10934 VDD.n10933 0.0434688
R19650 VDD.n10933 VDD.n10931 0.0434688
R19651 VDD.n10931 VDD.n10930 0.0434688
R19652 VDD.n10918 VDD.n10917 0.0434688
R19653 VDD.n10917 VDD.n10916 0.0434688
R19654 VDD.n10916 VDD.n10914 0.0434688
R19655 VDD.n10910 VDD.n10909 0.0434688
R19656 VDD.n10909 VDD.n10908 0.0434688
R19657 VDD.n10908 VDD.n9345 0.0434688
R19658 VDD.n9143 VDD.n9142 0.0434688
R19659 VDD.n9144 VDD.n9105 0.0434688
R19660 VDD.n9884 VDD.n9826 0.0434688
R19661 VDD.n9884 VDD.n9883 0.0434688
R19662 VDD.n9883 VDD.n9882 0.0434688
R19663 VDD.n9882 VDD.n9881 0.0434688
R19664 VDD.n9877 VDD.n9876 0.0434688
R19665 VDD.n9876 VDD.n9874 0.0434688
R19666 VDD.n9874 VDD.n9873 0.0434688
R19667 VDD.n9873 VDD.n9871 0.0434688
R19668 VDD.n9871 VDD.n9870 0.0434688
R19669 VDD.n9848 VDD.n9846 0.0434688
R19670 VDD.n9846 VDD.n9845 0.0434688
R19671 VDD.n9845 VDD.n9843 0.0434688
R19672 VDD.n9843 VDD.n9842 0.0434688
R19673 VDD.n9842 VDD.n9840 0.0434688
R19674 VDD.n9840 VDD.n9839 0.0434688
R19675 VDD.n9839 VDD.n9454 0.0434688
R19676 VDD.n9892 VDD.n9454 0.0434688
R19677 VDD.n9893 VDD.n9892 0.0434688
R19678 VDD.n9895 VDD.n9893 0.0434688
R19679 VDD.n9896 VDD.n9895 0.0434688
R19680 VDD.n9897 VDD.n9896 0.0434688
R19681 VDD.n9898 VDD.n9897 0.0434688
R19682 VDD.n10665 VDD.n9898 0.0434688
R19683 VDD.n12698 VDD.n12697 0.0433094
R19684 VDD.n10286 VDD.n10285 0.0433094
R19685 VDD.n10331 VDD.n10209 0.0433094
R19686 VDD.n10384 VDD.n10383 0.0433094
R19687 VDD.n9525 VDD.n9522 0.0430273
R19688 VDD.n9482 VDD.n9479 0.0430273
R19689 VDD.n8819 VDD.n8803 0.0429751
R19690 VDD.n8930 VDD.n8768 0.0429751
R19691 VDD.n10059 VDD.n10016 0.042958
R19692 VDD.n10086 VDD.n10003 0.042958
R19693 VDD.n10583 VDD.n10132 0.042958
R19694 VDD.n10559 VDD.n10558 0.042958
R19695 VDD.n10897 VDD.n10671 0.0428604
R19696 VDD.n9596 VDD.n9577 0.0426869
R19697 VDD.n9731 VDD.n9556 0.0426869
R19698 VDD.n9759 VDD.n9752 0.0426869
R19699 VDD.n9780 VDD.n9514 0.0426869
R19700 VDD.n9806 VDD.n9798 0.0426869
R19701 VDD.n10771 VDD.n10695 0.0426869
R19702 VDD.n10767 VDD.n10700 0.0426869
R19703 VDD.n8938 VDD.n8884 0.0420568
R19704 VDD.n8841 VDD.n8783 0.0420568
R19705 VDD.n9028 VDD.n8791 0.0420568
R19706 VDD.n9270 VDD.n9260 0.0420568
R19707 VDD.n9147 VDD.n9095 0.0415156
R19708 VDD.n9133 VDD.n9132 0.0415156
R19709 VDD.n9146 VDD.n9145 0.0415156
R19710 VDD.n9654 VDD.n9644 0.0412609
R19711 VDD.n9672 VDD.n9660 0.0412609
R19712 VDD.n10797 VDD.n10787 0.0412609
R19713 VDD.n10815 VDD.n10803 0.0412609
R19714 VDD.n8873 VDD.n8863 0.0412609
R19715 VDD.n8957 VDD.n8956 0.0412609
R19716 VDD.n8971 VDD.n8856 0.0412609
R19717 VDD.n8980 VDD.n8979 0.0412609
R19718 VDD.n8993 VDD.n8828 0.0412609
R19719 VDD.n9011 VDD.n8999 0.0412609
R19720 VDD.n9284 VDD.n9274 0.0412609
R19721 VDD.n9414 VDD.n9404 0.0412609
R19722 VDD VDD.n2473 0.0412609
R19723 VDD VDD.n833 0.0412609
R19724 VDD.n10576 VDD.n10573 0.041125
R19725 VDD.n10939 VDD.n10938 0.041125
R19726 VDD.n10712 VDD 0.041125
R19727 VDD.n10630 VDD.n10582 0.0403437
R19728 VDD.n10930 VDD.n10928 0.0403437
R19729 VDD.n9849 VDD.n9848 0.0403437
R19730 VDD.n10922 VDD.n9324 0.0398734
R19731 VDD.n9104 VDD.n9097 0.0395625
R19732 VDD.n12444 VDD.n12443 0.0385435
R19733 VDD.n10036 VDD.n10035 0.0385435
R19734 VDD.n10595 VDD.n10594 0.0385435
R19735 VDD.n10557 VDD.n10532 0.0385435
R19736 VDD.n9619 VDD.n9567 0.0385435
R19737 VDD.n9689 VDD.n9683 0.0385435
R19738 VDD.n9708 VDD.n9680 0.0385435
R19739 VDD.n10858 VDD.n10779 0.0385435
R19740 VDD.n10839 VDD.n10782 0.0385435
R19741 VDD.n10743 VDD.n10742 0.0385435
R19742 VDD.n9937 VDD.n9936 0.0385068
R19743 VDD.n5735 VDD.n5718 0.0385068
R19744 VDD.n5768 VDD 0.0385068
R19745 VDD.n5712 VDD 0.0385068
R19746 VDD.n4095 VDD.n4078 0.0385068
R19747 VDD.n4128 VDD 0.0385068
R19748 VDD.n4072 VDD 0.0385068
R19749 VDD.n2454 VDD.n2437 0.0385068
R19750 VDD.n2488 VDD 0.0385068
R19751 VDD.n2431 VDD 0.0385068
R19752 VDD.n814 VDD.n797 0.0385068
R19753 VDD.n848 VDD 0.0385068
R19754 VDD.n791 VDD 0.0385068
R19755 VDD.n10439 VDD.n10155 0.0380981
R19756 VDD.n10019 VDD.n10018 0.0380882
R19757 VDD.n10088 VDD.n10087 0.0380882
R19758 VDD.n10138 VDD.n10137 0.0380882
R19759 VDD.n10530 VDD.n10513 0.0380882
R19760 VDD.n9826 VDD.n9825 0.038
R19761 VDD.n10666 VDD.n10665 0.038
R19762 VDD VDD.n9956 0.0377706
R19763 VDD.n9153 VDD.n9085 0.0376094
R19764 VDD.n9096 VDD.n9087 0.0376094
R19765 VDD.n9099 VDD.n9098 0.0356562
R19766 VDD.n10948 VDD.n10946 0.035222
R19767 VDD.n9394 VDD.n9352 0.0351381
R19768 VDD.n10440 VDD.n10439 0.0345604
R19769 VDD.n5754 VDD.n5753 0.0343645
R19770 VDD.n12777 VDD.n6570 0.034112
R19771 VDD.n9930 VDD.n9927 0.033866
R19772 VDD.n10956 VDD.n9225 0.0338623
R19773 VDD.n9137 VDD.n9107 0.0337031
R19774 VDD.n9136 VDD.n9135 0.0337031
R19775 VDD.n12495 VDD.n6908 0.0331087
R19776 VDD.n12449 VDD.n12448 0.0331087
R19777 VDD.n9612 VDD.n9571 0.0331087
R19778 VDD.n9685 VDD.n9684 0.0331087
R19779 VDD.n9713 VDD.n9679 0.0331087
R19780 VDD.n10863 VDD.n10778 0.0331087
R19781 VDD.n10834 VDD.n10783 0.0331087
R19782 VDD.n10752 VDD.n10713 0.0331087
R19783 VDD.n10676 VDD.n10669 0.0330948
R19784 VDD.n9861 VDD.n9831 0.0322427
R19785 VDD.n9447 VDD.n9446 0.0319008
R19786 VDD.n9929 VDD 0.03175
R19787 VDD.n9086 VDD.n9081 0.03175
R19788 VDD.n12780 VDD 0.0315923
R19789 VDD.n10085 VDD.n10002 0.0314198
R19790 VDD.n8839 VDD.n8780 0.0312849
R19791 VDD.n9269 VDD.n9268 0.0312849
R19792 VDD VDD.n12780 0.0311212
R19793 VDD.n9357 VDD.n9350 0.0311134
R19794 VDD.n9947 VDD.n9946 0.0309412
R19795 VDD.n8936 VDD.n8885 0.0308558
R19796 VDD.n9726 VDD.n9725 0.0303913
R19797 VDD.n10823 VDD.n10786 0.0303913
R19798 VDD.n8850 VDD.n8836 0.0303913
R19799 VDD.n9019 VDD.n8827 0.0303913
R19800 VDD.n8947 VDD.n8879 0.0303913
R19801 VDD.n9294 VDD.n9273 0.0303913
R19802 VDD.n9425 VDD.n9399 0.0303913
R19803 VDD.n8926 VDD.n8925 0.0303633
R19804 VDD.n9044 VDD.n8785 0.0303633
R19805 VDD.n8806 VDD.n8792 0.0303633
R19806 VDD.n9315 VDD.n9257 0.0303633
R19807 VDD.n10925 VDD.n9329 0.0303633
R19808 VDD.n10122 VDD.n10119 0.0301875
R19809 VDD.n10571 VDD.n10569 0.0301875
R19810 VDD.n9320 VDD.n9319 0.0301875
R19811 VDD.n10511 VDD.n10152 0.0301381
R19812 VDD.n9055 VDD.n8772 0.0301368
R19813 VDD.n8759 VDD.n8756 0.0301368
R19814 VDD.n9043 VDD.n8775 0.0301368
R19815 VDD.n9252 VDD.n9251 0.0301368
R19816 VDD.n10474 VDD.n10454 0.0299811
R19817 VDD.n10475 VDD.n10452 0.0299811
R19818 VDD.n10079 VDD.n10020 0.0297969
R19819 VDD.n10113 VDD.n10112 0.0297969
R19820 VDD.n10639 VDD.n10638 0.0297969
R19821 VDD.n10526 VDD.n10510 0.0297969
R19822 VDD.n9115 VDD.n9113 0.0297969
R19823 VDD.n10012 VDD.n10009 0.0297952
R19824 VDD.n9041 VDD.n8777 0.0291557
R19825 VDD.n8894 VDD.n8757 0.0291557
R19826 VDD.n9262 VDD.n9249 0.0291557
R19827 VDD.n10465 VDD.n10443 0.0288019
R19828 VDD.n10463 VDD.n10462 0.0288019
R19829 VDD.n10464 VDD.n10444 0.0288019
R19830 VDD.n6608 VDD.n6574 0.0280588
R19831 VDD.n9954 VDD 0.0280229
R19832 VDD.n5706 VDD 0.0280227
R19833 VDD.n4066 VDD 0.0280227
R19834 VDD.n2425 VDD 0.0280227
R19835 VDD.n784 VDD 0.0280227
R19836 VDD.n10426 VDD.n10159 0.0279836
R19837 VDD.n9611 VDD.n9575 0.0278438
R19838 VDD.n9741 VDD.n9554 0.0278438
R19839 VDD.n9546 VDD.n9543 0.0278438
R19840 VDD.n9532 VDD.n9527 0.0278438
R19841 VDD.n9786 VDD.n9513 0.0278438
R19842 VDD.n9813 VDD.n9502 0.0278438
R19843 VDD.n9489 VDD.n9484 0.0278438
R19844 VDD.n10880 VDD.n10669 0.0278438
R19845 VDD.n10865 VDD.n10864 0.0278438
R19846 VDD.n10754 VDD.n10753 0.0278438
R19847 VDD.n9718 VDD.n9678 0.0276739
R19848 VDD.n10829 VDD.n10784 0.0276739
R19849 VDD.n10468 VDD.n10467 0.0276226
R19850 VDD.n5734 VDD.n5722 0.027527
R19851 VDD.n5722 VDD.n5721 0.027527
R19852 VDD.n4094 VDD.n4082 0.027527
R19853 VDD.n4082 VDD.n4081 0.027527
R19854 VDD.n2453 VDD.n2441 0.027527
R19855 VDD.n2441 VDD.n2440 0.027527
R19856 VDD.n813 VDD.n801 0.027527
R19857 VDD.n801 VDD.n800 0.027527
R19858 VDD.n6572 VDD.n6571 0.0273817
R19859 VDD.n12775 VDD.n6572 0.0273817
R19860 VDD.n12774 VDD.n6574 0.0273817
R19861 VDD.n10130 VDD.n10129 0.0270625
R19862 VDD.n10471 VDD.n10460 0.0264434
R19863 VDD.n10470 VDD.n10468 0.0264434
R19864 VDD.n9155 VDD.n9083 0.0258906
R19865 VDD.n9128 VDD.n9109 0.0258906
R19866 VDD.n9127 VDD.n9126 0.0258906
R19867 VDD.n9126 VDD.n9111 0.0258906
R19868 VDD.n9125 VDD.n9108 0.0258906
R19869 VDD.n9125 VDD.n9124 0.0258906
R19870 VDD.n9953 VDD.n9952 0.025386
R19871 VDD.n10471 VDD.n10459 0.0252642
R19872 VDD.n10470 VDD.n10463 0.0252642
R19873 VDD.n9719 VDD.n9677 0.0249565
R19874 VDD.n10828 VDD.n10785 0.0249565
R19875 VDD.n8840 VDD.n8838 0.0249565
R19876 VDD.n8845 VDD.n8837 0.0249565
R19877 VDD.n9029 VDD.n8825 0.0249565
R19878 VDD.n9024 VDD.n8826 0.0249565
R19879 VDD.n8937 VDD.n8883 0.0249565
R19880 VDD.n8942 VDD.n8881 0.0249565
R19881 VDD.n9272 VDD.n9271 0.0249565
R19882 VDD.n9299 VDD.n9298 0.0249565
R19883 VDD.n9437 VDD.n9436 0.0249565
R19884 VDD.n9427 VDD.n9395 0.0249565
R19885 VDD.n9878 VDD.n9877 0.0247187
R19886 VDD.n5768 VDD.n5711 0.024466
R19887 VDD.n4128 VDD.n4071 0.024466
R19888 VDD.n2488 VDD.n2430 0.024466
R19889 VDD.n848 VDD.n790 0.024466
R19890 VDD VDD.n6563 0.024
R19891 VDD.n10070 VDD.n10010 0.0239375
R19892 VDD.n10117 VDD.n10007 0.0239375
R19893 VDD.n10631 VDD.n10147 0.0239375
R19894 VDD.n10517 VDD.n10150 0.0239375
R19895 VDD.n9052 VDD.n8778 0.0239375
R19896 VDD.n8804 VDD.n8800 0.0239375
R19897 VDD.n8923 VDD.n8769 0.0239375
R19898 VDD.n9058 VDD.n8762 0.0239375
R19899 VDD.n9256 VDD.n9250 0.0239375
R19900 VDD.n9338 VDD.n9322 0.0239375
R19901 VDD.n9444 VDD.n9358 0.0239375
R19902 VDD.n9160 VDD.n9159 0.0239375
R19903 VDD.n9103 VDD.n9102 0.0239375
R19904 VDD VDD.n5751 0.0235263
R19905 VDD.n4112 VDD 0.0235263
R19906 VDD.n10913 VDD.n10910 0.0231563
R19907 VDD.n9356 VDD.n9227 0.022375
R19908 VDD.n9723 VDD.n9677 0.0222391
R19909 VDD.n10824 VDD.n10785 0.0222391
R19910 VDD.n8844 VDD.n8838 0.0222391
R19911 VDD.n8849 VDD.n8837 0.0222391
R19912 VDD.n9025 VDD.n8825 0.0222391
R19913 VDD.n9020 VDD.n8826 0.0222391
R19914 VDD.n8941 VDD.n8883 0.0222391
R19915 VDD.n8946 VDD.n8881 0.0222391
R19916 VDD.n9300 VDD.n9272 0.0222391
R19917 VDD.n9298 VDD.n9295 0.0222391
R19918 VDD.n9436 VDD.n9435 0.0222391
R19919 VDD.n9427 VDD.n9426 0.0222391
R19920 VDD.n10060 VDD.n10058 0.0219844
R19921 VDD.n10105 VDD.n10104 0.0219844
R19922 VDD.n10621 VDD.n10620 0.0219844
R19923 VDD.n10560 VDD.n10509 0.0219844
R19924 VDD.n9037 VDD.n9036 0.0219844
R19925 VDD.n8818 VDD.n8814 0.0219844
R19926 VDD.n8919 VDD.n8918 0.0219844
R19927 VDD.n8899 VDD.n8898 0.0219844
R19928 VDD.n9306 VDD.n9305 0.0219844
R19929 VDD.n9335 VDD.n9334 0.0219844
R19930 VDD.n9382 VDD.n9381 0.0219844
R19931 VDD.n9119 VDD.n9118 0.0219844
R19932 VDD.n5775 VDD.n5708 0.0218675
R19933 VDD.n4135 VDD.n4068 0.0218675
R19934 VDD.n2495 VDD.n2427 0.0218675
R19935 VDD.n10461 VDD.n10458 0.0217264
R19936 VDD.n10466 VDD.n10457 0.0217264
R19937 VDD.n10483 VDD.n10445 0.0217264
R19938 VDD VDD.n9953 0.0217156
R19939 VDD.n9956 VDD 0.0217156
R19940 VDD.n9937 VDD.n9922 0.0215953
R19941 VDD.n5720 VDD.n5711 0.0215953
R19942 VDD.n4080 VDD.n4071 0.0215953
R19943 VDD.n2439 VDD.n2430 0.0215953
R19944 VDD.n799 VDD.n790 0.0215953
R19945 VDD.n12778 VDD.n6569 0.0211408
R19946 VDD.n10901 VDD.n10659 0.0210308
R19947 VDD.n10914 VDD.n10913 0.0208125
R19948 VDD.n9858 VDD.n9828 0.0205059
R19949 VDD.n10886 VDD.n10885 0.0205059
R19950 VDD.n9861 VDD.n9830 0.0200312
R19951 VDD.n10675 VDD.n10672 0.0200312
R19952 VDD.n9161 VDD.n9160 0.0200312
R19953 VDD.n9162 VDD.n9081 0.0200312
R19954 VDD.n8755 VDD.n8752 0.0198977
R19955 VDD.n11018 VDD.n11017 0.0197278
R19956 VDD.n9030 VDD.n8824 0.0196275
R19957 VDD.n9714 VDD.n9678 0.0195217
R19958 VDD.n10833 VDD.n10784 0.0195217
R19959 VDD.n10488 VDD.n10156 0.0193679
R19960 VDD.n5776 VDD.n5774 0.0193464
R19961 VDD.n4136 VDD.n4134 0.0193464
R19962 VDD.n2496 VDD.n2494 0.0193464
R19963 VDD.n9881 VDD.n9878 0.01925
R19964 VDD.n8921 VDD.n8920 0.0186403
R19965 VDD.n9035 VDD.n8786 0.0186403
R19966 VDD.n8817 VDD.n8793 0.0186403
R19967 VDD.n9304 VDD.n9259 0.0186403
R19968 VDD.n9337 VDD.n9336 0.0186403
R19969 VDD.n9601 VDD.n9578 0.0185773
R19970 VDD.n9537 VDD.n9536 0.0185773
R19971 VDD.n9790 VDD.n9515 0.0185773
R19972 VDD.n9494 VDD.n9493 0.0185773
R19973 VDD.n10491 VDD.n10438 0.0181887
R19974 VDD.n9141 VDD.n9106 0.0180781
R19975 VDD.n9133 VDD.n9107 0.0180781
R19976 VDD.n9122 VDD.n9114 0.0180781
R19977 VDD.n9135 VDD.n9134 0.0180781
R19978 VDD.n9123 VDD.n9112 0.0180781
R19979 VDD.n9042 VDD.n8779 0.0176875
R19980 VDD.n9318 VDD.n9248 0.0176875
R19981 VDD.n9187 VDD.n9080 0.0176875
R19982 VDD.n4114 VDD.n4113 0.0174323
R19983 VDD.n10649 VDD.n10130 0.0169062
R19984 VDD.n10498 VDD.n10156 0.0169062
R19985 VDD.n11006 VDD.n8754 0.0169062
R19986 VDD.n9080 VDD.n9079 0.0169062
R19987 VDD.n11019 VDD.n8738 0.0169062
R19988 VDD.n8840 VDD.n8839 0.0168893
R19989 VDD.n9030 VDD.n9029 0.0168893
R19990 VDD.n8937 VDD.n8936 0.0168893
R19991 VDD.n9271 VDD.n9269 0.0168893
R19992 VDD.n9437 VDD.n9394 0.0168893
R19993 VDD.n12485 VDD.n6567 0.0168043
R19994 VDD.n9727 VDD.n9726 0.0168043
R19995 VDD.n10819 VDD.n10786 0.0168043
R19996 VDD.n8854 VDD.n8836 0.0168043
R19997 VDD.n9015 VDD.n8827 0.0168043
R19998 VDD.n8951 VDD.n8879 0.0168043
R19999 VDD.n9290 VDD.n9273 0.0168043
R20000 VDD.n9420 VDD.n9399 0.0168043
R20001 VDD.n5774 VDD 0.0166045
R20002 VDD.n4134 VDD 0.0166045
R20003 VDD.n2494 VDD 0.0166045
R20004 VDD.n786 VDD 0.0166045
R20005 VDD.n5735 VDD.n5734 0.0165473
R20006 VDD.n4095 VDD.n4094 0.0165473
R20007 VDD.n2454 VDD.n2453 0.0165473
R20008 VDD.n814 VDD.n813 0.0165473
R20009 VDD.n9597 VDD.n9596 0.016125
R20010 VDD.n9590 VDD.n9581 0.016125
R20011 VDD.n9731 VDD.n9552 0.016125
R20012 VDD.n9736 VDD.n9551 0.016125
R20013 VDD.n9746 VDD.n9745 0.016125
R20014 VDD.n9752 VDD.n9751 0.016125
R20015 VDD.n9760 VDD.n9541 0.016125
R20016 VDD.n9753 VDD.n9542 0.016125
R20017 VDD.n9776 VDD.n9522 0.016125
R20018 VDD.n9771 VDD.n9770 0.016125
R20019 VDD.n9780 VDD.n9779 0.016125
R20020 VDD.n9794 VDD.n9509 0.016125
R20021 VDD.n9798 VDD.n9797 0.016125
R20022 VDD.n9807 VDD.n9498 0.016125
R20023 VDD.n9803 VDD.n9499 0.016125
R20024 VDD.n9823 VDD.n9479 0.016125
R20025 VDD.n9818 VDD.n9817 0.016125
R20026 VDD.n9851 VDD.n9850 0.016125
R20027 VDD.n9853 VDD.n9835 0.016125
R20028 VDD.n10880 VDD.n10673 0.016125
R20029 VDD.n10894 VDD.n10677 0.016125
R20030 VDD.n10772 VDD.n10771 0.016125
R20031 VDD.n10875 VDD.n10874 0.016125
R20032 VDD.n10869 VDD.n10775 0.016125
R20033 VDD.n10768 VDD.n10767 0.016125
R20034 VDD.n10703 VDD.n10696 0.016125
R20035 VDD.n10758 VDD.n10709 0.016125
R20036 VDD.n9448 VDD.n9351 0.016125
R20037 VDD.n9147 VDD.n9094 0.016125
R20038 VDD.n9142 VDD.n9141 0.016125
R20039 VDD.n9163 VDD.n9162 0.016125
R20040 VDD.n11022 VDD.n8739 0.016125
R20041 VDD.n5726 VDD.n5723 0.0157415
R20042 VDD.n4086 VDD.n4083 0.0157415
R20043 VDD.n2445 VDD.n2442 0.0157415
R20044 VDD.n805 VDD.n802 0.0157415
R20045 VDD.n6561 VDD 0.0146
R20046 VDD.n4921 VDD 0.0146
R20047 VDD.n3281 VDD 0.0146
R20048 VDD.n1640 VDD 0.0146
R20049 VDD.n10640 VDD.n10135 0.0145625
R20050 VDD.n9867 VDD.n9832 0.0145625
R20051 VDD.n10942 VDD.n9242 0.0143978
R20052 VDD.n10942 VDD.n9245 0.0143978
R20053 VDD.n9245 VDD.n9241 0.0143978
R20054 VDD.n10936 VDD.n9233 0.0143978
R20055 VDD.n10932 VDD.n9233 0.0143978
R20056 VDD.n10932 VDD.n9240 0.0143978
R20057 VDD.n10929 VDD.n9240 0.0143978
R20058 VDD.n10929 VDD.n9234 0.0143978
R20059 VDD.n10919 VDD.n9239 0.0143978
R20060 VDD.n10915 VDD.n9239 0.0143978
R20061 VDD.n10915 VDD.n9235 0.0143978
R20062 VDD.n10911 VDD.n9238 0.0143978
R20063 VDD.n10907 VDD.n9238 0.0143978
R20064 VDD.n10907 VDD.n10906 0.0143978
R20065 VDD.n9885 VDD.n9472 0.0143978
R20066 VDD.n9885 VDD.n9473 0.0143978
R20067 VDD.n9473 VDD.n9467 0.0143978
R20068 VDD.n9880 VDD.n9467 0.0143978
R20069 VDD.n9875 VDD.n9460 0.0143978
R20070 VDD.n9875 VDD.n9466 0.0143978
R20071 VDD.n9872 VDD.n9466 0.0143978
R20072 VDD.n9872 VDD.n9461 0.0143978
R20073 VDD.n9869 VDD.n9461 0.0143978
R20074 VDD.n9847 VDD.n9465 0.0143978
R20075 VDD.n9847 VDD.n9462 0.0143978
R20076 VDD.n9844 VDD.n9462 0.0143978
R20077 VDD.n9844 VDD.n9464 0.0143978
R20078 VDD.n9841 VDD.n9464 0.0143978
R20079 VDD.n9841 VDD.n9463 0.0143978
R20080 VDD.n9463 VDD.n9455 0.0143978
R20081 VDD.n9890 VDD.n9455 0.0143978
R20082 VDD.n9891 VDD.n9890 0.0143978
R20083 VDD.n9891 VDD.n9452 0.0143978
R20084 VDD.n9894 VDD.n9452 0.0143978
R20085 VDD.n9894 VDD.n9451 0.0143978
R20086 VDD.n9453 VDD.n9451 0.0143978
R20087 VDD.n10902 VDD.n9453 0.0143978
R20088 VDD.n10902 VDD.n9901 0.0143978
R20089 VDD.n10121 VDD.n9987 0.0143978
R20090 VDD.n10125 VDD.n9987 0.0143978
R20091 VDD.n10128 VDD.n9991 0.0143978
R20092 VDD.n10650 VDD.n10000 0.0143978
R20093 VDD.n10000 VDD.n9990 0.0143978
R20094 VDD.n10645 VDD.n9990 0.0143978
R20095 VDD.n10645 VDD.n9988 0.0143978
R20096 VDD.n10642 VDD.n9988 0.0143978
R20097 VDD.n10581 VDD.n9989 0.0143978
R20098 VDD.n10581 VDD.n9986 0.0143978
R20099 VDD.n10578 VDD.n9986 0.0143978
R20100 VDD.n10578 VDD.n9993 0.0143978
R20101 VDD.n10574 VDD.n9985 0.0143978
R20102 VDD.n10570 VDD.n9985 0.0143978
R20103 VDD.n10022 VDD.n10011 0.0141719
R20104 VDD.n10090 VDD.n10004 0.0141719
R20105 VDD.n10629 VDD.n10140 0.0141719
R20106 VDD.n10525 VDD.n10152 0.0141719
R20107 VDD.n9599 VDD.n9575 0.0141719
R20108 VDD.n9741 VDD.n9553 0.0141719
R20109 VDD.n9767 VDD.n9543 0.0141719
R20110 VDD.n9532 VDD.n9520 0.0141719
R20111 VDD.n9786 VDD.n9508 0.0141719
R20112 VDD.n9814 VDD.n9813 0.0141719
R20113 VDD.n9489 VDD.n9477 0.0141719
R20114 VDD.n9858 VDD.n9830 0.0141719
R20115 VDD.n10886 VDD.n10675 0.0141719
R20116 VDD.n10866 VDD.n10865 0.0141719
R20117 VDD.n10755 VDD.n10754 0.0141719
R20118 VDD.n9154 VDD.n9153 0.0141719
R20119 VDD.n6911 VDD.n6908 0.014087
R20120 VDD.n12448 VDD.n12445 0.014087
R20121 VDD.n9618 VDD.n9571 0.014087
R20122 VDD.n9688 VDD.n9685 0.014087
R20123 VDD.n9709 VDD.n9679 0.014087
R20124 VDD.n10859 VDD.n10778 0.014087
R20125 VDD.n10838 VDD.n10783 0.014087
R20126 VDD.n10716 VDD.n10713 0.014087
R20127 VDD.n10125 VDD.n10124 0.0138925
R20128 VDD.n10921 VDD.n9323 0.0137813
R20129 VDD.n9957 VDD 0.0136881
R20130 VDD.n10937 VDD.n9241 0.0136398
R20131 VDD.n10575 VDD.n10574 0.0136398
R20132 VDD.n10643 VDD.n10131 0.013
R20133 VDD.n10918 VDD.n9326 0.013
R20134 VDD.n9870 VDD.n9827 0.013
R20135 VDD.n11014 VDD.n8743 0.0128788
R20136 VDD.n9067 VDD.n8751 0.0128788
R20137 VDD.n11004 VDD.n8751 0.0128788
R20138 VDD.n11015 VDD.n11014 0.0128788
R20139 VDD.n6560 VDD.n6559 0.0127863
R20140 VDD.n4920 VDD.n4919 0.0127863
R20141 VDD.n3280 VDD.n3279 0.0127863
R20142 VDD.n9733 VDD.n9558 0.0127111
R20143 VDD.n9757 VDD.n9756 0.0127111
R20144 VDD.n9801 VDD.n9799 0.0127111
R20145 VDD.n10873 VDD.n10872 0.0127111
R20146 VDD.n10760 VDD.n10707 0.0127111
R20147 VDD.n9472 VDD.n9471 0.012629
R20148 VDD.n10661 VDD.n9901 0.012629
R20149 VDD.n10485 VDD.n10441 0.0122925
R20150 VDD.n10489 VDD.n10488 0.0122925
R20151 VDD.n10490 VDD.n10440 0.0122925
R20152 VDD.n10069 VDD.n10009 0.0122188
R20153 VDD.n10058 VDD.n10014 0.0122188
R20154 VDD.n10093 VDD.n10084 0.0122188
R20155 VDD.n10106 VDD.n10105 0.0122188
R20156 VDD.n10628 VDD.n10584 0.0122188
R20157 VDD.n10620 VDD.n10619 0.0122188
R20158 VDD.n10567 VDD.n10153 0.0122188
R20159 VDD.n10509 VDD.n10508 0.0122188
R20160 VDD.n9609 VDD.n9581 0.0122188
R20161 VDD.n9770 VDD.n9539 0.0122188
R20162 VDD.n9794 VDD.n9793 0.0122188
R20163 VDD.n9817 VDD.n9496 0.0122188
R20164 VDD.n9866 VDD.n9835 0.0122188
R20165 VDD.n10894 VDD.n10668 0.0122188
R20166 VDD.n9038 VDD.n9037 0.0122188
R20167 VDD.n9046 VDD.n9045 0.0122188
R20168 VDD.n8814 VDD.n8810 0.0122188
R20169 VDD.n8809 VDD.n8807 0.0122188
R20170 VDD.n8918 VDD.n8770 0.0122188
R20171 VDD.n8924 VDD.n8774 0.0122188
R20172 VDD.n8900 VDD.n8899 0.0122188
R20173 VDD.n9064 VDD.n9063 0.0122188
R20174 VDD.n9307 VDD.n9306 0.0122188
R20175 VDD.n9317 VDD.n9316 0.0122188
R20176 VDD.n9334 VDD.n9333 0.0122188
R20177 VDD.n10927 VDD.n9327 0.0122188
R20178 VDD.n9381 VDD.n9354 0.0122188
R20179 VDD.n9389 VDD.n9353 0.0122188
R20180 VDD.n9098 VDD.n9085 0.0122188
R20181 VDD.n9137 VDD.n9106 0.0122188
R20182 VDD.n9119 VDD.n9114 0.0122188
R20183 VDD.n9097 VDD.n9096 0.0122188
R20184 VDD.n5770 VDD 0.0121071
R20185 VDD.n4130 VDD 0.0121071
R20186 VDD.n2490 VDD 0.0121071
R20187 VDD.n850 VDD 0.0121071
R20188 VDD.n6558 VDD.n5772 0.0115787
R20189 VDD.n4918 VDD.n4132 0.0115787
R20190 VDD.n3278 VDD.n2492 0.0115787
R20191 VDD.n1638 VDD.n1227 0.0115787
R20192 VDD.n5730 VDD.n5729 0.0114797
R20193 VDD.n5721 VDD.n5720 0.0114797
R20194 VDD.n4090 VDD.n4089 0.0114797
R20195 VDD.n4081 VDD.n4080 0.0114797
R20196 VDD.n2449 VDD.n2448 0.0114797
R20197 VDD.n2440 VDD.n2439 0.0114797
R20198 VDD.n809 VDD.n808 0.0114797
R20199 VDD.n800 VDD.n799 0.0114797
R20200 VDD.n9445 VDD.n9345 0.0114375
R20201 VDD.n10456 VDD.n10450 0.0111132
R20202 VDD.n10487 VDD.n10441 0.0111132
R20203 VDD.n10898 VDD.n10670 0.0106562
R20204 VDD.n10896 VDD.n10670 0.0106562
R20205 VDD.n10070 VDD.n10069 0.0102656
R20206 VDD.n10093 VDD.n10007 0.0102656
R20207 VDD.n10584 VDD.n10147 0.0102656
R20208 VDD.n10517 VDD.n10153 0.0102656
R20209 VDD.n9045 VDD.n8778 0.0102656
R20210 VDD.n8807 VDD.n8804 0.0102656
R20211 VDD.n8924 VDD.n8923 0.0102656
R20212 VDD.n9063 VDD.n8762 0.0102656
R20213 VDD.n9316 VDD.n9256 0.0102656
R20214 VDD.n9338 VDD.n9327 0.0102656
R20215 VDD.n9389 VDD.n9358 0.0102656
R20216 VDD.n9242 VDD.n9236 0.0101021
R20217 VDD.n10920 VDD.n10919 0.0101021
R20218 VDD.n10121 VDD.n10120 0.0101021
R20219 VDD.n10570 VDD.n9994 0.0101021
R20220 VDD.n10456 VDD.n10451 0.00993396
R20221 VDD.n10485 VDD.n10484 0.00993396
R20222 VDD.n9869 VDD.n9868 0.00984946
R20223 VDD.n10642 VDD.n10641 0.00984946
R20224 VDD.n9930 VDD.n9929 0.00979054
R20225 VDD.n10083 VDD.n10008 0.00957737
R20226 VDD.n10118 VDD.n10001 0.00957737
R20227 VDD.n10512 VDD.n10499 0.00957737
R20228 VDD.n10158 VDD.n10156 0.00957737
R20229 VDD.n10080 VDD.n10008 0.00957737
R20230 VDD.n10114 VDD.n10001 0.00957737
R20231 VDD.n10531 VDD.n10512 0.00957737
R20232 VDD.n8893 VDD.n8761 0.00957737
R20233 VDD.n9054 VDD.n8773 0.00957737
R20234 VDD.n8820 VDD.n8802 0.00957737
R20235 VDD.n9057 VDD.n8761 0.00957737
R20236 VDD.n8929 VDD.n8773 0.00957737
R20237 VDD.n8823 VDD.n8802 0.00957737
R20238 VDD.n9344 VDD.n9326 0.00957737
R20239 VDD.n10949 VDD.n9226 0.00957737
R20240 VDD.n10921 VDD.n9344 0.00957737
R20241 VDD.n10949 VDD.n10947 0.00957737
R20242 VDD.n9610 VDD.n9579 0.00957737
R20243 VDD.n9748 VDD.n9747 0.00957737
R20244 VDD.n9768 VDD.n9540 0.00957737
R20245 VDD.n9777 VDD.n9519 0.00957737
R20246 VDD.n9792 VDD.n9507 0.00957737
R20247 VDD.n9815 VDD.n9497 0.00957737
R20248 VDD.n9824 VDD.n9476 0.00957737
R20249 VDD.n10777 VDD.n10774 0.00957737
R20250 VDD.n10712 VDD.n10698 0.00957737
R20251 VDD.n10970 VDD.n10969 0.00957737
R20252 VDD.n10708 VDD.n10698 0.00957737
R20253 VDD.n9495 VDD.n9476 0.00957737
R20254 VDD.n9805 VDD.n9497 0.00957737
R20255 VDD.n9538 VDD.n9519 0.00957737
R20256 VDD.n9795 VDD.n9507 0.00957737
R20257 VDD.n9758 VDD.n9540 0.00957737
R20258 VDD.n9588 VDD.n9579 0.00957737
R20259 VDD.n9749 VDD.n9748 0.00957737
R20260 VDD.n10777 VDD.n10770 0.00957737
R20261 VDD.n10970 VDD.n9213 0.00957737
R20262 VDD.n11007 VDD.n8748 0.00955797
R20263 VDD.n11013 VDD.n11012 0.00955797
R20264 VDD.n10906 VDD.n9449 0.00934409
R20265 VDD.n5753 VDD.n5752 0.00927193
R20266 VDD.n4113 VDD.n4111 0.00927193
R20267 VDD.n9213 VDD.n9211 0.00923422
R20268 VDD.n10081 VDD.n10015 0.0091882
R20269 VDD.n10116 VDD.n10115 0.0091882
R20270 VDD.n10134 VDD.n10131 0.0091882
R20271 VDD.n10568 VDD.n10151 0.0091882
R20272 VDD.n10640 VDD.n10134 0.0091882
R20273 VDD.n10081 VDD.n10080 0.0091882
R20274 VDD.n10115 VDD.n10114 0.0091882
R20275 VDD.n10531 VDD.n10151 0.0091882
R20276 VDD.n11007 VDD.n8749 0.0091882
R20277 VDD.n9065 VDD.n8758 0.0091882
R20278 VDD.n8929 VDD.n8767 0.0091882
R20279 VDD.n9042 VDD.n8776 0.0091882
R20280 VDD.n8823 VDD.n8801 0.0091882
R20281 VDD.n8893 VDD.n8758 0.0091882
R20282 VDD.n8812 VDD.n8801 0.0091882
R20283 VDD.n9053 VDD.n8776 0.0091882
R20284 VDD.n9056 VDD.n8767 0.0091882
R20285 VDD.n11002 VDD.n8749 0.0091882
R20286 VDD.n9255 VDD.n9248 0.0091882
R20287 VDD.n9448 VDD.n9349 0.0091882
R20288 VDD.n10955 VDD.n10954 0.0091882
R20289 VDD.n9445 VDD.n9349 0.0091882
R20290 VDD.n10954 VDD.n10947 0.0091882
R20291 VDD.n9255 VDD.n9254 0.0091882
R20292 VDD.n9610 VDD.n9576 0.0091882
R20293 VDD.n9747 VDD.n9555 0.0091882
R20294 VDD.n9750 VDD.n9544 0.0091882
R20295 VDD.n9769 VDD.n9521 0.0091882
R20296 VDD.n9792 VDD.n9511 0.0091882
R20297 VDD.n9805 VDD.n9501 0.0091882
R20298 VDD.n9816 VDD.n9478 0.0091882
R20299 VDD.n9834 VDD.n9827 0.0091882
R20300 VDD.n10774 VDD.n10773 0.0091882
R20301 VDD.n10769 VDD.n10697 0.0091882
R20302 VDD.n9495 VDD.n9478 0.0091882
R20303 VDD.n10773 VDD.n10674 0.0091882
R20304 VDD.n10708 VDD.n10697 0.0091882
R20305 VDD.n9867 VDD.n9834 0.0091882
R20306 VDD.n9796 VDD.n9501 0.0091882
R20307 VDD.n9778 VDD.n9511 0.0091882
R20308 VDD.n9538 VDD.n9521 0.0091882
R20309 VDD.n9598 VDD.n9576 0.0091882
R20310 VDD.n9587 VDD.n9555 0.0091882
R20311 VDD.n9758 VDD.n9544 0.0091882
R20312 VDD.n9215 VDD.n9211 0.00914234
R20313 VDD.n10128 VDD.n9999 0.0090914
R20314 VDD.n5730 VDD.n5728 0.00894595
R20315 VDD.n4090 VDD.n4088 0.00894595
R20316 VDD.n2449 VDD.n2447 0.00894595
R20317 VDD.n809 VDD.n807 0.00894595
R20318 VDD.n2473 VDD.n2470 0.00887321
R20319 VDD.n2473 VDD.n2472 0.00887321
R20320 VDD.n833 VDD.n830 0.00887321
R20321 VDD.n833 VDD.n832 0.00887321
R20322 VDD.n11011 VDD.n8744 0.00867391
R20323 VDD.n12443 VDD.n12441 0.00865217
R20324 VDD.n10051 VDD.n10036 0.00865217
R20325 VDD.n10610 VDD.n10595 0.00865217
R20326 VDD.n10536 VDD.n10532 0.00865217
R20327 VDD.n9625 VDD.n9567 0.00865217
R20328 VDD.n9693 VDD.n9683 0.00865217
R20329 VDD.n9704 VDD.n9680 0.00865217
R20330 VDD.n10854 VDD.n10779 0.00865217
R20331 VDD.n10843 VDD.n10782 0.00865217
R20332 VDD.n10742 VDD.n10741 0.00865217
R20333 VDD.n11016 VDD.n11013 0.00865217
R20334 VDD.n9879 VDD.n9460 0.00833333
R20335 VDD.n10060 VDD.n10059 0.0083125
R20336 VDD.n10104 VDD.n10003 0.0083125
R20337 VDD.n10621 VDD.n10583 0.0083125
R20338 VDD.n10560 VDD.n10559 0.0083125
R20339 VDD.n9036 VDD.n8777 0.0083125
R20340 VDD.n8819 VDD.n8818 0.0083125
R20341 VDD.n8919 VDD.n8768 0.0083125
R20342 VDD.n8898 VDD.n8757 0.0083125
R20343 VDD.n9305 VDD.n9249 0.0083125
R20344 VDD.n9335 VDD.n9324 0.0083125
R20345 VDD.n9382 VDD.n9357 0.0083125
R20346 VDD.n9159 VDD.n9083 0.0083125
R20347 VDD.n9132 VDD.n9109 0.0083125
R20348 VDD.n9128 VDD.n9127 0.0083125
R20349 VDD.n10453 VDD.n10442 0.0081375
R20350 VDD.n9348 VDD.n9228 0.00808064
R20351 VDD.n4923 VDD.n4922 0.00794492
R20352 VDD.n3283 VDD.n3282 0.00794492
R20353 VDD.n1642 VDD.n1641 0.00794492
R20354 VDD.n10912 VDD.n10911 0.00782796
R20355 VDD.n11007 VDD.n8746 0.00774638
R20356 VDD.n10459 VDD.n10458 0.00757547
R20357 VDD.n10896 VDD.n10895 0.00753125
R20358 VDD.n6559 VDD.n5773 0.00744444
R20359 VDD.n4919 VDD.n4133 0.00744444
R20360 VDD.n3279 VDD.n2493 0.00744444
R20361 VDD.n10912 VDD.n9235 0.00706989
R20362 VDD.n10472 VDD.n10455 0.00694587
R20363 VDD.n10707 VDD.n10696 0.00685176
R20364 VDD.n10874 VDD.n10873 0.00685176
R20365 VDD.n9799 VDD.n9498 0.00685176
R20366 VDD.n9757 VDD.n9541 0.00685176
R20367 VDD.n9558 VDD.n9551 0.00685176
R20368 VDD.n9887 VDD.n9468 0.0068172
R20369 VDD.n11017 VDD.n11015 0.00678574
R20370 VDD.n10945 VDD.n9227 0.00675
R20371 VDD.n10898 VDD.n10667 0.00675
R20372 VDD.n9067 VDD.n8755 0.00661507
R20373 VDD.n9880 VDD.n9879 0.00656452
R20374 VDD.n9949 VDD.n9948 0.00641216
R20375 VDD.n10460 VDD.n10457 0.00639623
R20376 VDD.n6558 VDD.n5777 0.00638768
R20377 VDD.n5705 VDD.n5704 0.00638768
R20378 VDD.n4918 VDD.n4137 0.00638768
R20379 VDD.n4065 VDD.n4064 0.00638768
R20380 VDD.n3278 VDD.n2497 0.00638768
R20381 VDD.n2424 VDD.n2423 0.00638768
R20382 VDD.n1227 VDD.n855 0.00638768
R20383 VDD.n782 VDD.n781 0.00638768
R20384 VDD.n9609 VDD.n9608 0.00635938
R20385 VDD.n9539 VDD.n9526 0.00635938
R20386 VDD.n9793 VDD.n9512 0.00635938
R20387 VDD.n9496 VDD.n9483 0.00635938
R20388 VDD.n9866 VDD.n9865 0.00635938
R20389 VDD.n10891 VDD.n10668 0.00635938
R20390 VDD.n10897 VDD.n10672 0.00635938
R20391 VDD.n11008 VDD.n8747 0.00635938
R20392 VDD.n9155 VDD.n9154 0.00635938
R20393 VDD.n9102 VDD.n9094 0.00635938
R20394 VDD.n9654 VDD.n9653 0.00593478
R20395 VDD.n9662 VDD.n9660 0.00593478
R20396 VDD.n10797 VDD.n10796 0.00593478
R20397 VDD.n10805 VDD.n10803 0.00593478
R20398 VDD.n8873 VDD.n8872 0.00593478
R20399 VDD.n8957 VDD.n8859 0.00593478
R20400 VDD.n8971 VDD.n8970 0.00593478
R20401 VDD.n8980 VDD.n8831 0.00593478
R20402 VDD.n8993 VDD.n8992 0.00593478
R20403 VDD.n9001 VDD.n8999 0.00593478
R20404 VDD.n9284 VDD.n9283 0.00593478
R20405 VDD.n9414 VDD.n9413 0.00593478
R20406 VDD.n10650 VDD.n9999 0.00580645
R20407 VDD.n11010 VDD.n8745 0.0056087
R20408 VDD.n9449 VDD.n9348 0.00555376
R20409 VDD.n9066 VDD.n8754 0.0051875
R20410 VDD.n11022 VDD.n8741 0.0051875
R20411 VDD.n9868 VDD.n9465 0.00504839
R20412 VDD.n10641 VDD.n9989 0.00504839
R20413 VDD.n8752 VDD.n8745 0.00492754
R20414 VDD.n10679 VDD.n10673 0.00490286
R20415 VDD.n9850 VDD.n9833 0.00490286
R20416 VDD.n10904 VDD.n9236 0.0047957
R20417 VDD.n10920 VDD.n9234 0.0047957
R20418 VDD.n10944 VDD.n9230 0.0047957
R20419 VDD.n10120 VDD.n9992 0.0047957
R20420 VDD.n10657 VDD.n9994 0.0047957
R20421 VDD.n10486 VDD.n10442 0.00449057
R20422 VDD.n10079 VDD.n10019 0.00440625
R20423 VDD.n10082 VDD.n10014 0.00440625
R20424 VDD.n10113 VDD.n10088 0.00440625
R20425 VDD.n10106 VDD.n10002 0.00440625
R20426 VDD.n10639 VDD.n10138 0.00440625
R20427 VDD.n10619 VDD.n10148 0.00440625
R20428 VDD.n10513 VDD.n10510 0.00440625
R20429 VDD.n10508 VDD.n10149 0.00440625
R20430 VDD.n9746 VDD.n9553 0.00440625
R20431 VDD.n9767 VDD.n9542 0.00440625
R20432 VDD.n9814 VDD.n9499 0.00440625
R20433 VDD.n10866 VDD.n10775 0.00440625
R20434 VDD.n10755 VDD.n10709 0.00440625
R20435 VDD.n9038 VDD.n8775 0.00440625
R20436 VDD.n8821 VDD.n8810 0.00440625
R20437 VDD.n9055 VDD.n8770 0.00440625
R20438 VDD.n8900 VDD.n8756 0.00440625
R20439 VDD.n11003 VDD.n11002 0.00440625
R20440 VDD.n9307 VDD.n9251 0.00440625
R20441 VDD.n9333 VDD.n9321 0.00440625
R20442 VDD.n9446 VDD.n9354 0.00440625
R20443 VDD.n9103 VDD.n9099 0.00440625
R20444 VDD.n9143 VDD.n9095 0.00440625
R20445 VDD.n9122 VDD.n9113 0.00440625
R20446 VDD.n9145 VDD.n9144 0.00440625
R20447 VDD.n11023 VDD.n8736 0.00433093
R20448 VDD.n9232 VDD.n9230 0.00429032
R20449 VDD.n10653 VDD.n9992 0.00429032
R20450 VDD.n10657 VDD.n9997 0.00429032
R20451 VDD.n10473 VDD.n10472 0.00397228
R20452 VDD VDD.n12782 0.00363333
R20453 VDD.n10630 VDD.n10135 0.003625
R20454 VDD.n10928 VDD.n9323 0.003625
R20455 VDD.n9849 VDD.n9832 0.003625
R20456 VDD.n10667 VDD.n10666 0.003625
R20457 VDD.n10040 VDD.n10037 0.00321739
R20458 VDD.n10599 VDD.n10596 0.00321739
R20459 VDD.n10547 VDD.n10546 0.00321739
R20460 VDD.n9626 VDD.n9562 0.00321739
R20461 VDD.n9698 VDD.n9682 0.00321739
R20462 VDD.n9699 VDD.n9681 0.00321739
R20463 VDD.n10849 VDD.n10780 0.00321739
R20464 VDD.n10848 VDD.n10781 0.00321739
R20465 VDD.n10734 VDD.n10730 0.00321739
R20466 VDD.n8892 VDD.n8890 0.00321739
R20467 VDD.n9372 VDD.n9371 0.00321739
R20468 VDD.n9925 VDD.n9924 0.00303378
R20469 VDD VDD.n5712 0.00303378
R20470 VDD VDD.n4072 0.00303378
R20471 VDD VDD.n2431 0.00303378
R20472 VDD VDD.n791 0.00303378
R20473 VDD.n9599 VDD.n9578 0.00295228
R20474 VDD.n9537 VDD.n9520 0.00295228
R20475 VDD.n9515 VDD.n9508 0.00295228
R20476 VDD.n9494 VDD.n9477 0.00295228
R20477 VDD.n10466 VDD.n10465 0.00285849
R20478 VDD.n10467 VDD.n10464 0.00285849
R20479 VDD.n10491 VDD.n10490 0.00285849
R20480 VDD.n10577 VDD.n10576 0.00284375
R20481 VDD.n10938 VDD.n10935 0.00284375
R20482 VDD.n10654 VDD.n9998 0.00278115
R20483 VDD.n10652 VDD.n9998 0.00278115
R20484 VDD.n5775 VDD.n5773 0.00263675
R20485 VDD.n4135 VDD.n4133 0.00263675
R20486 VDD.n2495 VDD.n2493 0.00263675
R20487 VDD.n854 VDD.n853 0.00263675
R20488 VDD.n9474 VDD.n9457 0.00262546
R20489 VDD.n9470 VDD.n9457 0.00262546
R20490 VDD.n10944 VDD.n9228 0.00252151
R20491 VDD.n12700 VDD.n6609 0.00251613
R20492 VDD.n10022 VDD.n10020 0.00245312
R20493 VDD.n10112 VDD.n10090 0.00245312
R20494 VDD.n10638 VDD.n10140 0.00245312
R20495 VDD.n10526 VDD.n10525 0.00245312
R20496 VDD.n10163 VDD.n6918 0.00244542
R20497 VDD.n10664 VDD.n9899 0.00243946
R20498 VDD.n10943 VDD.n9231 0.00243946
R20499 VDD.n9231 VDD.n9229 0.00243946
R20500 VDD.n10664 VDD.n10663 0.00243946
R20501 VDD.n5777 VDD.n5776 0.00231159
R20502 VDD.n4137 VDD.n4136 0.00231159
R20503 VDD.n2497 VDD.n2496 0.00231159
R20504 VDD.n855 VDD.n852 0.00231159
R20505 VDD.n9887 VDD.n9471 0.00226882
R20506 VDD.n10900 VDD.n10661 0.00226882
R20507 VDD.n9957 VDD.n9954 0.00222018
R20508 VDD.n11005 VDD.n11004 0.0022029
R20509 VDD.n10433 VDD.n6916 0.00207156
R20510 VDD.n10421 VDD.n6917 0.00207156
R20511 VDD.n9171 VDD.n9170 0.00207156
R20512 VDD.n9175 VDD.n9167 0.00207156
R20513 VDD.n10950 VDD.n9202 0.00207156
R20514 VDD.n9223 VDD.n9203 0.00207156
R20515 VDD.n10998 VDD.n10997 0.00207156
R20516 VDD.n9356 VDD.n9351 0.0020625
R20517 VDD.n9171 VDD.n9077 0.00194557
R20518 VDD.n9175 VDD.n9166 0.00194557
R20519 VDD.n10951 VDD.n10950 0.00194557
R20520 VDD.n9224 VDD.n9223 0.00194557
R20521 VDD.n10966 VDD.n9206 0.00194557
R20522 VDD.n10978 VDD.n9206 0.00194557
R20523 VDD.n9210 VDD.n9200 0.00194557
R20524 VDD.n10978 VDD.n9200 0.00194557
R20525 VDD.n10999 VDD.n10998 0.00194557
R20526 VDD.n10986 VDD.n9068 0.00194557
R20527 VDD.n10996 VDD.n10986 0.00194557
R20528 VDD.n10995 VDD.n10994 0.00194557
R20529 VDD.n10996 VDD.n10995 0.00194557
R20530 VDD.n8735 VDD.n8733 0.00194557
R20531 VDD.n10996 VDD.n8733 0.00194557
R20532 VDD.n10163 VDD.n10161 0.00194557
R20533 VDD.n10421 VDD.n10160 0.00194557
R20534 VDD.n10436 VDD.n10433 0.00194557
R20535 VDD.n10446 VDD.n6922 0.00194557
R20536 VDD.n12421 VDD.n6922 0.00194557
R20537 VDD.n10449 VDD.n6914 0.00194557
R20538 VDD.n12421 VDD.n6914 0.00194557
R20539 VDD.n8744 VDD.n8743 0.00186232
R20540 VDD.n10900 VDD.n10899 0.00176344
R20541 VDD.n10474 VDD.n10451 0.00167925
R20542 VDD.n10461 VDD.n10454 0.00167925
R20543 VDD.n10484 VDD.n10443 0.00167925
R20544 VDD.n10476 VDD.n10475 0.00167925
R20545 VDD.n10462 VDD.n10452 0.00167925
R20546 VDD.n10483 VDD.n10444 0.00167925
R20547 VDD.n5706 VDD.n5705 0.00145339
R20548 VDD.n4066 VDD.n4065 0.00145339
R20549 VDD.n2425 VDD.n2424 0.00145339
R20550 VDD.n10658 VDD.n9984 0.00145036
R20551 VDD.n10656 VDD.n9984 0.00145036
R20552 VDD.n9996 VDD.n9995 0.00143078
R20553 VDD.n9995 VDD.n6569 0.00143078
R20554 VDD.n9889 VDD.n9458 0.00141098
R20555 VDD.n9889 VDD.n9888 0.00141098
R20556 VDD.n11009 VDD.n8746 0.0014058
R20557 VDD.n9886 VDD.n9456 0.00139311
R20558 VDD.n9469 VDD.n9456 0.00139311
R20559 VDD.n9170 VDD.n7736 0.00137395
R20560 VDD.n9167 VDD.n7736 0.00137395
R20561 VDD.n10978 VDD.n9203 0.00137395
R20562 VDD.n10978 VDD.n9202 0.00137395
R20563 VDD.n10997 VDD.n10996 0.00137395
R20564 VDD.n12421 VDD.n6917 0.00137395
R20565 VDD.n12421 VDD.n6916 0.00137395
R20566 VDD.n10903 VDD.n9450 0.00136393
R20567 VDD.n9247 VDD.n9246 0.00136393
R20568 VDD.n9903 VDD.n9450 0.00136393
R20569 VDD.n9246 VDD.n9243 0.00136393
R20570 VDD.n10662 VDD.n10660 0.00134811
R20571 VDD.n9347 VDD.n9244 0.00134811
R20572 VDD.n10905 VDD.n9244 0.00134811
R20573 VDD.n10901 VDD.n10660 0.00134811
R20574 VDD.n11007 VDD.n11006 0.00128125
R20575 VDD.n11019 VDD.n11013 0.00128125
R20576 VDD.n11013 VDD.n8739 0.00128125
R20577 VDD.n10937 VDD.n10936 0.00125806
R20578 VDD.n10575 VDD.n9993 0.00125806
R20579 VDD.n10652 VDD.n10651 0.00119582
R20580 VDD.n10651 VDD.n9996 0.00119582
R20581 VDD.n6560 VDD.n5772 0.00119132
R20582 VDD.n4920 VDD.n4132 0.00119132
R20583 VDD.n3280 VDD.n2492 0.00119132
R20584 VDD.n1639 VDD.n1638 0.00119132
R20585 VDD.n9475 VDD.n9474 0.0011787
R20586 VDD.n9475 VDD.n9469 0.0011787
R20587 VDD.n6608 VDD.n6571 0.00117707
R20588 VDD.n10656 VDD.n10655 0.00117624
R20589 VDD.n10655 VDD.n10654 0.00117624
R20590 VDD.n9888 VDD.n9459 0.00116083
R20591 VDD.n9470 VDD.n9459 0.00116083
R20592 VDD.n10662 VDD.n9900 0.00115824
R20593 VDD.n9346 VDD.n9229 0.00115824
R20594 VDD.n9347 VDD.n9346 0.00115824
R20595 VDD.n10663 VDD.n9900 0.00115824
R20596 VDD.n9903 VDD.n9902 0.00114242
R20597 VDD.n10943 VDD.n9237 0.00114242
R20598 VDD.n9247 VDD.n9237 0.00114242
R20599 VDD.n9902 VDD.n9899 0.00114242
R20600 VDD.n5774 VDD.n5708 0.00112276
R20601 VDD.n4134 VDD.n4068 0.00112276
R20602 VDD.n2494 VDD.n2427 0.00112276
R20603 VDD.n787 VDD.n786 0.00112276
R20604 VDD.n10977 VDD.n9207 0.00105433
R20605 VDD.n10985 VDD.n10984 0.00104275
R20606 VDD.n10977 VDD.n10976 0.00104275
R20607 VDD.n12421 VDD.n12420 0.00103737
R20608 VDD.n5707 VDD.n4922 0.00103419
R20609 VDD.n4067 VDD.n3282 0.00103419
R20610 VDD.n2426 VDD.n1641 0.00103419
R20611 VDD.n785 VDD.n783 0.00103419
R20612 VDD.n10985 VDD.n9072 0.00101611
R20613 VDD.n10480 VDD.n6915 0.00101576
R20614 VDD.n9204 VDD.n9198 0.00101522
R20615 VDD.n10428 VDD.n6919 0.00100772
R20616 VDD.n12420 VDD.n12419 0.00100538
R20617 VDD.n10124 VDD.n9991 0.00100538
R20618 VDD.n10991 VDD.n9071 0.00100409
R20619 VDD.n10963 VDD.n9201 0.00100409
R20620 VDD.n10423 VDD.n6918 0.00100372
R20621 VDD.n9193 VDD.n9192 0.00100292
R20622 VDD.n9192 VDD.n9191 0.00100251
R20623 VDD.n10961 VDD.n9201 0.00100251
R20624 VDD.n10989 VDD.n9071 0.00100251
R20625 VDD.n12421 VDD.n6915 0.00100095
R20626 VDD.n10978 VDD.n9204 0.00100089
R20627 VDD.n6701 VDD.n6700 0.00100055
R20628 VDD.n5704 VDD.n4923 0.00100041
R20629 VDD.n4064 VDD.n3283 0.00100041
R20630 VDD.n2423 VDD.n1642 0.00100041
R20631 VDD.n781 VDD.n410 0.00100041
R20632 VDD.n5707 VDD.n5706 0.00100036
R20633 VDD.n4067 VDD.n4066 0.00100036
R20634 VDD.n2426 VDD.n2425 0.00100036
R20635 VDD.n785 VDD.n784 0.00100036
R20636 VDD.n12421 VDD.n6919 0.00100024
R20637 VDD.n12773 VDD.n6573 0.00100002
R20638 VDD.n12421 VDD.n6918 0.001
R20639 VDD.n9192 VDD.n7736 0.001
R20640 VDD.n10978 VDD.n9201 0.001
R20641 VDD.n10978 VDD.n10977 0.001
R20642 VDD.n10996 VDD.n10985 0.001
R20643 VDD.n10996 VDD.n9071 0.001
R20644 VDD.n12776 VDD.n12775 0.000855023
R20645 VDD.n12776 VDD.n6571 0.000855023
R20646 VDD.n6561 VDD.n5708 0.000855023
R20647 VDD.n6561 VDD.n6560 0.000855023
R20648 VDD.n4921 VDD.n4068 0.000855023
R20649 VDD.n4921 VDD.n4920 0.000855023
R20650 VDD.n3281 VDD.n2427 0.000855023
R20651 VDD.n3281 VDD.n3280 0.000855023
R20652 VDD.n1640 VDD.n787 0.000855023
R20653 VDD.n1640 VDD.n1639 0.000855023
R20654 VDD.n12775 VDD.n12774 0.000855004
R20655 VDD.n10473 VDD.n10442 0.00079375
R20656 VDD.n10973 VDD.n9207 0.000554326
R20657 VDD.n10976 VDD.n10975 0.000542748
R20658 VDD.n10980 VDD.n10979 0.000542748
R20659 VDD.n10979 VDD.n10978 0.000542748
R20660 VDD.n10984 VDD.n10983 0.000542748
R20661 VDD.n9195 VDD.n9194 0.000542748
R20662 VDD.n9194 VDD.n7736 0.000542748
R20663 VDD.n12771 VDD.n6577 0.000542748
R20664 VDD.n6632 VDD.n6621 0.000542748
R20665 VDD.n12693 VDD.n6621 0.000542748
R20666 VDD.n12419 VDD.n12418 0.000542748
R20667 VDD.n12421 VDD.n6921 0.000542748
R20668 VDD.n10427 VDD.n6921 0.000542748
R20669 VDD.n9173 VDD.n7736 0.000523923
R20670 VDD.n10996 VDD.n8732 0.000523923
R20671 VDD.n8734 VDD.n8732 0.000523923
R20672 VDD.n9180 VDD.n9173 0.000523923
R20673 VDD.n10480 VDD.n10447 0.000516711
R20674 VDD.n9198 VDD.n9197 0.000516107
R20675 VDD.n10982 VDD.n9072 0.000516107
R20676 VDD.n10429 VDD.n10428 0.000507966
R20677 VDD.n10964 VDD.n10963 0.000504095
R20678 VDD.n10992 VDD.n10991 0.000504095
R20679 VDD.n10424 VDD.n10423 0.000503718
R20680 VDD.n9193 VDD.n9075 0.000502918
R20681 VDD.n9177 VDD.n9073 0.000502851
R20682 VDD.n9196 VDD.n9073 0.000502851
R20683 VDD.n9191 VDD.n9190 0.000502515
R20684 VDD.n10962 VDD.n10961 0.000502515
R20685 VDD.n10990 VDD.n10989 0.000502515
R20686 VDD.n6700 VDD.n6699 0.000501859
R20687 VDD.n9179 VDD.n9178 0.000501425
R20688 VDD.n9178 VDD.n9177 0.000501425
R20689 VDD.n6559 VDD.n6558 0.000500887
R20690 VDD.n6558 VDD.n6557 0.000500887
R20691 VDD.n5704 VDD.n5703 0.000500887
R20692 VDD.n4919 VDD.n4918 0.000500887
R20693 VDD.n4918 VDD.n4917 0.000500887
R20694 VDD.n4064 VDD.n4063 0.000500887
R20695 VDD.n3279 VDD.n3278 0.000500887
R20696 VDD.n3278 VDD.n3277 0.000500887
R20697 VDD.n2423 VDD.n2422 0.000500887
R20698 VDD.n1227 VDD.n856 0.000500887
R20699 VDD.n1227 VDD.n1226 0.000500887
R20700 VDD.n781 VDD.n780 0.000500887
R20701 VDD.n5705 VDD.n4922 0.000500755
R20702 VDD.n4065 VDD.n3282 0.000500755
R20703 VDD.n2424 VDD.n1641 0.000500755
R20704 VDD.n783 VDD.n782 0.000500755
R20705 VDD.n10326 VDD.n6924 0.000500648
R20706 VDD.t148 VDD.n6924 0.000500648
R20707 VDD.t148 VDD.n10210 0.000500648
R20708 VDD.n10210 VDD.n6576 0.000500648
R20709 VDD.n5777 VDD.n5773 0.000500446
R20710 VDD.n4137 VDD.n4133 0.000500446
R20711 VDD.n2497 VDD.n2493 0.000500446
R20712 VDD.n855 VDD.n854 0.000500446
R20713 VDD.n10974 VDD.n9208 0.000500389
R20714 VDD.n9220 VDD.n9208 0.000500389
R20715 VDD.n10981 VDD.n9074 0.000500389
R20716 VDD.n9220 VDD.n9074 0.000500389
R20717 VDD.n6013 VDD.n6012 0.000500314
R20718 VDD.n5159 VDD.n5158 0.000500314
R20719 VDD.n4373 VDD.n4372 0.000500314
R20720 VDD.n3519 VDD.n3518 0.000500314
R20721 VDD.n2733 VDD.n2732 0.000500314
R20722 VDD.n1878 VDD.n1877 0.000500314
R20723 VDD.n1610 VDD.n1609 0.000500314
R20724 VDD.n382 VDD.n381 0.000500314
R20725 VDD.n6017 VDD.n6016 0.000500201
R20726 VDD.n5163 VDD.n5162 0.000500201
R20727 VDD.n4377 VDD.n4376 0.000500201
R20728 VDD.n3523 VDD.n3522 0.000500201
R20729 VDD.n2737 VDD.n2736 0.000500201
R20730 VDD.n1882 VDD.n1881 0.000500201
R20731 VDD.n1636 VDD.n1635 0.000500201
R20732 VDD.n408 VDD.n407 0.000500201
R20733 VDD.n12773 VDD.n12772 0.000500031
R20734 EF_R2RVCE_0.comparator_0.VBN.n263 EF_R2RVCE_0.comparator_0.VBN.t2 60.2505
R20735 EF_R2RVCE_0.comparator_0.VBN.n284 EF_R2RVCE_0.comparator_0.VBN.t11 60.2505
R20736 EF_R2RVCE_0.comparator_0.VBN.n304 EF_R2RVCE_0.comparator_0.VBN.t10 60.2505
R20737 EF_R2RVCE_0.comparator_0.VBN.n306 EF_R2RVCE_0.comparator_0.VBN.t12 60.2505
R20738 EF_R2RVCE_0.comparator_0.VBN.n318 EF_R2RVCE_0.comparator_0.VBN.t9 60.2505
R20739 EF_R2RVCE_0.comparator_0.VBN.n97 EF_R2RVCE_0.comparator_0.VBN.n95 41.8847
R20740 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.t1 35.1154
R20741 EF_R2RVCE_0.comparator_0.VBN.n105 EF_R2RVCE_0.comparator_0.VBN.n102 26.3366
R20742 EF_R2RVCE_0.comparator_0.VBN.n52 EF_R2RVCE_0.comparator_0.VBN.n51 26.3366
R20743 EF_R2RVCE_0.comparator_0.VBN.n38 EF_R2RVCE_0.comparator_0.VBN.n35 26.3366
R20744 EF_R2RVCE_0.comparator_0.VBN.n97 EF_R2RVCE_0.comparator_0.VBN.n96 15.9528
R20745 EF_R2RVCE_0.comparator_0.VBN.n44 EF_R2RVCE_0.comparator_0.VBN.n42 12.8005
R20746 EF_R2RVCE_0.comparator_0.VBN.n44 EF_R2RVCE_0.comparator_0.VBN.n43 12.8005
R20747 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n267 9.3005
R20748 EF_R2RVCE_0.comparator_0.VBN.n273 EF_R2RVCE_0.comparator_0.VBN.n272 9.3005
R20749 EF_R2RVCE_0.comparator_0.VBN.n282 EF_R2RVCE_0.comparator_0.VBN.n281 9.3005
R20750 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n276 9.3005
R20751 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n287 9.3005
R20752 EF_R2RVCE_0.comparator_0.VBN.n302 EF_R2RVCE_0.comparator_0.VBN.n301 9.3005
R20753 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n296 9.3005
R20754 EF_R2RVCE_0.comparator_0.VBN.n293 EF_R2RVCE_0.comparator_0.VBN.n292 9.3005
R20755 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.n23 9.3005
R20756 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.n31 9.3005
R20757 EF_R2RVCE_0.comparator_0.VBN.n11 EF_R2RVCE_0.comparator_0.VBN.n40 9.3005
R20758 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n46 9.3005
R20759 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n55 9.3005
R20760 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n63 9.3005
R20761 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n71 9.3005
R20762 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n79 9.3005
R20763 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n87 9.3005
R20764 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n86 9.3005
R20765 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n85 9.3005
R20766 EF_R2RVCE_0.comparator_0.VBN.n85 EF_R2RVCE_0.comparator_0.VBN.n84 9.3005
R20767 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n78 9.3005
R20768 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n77 9.3005
R20769 EF_R2RVCE_0.comparator_0.VBN.n77 EF_R2RVCE_0.comparator_0.VBN.n76 9.3005
R20770 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n70 9.3005
R20771 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n69 9.3005
R20772 EF_R2RVCE_0.comparator_0.VBN.n69 EF_R2RVCE_0.comparator_0.VBN.n68 9.3005
R20773 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n62 9.3005
R20774 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n61 9.3005
R20775 EF_R2RVCE_0.comparator_0.VBN.n61 EF_R2RVCE_0.comparator_0.VBN.n60 9.3005
R20776 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n54 9.3005
R20777 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n53 9.3005
R20778 EF_R2RVCE_0.comparator_0.VBN.n53 EF_R2RVCE_0.comparator_0.VBN.n52 9.3005
R20779 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n45 9.3005
R20780 EF_R2RVCE_0.comparator_0.VBN.n11 EF_R2RVCE_0.comparator_0.VBN.n41 9.3005
R20781 EF_R2RVCE_0.comparator_0.VBN.n11 EF_R2RVCE_0.comparator_0.VBN.n39 9.3005
R20782 EF_R2RVCE_0.comparator_0.VBN.n39 EF_R2RVCE_0.comparator_0.VBN.n38 9.3005
R20783 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.n32 9.3005
R20784 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.n30 9.3005
R20785 EF_R2RVCE_0.comparator_0.VBN.n30 EF_R2RVCE_0.comparator_0.VBN.n29 9.3005
R20786 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.n24 9.3005
R20787 EF_R2RVCE_0.comparator_0.VBN.n14 EF_R2RVCE_0.comparator_0.VBN.n22 9.3005
R20788 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n155 9.3005
R20789 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n147 9.3005
R20790 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n139 9.3005
R20791 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n131 9.3005
R20792 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n123 9.3005
R20793 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n115 9.3005
R20794 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n107 9.3005
R20795 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n98 9.3005
R20796 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n106 9.3005
R20797 EF_R2RVCE_0.comparator_0.VBN.n106 EF_R2RVCE_0.comparator_0.VBN.n105 9.3005
R20798 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n99 9.3005
R20799 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n108 9.3005
R20800 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n114 9.3005
R20801 EF_R2RVCE_0.comparator_0.VBN.n114 EF_R2RVCE_0.comparator_0.VBN.n113 9.3005
R20802 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n122 9.3005
R20803 EF_R2RVCE_0.comparator_0.VBN.n122 EF_R2RVCE_0.comparator_0.VBN.n121 9.3005
R20804 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n116 9.3005
R20805 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n124 9.3005
R20806 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n130 9.3005
R20807 EF_R2RVCE_0.comparator_0.VBN.n130 EF_R2RVCE_0.comparator_0.VBN.n129 9.3005
R20808 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n138 9.3005
R20809 EF_R2RVCE_0.comparator_0.VBN.n138 EF_R2RVCE_0.comparator_0.VBN.n137 9.3005
R20810 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n132 9.3005
R20811 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n140 9.3005
R20812 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n146 9.3005
R20813 EF_R2RVCE_0.comparator_0.VBN.n146 EF_R2RVCE_0.comparator_0.VBN.n145 9.3005
R20814 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n154 9.3005
R20815 EF_R2RVCE_0.comparator_0.VBN.n154 EF_R2RVCE_0.comparator_0.VBN.n153 9.3005
R20816 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n148 9.3005
R20817 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n156 9.3005
R20818 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n162 9.3005
R20819 EF_R2RVCE_0.comparator_0.VBN.n162 EF_R2RVCE_0.comparator_0.VBN.n161 9.3005
R20820 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n170 9.3005
R20821 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n171 9.3005
R20822 EF_R2RVCE_0.comparator_0.VBN.n177 EF_R2RVCE_0.comparator_0.VBN.n176 9.3005
R20823 EF_R2RVCE_0.comparator_0.VBN.n92 EF_R2RVCE_0.comparator_0.VBN.n91 9.3005
R20824 EF_R2RVCE_0.comparator_0.VBN.n167 EF_R2RVCE_0.comparator_0.VBN.n166 9.3005
R20825 EF_R2RVCE_0.comparator_0.VBN.n20 EF_R2RVCE_0.comparator_0.VBN.n315 9.3005
R20826 EF_R2RVCE_0.comparator_0.VBN.n20 EF_R2RVCE_0.comparator_0.VBN.n313 9.3005
R20827 EF_R2RVCE_0.comparator_0.VBN.n313 EF_R2RVCE_0.comparator_0.VBN.n312 9.3005
R20828 EF_R2RVCE_0.comparator_0.VBN.n20 EF_R2RVCE_0.comparator_0.VBN.n314 9.3005
R20829 EF_R2RVCE_0.comparator_0.VBN.n17 EF_R2RVCE_0.comparator_0.VBN.n327 9.3005
R20830 EF_R2RVCE_0.comparator_0.VBN.n17 EF_R2RVCE_0.comparator_0.VBN.n326 9.3005
R20831 EF_R2RVCE_0.comparator_0.VBN.n17 EF_R2RVCE_0.comparator_0.VBN.n325 9.3005
R20832 EF_R2RVCE_0.comparator_0.VBN.n325 EF_R2RVCE_0.comparator_0.VBN.n324 9.3005
R20833 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n246 9.3005
R20834 EF_R2RVCE_0.comparator_0.VBN.n252 EF_R2RVCE_0.comparator_0.VBN.n251 9.3005
R20835 EF_R2RVCE_0.comparator_0.VBN.n261 EF_R2RVCE_0.comparator_0.VBN.n260 9.3005
R20836 EF_R2RVCE_0.comparator_0.VBN.n18 EF_R2RVCE_0.comparator_0.VBN.n255 9.3005
R20837 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n242 9.3005
R20838 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n197 9.3005
R20839 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n192 9.3005
R20840 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n243 9.3005
R20841 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n241 9.3005
R20842 EF_R2RVCE_0.comparator_0.VBN.n285 EF_R2RVCE_0.comparator_0.VBN.n284 8.76429
R20843 EF_R2RVCE_0.comparator_0.VBN.n305 EF_R2RVCE_0.comparator_0.VBN.n304 8.76429
R20844 EF_R2RVCE_0.comparator_0.VBN.n264 EF_R2RVCE_0.comparator_0.VBN.n263 8.76429
R20845 EF_R2RVCE_0.comparator_0.VBN.n271 EF_R2RVCE_0.comparator_0.VBN.n270 8.21641
R20846 EF_R2RVCE_0.comparator_0.VBN.n280 EF_R2RVCE_0.comparator_0.VBN.n279 8.21641
R20847 EF_R2RVCE_0.comparator_0.VBN.n291 EF_R2RVCE_0.comparator_0.VBN.n290 8.21641
R20848 EF_R2RVCE_0.comparator_0.VBN.n300 EF_R2RVCE_0.comparator_0.VBN.n299 8.21641
R20849 EF_R2RVCE_0.comparator_0.VBN.n311 EF_R2RVCE_0.comparator_0.VBN.n310 8.21641
R20850 EF_R2RVCE_0.comparator_0.VBN.n323 EF_R2RVCE_0.comparator_0.VBN.n322 8.21641
R20851 EF_R2RVCE_0.comparator_0.VBN.n250 EF_R2RVCE_0.comparator_0.VBN.n249 8.21641
R20852 EF_R2RVCE_0.comparator_0.VBN.n259 EF_R2RVCE_0.comparator_0.VBN.n258 8.21641
R20853 EF_R2RVCE_0.comparator_0.VBN.n160 EF_R2RVCE_0.comparator_0.VBN.n159 7.95102
R20854 EF_R2RVCE_0.comparator_0.VBN.n165 EF_R2RVCE_0.comparator_0.VBN.n164 7.95102
R20855 EF_R2RVCE_0.comparator_0.VBN.n105 EF_R2RVCE_0.comparator_0.VBN.n104 7.45411
R20856 EF_R2RVCE_0.comparator_0.VBN.n52 EF_R2RVCE_0.comparator_0.VBN.n50 7.45411
R20857 EF_R2RVCE_0.comparator_0.VBN.n38 EF_R2RVCE_0.comparator_0.VBN.n37 7.45411
R20858 EF_R2RVCE_0.comparator_0.VBN.n152 EF_R2RVCE_0.comparator_0.VBN.n151 6.9572
R20859 EF_R2RVCE_0.comparator_0.VBN.n175 EF_R2RVCE_0.comparator_0.VBN.n174 6.9572
R20860 EF_R2RVCE_0.comparator_0.VBN.n319 EF_R2RVCE_0.comparator_0.VBN.n318 6.92242
R20861 EF_R2RVCE_0.comparator_0.VBN.n307 EF_R2RVCE_0.comparator_0.VBN.n306 6.92012
R20862 EF_R2RVCE_0.comparator_0.VBN.n113 EF_R2RVCE_0.comparator_0.VBN.n112 6.46029
R20863 EF_R2RVCE_0.comparator_0.VBN.n60 EF_R2RVCE_0.comparator_0.VBN.n59 6.46029
R20864 EF_R2RVCE_0.comparator_0.VBN.n29 EF_R2RVCE_0.comparator_0.VBN.n28 6.46029
R20865 EF_R2RVCE_0.comparator_0.VBN.n158 EF_R2RVCE_0.comparator_0.VBN.n157 6.02403
R20866 EF_R2RVCE_0.comparator_0.VBN.n144 EF_R2RVCE_0.comparator_0.VBN.n143 5.96339
R20867 EF_R2RVCE_0.comparator_0.VBN.n90 EF_R2RVCE_0.comparator_0.VBN.n89 5.96339
R20868 EF_R2RVCE_0.comparator_0.VBN.n269 EF_R2RVCE_0.comparator_0.VBN.n268 5.64756
R20869 EF_R2RVCE_0.comparator_0.VBN.n278 EF_R2RVCE_0.comparator_0.VBN.n277 5.64756
R20870 EF_R2RVCE_0.comparator_0.VBN.n289 EF_R2RVCE_0.comparator_0.VBN.n288 5.64756
R20871 EF_R2RVCE_0.comparator_0.VBN.n298 EF_R2RVCE_0.comparator_0.VBN.n297 5.64756
R20872 EF_R2RVCE_0.comparator_0.VBN.n106 EF_R2RVCE_0.comparator_0.VBN.n101 5.64756
R20873 EF_R2RVCE_0.comparator_0.VBN.n53 EF_R2RVCE_0.comparator_0.VBN.n48 5.64756
R20874 EF_R2RVCE_0.comparator_0.VBN.n39 EF_R2RVCE_0.comparator_0.VBN.n34 5.64756
R20875 EF_R2RVCE_0.comparator_0.VBN.n309 EF_R2RVCE_0.comparator_0.VBN.n308 5.64756
R20876 EF_R2RVCE_0.comparator_0.VBN.n321 EF_R2RVCE_0.comparator_0.VBN.n320 5.64756
R20877 EF_R2RVCE_0.comparator_0.VBN.n248 EF_R2RVCE_0.comparator_0.VBN.n247 5.64756
R20878 EF_R2RVCE_0.comparator_0.VBN.n257 EF_R2RVCE_0.comparator_0.VBN.n256 5.64756
R20879 EF_R2RVCE_0.comparator_0.VBN.n225 EF_R2RVCE_0.comparator_0.VBN.t8 5.5395
R20880 EF_R2RVCE_0.comparator_0.VBN.n225 EF_R2RVCE_0.comparator_0.VBN.t5 5.5395
R20881 EF_R2RVCE_0.comparator_0.VBN.n210 EF_R2RVCE_0.comparator_0.VBN.t6 5.5395
R20882 EF_R2RVCE_0.comparator_0.VBN.n210 EF_R2RVCE_0.comparator_0.VBN.t7 5.5395
R20883 EF_R2RVCE_0.comparator_0.VBN.n121 EF_R2RVCE_0.comparator_0.VBN.n120 5.46648
R20884 EF_R2RVCE_0.comparator_0.VBN.n68 EF_R2RVCE_0.comparator_0.VBN.n67 5.46648
R20885 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n244 5.28613
R20886 EF_R2RVCE_0.comparator_0.VBN.n150 EF_R2RVCE_0.comparator_0.VBN.n149 5.27109
R20887 EF_R2RVCE_0.comparator_0.VBN.n136 EF_R2RVCE_0.comparator_0.VBN.n135 4.96957
R20888 EF_R2RVCE_0.comparator_0.VBN.n83 EF_R2RVCE_0.comparator_0.VBN.n82 4.96957
R20889 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n266 4.911
R20890 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n286 4.911
R20891 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n275 4.91005
R20892 EF_R2RVCE_0.comparator_0.VBN.n18 EF_R2RVCE_0.comparator_0.VBN.n254 4.91005
R20893 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n295 4.90905
R20894 EF_R2RVCE_0.comparator_0.VBN.n114 EF_R2RVCE_0.comparator_0.VBN.n110 4.89462
R20895 EF_R2RVCE_0.comparator_0.VBN.n61 EF_R2RVCE_0.comparator_0.VBN.n57 4.89462
R20896 EF_R2RVCE_0.comparator_0.VBN.n30 EF_R2RVCE_0.comparator_0.VBN.n26 4.89462
R20897 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n245 4.76425
R20898 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n44 4.6505
R20899 EF_R2RVCE_0.comparator_0.VBN.n219 EF_R2RVCE_0.comparator_0.VBN.n218 4.51815
R20900 EF_R2RVCE_0.comparator_0.VBN.n206 EF_R2RVCE_0.comparator_0.VBN.n205 4.51815
R20901 EF_R2RVCE_0.comparator_0.VBN.n142 EF_R2RVCE_0.comparator_0.VBN.n141 4.51815
R20902 EF_R2RVCE_0.comparator_0.VBN.n169 EF_R2RVCE_0.comparator_0.VBN.n163 4.51815
R20903 EF_R2RVCE_0.comparator_0.VBN.n195 EF_R2RVCE_0.comparator_0.VBN.n194 4.51815
R20904 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n232 4.5005
R20905 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n200 4.5005
R20906 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n224 4.5005
R20907 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n222 4.5005
R20908 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n229 4.5005
R20909 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n216 4.5005
R20910 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n204 4.5005
R20911 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n236 4.5005
R20912 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n213 4.5005
R20913 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n209 4.5005
R20914 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n94 4.5005
R20915 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n182 4.5005
R20916 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n179 4.5005
R20917 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n169 4.5005
R20918 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n274 4.5005
R20919 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n283 4.5005
R20920 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n303 4.5005
R20921 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n294 4.5005
R20922 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n253 4.5005
R20923 EF_R2RVCE_0.comparator_0.VBN.n18 EF_R2RVCE_0.comparator_0.VBN.n262 4.5005
R20924 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n195 4.5005
R20925 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n188 4.5005
R20926 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n190 4.5005
R20927 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n239 4.5005
R20928 EF_R2RVCE_0.comparator_0.VBN.n129 EF_R2RVCE_0.comparator_0.VBN.n128 4.47267
R20929 EF_R2RVCE_0.comparator_0.VBN.n76 EF_R2RVCE_0.comparator_0.VBN.n75 4.47267
R20930 EF_R2RVCE_0.comparator_0.VBN.n21 EF_R2RVCE_0.comparator_0.VBN.n7 4.44875
R20931 EF_R2RVCE_0.comparator_0.VBN.n7 EF_R2RVCE_0.comparator_0.VBN.n316 7.3305
R20932 EF_R2RVCE_0.comparator_0.VBN.n17 EF_R2RVCE_0.comparator_0.VBN.n329 4.24504
R20933 EF_R2RVCE_0.comparator_0.VBN.n122 EF_R2RVCE_0.comparator_0.VBN.n118 4.14168
R20934 EF_R2RVCE_0.comparator_0.VBN.n69 EF_R2RVCE_0.comparator_0.VBN.n65 4.14168
R20935 EF_R2RVCE_0.comparator_0.VBN.n128 EF_R2RVCE_0.comparator_0.VBN.n127 3.97576
R20936 EF_R2RVCE_0.comparator_0.VBN.n75 EF_R2RVCE_0.comparator_0.VBN.n74 3.97576
R20937 EF_R2RVCE_0.comparator_0.VBN.n134 EF_R2RVCE_0.comparator_0.VBN.n133 3.76521
R20938 EF_R2RVCE_0.comparator_0.VBN.n179 EF_R2RVCE_0.comparator_0.VBN.n173 3.76521
R20939 EF_R2RVCE_0.comparator_0.VBN.n182 EF_R2RVCE_0.comparator_0.VBN.n180 3.76521
R20940 EF_R2RVCE_0.comparator_0.VBN.n81 EF_R2RVCE_0.comparator_0.VBN.n80 3.76521
R20941 EF_R2RVCE_0.comparator_0.VBN.n239 EF_R2RVCE_0.comparator_0.VBN.n238 3.76521
R20942 EF_R2RVCE_0.comparator_0.VBN.n137 EF_R2RVCE_0.comparator_0.VBN.n136 3.47885
R20943 EF_R2RVCE_0.comparator_0.VBN.n84 EF_R2RVCE_0.comparator_0.VBN.n83 3.47885
R20944 EF_R2RVCE_0.comparator_0.VBN.n20 EF_R2RVCE_0.comparator_0.VBN.n307 3.47756
R20945 EF_R2RVCE_0.comparator_0.VBN.n17 EF_R2RVCE_0.comparator_0.VBN.n319 3.4767
R20946 EF_R2RVCE_0.comparator_0.VBN.n130 EF_R2RVCE_0.comparator_0.VBN.n126 3.38874
R20947 EF_R2RVCE_0.comparator_0.VBN.n77 EF_R2RVCE_0.comparator_0.VBN.n73 3.38874
R20948 EF_R2RVCE_0.comparator_0.VBN.n184 EF_R2RVCE_0.comparator_0.VBN.t4 3.3065
R20949 EF_R2RVCE_0.comparator_0.VBN.n184 EF_R2RVCE_0.comparator_0.VBN.t3 3.3065
R20950 EF_R2RVCE_0.comparator_0.VBN.n188 EF_R2RVCE_0.comparator_0.VBN.n186 3.74814
R20951 EF_R2RVCE_0.comparator_0.VBN.n15 EF_R2RVCE_0.comparator_0.VBN.n185 3.15814
R20952 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n219 3.03311
R20953 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n206 3.03311
R20954 EF_R2RVCE_0.comparator_0.VBN.n3 EF_R2RVCE_0.comparator_0.VBN.n285 3.03311
R20955 EF_R2RVCE_0.comparator_0.VBN.n2 EF_R2RVCE_0.comparator_0.VBN.n305 3.03311
R20956 EF_R2RVCE_0.comparator_0.VBN.n18 EF_R2RVCE_0.comparator_0.VBN.n264 3.03311
R20957 EF_R2RVCE_0.comparator_0.VBN.n126 EF_R2RVCE_0.comparator_0.VBN.n125 3.01226
R20958 EF_R2RVCE_0.comparator_0.VBN.n94 EF_R2RVCE_0.comparator_0.VBN.n88 3.01226
R20959 EF_R2RVCE_0.comparator_0.VBN.n73 EF_R2RVCE_0.comparator_0.VBN.n72 3.01226
R20960 EF_R2RVCE_0.comparator_0.VBN.n188 EF_R2RVCE_0.comparator_0.VBN.n187 3.01226
R20961 EF_R2RVCE_0.comparator_0.VBN.n120 EF_R2RVCE_0.comparator_0.VBN.n119 2.98194
R20962 EF_R2RVCE_0.comparator_0.VBN.n67 EF_R2RVCE_0.comparator_0.VBN.n66 2.98194
R20963 EF_R2RVCE_0.comparator_0.VBN.n236 EF_R2RVCE_0.comparator_0.VBN.n234 2.63579
R20964 EF_R2RVCE_0.comparator_0.VBN.n204 EF_R2RVCE_0.comparator_0.VBN.n202 2.63579
R20965 EF_R2RVCE_0.comparator_0.VBN.n138 EF_R2RVCE_0.comparator_0.VBN.n134 2.63579
R20966 EF_R2RVCE_0.comparator_0.VBN.n85 EF_R2RVCE_0.comparator_0.VBN.n81 2.63579
R20967 EF_R2RVCE_0.comparator_0.VBN.n239 EF_R2RVCE_0.comparator_0.VBN.n237 2.63579
R20968 EF_R2RVCE_0.comparator_0.VBN.n192 EF_R2RVCE_0.comparator_0.VBN.n191 2.61733
R20969 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n198 2.60826
R20970 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n230 2.60826
R20971 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n183 2.53421
R20972 EF_R2RVCE_0.comparator_0.VBN.n145 EF_R2RVCE_0.comparator_0.VBN.n144 2.48504
R20973 EF_R2RVCE_0.comparator_0.VBN.n91 EF_R2RVCE_0.comparator_0.VBN.n90 2.48504
R20974 EF_R2RVCE_0.comparator_0.VBN.n7 EF_R2RVCE_0.comparator_0.VBN.n17 2.42663
R20975 EF_R2RVCE_0.comparator_0.VBN.n7 EF_R2RVCE_0.comparator_0.VBN.n20 2.39724
R20976 EF_R2RVCE_0.comparator_0.VBN.n229 EF_R2RVCE_0.comparator_0.VBN.n227 2.25932
R20977 EF_R2RVCE_0.comparator_0.VBN.n221 EF_R2RVCE_0.comparator_0.VBN.n220 2.25932
R20978 EF_R2RVCE_0.comparator_0.VBN.n216 EF_R2RVCE_0.comparator_0.VBN.n214 2.25932
R20979 EF_R2RVCE_0.comparator_0.VBN.n208 EF_R2RVCE_0.comparator_0.VBN.n207 2.25932
R20980 EF_R2RVCE_0.comparator_0.VBN.n118 EF_R2RVCE_0.comparator_0.VBN.n117 2.25932
R20981 EF_R2RVCE_0.comparator_0.VBN.n65 EF_R2RVCE_0.comparator_0.VBN.n64 2.25932
R20982 EF_R2RVCE_0.comparator_0.VBN.n229 EF_R2RVCE_0.comparator_0.VBN.n228 2.25379
R20983 EF_R2RVCE_0.comparator_0.VBN.n216 EF_R2RVCE_0.comparator_0.VBN.n215 2.25379
R20984 EF_R2RVCE_0.comparator_0.VBN.n7 EF_R2RVCE_0.comparator_0.VBN.n317 2.2505
R20985 EF_R2RVCE_0.comparator_0.VBN.n197 EF_R2RVCE_0.comparator_0.VBN.n196 2.24766
R20986 EF_R2RVCE_0.comparator_0.VBN.n265 EF_R2RVCE_0.comparator_0.VBN.n18 2.073
R20987 EF_R2RVCE_0.comparator_0.VBN EF_R2RVCE_0.comparator_0.VBN.n19 2.06925
R20988 EF_R2RVCE_0.comparator_0.VBN.n112 EF_R2RVCE_0.comparator_0.VBN.n111 1.98813
R20989 EF_R2RVCE_0.comparator_0.VBN.n59 EF_R2RVCE_0.comparator_0.VBN.n58 1.98813
R20990 EF_R2RVCE_0.comparator_0.VBN.n28 EF_R2RVCE_0.comparator_0.VBN.n27 1.98813
R20991 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n172 1.94045
R20992 EF_R2RVCE_0.comparator_0.VBN.n146 EF_R2RVCE_0.comparator_0.VBN.n142 1.88285
R20993 EF_R2RVCE_0.comparator_0.VBN.n93 EF_R2RVCE_0.comparator_0.VBN.n92 1.88285
R20994 EF_R2RVCE_0.comparator_0.VBN.n195 EF_R2RVCE_0.comparator_0.VBN.n193 1.88285
R20995 EF_R2RVCE_0.comparator_0.VBN.n236 EF_R2RVCE_0.comparator_0.VBN.n235 1.87949
R20996 EF_R2RVCE_0.comparator_0.VBN.n204 EF_R2RVCE_0.comparator_0.VBN.n203 1.87949
R20997 EF_R2RVCE_0.comparator_0.VBN.n265 EF_R2RVCE_0.comparator_0.VBN.n3 1.85011
R20998 EF_R2RVCE_0.comparator_0.VBN.n217 EF_R2RVCE_0.comparator_0.VBN.n1 1.73899
R20999 EF_R2RVCE_0.comparator_0.VBN.n21 EF_R2RVCE_0.comparator_0.VBN.n172 1.70776
R21000 EF_R2RVCE_0.comparator_0.VBN.n19 EF_R2RVCE_0.comparator_0.VBN.n2 1.70567
R21001 EF_R2RVCE_0.comparator_0.VBN.n15 EF_R2RVCE_0.comparator_0.VBN.n184 1.61775
R21002 EF_R2RVCE_0.comparator_0.VBN.n95 EF_R2RVCE_0.comparator_0.VBN.t0 1.60717
R21003 EF_R2RVCE_0.comparator_0.VBN.n7 EF_R2RVCE_0.comparator_0.VBN 1.60425
R21004 EF_R2RVCE_0.comparator_0.VBN.n224 EF_R2RVCE_0.comparator_0.VBN.n223 1.50638
R21005 EF_R2RVCE_0.comparator_0.VBN.n213 EF_R2RVCE_0.comparator_0.VBN.n212 1.50638
R21006 EF_R2RVCE_0.comparator_0.VBN.n110 EF_R2RVCE_0.comparator_0.VBN.n109 1.50638
R21007 EF_R2RVCE_0.comparator_0.VBN.n169 EF_R2RVCE_0.comparator_0.VBN.n168 1.50638
R21008 EF_R2RVCE_0.comparator_0.VBN.n179 EF_R2RVCE_0.comparator_0.VBN.n178 1.50638
R21009 EF_R2RVCE_0.comparator_0.VBN.n94 EF_R2RVCE_0.comparator_0.VBN.n93 1.50638
R21010 EF_R2RVCE_0.comparator_0.VBN.n57 EF_R2RVCE_0.comparator_0.VBN.n56 1.50638
R21011 EF_R2RVCE_0.comparator_0.VBN.n26 EF_R2RVCE_0.comparator_0.VBN.n25 1.50638
R21012 EF_R2RVCE_0.comparator_0.VBN.n226 EF_R2RVCE_0.comparator_0.VBN.n225 1.50151
R21013 EF_R2RVCE_0.comparator_0.VBN.n211 EF_R2RVCE_0.comparator_0.VBN.n210 1.50148
R21014 EF_R2RVCE_0.comparator_0.VBN.n153 EF_R2RVCE_0.comparator_0.VBN.n152 1.49122
R21015 EF_R2RVCE_0.comparator_0.VBN.n176 EF_R2RVCE_0.comparator_0.VBN.n175 1.49122
R21016 EF_R2RVCE_0.comparator_0.VBN.n19 EF_R2RVCE_0.comparator_0.VBN.n265 1.26925
R21017 EF_R2RVCE_0.comparator_0.VBN.n217 EF_R2RVCE_0.comparator_0.VBN.n0 1.19668
R21018 EF_R2RVCE_0.comparator_0.VBN.n19 EF_R2RVCE_0.comparator_0.VBN.n21 1.1545
R21019 EF_R2RVCE_0.comparator_0.VBN.n154 EF_R2RVCE_0.comparator_0.VBN.n150 1.12991
R21020 EF_R2RVCE_0.comparator_0.VBN.n178 EF_R2RVCE_0.comparator_0.VBN.n177 1.12991
R21021 EF_R2RVCE_0.comparator_0.VBN.n190 EF_R2RVCE_0.comparator_0.VBN.n189 1.12991
R21022 EF_R2RVCE_0.comparator_0.VBN.n272 EF_R2RVCE_0.comparator_0.VBN.n271 1.09595
R21023 EF_R2RVCE_0.comparator_0.VBN.n281 EF_R2RVCE_0.comparator_0.VBN.n280 1.09595
R21024 EF_R2RVCE_0.comparator_0.VBN.n292 EF_R2RVCE_0.comparator_0.VBN.n291 1.09595
R21025 EF_R2RVCE_0.comparator_0.VBN.n301 EF_R2RVCE_0.comparator_0.VBN.n300 1.09595
R21026 EF_R2RVCE_0.comparator_0.VBN.n312 EF_R2RVCE_0.comparator_0.VBN.n311 1.09595
R21027 EF_R2RVCE_0.comparator_0.VBN.n324 EF_R2RVCE_0.comparator_0.VBN.n323 1.09595
R21028 EF_R2RVCE_0.comparator_0.VBN.n251 EF_R2RVCE_0.comparator_0.VBN.n250 1.09595
R21029 EF_R2RVCE_0.comparator_0.VBN.n260 EF_R2RVCE_0.comparator_0.VBN.n259 1.09595
R21030 EF_R2RVCE_0.comparator_0.VBN.n13 EF_R2RVCE_0.comparator_0.VBN.n97 1.03132
R21031 EF_R2RVCE_0.comparator_0.VBN.n104 EF_R2RVCE_0.comparator_0.VBN.n103 0.994314
R21032 EF_R2RVCE_0.comparator_0.VBN.n50 EF_R2RVCE_0.comparator_0.VBN.n49 0.994314
R21033 EF_R2RVCE_0.comparator_0.VBN.n37 EF_R2RVCE_0.comparator_0.VBN.n36 0.994314
R21034 EF_R2RVCE_0.comparator_0.VBN.n183 EF_R2RVCE_0.comparator_0.VBN.n217 0.890264
R21035 EF_R2RVCE_0.comparator_0.VBN.n0 EF_R2RVCE_0.comparator_0.VBN.n226 0.833636
R21036 EF_R2RVCE_0.comparator_0.VBN.n1 EF_R2RVCE_0.comparator_0.VBN.n211 0.833623
R21037 EF_R2RVCE_0.comparator_0.VBN.n6 EF_R2RVCE_0.comparator_0.VBN.n16 0.766876
R21038 EF_R2RVCE_0.comparator_0.VBN.n232 EF_R2RVCE_0.comparator_0.VBN.n231 0.753441
R21039 EF_R2RVCE_0.comparator_0.VBN.n222 EF_R2RVCE_0.comparator_0.VBN.n221 0.753441
R21040 EF_R2RVCE_0.comparator_0.VBN.n200 EF_R2RVCE_0.comparator_0.VBN.n199 0.753441
R21041 EF_R2RVCE_0.comparator_0.VBN.n209 EF_R2RVCE_0.comparator_0.VBN.n208 0.753441
R21042 EF_R2RVCE_0.comparator_0.VBN.n274 EF_R2RVCE_0.comparator_0.VBN.n273 0.753441
R21043 EF_R2RVCE_0.comparator_0.VBN.n273 EF_R2RVCE_0.comparator_0.VBN.n269 0.753441
R21044 EF_R2RVCE_0.comparator_0.VBN.n282 EF_R2RVCE_0.comparator_0.VBN.n278 0.753441
R21045 EF_R2RVCE_0.comparator_0.VBN.n283 EF_R2RVCE_0.comparator_0.VBN.n282 0.753441
R21046 EF_R2RVCE_0.comparator_0.VBN.n294 EF_R2RVCE_0.comparator_0.VBN.n293 0.753441
R21047 EF_R2RVCE_0.comparator_0.VBN.n293 EF_R2RVCE_0.comparator_0.VBN.n289 0.753441
R21048 EF_R2RVCE_0.comparator_0.VBN.n302 EF_R2RVCE_0.comparator_0.VBN.n298 0.753441
R21049 EF_R2RVCE_0.comparator_0.VBN.n303 EF_R2RVCE_0.comparator_0.VBN.n302 0.753441
R21050 EF_R2RVCE_0.comparator_0.VBN.n101 EF_R2RVCE_0.comparator_0.VBN.n100 0.753441
R21051 EF_R2RVCE_0.comparator_0.VBN.n48 EF_R2RVCE_0.comparator_0.VBN.n47 0.753441
R21052 EF_R2RVCE_0.comparator_0.VBN.n34 EF_R2RVCE_0.comparator_0.VBN.n33 0.753441
R21053 EF_R2RVCE_0.comparator_0.VBN.n313 EF_R2RVCE_0.comparator_0.VBN.n309 0.753441
R21054 EF_R2RVCE_0.comparator_0.VBN.n325 EF_R2RVCE_0.comparator_0.VBN.n321 0.753441
R21055 EF_R2RVCE_0.comparator_0.VBN.n253 EF_R2RVCE_0.comparator_0.VBN.n252 0.753441
R21056 EF_R2RVCE_0.comparator_0.VBN.n252 EF_R2RVCE_0.comparator_0.VBN.n248 0.753441
R21057 EF_R2RVCE_0.comparator_0.VBN.n261 EF_R2RVCE_0.comparator_0.VBN.n257 0.753441
R21058 EF_R2RVCE_0.comparator_0.VBN.n262 EF_R2RVCE_0.comparator_0.VBN.n261 0.753441
R21059 EF_R2RVCE_0.comparator_0.VBN.n329 EF_R2RVCE_0.comparator_0.VBN.n328 0.738413
R21060 EF_R2RVCE_0.comparator_0.VBN.n5 EF_R2RVCE_0.comparator_0.VBN.n4 0.700653
R21061 EF_R2RVCE_0.comparator_0.VBN.n4 EF_R2RVCE_0.comparator_0.VBN.n10 0.571152
R21062 EF_R2RVCE_0.comparator_0.VBN.n18 EF_R2RVCE_0.comparator_0.VBN.n6 0.498175
R21063 EF_R2RVCE_0.comparator_0.VBN.n161 EF_R2RVCE_0.comparator_0.VBN.n160 0.497407
R21064 EF_R2RVCE_0.comparator_0.VBN.n166 EF_R2RVCE_0.comparator_0.VBN.n165 0.497407
R21065 EF_R2RVCE_0.comparator_0.VBN.n16 EF_R2RVCE_0.comparator_0.VBN.n15 0.489854
R21066 EF_R2RVCE_0.comparator_0.VBN.n241 EF_R2RVCE_0.comparator_0.VBN.n240 0.461175
R21067 EF_R2RVCE_0.comparator_0.VBN.n12 EF_R2RVCE_0.comparator_0.VBN.n11 0.42713
R21068 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n5 0.387304
R21069 EF_R2RVCE_0.comparator_0.VBN.n11 EF_R2RVCE_0.comparator_0.VBN.n14 0.380935
R21070 EF_R2RVCE_0.comparator_0.VBN.n9 EF_R2RVCE_0.comparator_0.VBN.n8 0.380935
R21071 EF_R2RVCE_0.comparator_0.VBN.n10 EF_R2RVCE_0.comparator_0.VBN.n13 0.380935
R21072 EF_R2RVCE_0.comparator_0.VBN.n8 EF_R2RVCE_0.comparator_0.VBN.n12 0.380935
R21073 EF_R2RVCE_0.comparator_0.VBN.n234 EF_R2RVCE_0.comparator_0.VBN.n233 0.376971
R21074 EF_R2RVCE_0.comparator_0.VBN.n202 EF_R2RVCE_0.comparator_0.VBN.n201 0.376971
R21075 EF_R2RVCE_0.comparator_0.VBN.n162 EF_R2RVCE_0.comparator_0.VBN.n158 0.376971
R21076 EF_R2RVCE_0.comparator_0.VBN.n168 EF_R2RVCE_0.comparator_0.VBN.n167 0.376971
R21077 EF_R2RVCE_0.comparator_0.VBN.n182 EF_R2RVCE_0.comparator_0.VBN.n181 0.376971
R21078 a_1297_2982.n76 a_1297_2982.n74 8.05594
R21079 a_1297_2982.n76 a_1297_2982.n75 8.02924
R21080 a_1297_2982.n72 a_1297_2982.n71 6.13632
R21081 a_1297_2982.n10 a_1297_2982.n66 5.61043
R21082 a_1297_2982.n8 a_1297_2982.n35 5.61041
R21083 a_1297_2982.n6 a_1297_2982.n37 5.61041
R21084 a_1297_2982.n2 a_1297_2982.n65 5.61041
R21085 a_1297_2982.n0 a_1297_2982.n17 5.61037
R21086 a_1297_2982.n4 a_1297_2982.n47 5.61037
R21087 a_1297_2982.n3 a_1297_2982.n59 4.5005
R21088 a_1297_2982.n5 a_1297_2982.n55 4.5005
R21089 a_1297_2982.n5 a_1297_2982.n51 4.5005
R21090 a_1297_2982.n3 a_1297_2982.n63 4.5005
R21091 a_1297_2982.n7 a_1297_2982.n45 4.5005
R21092 a_1297_2982.n7 a_1297_2982.n41 4.5005
R21093 a_1297_2982.n9 a_1297_2982.n29 4.5005
R21094 a_1297_2982.n1 a_1297_2982.n25 4.5005
R21095 a_1297_2982.n1 a_1297_2982.n21 4.5005
R21096 a_1297_2982.n9 a_1297_2982.n33 4.5005
R21097 a_1297_2982.n11 a_1297_2982.n68 4.5005
R21098 a_1297_2982.n11 a_1297_2982.n70 4.5005
R21099 a_1297_2982.n25 a_1297_2982.n24 3.76521
R21100 a_1297_2982.n29 a_1297_2982.n28 3.76521
R21101 a_1297_2982.n41 a_1297_2982.n40 3.76521
R21102 a_1297_2982.n55 a_1297_2982.n54 3.76521
R21103 a_1297_2982.n59 a_1297_2982.n58 3.76521
R21104 a_1297_2982.n70 a_1297_2982.n69 3.76521
R21105 a_1297_2982.n21 a_1297_2982.n19 3.38874
R21106 a_1297_2982.n33 a_1297_2982.n31 3.38874
R21107 a_1297_2982.n45 a_1297_2982.n43 3.38874
R21108 a_1297_2982.n51 a_1297_2982.n49 3.38874
R21109 a_1297_2982.n63 a_1297_2982.n61 3.38874
R21110 a_1297_2982.n22 a_1297_2982.t6 3.3065
R21111 a_1297_2982.n22 a_1297_2982.t2 3.3065
R21112 a_1297_2982.n26 a_1297_2982.t5 3.3065
R21113 a_1297_2982.n26 a_1297_2982.t4 3.3065
R21114 a_1297_2982.n38 a_1297_2982.t3 3.3065
R21115 a_1297_2982.n38 a_1297_2982.t10 3.3065
R21116 a_1297_2982.n52 a_1297_2982.t7 3.3065
R21117 a_1297_2982.n52 a_1297_2982.t8 3.3065
R21118 a_1297_2982.n56 a_1297_2982.t9 3.3065
R21119 a_1297_2982.n56 a_1297_2982.t11 3.3065
R21120 a_1297_2982.t0 a_1297_2982.n76 3.3065
R21121 a_1297_2982.n76 a_1297_2982.t1 3.3065
R21122 a_1297_2982.n21 a_1297_2982.n20 3.01226
R21123 a_1297_2982.n33 a_1297_2982.n32 3.01226
R21124 a_1297_2982.n45 a_1297_2982.n44 3.01226
R21125 a_1297_2982.n51 a_1297_2982.n50 3.01226
R21126 a_1297_2982.n63 a_1297_2982.n62 3.01226
R21127 a_1297_2982.n68 a_1297_2982.n67 3.01226
R21128 a_1297_2982.n25 a_1297_2982.n23 2.63579
R21129 a_1297_2982.n29 a_1297_2982.n27 2.63579
R21130 a_1297_2982.n41 a_1297_2982.n39 2.63579
R21131 a_1297_2982.n55 a_1297_2982.n53 2.63579
R21132 a_1297_2982.n59 a_1297_2982.n57 2.63579
R21133 a_1297_2982.n11 a_1297_2982.n15 2.2019
R21134 a_1297_2982.n13 a_1297_2982.n1 2.18356
R21135 a_1297_2982.n9 a_1297_2982.n26 1.85087
R21136 a_1297_2982.n3 a_1297_2982.n56 1.85087
R21137 a_1297_2982.n1 a_1297_2982.n22 1.85087
R21138 a_1297_2982.n7 a_1297_2982.n38 1.85087
R21139 a_1297_2982.n5 a_1297_2982.n52 1.85087
R21140 a_1297_2982.n72 a_1297_2982.n11 1.48738
R21141 a_1297_2982.n12 a_1297_2982.n7 1.48434
R21142 a_1297_2982.n13 a_1297_2982.n9 1.48434
R21143 a_1297_2982.n14 a_1297_2982.n5 1.48434
R21144 a_1297_2982.n15 a_1297_2982.n3 1.48434
R21145 a_1297_2982.n14 a_1297_2982.n12 0.735439
R21146 a_1297_2982.n15 a_1297_2982.n14 0.718062
R21147 a_1297_2982.n12 a_1297_2982.n13 0.718062
R21148 a_1297_2982.n1 a_1297_2982.n0 0.577306
R21149 a_1297_2982.n5 a_1297_2982.n4 0.576306
R21150 a_1297_2982.n9 a_1297_2982.n8 0.576265
R21151 a_1297_2982.n7 a_1297_2982.n6 0.576265
R21152 a_1297_2982.n3 a_1297_2982.n2 0.576265
R21153 a_1297_2982.n11 a_1297_2982.n10 0.576237
R21154 a_1297_2982.n17 a_1297_2982.n16 0.461175
R21155 a_1297_2982.n35 a_1297_2982.n34 0.461175
R21156 a_1297_2982.n37 a_1297_2982.n36 0.461175
R21157 a_1297_2982.n47 a_1297_2982.n46 0.461175
R21158 a_1297_2982.n65 a_1297_2982.n64 0.461175
R21159 a_1297_2982.n19 a_1297_2982.n18 0.430121
R21160 a_1297_2982.n31 a_1297_2982.n30 0.430121
R21161 a_1297_2982.n43 a_1297_2982.n42 0.430121
R21162 a_1297_2982.n49 a_1297_2982.n48 0.430121
R21163 a_1297_2982.n61 a_1297_2982.n60 0.430121
R21164 a_1297_2982.n74 a_1297_2982.n73 0.429625
R21165 a_1297_2982.n76 a_1297_2982.n72 0.363995
R21166 VSS.n1033 VSS.t52 1049.46
R21167 VSS.n859 VSS.t37 1045.16
R21168 VSS.t4 VSS.t0 984.947
R21169 VSS.t49 VSS.t6 984.947
R21170 VSS.n1044 VSS.t4 492.474
R21171 VSS.n1044 VSS.t49 492.474
R21172 VSS.n1757 VSS.n1756 292.5
R21173 VSS.n1755 VSS.n1754 292.5
R21174 VSS.n1753 VSS.n1752 292.5
R21175 VSS.n1751 VSS.n1750 292.5
R21176 VSS.n1749 VSS.n1748 292.5
R21177 VSS.n98 VSS.n97 292.5
R21178 VSS.n101 VSS.n100 292.5
R21179 VSS.n101 VSS.n99 292.5
R21180 VSS.n98 VSS.n96 292.5
R21181 VSS.n1949 VSS.n1948 292.5
R21182 VSS.n1951 VSS.n1950 292.5
R21183 VSS.n1953 VSS.n1952 292.5
R21184 VSS.n1955 VSS.n1954 292.5
R21185 VSS.n1957 VSS.n1956 292.5
R21186 VSS.n1959 VSS.n1958 292.5
R21187 VSS.n1759 VSS.n1758 292.5
R21188 VSS.n2115 VSS.n2111 174.535
R21189 VSS.n1802 VSS.n1801 155.356
R21190 VSS.n1046 VSS.n1041 142.119
R21191 VSS.n1054 VSS.n1046 142.119
R21192 VSS.n1919 VSS.n1918 132.803
R21193 VSS.n129 VSS.n128 105.766
R21194 VSS.n129 VSS.n125 105.766
R21195 VSS.n129 VSS.n122 105.766
R21196 VSS.n129 VSS.n119 105.766
R21197 VSS.n129 VSS.n116 105.766
R21198 VSS.n129 VSS.n113 105.766
R21199 VSS.n129 VSS.n110 105.766
R21200 VSS.n129 VSS.n107 105.766
R21201 VSS.n129 VSS.n104 105.766
R21202 VSS.n1746 VSS.n1745 83.9534
R21203 VSS.n1946 VSS.n1945 83.9534
R21204 VSS.n130 VSS.n129 81.2519
R21205 VSS.n128 VSS.n127 80.9725
R21206 VSS.n128 VSS.n126 80.9721
R21207 VSS.n125 VSS.n123 80.9719
R21208 VSS.n122 VSS.n120 80.9719
R21209 VSS.n119 VSS.n117 80.9719
R21210 VSS.n116 VSS.n114 80.9719
R21211 VSS.n113 VSS.n111 80.9719
R21212 VSS.n110 VSS.n108 80.9719
R21213 VSS.n107 VSS.n105 80.9719
R21214 VSS.n104 VSS.n102 80.9719
R21215 VSS.n125 VSS.n124 80.9719
R21216 VSS.n122 VSS.n121 80.9719
R21217 VSS.n119 VSS.n118 80.9719
R21218 VSS.n116 VSS.n115 80.9719
R21219 VSS.n113 VSS.n112 80.9719
R21220 VSS.n110 VSS.n109 80.9719
R21221 VSS.n107 VSS.n106 80.9719
R21222 VSS.n104 VSS.n103 80.9719
R21223 VSS.n2434 VSS.t47 68.2323
R21224 VSS.n1394 VSS.t33 68.2319
R21225 VSS.n2313 VSS.t45 60.2505
R21226 VSS.n2297 VSS.t54 60.2505
R21227 VSS.n259 VSS.t27 60.2505
R21228 VSS.n243 VSS.t41 60.2505
R21229 VSS.n1542 VSS.t39 60.2505
R21230 VSS.n1433 VSS.t31 60.2505
R21231 VSS.n465 VSS.t43 60.2505
R21232 VSS.n449 VSS.t25 60.2505
R21233 VSS.n1140 VSS.t29 60.2505
R21234 VSS.n1221 VSS.t34 60.2505
R21235 VSS.n897 VSS.t51 60.2505
R21236 VSS.n622 VSS.t48 60.2505
R21237 VSS.n735 VSS.t36 60.2505
R21238 VSS.n129 VSS.n101 59.7441
R21239 VSS.n1802 VSS.n1800 59.7441
R21240 VSS.n1760 VSS.n1759 57.6005
R21241 VSS.n1960 VSS.n1959 57.6005
R21242 VSS.n1920 VSS.n1917 49.397
R21243 VSS.n2115 VSS.n2114 49.397
R21244 VSS.n1777 VSS.n1776 46.104
R21245 VSS.n1977 VSS.n1976 46.104
R21246 VSS.n1896 VSS.n1894 42.8108
R21247 VSS.n2091 VSS.n2090 42.8108
R21248 VSS.n1795 VSS.n1794 39.5177
R21249 VSS.n1349 VSS.t2 36.3246
R21250 VSS.n1873 VSS.n1871 36.2246
R21251 VSS.n2068 VSS.n2067 36.2246
R21252 VSS.t42 VSS.n372 35.3798
R21253 VSS.n981 VSS.t53 35.3798
R21254 VSS.n820 VSS.t38 35.3798
R21255 VSS.t26 VSS.n513 35.3798
R21256 VSS.n1930 VSS.t10 35.3798
R21257 VSS.n1825 VSS.n1824 32.9315
R21258 VSS.n101 VSS.n98 32.501
R21259 VSS.n98 VSS.n95 32.501
R21260 VSS.n1798 VSS.n1797 32.501
R21261 VSS.n1799 VSS.n1798 32.501
R21262 VSS.n1800 VSS.n1799 32.501
R21263 VSS.n2438 VSS.n2437 31.4488
R21264 VSS.n1398 VSS.n1397 31.4488
R21265 VSS.n975 VSS.n974 31.4488
R21266 VSS.n982 VSS.n981 31.4488
R21267 VSS.n814 VSS.n813 31.4488
R21268 VSS.n821 VSS.n820 31.4488
R21269 VSS.n1931 VSS.n1930 31.4488
R21270 VSS.n2124 VSS.n2123 31.4488
R21271 VSS.n866 VSS.n862 30.0212
R21272 VSS.n857 VSS.n856 30.0212
R21273 VSS.n1850 VSS.n1848 29.6384
R21274 VSS.n2045 VSS.n2044 29.6384
R21275 VSS.n2449 VSS.n2448 27.5177
R21276 VSS.n187 VSS.n186 27.5177
R21277 VSS.n1408 VSS.n1407 27.5177
R21278 VSS.n964 VSS.n963 27.5177
R21279 VSS.n993 VSS.n992 27.5177
R21280 VSS.n803 VSS.n802 27.5177
R21281 VSS.n832 VSS.n831 27.5177
R21282 VSS.n1306 VSS.n1305 27.5177
R21283 VSS.n1907 VSS.n1906 27.5177
R21284 VSS.n2100 VSS.n2099 27.5177
R21285 VSS.n1848 VSS.n1847 26.3453
R21286 VSS.n80 VSS.t11 26.289
R21287 VSS.n1747 VSS.n1746 25.6005
R21288 VSS.n1749 VSS.n1747 25.6005
R21289 VSS.n1751 VSS.n1749 25.6005
R21290 VSS.n1753 VSS.n1751 25.6005
R21291 VSS.n1755 VSS.n1753 25.6005
R21292 VSS.n1757 VSS.n1755 25.6005
R21293 VSS.n1759 VSS.n1757 25.6005
R21294 VSS.n1745 VSS.n1744 25.6005
R21295 VSS.n1744 VSS.n1743 25.6005
R21296 VSS.n1743 VSS.n1742 25.6005
R21297 VSS.n1742 VSS.n1741 25.6005
R21298 VSS.n1741 VSS.n1740 25.6005
R21299 VSS.n1740 VSS.n1739 25.6005
R21300 VSS.n1739 VSS.n1738 25.6005
R21301 VSS.n1738 VSS.n1737 25.6005
R21302 VSS.n1938 VSS.n1937 25.6005
R21303 VSS.n1939 VSS.n1938 25.6005
R21304 VSS.n1940 VSS.n1939 25.6005
R21305 VSS.n1941 VSS.n1940 25.6005
R21306 VSS.n1942 VSS.n1941 25.6005
R21307 VSS.n1943 VSS.n1942 25.6005
R21308 VSS.n1944 VSS.n1943 25.6005
R21309 VSS.n1945 VSS.n1944 25.6005
R21310 VSS.n1947 VSS.n1946 25.6005
R21311 VSS.n1949 VSS.n1947 25.6005
R21312 VSS.n1951 VSS.n1949 25.6005
R21313 VSS.n1953 VSS.n1951 25.6005
R21314 VSS.n1955 VSS.n1953 25.6005
R21315 VSS.n1957 VSS.n1955 25.6005
R21316 VSS.n1959 VSS.n1957 25.6005
R21317 VSS.n1764 VSS.n1763 25.2105
R21318 VSS.n1964 VSS.n1963 25.2105
R21319 VSS.n1965 VSS.n1964 25.2105
R21320 VSS.n1765 VSS.n1764 25.2105
R21321 VSS.n2460 VSS.n2459 23.5867
R21322 VSS.n198 VSS.n197 23.5867
R21323 VSS.n1421 VSS.n1420 23.5867
R21324 VSS.n953 VSS.n952 23.5867
R21325 VSS.n1006 VSS.n1005 23.5867
R21326 VSS.n792 VSS.n791 23.5867
R21327 VSS.n845 VSS.n844 23.5867
R21328 VSS.n1331 VSS.n1330 23.5867
R21329 VSS.n1884 VSS.n1883 23.5867
R21330 VSS.n2077 VSS.n2076 23.5867
R21331 VSS.n1827 VSS.n1825 23.0522
R21332 VSS.n2022 VSS.n2021 23.0522
R21333 VSS.n1367 VSS.n1366 22.9106
R21334 VSS.n1371 VSS.n1361 22.9106
R21335 VSS.n2422 VSS.n2421 21.6212
R21336 VSS.n158 VSS.n157 21.6212
R21337 VSS.n1457 VSS.n1456 21.6212
R21338 VSS.n921 VSS.n920 21.6212
R21339 VSS.n760 VSS.n759 21.6212
R21340 VSS.n1816 VSS.n1815 21.6212
R21341 VSS.n2009 VSS.n2008 21.6212
R21342 VSS.n1871 VSS.n1870 19.7591
R21343 VSS.n2473 VSS.n2472 19.6557
R21344 VSS.n211 VSS.n210 19.6557
R21345 VSS.n1477 VSS.n1476 19.6557
R21346 VSS.n942 VSS.n941 19.6557
R21347 VSS.n887 VSS.n886 19.6557
R21348 VSS.n781 VSS.n780 19.6557
R21349 VSS.n726 VSS.n725 19.6557
R21350 VSS.n1861 VSS.n1860 19.6557
R21351 VSS.n2054 VSS.n2053 19.6557
R21352 VSS.n1374 VSS.n1371 19.4788
R21353 VSS.n1997 VSS.n1996 19.1141
R21354 VSS.n1998 VSS.n1997 19.1141
R21355 VSS.n2411 VSS.n2410 17.6902
R21356 VSS.n150 VSS.n149 17.6902
R21357 VSS.n1468 VSS.n1467 17.6902
R21358 VSS.n932 VSS.n931 17.6902
R21359 VSS.n872 VSS.n871 17.6902
R21360 VSS.n771 VSS.n770 17.6902
R21361 VSS.n714 VSS.n713 17.6902
R21362 VSS.n1839 VSS.n1838 17.6902
R21363 VSS.n2032 VSS.n2031 17.6902
R21364 VSS.n1804 VSS.n1795 16.466
R21365 VSS.n1999 VSS.n1998 16.466
R21366 VSS.t9 VSS.n1796 16.2508
R21367 VSS.n1797 VSS.t9 16.2508
R21368 VSS.n2021 VSS.n2020 16.0158
R21369 VSS.n2020 VSS.n2019 16.0158
R21370 VSS.n2410 VSS.n2409 15.7246
R21371 VSS.n149 VSS.n148 15.7246
R21372 VSS.n1467 VSS.n1466 15.7246
R21373 VSS.n931 VSS.n930 15.7246
R21374 VSS.n871 VSS.n870 15.7246
R21375 VSS.n770 VSS.n769 15.7246
R21376 VSS.n713 VSS.n712 15.7246
R21377 VSS.n1838 VSS.n1837 15.7246
R21378 VSS.n2031 VSS.n2030 15.7246
R21379 VSS.n2474 VSS.n2473 13.7591
R21380 VSS.n212 VSS.n211 13.7591
R21381 VSS.n1478 VSS.n1477 13.7591
R21382 VSS.n943 VSS.n942 13.7591
R21383 VSS.n888 VSS.n887 13.7591
R21384 VSS.n782 VSS.n781 13.7591
R21385 VSS.n727 VSS.n726 13.7591
R21386 VSS.n1862 VSS.n1861 13.7591
R21387 VSS.n2055 VSS.n2054 13.7591
R21388 VSS.n1894 VSS.n1893 13.1729
R21389 VSS.n2043 VSS.n2042 12.8833
R21390 VSS.n2044 VSS.n2043 12.8833
R21391 VSS.n2133 VSS.n2131 12.8005
R21392 VSS.n2133 VSS.n2132 12.8005
R21393 VSS.n705 VSS.n702 12.0077
R21394 VSS.n2421 VSS.n2420 11.7936
R21395 VSS.n157 VSS.n156 11.7936
R21396 VSS.n1456 VSS.n1455 11.7936
R21397 VSS.n920 VSS.n919 11.7936
R21398 VSS.n862 VSS.n861 11.7936
R21399 VSS.n759 VSS.n758 11.7936
R21400 VSS.n856 VSS.n855 11.7936
R21401 VSS.n1815 VSS.n1814 11.7936
R21402 VSS.n2008 VSS.n2007 11.7936
R21403 VSS.n1779 VSS.n1777 9.87981
R21404 VSS.n2461 VSS.n2460 9.82809
R21405 VSS.n199 VSS.n198 9.82809
R21406 VSS.n1422 VSS.n1421 9.82809
R21407 VSS.n954 VSS.n953 9.82809
R21408 VSS.n1007 VSS.n1006 9.82809
R21409 VSS.n793 VSS.n792 9.82809
R21410 VSS.n846 VSS.n845 9.82809
R21411 VSS.n1332 VSS.n1331 9.82809
R21412 VSS.n1885 VSS.n1884 9.82809
R21413 VSS.n2078 VSS.n2077 9.82809
R21414 VSS.n2067 VSS.n2066 9.71624
R21415 VSS.n2066 VSS.n2065 9.71624
R21416 VSS.n1978 VSS.n1977 9.5667
R21417 VSS.n2309 VSS.n2308 9.3005
R21418 VSS.n2307 VSS.n2306 9.3005
R21419 VSS.n2305 VSS.n2304 9.3005
R21420 VSS.n2304 VSS.n2303 9.3005
R21421 VSS.n2325 VSS.n2324 9.3005
R21422 VSS.n2321 VSS.n2320 9.3005
R21423 VSS.n2320 VSS.n2319 9.3005
R21424 VSS.n2323 VSS.n2322 9.3005
R21425 VSS.n2333 VSS.n2332 9.3005
R21426 VSS.n2340 VSS.n2339 9.3005
R21427 VSS.n2347 VSS.n2346 9.3005
R21428 VSS.n2354 VSS.n2353 9.3005
R21429 VSS.n2361 VSS.n2360 9.3005
R21430 VSS.n2368 VSS.n2367 9.3005
R21431 VSS.n2374 VSS.n2373 9.3005
R21432 VSS.n2381 VSS.n2380 9.3005
R21433 VSS.n2388 VSS.n2387 9.3005
R21434 VSS.n2390 VSS.n2389 9.3005
R21435 VSS.n2386 VSS.n2385 9.3005
R21436 VSS.n2383 VSS.n2382 9.3005
R21437 VSS.n2379 VSS.n2378 9.3005
R21438 VSS.n2376 VSS.n2375 9.3005
R21439 VSS.n2372 VSS.n2371 9.3005
R21440 VSS.n2370 VSS.n2369 9.3005
R21441 VSS.n2366 VSS.n2365 9.3005
R21442 VSS.n2364 VSS.n2363 9.3005
R21443 VSS.n2359 VSS.n2358 9.3005
R21444 VSS.n2357 VSS.n2356 9.3005
R21445 VSS.n2352 VSS.n2351 9.3005
R21446 VSS.n2350 VSS.n2349 9.3005
R21447 VSS.n2345 VSS.n2344 9.3005
R21448 VSS.n2343 VSS.n2342 9.3005
R21449 VSS.n2338 VSS.n2337 9.3005
R21450 VSS.n2336 VSS.n2335 9.3005
R21451 VSS.n2331 VSS.n2330 9.3005
R21452 VSS.n2393 VSS.n2392 9.3005
R21453 VSS.n2443 VSS.n2442 9.3005
R21454 VSS.n2454 VSS.n2453 9.3005
R21455 VSS.n2441 VSS.n2440 9.3005
R21456 VSS.n2440 VSS.n2439 9.3005
R21457 VSS.n2445 VSS.n2444 9.3005
R21458 VSS.n2452 VSS.n2451 9.3005
R21459 VSS.n2451 VSS.n2450 9.3005
R21460 VSS.n2456 VSS.n2455 9.3005
R21461 VSS.n2463 VSS.n2462 9.3005
R21462 VSS.n2462 VSS.n2461 9.3005
R21463 VSS.n2467 VSS.n2466 9.3005
R21464 VSS.n2465 VSS.n2464 9.3005
R21465 VSS.n2423 VSS.n2422 9.3005
R21466 VSS.n2412 VSS.n2411 9.3005
R21467 VSS.n2475 VSS.n2474 9.3005
R21468 VSS.n2470 VSS.n2469 9.3005
R21469 VSS.n181 VSS.n180 9.3005
R21470 VSS.n192 VSS.n191 9.3005
R21471 VSS.n179 VSS.n178 9.3005
R21472 VSS.n178 VSS.n177 9.3005
R21473 VSS.n183 VSS.n182 9.3005
R21474 VSS.n190 VSS.n189 9.3005
R21475 VSS.n189 VSS.n188 9.3005
R21476 VSS.n194 VSS.n193 9.3005
R21477 VSS.n201 VSS.n200 9.3005
R21478 VSS.n200 VSS.n199 9.3005
R21479 VSS.n205 VSS.n204 9.3005
R21480 VSS.n203 VSS.n202 9.3005
R21481 VSS.n151 VSS.n150 9.3005
R21482 VSS.n159 VSS.n158 9.3005
R21483 VSS.n213 VSS.n212 9.3005
R21484 VSS.n208 VSS.n207 9.3005
R21485 VSS.n255 VSS.n254 9.3005
R21486 VSS.n253 VSS.n252 9.3005
R21487 VSS.n251 VSS.n250 9.3005
R21488 VSS.n250 VSS.n249 9.3005
R21489 VSS.n271 VSS.n270 9.3005
R21490 VSS.n267 VSS.n266 9.3005
R21491 VSS.n266 VSS.n265 9.3005
R21492 VSS.n269 VSS.n268 9.3005
R21493 VSS.n279 VSS.n278 9.3005
R21494 VSS.n286 VSS.n285 9.3005
R21495 VSS.n293 VSS.n292 9.3005
R21496 VSS.n300 VSS.n299 9.3005
R21497 VSS.n307 VSS.n306 9.3005
R21498 VSS.n314 VSS.n313 9.3005
R21499 VSS.n320 VSS.n319 9.3005
R21500 VSS.n327 VSS.n326 9.3005
R21501 VSS.n334 VSS.n333 9.3005
R21502 VSS.n336 VSS.n335 9.3005
R21503 VSS.n332 VSS.n331 9.3005
R21504 VSS.n329 VSS.n328 9.3005
R21505 VSS.n325 VSS.n324 9.3005
R21506 VSS.n322 VSS.n321 9.3005
R21507 VSS.n318 VSS.n317 9.3005
R21508 VSS.n316 VSS.n315 9.3005
R21509 VSS.n312 VSS.n311 9.3005
R21510 VSS.n310 VSS.n309 9.3005
R21511 VSS.n305 VSS.n304 9.3005
R21512 VSS.n303 VSS.n302 9.3005
R21513 VSS.n298 VSS.n297 9.3005
R21514 VSS.n296 VSS.n295 9.3005
R21515 VSS.n291 VSS.n290 9.3005
R21516 VSS.n289 VSS.n288 9.3005
R21517 VSS.n284 VSS.n283 9.3005
R21518 VSS.n282 VSS.n281 9.3005
R21519 VSS.n277 VSS.n276 9.3005
R21520 VSS.n339 VSS.n338 9.3005
R21521 VSS.n1550 VSS.n1549 9.3005
R21522 VSS.n1549 VSS.n1548 9.3005
R21523 VSS.n1554 VSS.n1553 9.3005
R21524 VSS.n1552 VSS.n1551 9.3005
R21525 VSS.n1561 VSS.n1560 9.3005
R21526 VSS.n1568 VSS.n1567 9.3005
R21527 VSS.n1575 VSS.n1574 9.3005
R21528 VSS.n1573 VSS.n1572 9.3005
R21529 VSS.n1571 VSS.n1570 9.3005
R21530 VSS.n1566 VSS.n1565 9.3005
R21531 VSS.n1564 VSS.n1563 9.3005
R21532 VSS.n1559 VSS.n1558 9.3005
R21533 VSS.n1403 VSS.n1402 9.3005
R21534 VSS.n1401 VSS.n1400 9.3005
R21535 VSS.n1400 VSS.n1399 9.3005
R21536 VSS.n1441 VSS.n1440 9.3005
R21537 VSS.n1440 VSS.n1439 9.3005
R21538 VSS.n1445 VSS.n1444 9.3005
R21539 VSS.n1443 VSS.n1442 9.3005
R21540 VSS.n1452 VSS.n1451 9.3005
R21541 VSS.n1463 VSS.n1462 9.3005
R21542 VSS.n1474 VSS.n1473 9.3005
R21543 VSS.n1479 VSS.n1478 9.3005
R21544 VSS.n1472 VSS.n1471 9.3005
R21545 VSS.n1470 VSS.n1469 9.3005
R21546 VSS.n1469 VSS.n1468 9.3005
R21547 VSS.n1461 VSS.n1460 9.3005
R21548 VSS.n1459 VSS.n1458 9.3005
R21549 VSS.n1458 VSS.n1457 9.3005
R21550 VSS.n1450 VSS.n1449 9.3005
R21551 VSS.n1405 VSS.n1404 9.3005
R21552 VSS.n1410 VSS.n1409 9.3005
R21553 VSS.n1423 VSS.n1422 9.3005
R21554 VSS.n1241 VSS.n1240 9.3005
R21555 VSS.n1248 VSS.n1247 9.3005
R21556 VSS.n1255 VSS.n1254 9.3005
R21557 VSS.n1253 VSS.n1252 9.3005
R21558 VSS.n1251 VSS.n1250 9.3005
R21559 VSS.n1246 VSS.n1245 9.3005
R21560 VSS.n1244 VSS.n1243 9.3005
R21561 VSS.n1239 VSS.n1238 9.3005
R21562 VSS.n1164 VSS.n1163 9.3005
R21563 VSS.n1168 VSS.n1167 9.3005
R21564 VSS.n1166 VSS.n1165 9.3005
R21565 VSS.n1171 VSS.n1170 9.3005
R21566 VSS.n1173 VSS.n1172 9.3005
R21567 VSS.n1175 VSS.n1174 9.3005
R21568 VSS.n1161 VSS.n1160 9.3005
R21569 VSS.n1159 VSS.n1158 9.3005
R21570 VSS.n1151 VSS.n1150 9.3005
R21571 VSS.n1132 VSS.n1131 9.3005
R21572 VSS.n1231 VSS.n1230 9.3005
R21573 VSS.n1233 VSS.n1232 9.3005
R21574 VSS.n1229 VSS.n1228 9.3005
R21575 VSS.n1228 VSS.n1227 9.3005
R21576 VSS.n1153 VSS.n1152 9.3005
R21577 VSS.n1149 VSS.n1148 9.3005
R21578 VSS.n1148 VSS.n1147 9.3005
R21579 VSS.n1139 VSS.n1138 9.3005
R21580 VSS.n1138 VSS.n1137 9.3005
R21581 VSS.n1218 VSS.n1217 9.3005
R21582 VSS.n461 VSS.n460 9.3005
R21583 VSS.n459 VSS.n458 9.3005
R21584 VSS.n457 VSS.n456 9.3005
R21585 VSS.n456 VSS.n455 9.3005
R21586 VSS.n478 VSS.n477 9.3005
R21587 VSS.n474 VSS.n473 9.3005
R21588 VSS.n473 VSS.n472 9.3005
R21589 VSS.n476 VSS.n475 9.3005
R21590 VSS.n1124 VSS.n1123 9.3005
R21591 VSS.n1123 VSS.n1122 9.3005
R21592 VSS.n1128 VSS.n1127 9.3005
R21593 VSS.n1126 VSS.n1125 9.3005
R21594 VSS.n486 VSS.n485 9.3005
R21595 VSS.n493 VSS.n492 9.3005
R21596 VSS.n500 VSS.n499 9.3005
R21597 VSS.n498 VSS.n497 9.3005
R21598 VSS.n496 VSS.n495 9.3005
R21599 VSS.n491 VSS.n490 9.3005
R21600 VSS.n489 VSS.n488 9.3005
R21601 VSS.n484 VSS.n483 9.3005
R21602 VSS.n907 VSS.n906 9.3005
R21603 VSS.n909 VSS.n908 9.3005
R21604 VSS.n905 VSS.n904 9.3005
R21605 VSS.n904 VSS.n903 9.3005
R21606 VSS.n998 VSS.n997 9.3005
R21607 VSS.n987 VSS.n986 9.3005
R21608 VSS.n971 VSS.n970 9.3005
R21609 VSS.n960 VSS.n959 9.3005
R21610 VSS.n949 VSS.n948 9.3005
R21611 VSS.n938 VSS.n937 9.3005
R21612 VSS.n927 VSS.n926 9.3005
R21613 VSS.n916 VSS.n915 9.3005
R21614 VSS.n914 VSS.n913 9.3005
R21615 VSS.n923 VSS.n922 9.3005
R21616 VSS.n922 VSS.n921 9.3005
R21617 VSS.n925 VSS.n924 9.3005
R21618 VSS.n934 VSS.n933 9.3005
R21619 VSS.n933 VSS.n932 9.3005
R21620 VSS.n936 VSS.n935 9.3005
R21621 VSS.n945 VSS.n944 9.3005
R21622 VSS.n944 VSS.n943 9.3005
R21623 VSS.n947 VSS.n946 9.3005
R21624 VSS.n956 VSS.n955 9.3005
R21625 VSS.n955 VSS.n954 9.3005
R21626 VSS.n958 VSS.n957 9.3005
R21627 VSS.n967 VSS.n966 9.3005
R21628 VSS.n966 VSS.n965 9.3005
R21629 VSS.n969 VSS.n968 9.3005
R21630 VSS.n978 VSS.n977 9.3005
R21631 VSS.n977 VSS.n976 9.3005
R21632 VSS.n985 VSS.n984 9.3005
R21633 VSS.n984 VSS.n983 9.3005
R21634 VSS.n989 VSS.n988 9.3005
R21635 VSS.n996 VSS.n995 9.3005
R21636 VSS.n995 VSS.n994 9.3005
R21637 VSS.n1000 VSS.n999 9.3005
R21638 VSS.n1008 VSS.n1007 9.3005
R21639 VSS.n889 VSS.n888 9.3005
R21640 VSS.n873 VSS.n872 9.3005
R21641 VSS.n632 VSS.n631 9.3005
R21642 VSS.n634 VSS.n633 9.3005
R21643 VSS.n630 VSS.n629 9.3005
R21644 VSS.n629 VSS.n628 9.3005
R21645 VSS.n690 VSS.n689 9.3005
R21646 VSS.n683 VSS.n682 9.3005
R21647 VSS.n677 VSS.n676 9.3005
R21648 VSS.n670 VSS.n669 9.3005
R21649 VSS.n663 VSS.n662 9.3005
R21650 VSS.n656 VSS.n655 9.3005
R21651 VSS.n649 VSS.n648 9.3005
R21652 VSS.n642 VSS.n641 9.3005
R21653 VSS.n640 VSS.n639 9.3005
R21654 VSS.n645 VSS.n644 9.3005
R21655 VSS.n647 VSS.n646 9.3005
R21656 VSS.n652 VSS.n651 9.3005
R21657 VSS.n654 VSS.n653 9.3005
R21658 VSS.n659 VSS.n658 9.3005
R21659 VSS.n661 VSS.n660 9.3005
R21660 VSS.n666 VSS.n665 9.3005
R21661 VSS.n668 VSS.n667 9.3005
R21662 VSS.n673 VSS.n672 9.3005
R21663 VSS.n675 VSS.n674 9.3005
R21664 VSS.n679 VSS.n678 9.3005
R21665 VSS.n681 VSS.n680 9.3005
R21666 VSS.n685 VSS.n684 9.3005
R21667 VSS.n688 VSS.n687 9.3005
R21668 VSS.n692 VSS.n691 9.3005
R21669 VSS.n745 VSS.n744 9.3005
R21670 VSS.n747 VSS.n746 9.3005
R21671 VSS.n743 VSS.n742 9.3005
R21672 VSS.n742 VSS.n741 9.3005
R21673 VSS.n837 VSS.n836 9.3005
R21674 VSS.n826 VSS.n825 9.3005
R21675 VSS.n810 VSS.n809 9.3005
R21676 VSS.n799 VSS.n798 9.3005
R21677 VSS.n788 VSS.n787 9.3005
R21678 VSS.n777 VSS.n776 9.3005
R21679 VSS.n766 VSS.n765 9.3005
R21680 VSS.n755 VSS.n754 9.3005
R21681 VSS.n753 VSS.n752 9.3005
R21682 VSS.n762 VSS.n761 9.3005
R21683 VSS.n761 VSS.n760 9.3005
R21684 VSS.n764 VSS.n763 9.3005
R21685 VSS.n773 VSS.n772 9.3005
R21686 VSS.n772 VSS.n771 9.3005
R21687 VSS.n775 VSS.n774 9.3005
R21688 VSS.n784 VSS.n783 9.3005
R21689 VSS.n783 VSS.n782 9.3005
R21690 VSS.n786 VSS.n785 9.3005
R21691 VSS.n795 VSS.n794 9.3005
R21692 VSS.n794 VSS.n793 9.3005
R21693 VSS.n797 VSS.n796 9.3005
R21694 VSS.n806 VSS.n805 9.3005
R21695 VSS.n805 VSS.n804 9.3005
R21696 VSS.n808 VSS.n807 9.3005
R21697 VSS.n817 VSS.n816 9.3005
R21698 VSS.n816 VSS.n815 9.3005
R21699 VSS.n824 VSS.n823 9.3005
R21700 VSS.n823 VSS.n822 9.3005
R21701 VSS.n828 VSS.n827 9.3005
R21702 VSS.n835 VSS.n834 9.3005
R21703 VSS.n834 VSS.n833 9.3005
R21704 VSS.n839 VSS.n838 9.3005
R21705 VSS.n715 VSS.n714 9.3005
R21706 VSS.n847 VSS.n846 9.3005
R21707 VSS.n728 VSS.n727 9.3005
R21708 VSS.n1318 VSS.n1317 9.3005
R21709 VSS.n1317 VSS.n1316 9.3005
R21710 VSS.n1320 VSS.n1319 9.3005
R21711 VSS.n1333 VSS.n1332 9.3005
R21712 VSS.n1322 VSS.n1321 9.3005
R21713 VSS.n1308 VSS.n1307 9.3005
R21714 VSS.n1817 VSS.n1816 9.3005
R21715 VSS.n1840 VSS.n1839 9.3005
R21716 VSS.n1863 VSS.n1862 9.3005
R21717 VSS.n1886 VSS.n1885 9.3005
R21718 VSS.n1909 VSS.n1908 9.3005
R21719 VSS.n1933 VSS.n1932 9.3005
R21720 VSS.n2126 VSS.n2125 9.3005
R21721 VSS.n2102 VSS.n2101 9.3005
R21722 VSS.n2079 VSS.n2078 9.3005
R21723 VSS.n2056 VSS.n2055 9.3005
R21724 VSS.n2033 VSS.n2032 9.3005
R21725 VSS.n2010 VSS.n2009 9.3005
R21726 VSS.n1785 VSS.n1784 9.3005
R21727 VSS.n1973 VSS.n1972 9.3005
R21728 VSS.n1985 VSS.n1984 9.3005
R21729 VSS.n1983 VSS.n1982 9.3005
R21730 VSS.n1971 VSS.n1970 9.3005
R21731 VSS.n1773 VSS.n1772 9.3005
R21732 VSS.n1771 VSS.n1770 9.3005
R21733 VSS.n1783 VSS.n1782 9.3005
R21734 VSS.n1981 VSS.n1980 9.3005
R21735 VSS.n1980 VSS.n1979 9.3005
R21736 VSS.n1969 VSS.n1968 9.3005
R21737 VSS.n1968 VSS.n1967 9.3005
R21738 VSS.n1769 VSS.n1768 9.3005
R21739 VSS.n1768 VSS.n1767 9.3005
R21740 VSS.n1781 VSS.n1780 9.3005
R21741 VSS.n1780 VSS.n1779 9.3005
R21742 VSS.n1805 VSS.n1804 9.3005
R21743 VSS.n1828 VSS.n1827 9.3005
R21744 VSS.n1851 VSS.n1850 9.3005
R21745 VSS.n1874 VSS.n1873 9.3005
R21746 VSS.n1897 VSS.n1896 9.3005
R21747 VSS.n1921 VSS.n1920 9.3005
R21748 VSS.n2116 VSS.n2115 9.3005
R21749 VSS.n2092 VSS.n2091 9.3005
R21750 VSS.n2069 VSS.n2068 9.3005
R21751 VSS.n2046 VSS.n2045 9.3005
R21752 VSS.n2023 VSS.n2022 9.3005
R21753 VSS.n2000 VSS.n1999 9.3005
R21754 VSS.n37 VSS.n36 9.3005
R21755 VSS.n1350 VSS.n1349 9.01392
R21756 VSS.n1612 VSS.n1611 9.01392
R21757 VSS.n1374 VSS.n1373 9.01392
R21758 VSS.n1373 VSS.n1372 9.01392
R21759 VSS.n1380 VSS.n1379 9.01392
R21760 VSS.n1351 VSS.n1350 9.01392
R21761 VSS.n1613 VSS.n1612 9.01392
R21762 VSS.n1605 VSS.n1604 9.01392
R21763 VSS.n1602 VSS.n1601 9.01392
R21764 VSS.n1141 VSS.n1140 8.76429
R21765 VSS.n466 VSS.n465 8.76429
R21766 VSS.n2302 VSS.n2301 8.21641
R21767 VSS.n2318 VSS.n2317 8.21641
R21768 VSS.n248 VSS.n247 8.21641
R21769 VSS.n264 VSS.n263 8.21641
R21770 VSS.n1547 VSS.n1546 8.21641
R21771 VSS.n1438 VSS.n1437 8.21641
R21772 VSS.n454 VSS.n453 8.21641
R21773 VSS.n1226 VSS.n1225 8.21641
R21774 VSS.n1146 VSS.n1145 8.21641
R21775 VSS.n1136 VSS.n1135 8.21641
R21776 VSS.n471 VSS.n470 8.21641
R21777 VSS.n1121 VSS.n1120 8.21641
R21778 VSS.n902 VSS.n901 8.21641
R21779 VSS.n627 VSS.n626 8.21641
R21780 VSS.n740 VSS.n739 8.21641
R21781 VSS.n136 VSS.n67 7.30029
R21782 VSS.n1803 VSS.n1802 7.0773
R21783 VSS.n87 VSS.n74 6.95702
R21784 VSS.n2298 VSS.n2297 6.92242
R21785 VSS.n244 VSS.n243 6.92242
R21786 VSS.n450 VSS.n449 6.92242
R21787 VSS.n623 VSS.n622 6.92012
R21788 VSS.n736 VSS.n735 6.92012
R21789 VSS.n1222 VSS.n1221 6.92012
R21790 VSS.n2314 VSS.n2313 6.92012
R21791 VSS.n260 VSS.n259 6.92012
R21792 VSS.n898 VSS.n897 6.92011
R21793 VSS.n1543 VSS.n1542 6.92007
R21794 VSS.n1434 VSS.n1433 6.92007
R21795 VSS.n2488 VSS.n2487 6.81049
R21796 VSS.n2492 VSS.n2491 6.81049
R21797 VSS.n2489 VSS.n2488 6.81049
R21798 VSS.n2500 VSS.n2499 6.81049
R21799 VSS.n2493 VSS.n2492 6.81049
R21800 VSS.n1917 VSS.n1916 6.58671
R21801 VSS.n2416 VSS.n2415 6.55106
R21802 VSS.n163 VSS.n162 6.55006
R21803 VSS.n2089 VSS.n2088 6.51388
R21804 VSS.n2090 VSS.n2089 6.51388
R21805 VSS.n1448 VSS.n1447 6.43466
R21806 VSS.n912 VSS.n911 6.43466
R21807 VSS.n751 VSS.n750 6.43466
R21808 VSS.n2436 VSS.n2435 6.02403
R21809 VSS.n175 VSS.n174 6.02403
R21810 VSS.n1396 VSS.n1395 6.02403
R21811 VSS.n973 VSS.n972 6.02403
R21812 VSS.n980 VSS.n979 6.02403
R21813 VSS.n812 VSS.n811 6.02403
R21814 VSS.n819 VSS.n818 6.02403
R21815 VSS.n1314 VSS.n1313 6.02403
R21816 VSS.n1934 VSS.n1927 6.02403
R21817 VSS.n1929 VSS.n1928 6.02403
R21818 VSS.n2122 VSS.n2121 6.02403
R21819 VSS.n2128 VSS.n2127 6.02403
R21820 VSS.n1762 VSS.n1761 6.02403
R21821 VSS.n1962 VSS.n1961 6.02403
R21822 VSS.n2450 VSS.n2449 5.89705
R21823 VSS.n188 VSS.n187 5.89705
R21824 VSS.n1409 VSS.n1408 5.89705
R21825 VSS.n965 VSS.n964 5.89705
R21826 VSS.n994 VSS.n993 5.89705
R21827 VSS.n804 VSS.n803 5.89705
R21828 VSS.n833 VSS.n832 5.89705
R21829 VSS.n1307 VSS.n1306 5.89705
R21830 VSS.n1908 VSS.n1907 5.89705
R21831 VSS.n2101 VSS.n2100 5.89705
R21832 VSS.n2300 VSS.n2299 5.64756
R21833 VSS.n2316 VSS.n2315 5.64756
R21834 VSS.n246 VSS.n245 5.64756
R21835 VSS.n262 VSS.n261 5.64756
R21836 VSS.n1545 VSS.n1544 5.64756
R21837 VSS.n1436 VSS.n1435 5.64756
R21838 VSS.n452 VSS.n451 5.64756
R21839 VSS.n1224 VSS.n1223 5.64756
R21840 VSS.n1144 VSS.n1143 5.64756
R21841 VSS.n1134 VSS.n1133 5.64756
R21842 VSS.n469 VSS.n468 5.64756
R21843 VSS.n1119 VSS.n1118 5.64756
R21844 VSS.n900 VSS.n899 5.64756
R21845 VSS.n625 VSS.n624 5.64756
R21846 VSS.n738 VSS.n737 5.64756
R21847 VSS.n1921 VSS.n1915 5.64756
R21848 VSS.n1923 VSS.n1921 5.64756
R21849 VSS.n2117 VSS.n2116 5.64756
R21850 VSS.n2116 VSS.n2110 5.64756
R21851 VSS.n600 VSS.n599 5.61038
R21852 VSS.n705 VSS.n704 5.61038
R21853 VSS.n1788 VSS.n1787 5.54695
R21854 VSS.n405 VSS.n404 5.39982
R21855 VSS.n2195 VSS.n2194 5.39151
R21856 VSS.n2279 VSS.n2278 5.39151
R21857 VSS.n225 VSS.n224 5.39151
R21858 VSS.n1706 VSS.n1705 5.39051
R21859 VSS.n2165 VSS.n2164 5.39051
R21860 VSS.n2225 VSS.n2224 5.39051
R21861 VSS.n2255 VSS.n2254 5.39051
R21862 VSS.n362 VSS.n361 5.39051
R21863 VSS.n62 VSS.n61 5.38802
R21864 VSS.n867 VSS.n866 5.3711
R21865 VSS.n858 VSS.n857 5.3711
R21866 VSS.n1557 VSS.n1556 5.28653
R21867 VSS.n638 VSS.n637 5.28613
R21868 VSS.n482 VSS.n481 5.2751
R21869 VSS.n1237 VSS.n1236 5.2751
R21870 VSS.n1157 VSS.n1156 5.2751
R21871 VSS.n2329 VSS.n2328 5.27461
R21872 VSS.n275 VSS.n274 5.27461
R21873 VSS.n2447 VSS.n2446 5.27109
R21874 VSS.n185 VSS.n184 5.27109
R21875 VSS.n962 VSS.n961 5.27109
R21876 VSS.n991 VSS.n990 5.27109
R21877 VSS.n801 VSS.n800 5.27109
R21878 VSS.n830 VSS.n829 5.27109
R21879 VSS.n1910 VSS.n1903 5.27109
R21880 VSS.n1905 VSS.n1904 5.27109
R21881 VSS.n2098 VSS.n2097 5.27109
R21882 VSS.n2104 VSS.n2103 5.27109
R21883 VSS.n1775 VSS.n1774 5.27109
R21884 VSS.n1975 VSS.n1974 5.27109
R21885 VSS.n1988 VSS.n1987 5.23535
R21886 VSS.n1718 VSS.n1717 5.13412
R21887 VSS.n2177 VSS.n2176 5.13412
R21888 VSS.n2207 VSS.n2206 5.13412
R21889 VSS.n2237 VSS.n2236 5.13412
R21890 VSS.n2269 VSS.n2268 5.13412
R21891 VSS.n377 VSS.n376 5.13412
R21892 VSS.n1897 VSS.n1892 4.89462
R21893 VSS.n1899 VSS.n1897 4.89462
R21894 VSS.n2093 VSS.n2092 4.89462
R21895 VSS.n2092 VSS.n2087 4.89462
R21896 VSS.n1969 VSS.n1960 4.84343
R21897 VSS.n1769 VSS.n1760 4.84343
R21898 VSS.n133 VSS.n132 4.83275
R21899 VSS.n2311 VSS.n2310 4.76425
R21900 VSS.n2326 VSS.n2312 4.76425
R21901 VSS.n257 VSS.n256 4.76425
R21902 VSS.n272 VSS.n258 4.76425
R21903 VSS.n1555 VSS.n1541 4.76425
R21904 VSS.n1446 VSS.n1432 4.76425
R21905 VSS.n463 VSS.n462 4.76425
R21906 VSS.n1234 VSS.n1220 4.76425
R21907 VSS.n1154 VSS.n1130 4.76425
R21908 VSS.n1219 VSS.n1216 4.76425
R21909 VSS.n479 VSS.n464 4.76425
R21910 VSS.n1129 VSS.n1117 4.76425
R21911 VSS.n910 VSS.n896 4.76425
R21912 VSS.n636 VSS.n635 4.76425
R21913 VSS.n749 VSS.n748 4.76425
R21914 VSS.n1401 VSS.n1394 4.68469
R21915 VSS.n2441 VSS.n2434 4.68392
R21916 VSS.n179 VSS.n173 4.68392
R21917 VSS.n1318 VSS.n1312 4.68392
R21918 VSS.n1142 VSS.n1141 4.6505
R21919 VSS.n467 VSS.n466 4.6505
R21920 VSS.n2152 VSS 4.60572
R21921 VSS.n2458 VSS.n2457 4.51815
R21922 VSS.n196 VSS.n195 4.51815
R21923 VSS.n1413 VSS.n1412 4.51815
R21924 VSS.n595 VSS.n594 4.51815
R21925 VSS.n951 VSS.n950 4.51815
R21926 VSS.n1004 VSS.n1003 4.51815
R21927 VSS.n1010 VSS.n1009 4.51815
R21928 VSS.n698 VSS.n697 4.51815
R21929 VSS.n790 VSS.n789 4.51815
R21930 VSS.n843 VSS.n842 4.51815
R21931 VSS.n849 VSS.n848 4.51815
R21932 VSS.n1311 VSS.n1310 4.51815
R21933 VSS.n1887 VSS.n1880 4.51815
R21934 VSS.n1882 VSS.n1881 4.51815
R21935 VSS.n2075 VSS.n2074 4.51815
R21936 VSS.n2081 VSS.n2080 4.51815
R21937 VSS.n1793 VSS.n1792 4.51815
R21938 VSS.n1807 VSS.n1806 4.51815
R21939 VSS.n2001 VSS.n1993 4.51815
R21940 VSS.n1995 VSS.n1994 4.51815
R21941 VSS.n1581 VSS.n1580 4.5005
R21942 VSS.n1483 VSS.n1482 4.5005
R21943 VSS.n1495 VSS.n1491 4.5005
R21944 VSS.n1499 VSS.n1488 4.5005
R21945 VSS.n1505 VSS.n1504 4.5005
R21946 VSS.n1511 VSS.n1510 4.5005
R21947 VSS.n1526 VSS.n1525 4.5005
R21948 VSS.n1530 VSS.n1519 4.5005
R21949 VSS.n1536 VSS.n1535 4.5005
R21950 VSS.n1539 VSS.n1516 4.5005
R21951 VSS.n1414 VSS.n1413 4.5005
R21952 VSS.n1418 VSS.n1393 4.5005
R21953 VSS.n1427 VSS.n1426 4.5005
R21954 VSS.n1430 VSS.n1390 4.5005
R21955 VSS.n1261 VSS.n1260 4.5005
R21956 VSS.n1181 VSS.n1180 4.5005
R21957 VSS.n506 VSS.n505 4.5005
R21958 VSS.n596 VSS.n595 4.5005
R21959 VSS.n1011 VSS.n1010 4.5005
R21960 VSS.n699 VSS.n698 4.5005
R21961 VSS.n850 VSS.n849 4.5005
R21962 VSS.n609 VSS.n605 4.5005
R21963 VSS.n618 VSS.n617 4.5005
R21964 VSS.n731 VSS.n730 4.5005
R21965 VSS.n879 VSS.n875 4.5005
R21966 VSS.n892 VSS.n891 4.5005
R21967 VSS.n576 VSS.n572 4.5005
R21968 VSS.n585 VSS.n584 4.5005
R21969 VSS.n718 VSS.n717 4.5005
R21970 VSS.n1324 VSS.n1311 4.5005
R21971 VSS.n1328 VSS.n1304 4.5005
R21972 VSS.n1337 VSS.n1336 4.5005
R21973 VSS.n1343 VSS.n1342 4.5005
R21974 VSS.n1207 VSS.n1184 4.5005
R21975 VSS.n1274 VSS.n1273 4.5005
R21976 VSS.n1278 VSS.n1267 4.5005
R21977 VSS.n1284 VSS.n1283 4.5005
R21978 VSS.n1287 VSS.n1264 4.5005
R21979 VSS.n533 VSS.n509 4.5005
R21980 VSS.n530 VSS.n529 4.5005
R21981 VSS.n520 VSS.n519 4.5005
R21982 VSS.n524 VSS.n512 4.5005
R21983 VSS.n1204 VSS.n1203 4.5005
R21984 VSS.n1194 VSS.n1193 4.5005
R21985 VSS.n1198 VSS.n1187 4.5005
R21986 VSS.n64 VSS.n60 4.5005
R21987 VSS.n52 VSS.n51 4.5005
R21988 VSS.n42 VSS.n41 4.5005
R21989 VSS.n31 VSS.n30 4.5005
R21990 VSS.n26 VSS.n25 4.5005
R21991 VSS.n416 VSS.n414 4.5005
R21992 VSS.n423 VSS.n422 4.5005
R21993 VSS.n231 VSS.n230 4.5005
R21994 VSS.n241 VSS.n240 4.5005
R21995 VSS.n216 VSS.n215 4.5005
R21996 VSS.n165 VSS.n161 4.5005
R21997 VSS.n2478 VSS.n2477 4.5005
R21998 VSS.n2285 VSS.n2284 4.5005
R21999 VSS.n2295 VSS.n2294 4.5005
R22000 VSS.n2257 VSS.n2253 4.5005
R22001 VSS.n2227 VSS.n2223 4.5005
R22002 VSS.n2233 VSS.n2219 4.5005
R22003 VSS.n2432 VSS.n2414 4.5005
R22004 VSS.n2426 VSS.n2425 4.5005
R22005 VSS.n2263 VSS.n2249 4.5005
R22006 VSS.n2203 VSS.n2189 4.5005
R22007 VSS.n2167 VSS.n2163 4.5005
R22008 VSS.n2197 VSS.n2193 4.5005
R22009 VSS.n364 VSS.n360 4.5005
R22010 VSS.n370 VSS.n356 4.5005
R22011 VSS.n171 VSS.n153 4.5005
R22012 VSS.n407 VSS.n403 4.5005
R22013 VSS.n1708 VSS.n1704 4.5005
R22014 VSS.n1714 VSS.n1700 4.5005
R22015 VSS.n2173 VSS.n2159 4.5005
R22016 VSS.n2399 VSS.n2398 4.5005
R22017 VSS.n345 VSS.n344 4.5005
R22018 VSS.n1704 VSS.n1702 4.14168
R22019 VSS.n2163 VSS.n2161 4.14168
R22020 VSS.n2193 VSS.n2191 4.14168
R22021 VSS.n2223 VSS.n2221 4.14168
R22022 VSS.n2253 VSS.n2251 4.14168
R22023 VSS.n2284 VSS.n2282 4.14168
R22024 VSS.n2423 VSS.n2419 4.14168
R22025 VSS.n2425 VSS.n2423 4.14168
R22026 VSS.n159 VSS.n155 4.14168
R22027 VSS.n161 VSS.n159 4.14168
R22028 VSS.n230 VSS.n228 4.14168
R22029 VSS.n360 VSS.n358 4.14168
R22030 VSS.n403 VSS.n401 4.14168
R22031 VSS.n1516 VSS.n1515 4.14168
R22032 VSS.n1510 VSS.n1509 4.14168
R22033 VSS.n1458 VSS.n1454 4.14168
R22034 VSS.n1390 VSS.n1389 4.14168
R22035 VSS.n509 VSS.n508 4.14168
R22036 VSS.n1264 VSS.n1263 4.14168
R22037 VSS.n1184 VSS.n1183 4.14168
R22038 VSS.n922 VSS.n918 4.14168
R22039 VSS.n865 VSS.n864 4.14168
R22040 VSS.n761 VSS.n757 4.14168
R22041 VSS.n854 VSS.n853 4.14168
R22042 VSS.n1342 VSS.n1341 4.14168
R22043 VSS.n1818 VSS.n1817 4.14168
R22044 VSS.n1817 VSS.n1813 4.14168
R22045 VSS.n2010 VSS.n2006 4.14168
R22046 VSS.n2012 VSS.n2010 4.14168
R22047 VSS.n1874 VSS.n1869 4.14168
R22048 VSS.n1876 VSS.n1874 4.14168
R22049 VSS.n2070 VSS.n2069 4.14168
R22050 VSS.n2069 VSS.n2064 4.14168
R22051 VSS.n41 VSS.n39 4.14168
R22052 VSS.n60 VSS.n58 4.14168
R22053 VSS.n1785 VSS.n1783 3.88788
R22054 VSS.n2392 VSS.n2391 3.76521
R22055 VSS.n2398 VSS.n2396 3.76521
R22056 VSS.n2469 VSS.n2468 3.76521
R22057 VSS.n2477 VSS.n2475 3.76521
R22058 VSS.n207 VSS.n206 3.76521
R22059 VSS.n215 VSS.n213 3.76521
R22060 VSS.n338 VSS.n337 3.76521
R22061 VSS.n344 VSS.n342 3.76521
R22062 VSS.n1535 VSS.n1534 3.76521
R22063 VSS.n1504 VSS.n1503 3.76521
R22064 VSS.n1426 VSS.n1425 3.76521
R22065 VSS.n529 VSS.n528 3.76521
R22066 VSS.n1283 VSS.n1282 3.76521
R22067 VSS.n1203 VSS.n1202 3.76521
R22068 VSS.n584 VSS.n583 3.76521
R22069 VSS.n940 VSS.n939 3.76521
R22070 VSS.n885 VSS.n884 3.76521
R22071 VSS.n891 VSS.n890 3.76521
R22072 VSS.n617 VSS.n616 3.76521
R22073 VSS.n779 VSS.n778 3.76521
R22074 VSS.n724 VSS.n723 3.76521
R22075 VSS.n730 VSS.n729 3.76521
R22076 VSS.n1336 VSS.n1335 3.76521
R22077 VSS.n1864 VSS.n1857 3.76521
R22078 VSS.n1859 VSS.n1858 3.76521
R22079 VSS.n2052 VSS.n2051 3.76521
R22080 VSS.n2058 VSS.n2057 3.76521
R22081 VSS.n1823 VSS.n1822 3.76521
R22082 VSS.n1830 VSS.n1829 3.76521
R22083 VSS.n2024 VSS.n2016 3.76521
R22084 VSS.n2018 VSS.n2017 3.76521
R22085 VSS.n16 VSS.n14 3.49117
R22086 VSS.n1550 VSS.n1543 3.47842
R22087 VSS.n1441 VSS.n1434 3.47842
R22088 VSS.n1229 VSS.n1222 3.47756
R22089 VSS.n630 VSS.n623 3.47756
R22090 VSS.n743 VSS.n736 3.47756
R22091 VSS.n2321 VSS.n2314 3.47756
R22092 VSS.n267 VSS.n260 3.47756
R22093 VSS.n905 VSS.n898 3.47753
R22094 VSS.n2305 VSS.n2298 3.4767
R22095 VSS.n251 VSS.n244 3.4767
R22096 VSS.n457 VSS.n450 3.4767
R22097 VSS.n1700 VSS.n1698 3.38874
R22098 VSS.n2159 VSS.n2157 3.38874
R22099 VSS.n2189 VSS.n2187 3.38874
R22100 VSS.n2219 VSS.n2217 3.38874
R22101 VSS.n2249 VSS.n2247 3.38874
R22102 VSS.n2294 VSS.n2292 3.38874
R22103 VSS.n2412 VSS.n2408 3.38874
R22104 VSS.n2414 VSS.n2412 3.38874
R22105 VSS.n151 VSS.n147 3.38874
R22106 VSS.n153 VSS.n151 3.38874
R22107 VSS.n240 VSS.n238 3.38874
R22108 VSS.n356 VSS.n354 3.38874
R22109 VSS.n414 VSS.n412 3.38874
R22110 VSS.n1469 VSS.n1465 3.38874
R22111 VSS.n572 VSS.n570 3.38874
R22112 VSS.n933 VSS.n929 3.38874
R22113 VSS.n873 VSS.n869 3.38874
R22114 VSS.n875 VSS.n873 3.38874
R22115 VSS.n605 VSS.n603 3.38874
R22116 VSS.n772 VSS.n768 3.38874
R22117 VSS.n715 VSS.n711 3.38874
R22118 VSS.n717 VSS.n715 3.38874
R22119 VSS.n1841 VSS.n1840 3.38874
R22120 VSS.n1840 VSS.n1836 3.38874
R22121 VSS.n2033 VSS.n2029 3.38874
R22122 VSS.n2035 VSS.n2033 3.38874
R22123 VSS.n1851 VSS.n1846 3.38874
R22124 VSS.n1853 VSS.n1851 3.38874
R22125 VSS.n2047 VSS.n2046 3.38874
R22126 VSS.n2046 VSS.n2041 3.38874
R22127 VSS.n51 VSS.n49 3.38874
R22128 VSS.n1381 VSS.n1380 3.33963
R22129 VSS.n1606 VSS.n1602 3.33963
R22130 VSS.n1606 VSS.n1605 3.33963
R22131 VSS.n2500 VSS.n2498 3.33963
R22132 VSS.n2489 VSS.n2486 3.33963
R22133 VSS.n1613 VSS.n1385 3.33963
R22134 VSS.n1613 VSS.n1610 3.33963
R22135 VSS.n1716 VSS.t22 3.3065
R22136 VSS.n1716 VSS.t15 3.3065
R22137 VSS.n2175 VSS.t24 3.3065
R22138 VSS.n2175 VSS.t23 3.3065
R22139 VSS.n2205 VSS.t56 3.3065
R22140 VSS.n2205 VSS.t16 3.3065
R22141 VSS.n2235 VSS.t14 3.3065
R22142 VSS.n2235 VSS.t18 3.3065
R22143 VSS.n2267 VSS.t12 3.3065
R22144 VSS.n2267 VSS.t55 3.3065
R22145 VSS.t55 VSS.n2266 3.3065
R22146 VSS.n2266 VSS.t46 3.3065
R22147 VSS.n374 VSS.t42 3.3065
R22148 VSS.t28 VSS.n374 3.3065
R22149 VSS.n375 VSS.t28 3.3065
R22150 VSS.n375 VSS.t20 3.3065
R22151 VSS.n418 VSS.t21 3.3065
R22152 VSS.n418 VSS.t19 3.3065
R22153 VSS.n1520 VSS.t40 3.3065
R22154 VSS.n1520 VSS.t8 3.3065
R22155 VSS.n1492 VSS.t3 3.3065
R22156 VSS.n1492 VSS.t32 3.3065
R22157 VSS.n514 VSS.t26 3.3065
R22158 VSS.n514 VSS.t44 3.3065
R22159 VSS.n1268 VSS.t35 3.3065
R22160 VSS.n1188 VSS.t30 3.3065
R22161 VSS.n589 VSS.t1 3.3065
R22162 VSS.n589 VSS.t5 3.3065
R22163 VSS.n702 VSS.t50 3.3065
R22164 VSS.n702 VSS.t7 3.3065
R22165 VSS.n15 VSS.t13 3.3065
R22166 VSS.n15 VSS.t17 3.3065
R22167 VSS.n1767 VSS.n1765 3.2936
R22168 VSS.n1967 VSS.n1965 3.2936
R22169 VSS.n2114 VSS.n2113 3.27567
R22170 VSS.n2113 VSS.n2112 3.27567
R22171 VSS.n1580 VSS.n1578 3.22952
R22172 VSS.n505 VSS.n503 3.22952
R22173 VSS.n1260 VSS.n1258 3.22952
R22174 VSS.n1180 VSS.n1178 3.22952
R22175 VSS.n1380 VSS.n1378 3.03311
R22176 VSS.n1375 VSS.n1374 3.03311
R22177 VSS.n1819 VSS.n1818 3.03311
R22178 VSS.n1842 VSS.n1841 3.03311
R22179 VSS.n1865 VSS.n1864 3.03311
R22180 VSS.n1888 VSS.n1887 3.03311
R22181 VSS.n1911 VSS.n1910 3.03311
R22182 VSS.n1935 VSS.n1934 3.03311
R22183 VSS.n2129 VSS.n2128 3.03311
R22184 VSS.n2105 VSS.n2104 3.03311
R22185 VSS.n2082 VSS.n2081 3.03311
R22186 VSS.n2059 VSS.n2058 3.03311
R22187 VSS.n2036 VSS.n2035 3.03311
R22188 VSS.n2013 VSS.n2012 3.03311
R22189 VSS.n2002 VSS.n2001 3.03311
R22190 VSS.n1808 VSS.n1807 3.03311
R22191 VSS.n1831 VSS.n1830 3.03311
R22192 VSS.n1854 VSS.n1853 3.03311
R22193 VSS.n1877 VSS.n1876 3.03311
R22194 VSS.n1900 VSS.n1899 3.03311
R22195 VSS.n1924 VSS.n1923 3.03311
R22196 VSS.n2118 VSS.n2117 3.03311
R22197 VSS.n2094 VSS.n2093 3.03311
R22198 VSS.n2071 VSS.n2070 3.03311
R22199 VSS.n2048 VSS.n2047 3.03311
R22200 VSS.n2025 VSS.n2024 3.03311
R22201 VSS.n1352 VSS.n1351 3.03311
R22202 VSS.n1614 VSS.n1613 3.03311
R22203 VSS.n2490 VSS.n2489 3.03311
R22204 VSS.n1605 VSS.n1603 3.03311
R22205 VSS.n1602 VSS.n1600 3.03311
R22206 VSS.n2501 VSS.n2500 3.03311
R22207 VSS.n2494 VSS.n2493 3.03311
R22208 VSS.n1700 VSS.n1699 3.01226
R22209 VSS.n2159 VSS.n2158 3.01226
R22210 VSS.n2189 VSS.n2188 3.01226
R22211 VSS.n2219 VSS.n2218 3.01226
R22212 VSS.n2249 VSS.n2248 3.01226
R22213 VSS.n2294 VSS.n2293 3.01226
R22214 VSS.n2408 VSS.n2407 3.01226
R22215 VSS.n2414 VSS.n2413 3.01226
R22216 VSS.n147 VSS.n146 3.01226
R22217 VSS.n153 VSS.n152 3.01226
R22218 VSS.n240 VSS.n239 3.01226
R22219 VSS.n356 VSS.n355 3.01226
R22220 VSS.n414 VSS.n413 3.01226
R22221 VSS.n1580 VSS.n1579 3.01226
R22222 VSS.n1465 VSS.n1464 3.01226
R22223 VSS.n1482 VSS.n1481 3.01226
R22224 VSS.n505 VSS.n504 3.01226
R22225 VSS.n1260 VSS.n1259 3.01226
R22226 VSS.n1180 VSS.n1179 3.01226
R22227 VSS.n572 VSS.n571 3.01226
R22228 VSS.n929 VSS.n928 3.01226
R22229 VSS.n869 VSS.n868 3.01226
R22230 VSS.n875 VSS.n874 3.01226
R22231 VSS.n605 VSS.n604 3.01226
R22232 VSS.n768 VSS.n767 3.01226
R22233 VSS.n711 VSS.n710 3.01226
R22234 VSS.n717 VSS.n716 3.01226
R22235 VSS.n1841 VSS.n1834 3.01226
R22236 VSS.n1836 VSS.n1835 3.01226
R22237 VSS.n2029 VSS.n2028 3.01226
R22238 VSS.n2035 VSS.n2034 3.01226
R22239 VSS.n1846 VSS.n1845 3.01226
R22240 VSS.n1853 VSS.n1852 3.01226
R22241 VSS.n2047 VSS.n2039 3.01226
R22242 VSS.n2041 VSS.n2040 3.01226
R22243 VSS.n51 VSS.n50 3.01226
R22244 VSS.n2152 VSS.n2151 2.94883
R22245 VSS.n2398 VSS.n2397 2.63579
R22246 VSS.n2477 VSS.n2476 2.63579
R22247 VSS.n215 VSS.n214 2.63579
R22248 VSS.n344 VSS.n343 2.63579
R22249 VSS.n422 VSS.n421 2.63579
R22250 VSS.n1480 VSS.n1479 2.63579
R22251 VSS.n584 VSS.n582 2.63579
R22252 VSS.n944 VSS.n940 2.63579
R22253 VSS.n889 VSS.n885 2.63579
R22254 VSS.n891 VSS.n889 2.63579
R22255 VSS.n617 VSS.n615 2.63579
R22256 VSS.n783 VSS.n779 2.63579
R22257 VSS.n728 VSS.n724 2.63579
R22258 VSS.n730 VSS.n728 2.63579
R22259 VSS.n1864 VSS.n1863 2.63579
R22260 VSS.n1863 VSS.n1859 2.63579
R22261 VSS.n2056 VSS.n2052 2.63579
R22262 VSS.n2058 VSS.n2056 2.63579
R22263 VSS.n1828 VSS.n1823 2.63579
R22264 VSS.n1830 VSS.n1828 2.63579
R22265 VSS.n2024 VSS.n2023 2.63579
R22266 VSS.n2023 VSS.n2018 2.63579
R22267 VSS.n25 VSS.n21 2.63579
R22268 VSS.n1535 VSS.n1533 2.529
R22269 VSS.n1504 VSS.n1502 2.529
R22270 VSS.n529 VSS.n527 2.529
R22271 VSS.n1283 VSS.n1281 2.529
R22272 VSS.n1203 VSS.n1201 2.529
R22273 VSS.n1346 VSS.n1345 2.35698
R22274 VSS.n2134 VSS.n2133 2.28739
R22275 VSS.n1704 VSS.n1703 2.25932
R22276 VSS.n2163 VSS.n2162 2.25932
R22277 VSS.n2193 VSS.n2192 2.25932
R22278 VSS.n2223 VSS.n2222 2.25932
R22279 VSS.n2253 VSS.n2252 2.25932
R22280 VSS.n2284 VSS.n2283 2.25932
R22281 VSS.n2419 VSS.n2418 2.25932
R22282 VSS.n2425 VSS.n2424 2.25932
R22283 VSS.n155 VSS.n154 2.25932
R22284 VSS.n161 VSS.n160 2.25932
R22285 VSS.n230 VSS.n229 2.25932
R22286 VSS.n360 VSS.n359 2.25932
R22287 VSS.n403 VSS.n402 2.25932
R22288 VSS.n1518 VSS.n1517 2.25932
R22289 VSS.n1487 VSS.n1486 2.25932
R22290 VSS.n1454 VSS.n1453 2.25932
R22291 VSS.n1392 VSS.n1391 2.25932
R22292 VSS.n511 VSS.n510 2.25932
R22293 VSS.n1266 VSS.n1265 2.25932
R22294 VSS.n1186 VSS.n1185 2.25932
R22295 VSS.n918 VSS.n917 2.25932
R22296 VSS.n864 VSS.n863 2.25932
R22297 VSS.n757 VSS.n756 2.25932
R22298 VSS.n853 VSS.n852 2.25932
R22299 VSS.n1303 VSS.n1302 2.25932
R22300 VSS.n1818 VSS.n1811 2.25932
R22301 VSS.n1813 VSS.n1812 2.25932
R22302 VSS.n2006 VSS.n2005 2.25932
R22303 VSS.n2012 VSS.n2011 2.25932
R22304 VSS.n1869 VSS.n1868 2.25932
R22305 VSS.n1876 VSS.n1875 2.25932
R22306 VSS.n2070 VSS.n2062 2.25932
R22307 VSS.n2064 VSS.n2063 2.25932
R22308 VSS.n41 VSS.n40 2.25932
R22309 VSS.n60 VSS.n59 2.25932
R22310 VSS.n1055 VSS.n1054 2.24394
R22311 VSS.n36 VSS.n35 2.24086
R22312 VSS.n1920 VSS.n1919 2.11221
R22313 VSS.n1967 VSS.n1966 2.11221
R22314 VSS.n1767 VSS.n1766 2.11221
R22315 VSS.n1779 VSS.n1778 2.11221
R22316 VSS.n1804 VSS.n1803 2.11221
R22317 VSS.n1827 VSS.n1826 2.11221
R22318 VSS.n1850 VSS.n1849 2.11221
R22319 VSS.n1873 VSS.n1872 2.11221
R22320 VSS.n1896 VSS.n1895 2.11221
R22321 VSS.n2439 VSS.n2438 1.96602
R22322 VSS.n177 VSS.n176 1.96602
R22323 VSS.n1399 VSS.n1398 1.96602
R22324 VSS.n976 VSS.n975 1.96602
R22325 VSS.n983 VSS.n982 1.96602
R22326 VSS.n815 VSS.n814 1.96602
R22327 VSS.n822 VSS.n821 1.96602
R22328 VSS.n1316 VSS.n1315 1.96602
R22329 VSS.n1932 VSS.n1931 1.96602
R22330 VSS.n2125 VSS.n2124 1.96602
R22331 VSS.n2462 VSS.n2458 1.88285
R22332 VSS.n200 VSS.n196 1.88285
R22333 VSS.n1424 VSS.n1423 1.88285
R22334 VSS.n595 VSS.n593 1.88285
R22335 VSS.n955 VSS.n951 1.88285
R22336 VSS.n1008 VSS.n1004 1.88285
R22337 VSS.n1010 VSS.n1008 1.88285
R22338 VSS.n698 VSS.n696 1.88285
R22339 VSS.n794 VSS.n790 1.88285
R22340 VSS.n847 VSS.n843 1.88285
R22341 VSS.n849 VSS.n847 1.88285
R22342 VSS.n1334 VSS.n1333 1.88285
R22343 VSS.n1887 VSS.n1886 1.88285
R22344 VSS.n1886 VSS.n1882 1.88285
R22345 VSS.n2079 VSS.n2075 1.88285
R22346 VSS.n2081 VSS.n2079 1.88285
R22347 VSS.n1805 VSS.n1793 1.88285
R22348 VSS.n1807 VSS.n1805 1.88285
R22349 VSS.n2001 VSS.n2000 1.88285
R22350 VSS.n2000 VSS.n1995 1.88285
R22351 VSS.n25 VSS.n24 1.88285
R22352 VSS.n1525 VSS.n1524 1.82308
R22353 VSS.n1491 VSS.n1490 1.82308
R22354 VSS.n519 VSS.n518 1.82308
R22355 VSS.n1273 VSS.n1272 1.82308
R22356 VSS.n1193 VSS.n1192 1.82308
R22357 VSS.n1299 VSS.n1298 1.71173
R22358 VSS.n1056 VSS.n1055 1.70717
R22359 VSS.n1647 VSS.n1646 1.70597
R22360 VSS.n1634 VSS.n1633 1.70597
R22361 VSS.n1647 VSS.n1641 1.70596
R22362 VSS.n1104 VSS.n1103 1.70592
R22363 VSS.n1636 VSS.n545 1.70592
R22364 VSS.n566 VSS.n565 1.70591
R22365 VSS.n1098 VSS.n1097 1.70577
R22366 VSS.n555 VSS.n554 1.70511
R22367 VSS.n546 VSS 1.68959
R22368 VSS.n143 VSS.n66 1.6655
R22369 VSS.n1787 VSS.n1786 1.65133
R22370 VSS.n1987 VSS.n1986 1.65133
R22371 VSS.n16 VSS.n15 1.60574
R22372 VSS.n2266 VSS.n2265 1.60111
R22373 VSS.n374 VSS.n373 1.60111
R22374 VSS.n702 VSS.n701 1.60111
R22375 VSS.n591 VSS.n590 1.52198
R22376 VSS.n1074 VSS.n601 1.51434
R22377 VSS.n1065 VSS.n706 1.51434
R22378 VSS.n1061 VSS.n858 1.51434
R22379 VSS.n1025 VSS.n867 1.51289
R22380 VSS.n1892 VSS.n1891 1.50638
R22381 VSS.n1899 VSS.n1898 1.50638
R22382 VSS.n2093 VSS.n2085 1.50638
R22383 VSS.n2087 VSS.n2086 1.50638
R22384 VSS.n30 VSS.n29 1.50638
R22385 VSS.n2481 VSS.n2480 1.48392
R22386 VSS.n2273 VSS.n2272 1.48392
R22387 VSS.n2241 VSS.n2240 1.48392
R22388 VSS.n381 VSS.n380 1.48392
R22389 VSS.n219 VSS.n218 1.48392
R22390 VSS.n1722 VSS.n1721 1.48392
R22391 VSS.n2181 VSS.n2180 1.48392
R22392 VSS.n348 VSS.n347 1.48392
R22393 VSS.n2402 VSS.n2401 1.48392
R22394 VSS.n2211 VSS.n2210 1.48392
R22395 VSS.n1521 VSS.n1520 1.46886
R22396 VSS.n1189 VSS.n1188 1.46886
R22397 VSS.n515 VSS.n514 1.46879
R22398 VSS.n1269 VSS.n1268 1.46879
R22399 VSS.n1493 VSS.n1492 1.46878
R22400 VSS.n85 VSS.n84 1.43435
R22401 VSS.n1718 VSS.n1716 1.41292
R22402 VSS.n2177 VSS.n2175 1.41292
R22403 VSS.n2207 VSS.n2205 1.41292
R22404 VSS.n2237 VSS.n2235 1.41292
R22405 VSS.n2269 VSS.n2267 1.41292
R22406 VSS.n377 VSS.n375 1.41292
R22407 VSS.n426 VSS.n425 1.34465
R22408 VSS.n426 VSS.n410 1.34235
R22409 VSS.n446 VSS.n445 1.13717
R22410 VSS.n440 VSS.n439 1.13717
R22411 VSS.n1296 VSS.n1295 1.13717
R22412 VSS.n1211 VSS.n1210 1.13717
R22413 VSS.n543 VSS.n542 1.13717
R22414 VSS.n1631 VSS.n1630 1.13717
R22415 VSS.n1074 VSS.n597 1.13083
R22416 VSS.n1065 VSS.n700 1.13027
R22417 VSS.n1061 VSS.n851 1.13027
R22418 VSS.n1025 VSS.n1012 1.13002
R22419 VSS.n2451 VSS.n2447 1.12991
R22420 VSS.n189 VSS.n185 1.12991
R22421 VSS.n1411 VSS.n1410 1.12991
R22422 VSS.n966 VSS.n962 1.12991
R22423 VSS.n995 VSS.n991 1.12991
R22424 VSS.n805 VSS.n801 1.12991
R22425 VSS.n834 VSS.n830 1.12991
R22426 VSS.n1309 VSS.n1308 1.12991
R22427 VSS.n1910 VSS.n1909 1.12991
R22428 VSS.n1909 VSS.n1905 1.12991
R22429 VSS.n2102 VSS.n2098 1.12991
R22430 VSS.n2104 VSS.n2102 1.12991
R22431 VSS.n1780 VSS.n1775 1.12991
R22432 VSS.n1980 VSS.n1975 1.12991
R22433 VSS.n23 VSS.n22 1.12991
R22434 VSS.n65 VSS.n64 1.1255
R22435 VSS.n2303 VSS.n2302 1.09595
R22436 VSS.n2319 VSS.n2318 1.09595
R22437 VSS.n249 VSS.n248 1.09595
R22438 VSS.n265 VSS.n264 1.09595
R22439 VSS.n1548 VSS.n1547 1.09595
R22440 VSS.n1439 VSS.n1438 1.09595
R22441 VSS.n455 VSS.n454 1.09595
R22442 VSS.n1227 VSS.n1226 1.09595
R22443 VSS.n1147 VSS.n1146 1.09595
R22444 VSS.n1137 VSS.n1136 1.09595
R22445 VSS.n472 VSS.n471 1.09595
R22446 VSS.n1122 VSS.n1121 1.09595
R22447 VSS.n903 VSS.n902 1.09595
R22448 VSS.n628 VSS.n627 1.09595
R22449 VSS.n741 VSS.n740 1.09595
R22450 VSS.n419 VSS.n418 1.0555
R22451 VSS.n1589 VSS.n1513 0.903813
R22452 VSS.n1291 VSS.n1289 0.903813
R22453 VSS.n1621 VSS.n1346 0.903541
R22454 VSS.n1585 VSS.n1582 0.90354
R22455 VSS.n1594 VSS.n1484 0.90354
R22456 VSS.n2153 VSS.n2152 0.790344
R22457 VSS.n1031 VSS.n1030 0.787987
R22458 VSS.n2304 VSS.n2300 0.753441
R22459 VSS.n2320 VSS.n2316 0.753441
R22460 VSS.n250 VSS.n246 0.753441
R22461 VSS.n266 VSS.n262 0.753441
R22462 VSS.n1549 VSS.n1545 0.753441
R22463 VSS.n1482 VSS.n1480 0.753441
R22464 VSS.n1426 VSS.n1424 0.753441
R22465 VSS.n1413 VSS.n1411 0.753441
R22466 VSS.n1440 VSS.n1436 0.753441
R22467 VSS.n456 VSS.n452 0.753441
R22468 VSS.n1228 VSS.n1224 0.753441
R22469 VSS.n1148 VSS.n1144 0.753441
R22470 VSS.n1138 VSS.n1134 0.753441
R22471 VSS.n473 VSS.n469 0.753441
R22472 VSS.n1123 VSS.n1119 0.753441
R22473 VSS.n904 VSS.n900 0.753441
R22474 VSS.n629 VSS.n625 0.753441
R22475 VSS.n742 VSS.n738 0.753441
R22476 VSS.n1336 VSS.n1334 0.753441
R22477 VSS.n1311 VSS.n1309 0.753441
R22478 VSS.n1915 VSS.n1914 0.753441
R22479 VSS.n1923 VSS.n1922 0.753441
R22480 VSS.n2117 VSS.n2108 0.753441
R22481 VSS.n2110 VSS.n2109 0.753441
R22482 VSS.n24 VSS.n23 0.753441
R22483 VSS.n1599 VSS.n1598 0.720975
R22484 VSS.n1616 VSS.n1615 0.720975
R22485 VSS.n1210 VSS.n1209 0.707257
R22486 VSS.n542 VSS.n535 0.707257
R22487 VSS.n1587 VSS.n1586 0.682531
R22488 VSS.n1063 VSS.n1062 0.682531
R22489 VSS.n2184 VSS.n2183 0.682531
R22490 VSS.n2214 VSS.n2213 0.682531
R22491 VSS.n2244 VSS.n2243 0.682531
R22492 VSS.n1679 VSS.n1678 0.6825
R22493 VSS.n420 VSS.n419 0.640088
R22494 VSS.n2505 VSS.n2502 0.614024
R22495 VSS.n1513 VSS.n1485 0.594417
R22496 VSS.n1522 VSS.n1521 0.575661
R22497 VSS.n1270 VSS.n1269 0.575335
R22498 VSS.n516 VSS.n515 0.574421
R22499 VSS.n1190 VSS.n1189 0.574409
R22500 VSS.n1083 VSS.n1082 0.568833
R22501 VSS.n1494 VSS.n1493 0.561441
R22502 VSS.n2153 VSS.n1724 0.541125
R22503 VSS.n1067 VSS.n1066 0.534875
R22504 VSS.n1702 VSS.n1701 0.461175
R22505 VSS.n2161 VSS.n2160 0.461175
R22506 VSS.n2191 VSS.n2190 0.461175
R22507 VSS.n2221 VSS.n2220 0.461175
R22508 VSS.n2251 VSS.n2250 0.461175
R22509 VSS.n2335 VSS.n2334 0.461175
R22510 VSS.n2282 VSS.n2281 0.461175
R22511 VSS.n281 VSS.n280 0.461175
R22512 VSS.n228 VSS.n227 0.461175
R22513 VSS.n358 VSS.n357 0.461175
R22514 VSS.n401 VSS.n400 0.461175
R22515 VSS.n1563 VSS.n1562 0.461175
R22516 VSS.n488 VSS.n487 0.461175
R22517 VSS.n1243 VSS.n1242 0.461175
R22518 VSS.n1163 VSS.n1162 0.461175
R22519 VSS.n599 VSS.n598 0.461175
R22520 VSS.n704 VSS.n703 0.461175
R22521 VSS.n58 VSS.n57 0.461175
R22522 VSS.n644 VSS.n643 0.460679
R22523 VSS.n141 VSS.n140 0.430441
R22524 VSS.n1698 VSS.n1697 0.430121
R22525 VSS.n2157 VSS.n2156 0.430121
R22526 VSS.n2187 VSS.n2186 0.430121
R22527 VSS.n2217 VSS.n2216 0.430121
R22528 VSS.n2247 VSS.n2246 0.430121
R22529 VSS.n2342 VSS.n2341 0.430121
R22530 VSS.n2292 VSS.n2291 0.430121
R22531 VSS.n288 VSS.n287 0.430121
R22532 VSS.n238 VSS.n237 0.430121
R22533 VSS.n354 VSS.n353 0.430121
R22534 VSS.n412 VSS.n411 0.430121
R22535 VSS.n1570 VSS.n1569 0.430121
R22536 VSS.n495 VSS.n494 0.430121
R22537 VSS.n1250 VSS.n1249 0.430121
R22538 VSS.n1170 VSS.n1169 0.430121
R22539 VSS.n570 VSS.n569 0.430121
R22540 VSS.n603 VSS.n602 0.430121
R22541 VSS.n49 VSS.n48 0.430121
R22542 VSS.n651 VSS.n650 0.429625
R22543 VSS.n1448 VSS.n1446 0.420318
R22544 VSS.n912 VSS.n910 0.420318
R22545 VSS.n751 VSS.n749 0.420318
R22546 VSS.n2349 VSS.n2348 0.398603
R22547 VSS.n295 VSS.n294 0.398603
R22548 VSS.n582 VSS.n581 0.398603
R22549 VSS.n615 VSS.n614 0.398603
R22550 VSS.n658 VSS.n657 0.398108
R22551 VSS.n1028 VSS.n1027 0.382531
R22552 VSS.n590 VSS.n589 0.378264
R22553 VSS.n2440 VSS.n2436 0.376971
R22554 VSS.n178 VSS.n175 0.376971
R22555 VSS.n1516 VSS.n1514 0.376971
R22556 VSS.n1519 VSS.n1518 0.376971
R22557 VSS.n1510 VSS.n1508 0.376971
R22558 VSS.n1488 VSS.n1487 0.376971
R22559 VSS.n1390 VSS.n1388 0.376971
R22560 VSS.n1393 VSS.n1392 0.376971
R22561 VSS.n1400 VSS.n1396 0.376971
R22562 VSS.n509 VSS.n507 0.376971
R22563 VSS.n512 VSS.n511 0.376971
R22564 VSS.n1264 VSS.n1262 0.376971
R22565 VSS.n1267 VSS.n1266 0.376971
R22566 VSS.n1184 VSS.n1182 0.376971
R22567 VSS.n1187 VSS.n1186 0.376971
R22568 VSS.n977 VSS.n973 0.376971
R22569 VSS.n984 VSS.n980 0.376971
R22570 VSS.n816 VSS.n812 0.376971
R22571 VSS.n823 VSS.n819 0.376971
R22572 VSS.n1342 VSS.n1340 0.376971
R22573 VSS.n1304 VSS.n1303 0.376971
R22574 VSS.n1317 VSS.n1314 0.376971
R22575 VSS.n1934 VSS.n1933 0.376971
R22576 VSS.n1933 VSS.n1929 0.376971
R22577 VSS.n2126 VSS.n2122 0.376971
R22578 VSS.n2128 VSS.n2126 0.376971
R22579 VSS.n1768 VSS.n1762 0.376971
R22580 VSS.n1968 VSS.n1962 0.376971
R22581 VSS.n2356 VSS.n2355 0.366615
R22582 VSS.n302 VSS.n301 0.366615
R22583 VSS.n696 VSS.n695 0.366615
R22584 VSS.n2385 VSS.n2384 0.366119
R22585 VSS.n331 VSS.n330 0.366119
R22586 VSS.n665 VSS.n664 0.366119
R22587 VSS.n866 VSS.n865 0.337513
R22588 VSS.n857 VSS.n854 0.337513
R22589 VSS.n2363 VSS.n2362 0.334147
R22590 VSS.n309 VSS.n308 0.334147
R22591 VSS.n687 VSS.n686 0.334147
R22592 VSS.n2378 VSS.n2377 0.333652
R22593 VSS.n324 VSS.n323 0.333652
R22594 VSS.n672 VSS.n671 0.333652
R22595 VSS.n1592 VSS.n1591 0.324719
R22596 VSS.n222 VSS.n221 0.324719
R22597 VSS.n351 VSS.n350 0.324719
R22598 VSS.n2276 VSS.n2275 0.324719
R22599 VSS.n2405 VSS.n2404 0.324719
R22600 VSS.n1557 VSS.n1555 0.316384
R22601 VSS.n638 VSS.n636 0.316384
R22602 VSS VSS.n1058 0.313
R22603 VSS.n144 VSS.n143 0.298156
R22604 VSS.n601 VSS.n600 0.297854
R22605 VSS.n706 VSS.n705 0.297854
R22606 VSS.n2178 VSS.n2177 0.251319
R22607 VSS.n2270 VSS.n2269 0.251319
R22608 VSS.n378 VSS.n377 0.251319
R22609 VSS.n2208 VSS.n2207 0.251319
R22610 VSS.n2238 VSS.n2237 0.251319
R22611 VSS.n1719 VSS.n1718 0.251319
R22612 VSS.n1294 VSS.n1293 0.234094
R22613 VSS.n17 VSS.n16 0.23152
R22614 VSS.n2327 VSS.n2311 0.229427
R22615 VSS.n2327 VSS.n2326 0.229427
R22616 VSS.n273 VSS.n257 0.229427
R22617 VSS.n273 VSS.n272 0.229427
R22618 VSS.n480 VSS.n463 0.229427
R22619 VSS.n480 VSS.n479 0.229427
R22620 VSS.n1155 VSS.n1129 0.229427
R22621 VSS.n1155 VSS.n1154 0.229427
R22622 VSS.n1235 VSS.n1219 0.229427
R22623 VSS.n1235 VSS.n1234 0.229427
R22624 VSS.n2329 VSS.n2327 0.191391
R22625 VSS.n275 VSS.n273 0.191391
R22626 VSS.n1237 VSS.n1235 0.191391
R22627 VSS.n1157 VSS.n1155 0.191391
R22628 VSS.n482 VSS.n480 0.191391
R22629 VSS.n2372 VSS.n2370 0.190717
R22630 VSS.n318 VSS.n316 0.190717
R22631 VSS.n474 VSS.n467 0.190717
R22632 VSS.n1149 VSS.n1142 0.190717
R22633 VSS.n1142 VSS.n1139 0.190717
R22634 VSS.n985 VSS.n978 0.190717
R22635 VSS.n681 VSS.n679 0.190717
R22636 VSS.n824 VSS.n817 0.190717
R22637 VSS.n2331 VSS.n2329 0.164777
R22638 VSS.n277 VSS.n275 0.164777
R22639 VSS.n1450 VSS.n1448 0.164777
R22640 VSS.n1239 VSS.n1237 0.164777
R22641 VSS.n1159 VSS.n1157 0.164777
R22642 VSS.n484 VSS.n482 0.164777
R22643 VSS.n914 VSS.n912 0.164777
R22644 VSS.n753 VSS.n751 0.164777
R22645 VSS.n2311 VSS.n2309 0.15935
R22646 VSS.n2326 VSS.n2325 0.15935
R22647 VSS.n257 VSS.n255 0.15935
R22648 VSS.n272 VSS.n271 0.15935
R22649 VSS.n1555 VSS.n1554 0.15935
R22650 VSS.n1446 VSS.n1445 0.15935
R22651 VSS.n463 VSS.n461 0.15935
R22652 VSS.n479 VSS.n478 0.15935
R22653 VSS.n1129 VSS.n1128 0.15935
R22654 VSS.n1154 VSS.n1153 0.15935
R22655 VSS.n1219 VSS.n1218 0.15935
R22656 VSS.n1234 VSS.n1233 0.15935
R22657 VSS.n910 VSS.n909 0.15935
R22658 VSS.n636 VSS.n634 0.15935
R22659 VSS.n749 VSS.n747 0.15935
R22660 VSS.n384 VSS.n383 0.15675
R22661 VSS.n1979 VSS.n1978 0.15307
R22662 VSS.n1100 VSS.n1099 0.148462
R22663 VSS.n2338 VSS.n2336 0.144522
R22664 VSS.n2345 VSS.n2343 0.144522
R22665 VSS.n2352 VSS.n2350 0.144522
R22666 VSS.n2359 VSS.n2357 0.144522
R22667 VSS.n2366 VSS.n2364 0.144522
R22668 VSS.n2379 VSS.n2376 0.144522
R22669 VSS.n2386 VSS.n2383 0.144522
R22670 VSS.n2452 VSS.n2445 0.144522
R22671 VSS.n2463 VSS.n2456 0.144522
R22672 VSS.n190 VSS.n183 0.144522
R22673 VSS.n201 VSS.n194 0.144522
R22674 VSS.n284 VSS.n282 0.144522
R22675 VSS.n291 VSS.n289 0.144522
R22676 VSS.n298 VSS.n296 0.144522
R22677 VSS.n305 VSS.n303 0.144522
R22678 VSS.n312 VSS.n310 0.144522
R22679 VSS.n325 VSS.n322 0.144522
R22680 VSS.n332 VSS.n329 0.144522
R22681 VSS.n1566 VSS.n1564 0.144522
R22682 VSS.n1573 VSS.n1571 0.144522
R22683 VSS.n1461 VSS.n1459 0.144522
R22684 VSS.n1472 VSS.n1470 0.144522
R22685 VSS.n1246 VSS.n1244 0.144522
R22686 VSS.n1253 VSS.n1251 0.144522
R22687 VSS.n1166 VSS.n1164 0.144522
R22688 VSS.n1173 VSS.n1171 0.144522
R22689 VSS.n491 VSS.n489 0.144522
R22690 VSS.n498 VSS.n496 0.144522
R22691 VSS.n925 VSS.n923 0.144522
R22692 VSS.n936 VSS.n934 0.144522
R22693 VSS.n947 VSS.n945 0.144522
R22694 VSS.n958 VSS.n956 0.144522
R22695 VSS.n969 VSS.n967 0.144522
R22696 VSS.n996 VSS.n989 0.144522
R22697 VSS.n647 VSS.n645 0.144522
R22698 VSS.n654 VSS.n652 0.144522
R22699 VSS.n661 VSS.n659 0.144522
R22700 VSS.n668 VSS.n666 0.144522
R22701 VSS.n675 VSS.n673 0.144522
R22702 VSS.n688 VSS.n685 0.144522
R22703 VSS.n764 VSS.n762 0.144522
R22704 VSS.n775 VSS.n773 0.144522
R22705 VSS.n786 VSS.n784 0.144522
R22706 VSS.n797 VSS.n795 0.144522
R22707 VSS.n808 VSS.n806 0.144522
R22708 VSS.n835 VSS.n828 0.144522
R22709 VSS.n1981 VSS.n1973 0.144522
R22710 VSS.n1781 VSS.n1773 0.144522
R22711 VSS.n2154 VSS.n2153 0.141906
R22712 VSS.n1559 VSS.n1557 0.141804
R22713 VSS.n640 VSS.n638 0.141804
R22714 VSS.n2396 VSS.n2395 0.125448
R22715 VSS.n342 VSS.n341 0.125448
R22716 VSS.n1578 VSS.n1577 0.125448
R22717 VSS.n503 VSS.n502 0.125448
R22718 VSS.n1258 VSS.n1257 0.125448
R22719 VSS.n1178 VSS.n1177 0.125448
R22720 VSS.n2393 VSS.n2390 0.122443
R22721 VSS.n2470 VSS.n2467 0.122443
R22722 VSS.n208 VSS.n205 0.122443
R22723 VSS.n339 VSS.n336 0.122443
R22724 VSS.n1596 VSS.n1595 0.113781
R22725 VSS.n1619 VSS.n1618 0.113781
R22726 VSS.n1001 VSS.n1000 0.106563
R22727 VSS.n693 VSS.n692 0.106563
R22728 VSS.n840 VSS.n839 0.106563
R22729 VSS.n1533 VSS.n1532 0.0902327
R22730 VSS.n1502 VSS.n1501 0.0902327
R22731 VSS.n527 VSS.n526 0.0902327
R22732 VSS.n1281 VSS.n1280 0.0902327
R22733 VSS.n1201 VSS.n1200 0.0902327
R22734 VSS.n2501 VSS.n2495 0.0861908
R22735 VSS.n1614 VSS.n1376 0.0861908
R22736 VSS.n2502 VSS.n2501 0.0777426
R22737 VSS.n410 VSS.n409 0.07529
R22738 VSS.n1615 VSS.n1352 0.0740544
R22739 VSS.n1582 VSS.n1540 0.0699908
R22740 VSS.n1484 VSS.n1431 0.0699908
R22741 VSS.n1346 VSS.n1344 0.0699908
R22742 VSS.n1289 VSS.n1288 0.0695895
R22743 VSS.n1513 VSS.n1512 0.0695894
R22744 VSS.n1600 VSS.n1599 0.0683603
R22745 VSS.n1615 VSS.n1614 0.0683603
R22746 VSS.n1406 VSS.n1405 0.0679423
R22747 VSS.n1323 VSS.n1322 0.0676044
R22748 VSS.n1059 VSS 0.066125
R22749 VSS VSS.n2507 0.066125
R22750 VSS.n1209 VSS.n1208 0.0638939
R22751 VSS.n535 VSS.n534 0.0638939
R22752 VSS.n2502 VSS.n2490 0.0636644
R22753 VSS.n575 VSS.n574 0.0618569
R22754 VSS.n608 VSS.n607 0.0618569
R22755 VSS.n709 VSS.n708 0.0618569
R22756 VSS.n878 VSS.n877 0.0615154
R22757 VSS.n2180 VSS.n2174 0.0611815
R22758 VSS.n2272 VSS.n2264 0.0611815
R22759 VSS.n2480 VSS.n2433 0.0611815
R22760 VSS.n218 VSS.n172 0.0611815
R22761 VSS.n380 VSS.n371 0.0611815
R22762 VSS.n2240 VSS.n2234 0.0611815
R22763 VSS.n1721 VSS.n1715 0.0611815
R22764 VSS.n2210 VSS.n2204 0.0608398
R22765 VSS.n2401 VSS.n2296 0.0608398
R22766 VSS.n347 VSS.n242 0.0608398
R22767 VSS.n1329 VSS.n1328 0.0604712
R22768 VSS.n1712 VSS.n1711 0.0584854
R22769 VSS.n2171 VSS.n2170 0.0584854
R22770 VSS.n2201 VSS.n2200 0.0584854
R22771 VSS.n2231 VSS.n2230 0.0584854
R22772 VSS.n2261 VSS.n2260 0.0584854
R22773 VSS.n2289 VSS.n2288 0.0584854
R22774 VSS.n2430 VSS.n2429 0.0584854
R22775 VSS.n169 VSS.n168 0.0584854
R22776 VSS.n235 VSS.n234 0.0584854
R22777 VSS.n368 VSS.n367 0.0584854
R22778 VSS.n2495 VSS.n2494 0.0566413
R22779 VSS.n1378 VSS.n1377 0.0566413
R22780 VSS.n1376 VSS.n1375 0.0566413
R22781 VSS.n579 VSS.n578 0.0565323
R22782 VSS.n882 VSS.n881 0.0565323
R22783 VSS.n612 VSS.n611 0.0565323
R22784 VSS.n721 VSS.n720 0.0565323
R22785 VSS.n425 VSS.n417 0.0558464
R22786 VSS.n1524 VSS.n1523 0.0547459
R22787 VSS.n1490 VSS.n1489 0.0547459
R22788 VSS.n518 VSS.n517 0.0547459
R22789 VSS.n1272 VSS.n1271 0.0547459
R22790 VSS.n1192 VSS.n1191 0.0547459
R22791 VSS.n6 VSS.n5 0.053
R22792 VSS.n588 VSS.n587 0.0526261
R22793 VSS.n587 VSS.n586 0.0526261
R22794 VSS.n895 VSS.n894 0.0526261
R22795 VSS.n894 VSS.n893 0.0526261
R22796 VSS.n621 VSS.n620 0.0526261
R22797 VSS.n620 VSS.n619 0.0526261
R22798 VSS.n734 VSS.n733 0.0526261
R22799 VSS.n733 VSS.n732 0.0526261
R22800 VSS.n425 VSS.n424 0.0502162
R22801 VSS.n1695 VSS.n1694 0.0497188
R22802 VSS.n37 VSS.n34 0.0493281
R22803 VSS.n46 VSS.n45 0.0493281
R22804 VSS.n55 VSS.n54 0.0493281
R22805 VSS VSS.n2483 0.0489375
R22806 VSS.n580 VSS.n579 0.0487198
R22807 VSS.n883 VSS.n882 0.0487198
R22808 VSS.n613 VSS.n612 0.0487198
R22809 VSS.n722 VSS.n721 0.0487198
R22810 VSS.n1624 VSS.n1623 0.0481562
R22811 VSS.n1711 VSS.n1710 0.0467667
R22812 VSS.n2170 VSS.n2169 0.0467667
R22813 VSS.n2200 VSS.n2199 0.0467667
R22814 VSS.n2230 VSS.n2229 0.0467667
R22815 VSS.n2260 VSS.n2259 0.0467667
R22816 VSS.n2288 VSS.n2287 0.0467667
R22817 VSS.n2429 VSS.n2428 0.0467667
R22818 VSS.n168 VSS.n167 0.0467667
R22819 VSS.n234 VSS.n233 0.0467667
R22820 VSS.n367 VSS.n366 0.0467667
R22821 VSS.n525 VSS.n524 0.0464244
R22822 VSS.n1199 VSS.n1198 0.0464244
R22823 VSS.n1500 VSS.n1499 0.0461141
R22824 VSS.n1531 VSS.n1530 0.0461141
R22825 VSS.n1419 VSS.n1418 0.0461141
R22826 VSS.n1279 VSS.n1278 0.045605
R22827 VSS.n1284 VSS.n1279 0.0454086
R22828 VSS.n2210 VSS.n2209 0.0449804
R22829 VSS.n2401 VSS.n2400 0.0449804
R22830 VSS.n347 VSS.n346 0.0449804
R22831 VSS.n1536 VSS.n1531 0.0448907
R22832 VSS.n1505 VSS.n1500 0.0448907
R22833 VSS.n1427 VSS.n1419 0.0448907
R22834 VSS.n1721 VSS.n1720 0.04464
R22835 VSS.n2180 VSS.n2179 0.04464
R22836 VSS.n2240 VSS.n2239 0.04464
R22837 VSS.n2272 VSS.n2271 0.04464
R22838 VSS.n2480 VSS.n2479 0.04464
R22839 VSS.n218 VSS.n217 0.04464
R22840 VSS.n380 VSS.n379 0.04464
R22841 VSS.n1204 VSS.n1199 0.0445792
R22842 VSS.n530 VSS.n525 0.0445792
R22843 VSS.n877 VSS.n876 0.0443642
R22844 VSS.n574 VSS.n573 0.0440244
R22845 VSS.n607 VSS.n606 0.0440244
R22846 VSS.n708 VSS.n707 0.0440244
R22847 VSS.n2368 VSS.n2366 0.0439783
R22848 VSS.n2376 VSS.n2374 0.0439783
R22849 VSS.n2445 VSS.n2443 0.0439783
R22850 VSS.n183 VSS.n181 0.0439783
R22851 VSS.n314 VSS.n312 0.0439783
R22852 VSS.n322 VSS.n320 0.0439783
R22853 VSS.n1405 VSS.n1403 0.0439783
R22854 VSS.n971 VSS.n969 0.0439783
R22855 VSS.n989 VSS.n987 0.0439783
R22856 VSS.n677 VSS.n675 0.0439783
R22857 VSS.n685 VSS.n683 0.0439783
R22858 VSS.n810 VSS.n808 0.0439783
R22859 VSS.n828 VSS.n826 0.0439783
R22860 VSS.n1322 VSS.n1320 0.0439783
R22861 VSS.n1973 VSS.n1971 0.0439783
R22862 VSS.n1773 VSS.n1771 0.0439783
R22863 VSS.n1021 VSS.n1020 0.0434688
R22864 VSS.n1020 VSS.n1019 0.0434688
R22865 VSS.n1019 VSS.n1018 0.0434688
R22866 VSS.n1018 VSS.n1017 0.0434688
R22867 VSS.n1017 VSS.n1016 0.0434688
R22868 VSS.n1016 VSS.n1015 0.0434688
R22869 VSS.n1013 VSS.n568 0.0434688
R22870 VSS.n1082 VSS.n568 0.0434688
R22871 VSS.n1082 VSS.n1081 0.0434688
R22872 VSS.n1081 VSS.n1080 0.0434688
R22873 VSS.n1080 VSS.n1079 0.0434688
R22874 VSS.n1079 VSS.n1078 0.0434688
R22875 VSS.n1078 VSS.n1077 0.0434688
R22876 VSS.n1071 VSS.n1070 0.0434688
R22877 VSS.n1626 VSS.n1625 0.0434688
R22878 VSS.n1627 VSS.n1626 0.0434688
R22879 VSS.n1629 VSS.n1628 0.0434688
R22880 VSS.n1112 VSS.n1111 0.0434688
R22881 VSS.n1215 VSS.n1214 0.0434688
R22882 VSS.n386 VSS.n385 0.0434688
R22883 VSS.n387 VSS.n386 0.0434688
R22884 VSS.n388 VSS.n387 0.0434688
R22885 VSS.n389 VSS.n388 0.0434688
R22886 VSS.n392 VSS.n391 0.0434688
R22887 VSS.n393 VSS.n392 0.0434688
R22888 VSS.n394 VSS.n393 0.0434688
R22889 VSS.n395 VSS.n394 0.0434688
R22890 VSS.n396 VSS.n395 0.0434688
R22891 VSS.n397 VSS.n396 0.0434688
R22892 VSS.n1680 VSS.n1679 0.0434688
R22893 VSS.n1681 VSS.n1680 0.0434688
R22894 VSS.n1682 VSS.n1681 0.0434688
R22895 VSS.n1683 VSS.n1682 0.0434688
R22896 VSS.n1684 VSS.n1683 0.0434688
R22897 VSS.n1685 VSS.n1684 0.0434688
R22898 VSS.n1688 VSS.n1687 0.0434688
R22899 VSS.n1689 VSS.n1688 0.0434688
R22900 VSS.n1690 VSS.n1689 0.0434688
R22901 VSS.n1691 VSS.n1690 0.0434688
R22902 VSS.n1692 VSS.n1691 0.0434688
R22903 VSS.n1693 VSS.n1692 0.0434688
R22904 VSS.n390 VSS.n389 0.0426875
R22905 VSS.n1495 VSS.n1494 0.0419945
R22906 VSS.n1113 VSS.n1112 0.0419063
R22907 VSS.n26 VSS.n20 0.0415156
R22908 VSS.n2309 VSS.n2307 0.0412609
R22909 VSS.n2325 VSS.n2323 0.0412609
R22910 VSS.n255 VSS.n253 0.0412609
R22911 VSS.n271 VSS.n269 0.0412609
R22912 VSS.n1554 VSS.n1552 0.0412609
R22913 VSS.n1445 VSS.n1443 0.0412609
R22914 VSS.n461 VSS.n459 0.0412609
R22915 VSS.n478 VSS.n476 0.0412609
R22916 VSS.n1128 VSS.n1126 0.0412609
R22917 VSS.n1153 VSS.n1151 0.0412609
R22918 VSS.n1233 VSS.n1231 0.0412609
R22919 VSS.n909 VSS.n907 0.0412609
R22920 VSS.n634 VSS.n632 0.0412609
R22921 VSS.n747 VSS.n745 0.0412609
R22922 VSS.n445 VSS.n444 0.041125
R22923 VSS.n2361 VSS.n2359 0.0385435
R22924 VSS.n2383 VSS.n2381 0.0385435
R22925 VSS.n2456 VSS.n2454 0.0385435
R22926 VSS.n194 VSS.n192 0.0385435
R22927 VSS.n307 VSS.n305 0.0385435
R22928 VSS.n329 VSS.n327 0.0385435
R22929 VSS.n960 VSS.n958 0.0385435
R22930 VSS.n1000 VSS.n998 0.0385435
R22931 VSS.n670 VSS.n668 0.0385435
R22932 VSS.n692 VSS.n690 0.0385435
R22933 VSS.n799 VSS.n797 0.0385435
R22934 VSS.n839 VSS.n837 0.0385435
R22935 VSS.n385 VSS.n384 0.038
R22936 VSS.n1694 VSS.n1693 0.038
R22937 VSS.n1069 VSS.n1068 0.0372187
R22938 VSS.n1679 VSS.n428 0.0372187
R22939 VSS.n1630 VSS.n1629 0.0356562
R22940 VSS.n439 VSS.n438 0.0356562
R22941 VSS.n19 VSS.n18 0.0356562
R22942 VSS.n54 VSS.n53 0.0356562
R22943 VSS.n1625 VSS.n1624 0.034875
R22944 VSS.n1295 VSS.n1294 0.034875
R22945 VSS.n1686 VSS.n1685 0.0340938
R22946 VSS.n2354 VSS.n2352 0.0331087
R22947 VSS.n2390 VSS.n2388 0.0331087
R22948 VSS.n2467 VSS.n2465 0.0331087
R22949 VSS.n205 VSS.n203 0.0331087
R22950 VSS.n300 VSS.n298 0.0331087
R22951 VSS.n336 VSS.n334 0.0331087
R22952 VSS.n949 VSS.n947 0.0331087
R22953 VSS.n663 VSS.n661 0.0331087
R22954 VSS.n788 VSS.n786 0.0331087
R22955 VSS.n1072 VSS.n1071 0.0325312
R22956 VSS.n63 VSS.n62 0.03175
R22957 VSS.n9 VSS.n8 0.03175
R22958 VSS.n13 VSS.n12 0.03175
R22959 VSS.n1023 VSS.n1022 0.0309688
R22960 VSS.n1015 VSS.n1014 0.0309688
R22961 VSS.n410 VSS.n408 0.0306452
R22962 VSS.n520 VSS.n516 0.0304205
R22963 VSS.n1194 VSS.n1190 0.0304205
R22964 VSS.n2336 VSS.n2333 0.0303913
R22965 VSS.n282 VSS.n279 0.0303913
R22966 VSS.n1564 VSS.n1561 0.0303913
R22967 VSS.n1459 VSS.n1452 0.0303913
R22968 VSS.n1244 VSS.n1241 0.0303913
R22969 VSS.n1164 VSS.n1161 0.0303913
R22970 VSS.n489 VSS.n486 0.0303913
R22971 VSS.n923 VSS.n916 0.0303913
R22972 VSS.n645 VSS.n642 0.0303913
R22973 VSS.n762 VSS.n755 0.0303913
R22974 VSS.n1022 VSS.n1021 0.0301875
R22975 VSS.n1068 VSS.n1067 0.0301875
R22976 VSS.n1337 VSS.n1329 0.0301368
R22977 VSS.n1707 VSS.n1706 0.0297969
R22978 VSS.n2166 VSS.n2165 0.0297969
R22979 VSS.n2196 VSS.n2195 0.0297969
R22980 VSS.n2226 VSS.n2225 0.0297969
R22981 VSS.n2256 VSS.n2255 0.0297969
R22982 VSS.n2280 VSS.n2279 0.0297969
R22983 VSS.n2417 VSS.n2416 0.0297969
R22984 VSS.n164 VSS.n163 0.0297969
R22985 VSS.n226 VSS.n225 0.0297969
R22986 VSS.n363 VSS.n362 0.0297969
R22987 VSS.n3 VSS.n2 0.02925
R22988 VSS.n1324 VSS.n1323 0.0288505
R22989 VSS.n1274 VSS.n1270 0.0288505
R22990 VSS.n1526 VSS.n1522 0.0285117
R22991 VSS.n1414 VSS.n1406 0.0285117
R22992 VSS.n1726 VSS.n1725 0.0282778
R22993 VSS.n1727 VSS.n1726 0.0282778
R22994 VSS.n1728 VSS.n1727 0.0282778
R22995 VSS.n1729 VSS.n1728 0.0282778
R22996 VSS.n1730 VSS.n1729 0.0282778
R22997 VSS.n1731 VSS.n1730 0.0282778
R22998 VSS.n1732 VSS.n1731 0.0282778
R22999 VSS.n1733 VSS.n1732 0.0282778
R23000 VSS.n1734 VSS.n1733 0.0282778
R23001 VSS.n1735 VSS.n1734 0.0282778
R23002 VSS.n1736 VSS.n1735 0.0282778
R23003 VSS.n2138 VSS.n2137 0.0282778
R23004 VSS.n2139 VSS.n2138 0.0282778
R23005 VSS.n2140 VSS.n2139 0.0282778
R23006 VSS.n2141 VSS.n2140 0.0282778
R23007 VSS.n2142 VSS.n2141 0.0282778
R23008 VSS.n2143 VSS.n2142 0.0282778
R23009 VSS.n2144 VSS.n2143 0.0282778
R23010 VSS.n2145 VSS.n2144 0.0282778
R23011 VSS.n2146 VSS.n2145 0.0282778
R23012 VSS.n2147 VSS.n2146 0.0282778
R23013 VSS.n2148 VSS.n2147 0.0282778
R23014 VSS.n2149 VSS.n2148 0.0282778
R23015 VSS.n66 VSS.n65 0.028
R23016 VSS.n537 VSS.n536 0.0278438
R23017 VSS.n45 VSS.n44 0.0278438
R23018 VSS.n2347 VSS.n2345 0.0276739
R23019 VSS.n293 VSS.n291 0.0276739
R23020 VSS.n938 VSS.n936 0.0276739
R23021 VSS.n656 VSS.n654 0.0276739
R23022 VSS.n777 VSS.n775 0.0276739
R23023 VSS.n2 VSS.n1 0.02675
R23024 VSS.n65 VSS.n13 0.02675
R23025 VSS.n2136 VSS.n1736 0.0267346
R23026 VSS.n31 VSS.n28 0.0258906
R23027 VSS.n540 VSS.n539 0.0255
R23028 VSS.n1209 VSS.n1181 0.0250149
R23029 VSS.n535 VSS.n506 0.0250149
R23030 VSS.n2343 VSS.n2340 0.0249565
R23031 VSS.n289 VSS.n286 0.0249565
R23032 VSS.n1571 VSS.n1568 0.0249565
R23033 VSS.n1575 VSS.n1573 0.0249565
R23034 VSS.n1470 VSS.n1463 0.0249565
R23035 VSS.n1474 VSS.n1472 0.0249565
R23036 VSS.n1251 VSS.n1248 0.0249565
R23037 VSS.n1255 VSS.n1253 0.0249565
R23038 VSS.n1171 VSS.n1168 0.0249565
R23039 VSS.n1175 VSS.n1173 0.0249565
R23040 VSS.n496 VSS.n493 0.0249565
R23041 VSS.n500 VSS.n498 0.0249565
R23042 VSS.n934 VSS.n927 0.0249565
R23043 VSS.n652 VSS.n649 0.0249565
R23044 VSS.n773 VSS.n766 0.0249565
R23045 VSS.n2134 VSS.n2130 0.0248056
R23046 VSS.n592 VSS.n591 0.0239375
R23047 VSS.n1002 VSS.n1001 0.0239375
R23048 VSS.n694 VSS.n693 0.0239375
R23049 VSS.n841 VSS.n840 0.0239375
R23050 VSS.n33 VSS.n32 0.0239375
R23051 VSS.n2135 VSS.n1936 0.0234167
R23052 VSS.n142 VSS.n139 0.0232776
R23053 VSS.n12 VSS.n11 0.023
R23054 VSS.n2150 VSS.n2149 0.0228765
R23055 VSS.n406 VSS.n405 0.022459
R23056 VSS.n1638 VSS.n1637 0.0223109
R23057 VSS.n2340 VSS.n2338 0.0222391
R23058 VSS.n286 VSS.n284 0.0222391
R23059 VSS.n1568 VSS.n1566 0.0222391
R23060 VSS.n1576 VSS.n1575 0.0222391
R23061 VSS.n1463 VSS.n1461 0.0222391
R23062 VSS.n1475 VSS.n1474 0.0222391
R23063 VSS.n1248 VSS.n1246 0.0222391
R23064 VSS.n1256 VSS.n1255 0.0222391
R23065 VSS.n1168 VSS.n1166 0.0222391
R23066 VSS.n1176 VSS.n1175 0.0222391
R23067 VSS.n493 VSS.n491 0.0222391
R23068 VSS.n501 VSS.n500 0.0222391
R23069 VSS.n927 VSS.n925 0.0222391
R23070 VSS.n649 VSS.n647 0.0222391
R23071 VSS.n766 VSS.n764 0.0222391
R23072 VSS.n408 VSS.n407 0.0219844
R23073 VSS.n1539 VSS.n1538 0.0219844
R23074 VSS.n1528 VSS.n1527 0.0219844
R23075 VSS.n1511 VSS.n1507 0.0219844
R23076 VSS.n1497 VSS.n1496 0.0219844
R23077 VSS.n1430 VSS.n1429 0.0219844
R23078 VSS.n1416 VSS.n1415 0.0219844
R23079 VSS.n1287 VSS.n1286 0.0219844
R23080 VSS.n1276 VSS.n1275 0.0219844
R23081 VSS.n1207 VSS.n1206 0.0219844
R23082 VSS.n1196 VSS.n1195 0.0219844
R23083 VSS.n533 VSS.n532 0.0219844
R23084 VSS.n522 VSS.n521 0.0219844
R23085 VSS.n1343 VSS.n1339 0.0219844
R23086 VSS.n1326 VSS.n1325 0.0219844
R23087 VSS.n42 VSS.n38 0.0219844
R23088 VSS.n64 VSS.n56 0.0219844
R23089 VSS.n10 VSS.n9 0.02175
R23090 VSS.n1077 VSS.n1076 0.0208125
R23091 VSS.n1710 VSS.n1709 0.0205304
R23092 VSS.n2199 VSS.n2198 0.0205304
R23093 VSS.n2229 VSS.n2228 0.0205304
R23094 VSS.n2287 VSS.n2286 0.0205304
R23095 VSS.n233 VSS.n232 0.0205304
R23096 VSS.n366 VSS.n365 0.0205304
R23097 VSS.n4 VSS.n3 0.0205
R23098 VSS.n1012 VSS.n895 0.0204768
R23099 VSS.n700 VSS.n621 0.0204759
R23100 VSS.n851 VSS.n734 0.0204759
R23101 VSS.n597 VSS.n588 0.020474
R23102 VSS.n2399 VSS.n2394 0.0200312
R23103 VSS.n2478 VSS.n2471 0.0200312
R23104 VSS.n216 VSS.n209 0.0200312
R23105 VSS.n345 VSS.n340 0.0200312
R23106 VSS.n585 VSS.n580 0.0200312
R23107 VSS.n892 VSS.n883 0.0200312
R23108 VSS.n618 VSS.n613 0.0200312
R23109 VSS.n731 VSS.n722 0.0200312
R23110 VSS.n34 VSS.n33 0.0200312
R23111 VSS.n56 VSS.n55 0.0200312
R23112 VSS.n2350 VSS.n2347 0.0195217
R23113 VSS.n296 VSS.n293 0.0195217
R23114 VSS.n945 VSS.n938 0.0195217
R23115 VSS.n659 VSS.n656 0.0195217
R23116 VSS.n784 VSS.n777 0.0195217
R23117 VSS.n1988 VSS.n1985 0.0191458
R23118 VSS.n1289 VSS.n1261 0.0188525
R23119 VSS.n1581 VSS.n1576 0.0188424
R23120 VSS.n1483 VSS.n1475 0.0188424
R23121 VSS.n1261 VSS.n1256 0.0188424
R23122 VSS.n1181 VSS.n1176 0.0188424
R23123 VSS.n506 VSS.n501 0.0188424
R23124 VSS.n1788 VSS.n1785 0.0185819
R23125 VSS.n1582 VSS.n1581 0.0184465
R23126 VSS.n1484 VSS.n1483 0.0184465
R23127 VSS.n1985 VSS.n1983 0.018314
R23128 VSS.n1715 VSS.n1714 0.0180781
R23129 VSS.n2174 VSS.n2173 0.0180781
R23130 VSS.n2169 VSS.n2168 0.0180781
R23131 VSS.n2204 VSS.n2203 0.0180781
R23132 VSS.n2234 VSS.n2233 0.0180781
R23133 VSS.n2264 VSS.n2263 0.0180781
R23134 VSS.n2259 VSS.n2258 0.0180781
R23135 VSS.n2296 VSS.n2295 0.0180781
R23136 VSS.n2433 VSS.n2432 0.0180781
R23137 VSS.n2428 VSS.n2427 0.0180781
R23138 VSS.n172 VSS.n171 0.0180781
R23139 VSS.n167 VSS.n166 0.0180781
R23140 VSS.n242 VSS.n241 0.0180781
R23141 VSS.n371 VSS.n370 0.0180781
R23142 VSS.n417 VSS.n416 0.0180781
R23143 VSS.n52 VSS.n47 0.0180781
R23144 VSS.n8 VSS.n7 0.018
R23145 VSS.n1586 VSS.n1585 0.0176875
R23146 VSS.n1595 VSS.n1594 0.0176875
R23147 VSS.n1291 VSS.n1290 0.0176875
R23148 VSS.n1066 VSS.n1065 0.0169062
R23149 VSS.n1062 VSS.n1061 0.0169062
R23150 VSS.n2333 VSS.n2331 0.0168043
R23151 VSS.n279 VSS.n277 0.0168043
R23152 VSS.n1561 VSS.n1559 0.0168043
R23153 VSS.n1452 VSS.n1450 0.0168043
R23154 VSS.n1241 VSS.n1239 0.0168043
R23155 VSS.n1161 VSS.n1159 0.0168043
R23156 VSS.n486 VSS.n484 0.0168043
R23157 VSS.n916 VSS.n914 0.0168043
R23158 VSS.n642 VSS.n640 0.0168043
R23159 VSS.n755 VSS.n753 0.0168043
R23160 VSS.n576 VSS.n575 0.016125
R23161 VSS.n879 VSS.n878 0.016125
R23162 VSS.n609 VSS.n608 0.016125
R23163 VSS.n718 VSS.n709 0.016125
R23164 VSS.n538 VSS.n537 0.016125
R23165 VSS.n47 VSS.n46 0.016125
R23166 VSS.n53 VSS.n52 0.016125
R23167 VSS.n398 VSS.n397 0.016125
R23168 VSS.n7 VSS.n6 0.0155
R23169 VSS.n1210 VSS.n1114 0.0153437
R23170 VSS.n1647 VSS.n431 0.0143978
R23171 VSS.n1648 VSS.n1647 0.0143978
R23172 VSS.n1649 VSS.n1648 0.0143978
R23173 VSS.n1650 VSS.n1649 0.0143978
R23174 VSS.n1653 VSS.n1652 0.0143978
R23175 VSS.n1654 VSS.n1653 0.0143978
R23176 VSS.n1655 VSS.n1654 0.0143978
R23177 VSS.n1656 VSS.n1655 0.0143978
R23178 VSS.n1657 VSS.n1656 0.0143978
R23179 VSS.n1658 VSS.n1657 0.0143978
R23180 VSS.n1678 VSS.n1660 0.0143978
R23181 VSS.n1678 VSS.n1677 0.0143978
R23182 VSS.n1677 VSS.n1676 0.0143978
R23183 VSS.n1676 VSS.n1675 0.0143978
R23184 VSS.n1675 VSS.n1674 0.0143978
R23185 VSS.n1674 VSS.n1673 0.0143978
R23186 VSS.n1673 VSS.n1672 0.0143978
R23187 VSS.n1670 VSS.n1669 0.0143978
R23188 VSS.n1669 VSS.n1668 0.0143978
R23189 VSS.n1668 VSS.n1667 0.0143978
R23190 VSS.n1667 VSS.n1666 0.0143978
R23191 VSS.n1666 VSS.n1665 0.0143978
R23192 VSS.n1665 VSS.n1664 0.0143978
R23193 VSS.n565 VSS.n564 0.0143978
R23194 VSS.n564 VSS.n563 0.0143978
R23195 VSS.n563 VSS.n562 0.0143978
R23196 VSS.n562 VSS.n561 0.0143978
R23197 VSS.n561 VSS.n560 0.0143978
R23198 VSS.n558 VSS.n557 0.0143978
R23199 VSS.n1084 VSS.n1083 0.0143978
R23200 VSS.n1085 VSS.n1084 0.0143978
R23201 VSS.n1086 VSS.n1085 0.0143978
R23202 VSS.n1087 VSS.n1086 0.0143978
R23203 VSS.n1088 VSS.n1087 0.0143978
R23204 VSS.n1091 VSS.n1090 0.0143978
R23205 VSS.n1097 VSS.n1091 0.0143978
R23206 VSS.n1633 VSS.n1301 0.0143978
R23207 VSS.n1633 VSS.n1632 0.0143978
R23208 VSS.n435 VSS.n434 0.0143978
R23209 VSS.n545 VSS.n435 0.0143978
R23210 VSS.n545 VSS.n544 0.0143978
R23211 VSS.n448 VSS.n447 0.0143978
R23212 VSS.n442 VSS.n441 0.0143978
R23213 VSS.n1109 VSS.n1108 0.0143978
R23214 VSS.n1110 VSS.n1109 0.0143978
R23215 VSS.n1213 VSS.n1212 0.0143978
R23216 VSS.n1720 VSS.n1719 0.0141719
R23217 VSS.n2179 VSS.n2178 0.0141719
R23218 VSS.n2209 VSS.n2208 0.0141719
R23219 VSS.n2239 VSS.n2238 0.0141719
R23220 VSS.n2271 VSS.n2270 0.0141719
R23221 VSS.n2394 VSS.n2393 0.0141719
R23222 VSS.n2400 VSS.n2399 0.0141719
R23223 VSS.n2471 VSS.n2470 0.0141719
R23224 VSS.n2479 VSS.n2478 0.0141719
R23225 VSS.n209 VSS.n208 0.0141719
R23226 VSS.n217 VSS.n216 0.0141719
R23227 VSS.n340 VSS.n339 0.0141719
R23228 VSS.n346 VSS.n345 0.0141719
R23229 VSS.n379 VSS.n378 0.0141719
R23230 VSS.n424 VSS.n423 0.0141719
R23231 VSS.n1537 VSS.n1536 0.0141719
R23232 VSS.n1506 VSS.n1505 0.0141719
R23233 VSS.n1428 VSS.n1427 0.0141719
R23234 VSS.n1285 VSS.n1284 0.0141719
R23235 VSS.n1205 VSS.n1204 0.0141719
R23236 VSS.n531 VSS.n530 0.0141719
R23237 VSS.n586 VSS.n585 0.0141719
R23238 VSS.n893 VSS.n892 0.0141719
R23239 VSS.n619 VSS.n618 0.0141719
R23240 VSS.n732 VSS.n731 0.0141719
R23241 VSS.n1338 VSS.n1337 0.0141719
R23242 VSS.n27 VSS.n26 0.0141719
R23243 VSS.n1651 VSS.n1650 0.0141452
R23244 VSS.n543 VSS.n448 0.0141452
R23245 VSS.n2357 VSS.n2354 0.014087
R23246 VSS.n2388 VSS.n2386 0.014087
R23247 VSS.n2465 VSS.n2463 0.014087
R23248 VSS.n203 VSS.n201 0.014087
R23249 VSS.n303 VSS.n300 0.014087
R23250 VSS.n334 VSS.n332 0.014087
R23251 VSS.n956 VSS.n949 0.014087
R23252 VSS.n666 VSS.n663 0.014087
R23253 VSS.n795 VSS.n788 0.014087
R23254 VSS.n446 VSS.n442 0.0136398
R23255 VSS.n1014 VSS.n1013 0.013
R23256 VSS.n1791 VSS.n1790 0.013
R23257 VSS.n1810 VSS.n1809 0.013
R23258 VSS.n1821 VSS.n1820 0.013
R23259 VSS.n1833 VSS.n1832 0.013
R23260 VSS.n1844 VSS.n1843 0.013
R23261 VSS.n1856 VSS.n1855 0.013
R23262 VSS.n1867 VSS.n1866 0.013
R23263 VSS.n1879 VSS.n1878 0.013
R23264 VSS.n1890 VSS.n1889 0.013
R23265 VSS.n1902 VSS.n1901 0.013
R23266 VSS.n1913 VSS.n1912 0.013
R23267 VSS.n1926 VSS.n1925 0.013
R23268 VSS.n2120 VSS.n2119 0.013
R23269 VSS.n2107 VSS.n2106 0.013
R23270 VSS.n2096 VSS.n2095 0.013
R23271 VSS.n2084 VSS.n2083 0.013
R23272 VSS.n2073 VSS.n2072 0.013
R23273 VSS.n2061 VSS.n2060 0.013
R23274 VSS.n2050 VSS.n2049 0.013
R23275 VSS.n2038 VSS.n2037 0.013
R23276 VSS.n2027 VSS.n2026 0.013
R23277 VSS.n2015 VSS.n2014 0.013
R23278 VSS.n2004 VSS.n2003 0.013
R23279 VSS.n1992 VSS.n1991 0.013
R23280 VSS.n5 VSS.n4 0.013
R23281 VSS.n431 VSS.n430 0.012629
R23282 VSS.n1664 VSS.n1663 0.012629
R23283 VSS.n1076 VSS.n1075 0.012435
R23284 VSS.n1060 VSS.n1059 0.0124292
R23285 VSS.n1064 VSS.n1063 0.0124292
R23286 VSS.n1089 VSS.n1088 0.0123763
R23287 VSS.n1096 VSS.n1095 0.0123763
R23288 VSS.n1714 VSS.n1713 0.0122188
R23289 VSS.n1708 VSS.n1707 0.0122188
R23290 VSS.n2167 VSS.n2166 0.0122188
R23291 VSS.n2203 VSS.n2202 0.0122188
R23292 VSS.n2197 VSS.n2196 0.0122188
R23293 VSS.n2233 VSS.n2232 0.0122188
R23294 VSS.n2227 VSS.n2226 0.0122188
R23295 VSS.n2257 VSS.n2256 0.0122188
R23296 VSS.n2295 VSS.n2290 0.0122188
R23297 VSS.n2285 VSS.n2280 0.0122188
R23298 VSS.n2426 VSS.n2417 0.0122188
R23299 VSS.n165 VSS.n164 0.0122188
R23300 VSS.n241 VSS.n236 0.0122188
R23301 VSS.n231 VSS.n226 0.0122188
R23302 VSS.n370 VSS.n369 0.0122188
R23303 VSS.n364 VSS.n363 0.0122188
R23304 VSS.n407 VSS.n406 0.0122188
R23305 VSS.n1529 VSS.n1528 0.0122188
R23306 VSS.n1498 VSS.n1497 0.0122188
R23307 VSS.n1417 VSS.n1416 0.0122188
R23308 VSS.n1277 VSS.n1276 0.0122188
R23309 VSS.n1197 VSS.n1196 0.0122188
R23310 VSS.n523 VSS.n522 0.0122188
R23311 VSS.n1327 VSS.n1326 0.0122188
R23312 VSS.n38 VSS.n37 0.0122188
R23313 VSS.n43 VSS.n42 0.0122188
R23314 VSS.n44 VSS.n43 0.0122188
R23315 VSS.n64 VSS.n63 0.0122188
R23316 VSS.n1597 VSS.n1596 0.0118907
R23317 VSS.n1348 VSS.n1347 0.0118907
R23318 VSS.n440 VSS.n436 0.011871
R23319 VSS.n1297 VSS.n1296 0.0116183
R23320 VSS.n1935 VSS.n1926 0.0116111
R23321 VSS.n2129 VSS.n2120 0.0116111
R23322 VSS.n1073 VSS.n1072 0.0114375
R23323 VSS.n427 VSS.n426 0.0114375
R23324 VSS.n1672 VSS.n1671 0.0113656
R23325 VSS.n1924 VSS.n1913 0.0109167
R23326 VSS.n2118 VSS.n2107 0.0109167
R23327 VSS.n1659 VSS.n1658 0.0108602
R23328 VSS.n2172 VSS.n2171 0.010758
R23329 VSS.n2262 VSS.n2261 0.010758
R23330 VSS.n2431 VSS.n2430 0.010758
R23331 VSS.n170 VSS.n169 0.010758
R23332 VSS.n881 VSS.n880 0.0107521
R23333 VSS.n611 VSS.n610 0.0107521
R23334 VSS.n720 VSS.n719 0.0107521
R23335 VSS.n11 VSS.n10 0.0105
R23336 VSS.n88 VSS.n87 0.0104225
R23337 VSS.n560 VSS.n559 0.0103548
R23338 VSS.n1538 VSS.n1537 0.0102656
R23339 VSS.n1527 VSS.n1526 0.0102656
R23340 VSS.n1507 VSS.n1506 0.0102656
R23341 VSS.n1496 VSS.n1495 0.0102656
R23342 VSS.n1429 VSS.n1428 0.0102656
R23343 VSS.n1415 VSS.n1414 0.0102656
R23344 VSS.n1286 VSS.n1285 0.0102656
R23345 VSS.n1275 VSS.n1274 0.0102656
R23346 VSS.n1206 VSS.n1205 0.0102656
R23347 VSS.n1195 VSS.n1194 0.0102656
R23348 VSS.n532 VSS.n531 0.0102656
R23349 VSS.n521 VSS.n520 0.0102656
R23350 VSS.n596 VSS.n592 0.0102656
R23351 VSS.n1011 VSS.n1002 0.0102656
R23352 VSS.n699 VSS.n694 0.0102656
R23353 VSS.n850 VSS.n841 0.0102656
R23354 VSS.n1339 VSS.n1338 0.0102656
R23355 VSS.n1325 VSS.n1324 0.0102656
R23356 VSS.n1911 VSS.n1902 0.0102222
R23357 VSS.n2105 VSS.n2096 0.0102222
R23358 VSS.n554 VSS.n553 0.0101021
R23359 VSS.n1095 VSS.n1094 0.0101021
R23360 VSS.n1687 VSS.n1686 0.009875
R23361 VSS.n577 VSS.n576 0.00987154
R23362 VSS.n578 VSS.n577 0.00967578
R23363 VSS.n1598 VSS.n1387 0.00962927
R23364 VSS.n1617 VSS.n1616 0.00962927
R23365 VSS.n1212 VSS.n1211 0.00959677
R23366 VSS.n1591 VSS.n1590 0.00957737
R23367 VSS.n1590 VSS.n1589 0.00957737
R23368 VSS.n1024 VSS.n1023 0.00957737
R23369 VSS.n1025 VSS.n1024 0.00957737
R23370 VSS.n1623 VSS.n1622 0.00957737
R23371 VSS.n542 VSS.n541 0.00957737
R23372 VSS.n1210 VSS.n1116 0.00957737
R23373 VSS.n1622 VSS.n1621 0.00957737
R23374 VSS.n1116 VSS.n1115 0.00957737
R23375 VSS.n541 VSS.n540 0.00957737
R23376 VSS.n221 VSS.n220 0.00957737
R23377 VSS.n349 VSS.n348 0.00957737
R23378 VSS.n383 VSS.n382 0.00957737
R23379 VSS.n1723 VSS.n1722 0.00957737
R23380 VSS.n2183 VSS.n2182 0.00957737
R23381 VSS.n2213 VSS.n2212 0.00957737
R23382 VSS.n2242 VSS.n2241 0.00957737
R23383 VSS.n2275 VSS.n2274 0.00957737
R23384 VSS.n2403 VSS.n2402 0.00957737
R23385 VSS.n2483 VSS.n2482 0.00957737
R23386 VSS.n2504 VSS.n2503 0.00957737
R23387 VSS.n382 VSS.n381 0.00957737
R23388 VSS.n350 VSS.n349 0.00957737
R23389 VSS.n220 VSS.n219 0.00957737
R23390 VSS.n2482 VSS.n2481 0.00957737
R23391 VSS.n2404 VSS.n2403 0.00957737
R23392 VSS.n2274 VSS.n2273 0.00957737
R23393 VSS.n2212 VSS.n2211 0.00957737
R23394 VSS.n2243 VSS.n2242 0.00957737
R23395 VSS.n2182 VSS.n2181 0.00957737
R23396 VSS.n1724 VSS.n1723 0.00957737
R23397 VSS.n2505 VSS.n2504 0.00957737
R23398 VSS.n1900 VSS.n1890 0.00952778
R23399 VSS.n2094 VSS.n2084 0.00952778
R23400 VSS.n1387 VSS.n1386 0.00952566
R23401 VSS.n1618 VSS.n1617 0.00952566
R23402 VSS.n2506 VSS.n2505 0.00923422
R23403 VSS.n1585 VSS.n1584 0.0091882
R23404 VSS.n1588 VSS.n1587 0.0091882
R23405 VSS.n1594 VSS.n1593 0.0091882
R23406 VSS.n1593 VSS.n1592 0.0091882
R23407 VSS.n1589 VSS.n1588 0.0091882
R23408 VSS.n1584 VSS.n1583 0.0091882
R23409 VSS.n1027 VSS.n1026 0.0091882
R23410 VSS.n1026 VSS.n1025 0.0091882
R23411 VSS.n1621 VSS.n1620 0.0091882
R23412 VSS.n1292 VSS.n1291 0.0091882
R23413 VSS.n1620 VSS.n1619 0.0091882
R23414 VSS.n1293 VSS.n1292 0.0091882
R23415 VSS.n219 VSS.n145 0.0091882
R23416 VSS.n348 VSS.n223 0.0091882
R23417 VSS.n352 VSS.n351 0.0091882
R23418 VSS.n426 VSS.n399 0.0091882
R23419 VSS.n1722 VSS.n1696 0.0091882
R23420 VSS.n2181 VSS.n2155 0.0091882
R23421 VSS.n2185 VSS.n2184 0.0091882
R23422 VSS.n2241 VSS.n2215 0.0091882
R23423 VSS.n2273 VSS.n2245 0.0091882
R23424 VSS.n2402 VSS.n2277 0.0091882
R23425 VSS.n2406 VSS.n2405 0.0091882
R23426 VSS.n223 VSS.n222 0.0091882
R23427 VSS.n145 VSS.n144 0.0091882
R23428 VSS.n2277 VSS.n2276 0.0091882
R23429 VSS.n2245 VSS.n2244 0.0091882
R23430 VSS.n2215 VSS.n2214 0.0091882
R23431 VSS.n2481 VSS.n2406 0.0091882
R23432 VSS.n2211 VSS.n2185 0.0091882
R23433 VSS.n2155 VSS.n2154 0.0091882
R23434 VSS.n381 VSS.n352 0.0091882
R23435 VSS.n399 VSS.n398 0.0091882
R23436 VSS.n1696 VSS.n1695 0.0091882
R23437 VSS.n2507 VSS.n2506 0.00914234
R23438 VSS.n1809 VSS.n1808 0.00883333
R23439 VSS.n1888 VSS.n1879 0.00883333
R23440 VSS.n2082 VSS.n2073 0.00883333
R23441 VSS.n2003 VSS.n2002 0.00883333
R23442 VSS.n880 VSS.n879 0.00879896
R23443 VSS.n610 VSS.n609 0.00879896
R23444 VSS.n719 VSS.n718 0.00879896
R23445 VSS.n2364 VSS.n2361 0.00865217
R23446 VSS.n2381 VSS.n2379 0.00865217
R23447 VSS.n2454 VSS.n2452 0.00865217
R23448 VSS.n192 VSS.n190 0.00865217
R23449 VSS.n310 VSS.n307 0.00865217
R23450 VSS.n327 VSS.n325 0.00865217
R23451 VSS.n967 VSS.n960 0.00865217
R23452 VSS.n998 VSS.n996 0.00865217
R23453 VSS.n673 VSS.n670 0.00865217
R23454 VSS.n690 VSS.n688 0.00865217
R23455 VSS.n806 VSS.n799 0.00865217
R23456 VSS.n837 VSS.n835 0.00865217
R23457 VSS.n1983 VSS.n1981 0.00865217
R23458 VSS.n1783 VSS.n1781 0.00865217
R23459 VSS.n1630 VSS.n1627 0.0083125
R23460 VSS.n439 VSS.n437 0.0083125
R23461 VSS.n20 VSS.n19 0.0083125
R23462 VSS.n32 VSS.n31 0.0083125
R23463 VSS.n1820 VSS.n1819 0.00813889
R23464 VSS.n1877 VSS.n1867 0.00813889
R23465 VSS.n2071 VSS.n2061 0.00813889
R23466 VSS.n2014 VSS.n2013 0.00813889
R23467 VSS.n416 VSS.n415 0.00765694
R23468 VSS.n1832 VSS.n1831 0.00744444
R23469 VSS.n1865 VSS.n1856 0.00744444
R23470 VSS.n2059 VSS.n2050 0.00744444
R23471 VSS.n2026 VSS.n2025 0.00744444
R23472 VSS.n2432 VSS.n2431 0.00685176
R23473 VSS.n2263 VSS.n2262 0.00685176
R23474 VSS.n171 VSS.n170 0.00685176
R23475 VSS.n2173 VSS.n2172 0.00685176
R23476 VSS.n1662 VSS.n1661 0.0068172
R23477 VSS.n1074 VSS.n1073 0.00675
R23478 VSS.n1070 VSS.n1069 0.00675
R23479 VSS.n1843 VSS.n1842 0.00675
R23480 VSS.n1854 VSS.n1844 0.00675
R23481 VSS.n2048 VSS.n2038 0.00675
R23482 VSS.n2037 VSS.n2036 0.00675
R23483 VSS.n428 VSS.n427 0.00675
R23484 VSS.n1065 VSS.n1064 0.00671462
R23485 VSS.n1061 VSS.n1060 0.00671462
R23486 VSS.n1598 VSS.n1597 0.00647588
R23487 VSS.n1616 VSS.n1348 0.00647588
R23488 VSS.n28 VSS.n27 0.00635938
R23489 VSS.n1790 VSS.n1789 0.00620828
R23490 VSS.n1842 VSS.n1833 0.00605556
R23491 VSS.n1855 VSS.n1854 0.00605556
R23492 VSS.n2049 VSS.n2048 0.00605556
R23493 VSS.n2036 VSS.n2027 0.00605556
R23494 VSS.n2307 VSS.n2305 0.00593478
R23495 VSS.n2323 VSS.n2321 0.00593478
R23496 VSS.n253 VSS.n251 0.00593478
R23497 VSS.n269 VSS.n267 0.00593478
R23498 VSS.n1552 VSS.n1550 0.00593478
R23499 VSS.n1443 VSS.n1441 0.00593478
R23500 VSS.n459 VSS.n457 0.00593478
R23501 VSS.n476 VSS.n474 0.00593478
R23502 VSS.n1126 VSS.n1124 0.00593478
R23503 VSS.n1151 VSS.n1149 0.00593478
R23504 VSS.n1139 VSS.n1132 0.00593478
R23505 VSS.n1231 VSS.n1229 0.00593478
R23506 VSS.n907 VSS.n905 0.00593478
R23507 VSS.n632 VSS.n630 0.00593478
R23508 VSS.n745 VSS.n743 0.00593478
R23509 VSS.n1075 VSS.n1074 0.00592961
R23510 VSS.n1103 VSS.n1101 0.00580645
R23511 VSS.n1 VSS.n0 0.0055
R23512 VSS.n1831 VSS.n1821 0.00536111
R23513 VSS.n1866 VSS.n1865 0.00536111
R23514 VSS.n2060 VSS.n2059 0.00536111
R23515 VSS.n2025 VSS.n2015 0.00536111
R23516 VSS.n1211 VSS.n1110 0.00530108
R23517 VSS.n1385 VSS.n1384 0.00507113
R23518 VSS.n1384 VSS.n1383 0.00507113
R23519 VSS.n1610 VSS.n1609 0.00507113
R23520 VSS.n1609 VSS.n1608 0.00507113
R23521 VSS.n2486 VSS.n2485 0.00507113
R23522 VSS.n2485 VSS.n2484 0.00507113
R23523 VSS.n2498 VSS.n2497 0.00507113
R23524 VSS.n2497 VSS.n2496 0.00507113
R23525 VSS.n1607 VSS.n1606 0.00507113
R23526 VSS.n1608 VSS.n1607 0.00507113
R23527 VSS.n1382 VSS.n1381 0.00507113
R23528 VSS.n1383 VSS.n1382 0.00507113
R23529 VSS.n1789 VSS.n1788 0.00500684
R23530 VSS.n597 VSS.n596 0.00492302
R23531 VSS.n700 VSS.n699 0.00492108
R23532 VSS.n851 VSS.n850 0.00492108
R23533 VSS.n1012 VSS.n1011 0.00492021
R23534 VSS.n423 VSS.n420 0.00490286
R23535 VSS.n554 VSS.n552 0.0047957
R23536 VSS.n1094 VSS.n1093 0.0047957
R23537 VSS.n1819 VSS.n1810 0.00466667
R23538 VSS.n1878 VSS.n1877 0.00466667
R23539 VSS.n2072 VSS.n2071 0.00466667
R23540 VSS.n2013 VSS.n2004 0.00466667
R23541 VSS.n1991 VSS.n1990 0.00466667
R23542 VSS.n559 VSS.n558 0.00454301
R23543 VSS.n1713 VSS.n1712 0.00440625
R23544 VSS.n2168 VSS.n2167 0.00440625
R23545 VSS.n2202 VSS.n2201 0.00440625
R23546 VSS.n2232 VSS.n2231 0.00440625
R23547 VSS.n2258 VSS.n2257 0.00440625
R23548 VSS.n2290 VSS.n2289 0.00440625
R23549 VSS.n2427 VSS.n2426 0.00440625
R23550 VSS.n166 VSS.n165 0.00440625
R23551 VSS.n236 VSS.n235 0.00440625
R23552 VSS.n369 VSS.n368 0.00440625
R23553 VSS.n18 VSS.n17 0.00440625
R23554 VSS.n552 VSS.n551 0.00429032
R23555 VSS.n1093 VSS.n1092 0.00429032
R23556 VSS.n1989 VSS.n1988 0.00428997
R23557 VSS.n1660 VSS.n1659 0.00403763
R23558 VSS.n1808 VSS.n1791 0.00397222
R23559 VSS.n1889 VSS.n1888 0.00397222
R23560 VSS.n2083 VSS.n2082 0.00397222
R23561 VSS.n2002 VSS.n1992 0.00397222
R23562 VSS.n1671 VSS.n1670 0.00353226
R23563 VSS.n1103 VSS.n1102 0.00327957
R23564 VSS.n1901 VSS.n1900 0.00327778
R23565 VSS.n2095 VSS.n2094 0.00327778
R23566 VSS.n2370 VSS.n2368 0.00321739
R23567 VSS.n2374 VSS.n2372 0.00321739
R23568 VSS.n2443 VSS.n2441 0.00321739
R23569 VSS.n181 VSS.n179 0.00321739
R23570 VSS.n316 VSS.n314 0.00321739
R23571 VSS.n320 VSS.n318 0.00321739
R23572 VSS.n1403 VSS.n1401 0.00321739
R23573 VSS.n978 VSS.n971 0.00321739
R23574 VSS.n987 VSS.n985 0.00321739
R23575 VSS.n679 VSS.n677 0.00321739
R23576 VSS.n683 VSS.n681 0.00321739
R23577 VSS.n817 VSS.n810 0.00321739
R23578 VSS.n826 VSS.n824 0.00321739
R23579 VSS.n1320 VSS.n1318 0.00321739
R23580 VSS.n1971 VSS.n1969 0.00321739
R23581 VSS.n1771 VSS.n1769 0.00321739
R23582 VSS.n1632 VSS.n1631 0.00302688
R23583 VSS.n441 VSS.n440 0.00302688
R23584 VSS.n1709 VSS.n1708 0.00295228
R23585 VSS.n2198 VSS.n2197 0.00295228
R23586 VSS.n2228 VSS.n2227 0.00295228
R23587 VSS.n2286 VSS.n2285 0.00295228
R23588 VSS.n232 VSS.n231 0.00295228
R23589 VSS.n365 VSS.n364 0.00295228
R23590 VSS.n445 VSS.n443 0.00284375
R23591 VSS.n1295 VSS.n1215 0.00284375
R23592 VSS.n556 VSS.n555 0.00278115
R23593 VSS.n555 VSS.n550 0.00278115
R23594 VSS.n1058 VSS.n1057 0.00269167
R23595 VSS.n1912 VSS.n1911 0.00258333
R23596 VSS.n2106 VSS.n2105 0.00258333
R23597 VSS.n1090 VSS.n1089 0.00252151
R23598 VSS.n1097 VSS.n1096 0.00252151
R23599 VSS.n1298 VSS.n1297 0.00252151
R23600 VSS.n1540 VSS.n1539 0.00245312
R23601 VSS.n1530 VSS.n1529 0.00245312
R23602 VSS.n1512 VSS.n1511 0.00245312
R23603 VSS.n1499 VSS.n1498 0.00245312
R23604 VSS.n1431 VSS.n1430 0.00245312
R23605 VSS.n1418 VSS.n1417 0.00245312
R23606 VSS.n1288 VSS.n1287 0.00245312
R23607 VSS.n1278 VSS.n1277 0.00245312
R23608 VSS.n1208 VSS.n1207 0.00245312
R23609 VSS.n1198 VSS.n1197 0.00245312
R23610 VSS.n534 VSS.n533 0.00245312
R23611 VSS.n524 VSS.n523 0.00245312
R23612 VSS.n1344 VSS.n1343 0.00245312
R23613 VSS.n1328 VSS.n1327 0.00245312
R23614 VSS.n430 VSS.n429 0.00226882
R23615 VSS.n1663 VSS.n1662 0.00226882
R23616 VSS.n1114 VSS.n1113 0.0020625
R23617 VSS.n2137 VSS.n2136 0.00204321
R23618 VSS.n1925 VSS.n1924 0.00188889
R23619 VSS.n2135 VSS.n2134 0.00188889
R23620 VSS.n2119 VSS.n2118 0.00188889
R23621 VSS.n94 VSS.n91 0.00175105
R23622 VSS.n1299 VSS.n1107 0.00166815
R23623 VSS.n433 VSS.n432 0.00166815
R23624 VSS.n1300 VSS.n1299 0.00166815
R23625 VSS.n860 VSS.n859 0.00149427
R23626 VSS.n1099 VSS.n1098 0.00145036
R23627 VSS.n1098 VSS.n567 0.00145036
R23628 VSS.n548 VSS.n547 0.00143078
R23629 VSS.n547 VSS.n546 0.00143078
R23630 VSS.n1057 VSS.n1056 0.00130794
R23631 VSS.n542 VSS.n538 0.00128125
R23632 VSS.n391 VSS.n390 0.00128125
R23633 VSS.n2151 VSS.n2150 0.00127161
R23634 VSS.n447 VSS.n446 0.00125806
R23635 VSS.n1296 VSS.n1213 0.00125806
R23636 VSS.n550 VSS.n549 0.00119582
R23637 VSS.n549 VSS.n548 0.00119582
R23638 VSS.n1936 VSS.n1935 0.00119444
R23639 VSS.n2130 VSS.n2129 0.00119444
R23640 VSS.n1990 VSS.n1989 0.00119444
R23641 VSS.n566 VSS.n556 0.00117624
R23642 VSS.n567 VSS.n566 0.00117624
R23643 VSS.n1637 VSS.n1636 0.0011689
R23644 VSS.n1644 VSS.n1643 0.0011689
R23645 VSS.n1645 VSS.n1644 0.0011689
R23646 VSS.n1636 VSS.n1635 0.0011689
R23647 VSS.n1105 VSS.n1104 0.00116156
R23648 VSS.n1639 VSS.n1638 0.00116156
R23649 VSS.n1640 VSS.n1639 0.00116156
R23650 VSS.n1104 VSS.n1100 0.00116156
R23651 VSS.n1365 VSS.n1364 0.00113518
R23652 VSS.n94 VSS.n93 0.00113518
R23653 VSS.n1355 VSS.n1354 0.00113518
R23654 VSS.n1360 VSS.n1359 0.00113518
R23655 VSS.n130 VSS.n94 0.00108774
R23656 VSS.n1107 VSS.n1106 0.00107344
R23657 VSS.n1641 VSS.n433 0.00107344
R23658 VSS.n1641 VSS.n1640 0.00107344
R23659 VSS.n1106 VSS.n1105 0.00107344
R23660 VSS.n1635 VSS.n1634 0.00106609
R23661 VSS.n1646 VSS.n1645 0.00106609
R23662 VSS.n1634 VSS.n1300 0.00106609
R23663 VSS.n1646 VSS.n1642 0.00106609
R23664 VSS.n1357 VSS.n1355 0.00101803
R23665 VSS.n1359 VSS.n1357 0.00101803
R23666 VSS.n83 VSS.n80 0.0010087
R23667 VSS.n1051 VSS.n1050 0.00100166
R23668 VSS.n1038 VSS.n1037 0.00100166
R23669 VSS.n1364 VSS.n1363 0.00100123
R23670 VSS.n1051 VSS.n1048 0.00100102
R23671 VSS.n1038 VSS.n1035 0.00100102
R23672 VSS.n137 VSS.n136 0.00100038
R23673 VSS.n1039 VSS.n1033 0.00100018
R23674 VSS.n136 VSS.n135 0.0010001
R23675 VSS.n139 VSS.n138 0.00100007
R23676 VSS.n1029 VSS.n1028 0.00100006
R23677 VSS.n142 VSS.n141 0.00100002
R23678 VSS.n1031 VSS.n1029 0.00100001
R23679 VSS.n1052 VSS.n1051 0.001
R23680 VSS.n1033 VSS.n1032 0.001
R23681 VSS.n1039 VSS.n1038 0.001
R23682 VSS.n1359 VSS.n1358 0.001
R23683 VSS.n1652 VSS.n1651 0.000752688
R23684 VSS.n544 VSS.n543 0.000752688
R23685 VSS.n79 VSS.n78 0.000670243
R23686 VSS.n85 VSS.n79 0.000670243
R23687 VSS.n86 VSS.n85 0.000670243
R23688 VSS.n1354 VSS.n1353 0.000635176
R23689 VSS.n1361 VSS.n1360 0.000635176
R23690 VSS.n1366 VSS.n1365 0.000635176
R23691 VSS.n93 VSS.n92 0.000635176
R23692 VSS.n132 VSS.n131 0.000635176
R23693 VSS.n131 VSS.n130 0.000635176
R23694 VSS.n89 VSS.n88 0.000631513
R23695 VSS.n135 VSS.n89 0.000631513
R23696 VSS.n1371 VSS.n1370 0.000552238
R23697 VSS.n1370 VSS.n1369 0.000552238
R23698 VSS.n1368 VSS.n1367 0.000552238
R23699 VSS.n1369 VSS.n1368 0.000552238
R23700 VSS.n76 VSS.n75 0.000512877
R23701 VSS.n77 VSS.n76 0.000512877
R23702 VSS.n86 VSS.n77 0.000512877
R23703 VSS.n134 VSS.n133 0.00051244
R23704 VSS.n135 VSS.n134 0.00051244
R23705 VSS.n87 VSS.n86 0.000511972
R23706 VSS.n84 VSS.n83 0.000510754
R23707 VSS.n1357 VSS.n1356 0.000509014
R23708 VSS.n74 VSS.n73 0.000507954
R23709 VSS.n73 VSS.n72 0.000507954
R23710 VSS.n69 VSS.n68 0.000507954
R23711 VSS.n72 VSS.n69 0.000507954
R23712 VSS.n1054 VSS.n1053 0.000505303
R23713 VSS.n1053 VSS.n1052 0.000505303
R23714 VSS.n1041 VSS.n1040 0.000505303
R23715 VSS.n1040 VSS.n1039 0.000505303
R23716 VSS.n71 VSS.n70 0.000503977
R23717 VSS.n72 VSS.n71 0.000503977
R23718 VSS.n1046 VSS.n1045 0.000503145
R23719 VSS.n1045 VSS.n1044 0.000503145
R23720 VSS.n1044 VSS.n1043 0.000503145
R23721 VSS.n1043 VSS.n1042 0.000503145
R23722 VSS.n1050 VSS.n1049 0.000501661
R23723 VSS.n1037 VSS.n1036 0.000501661
R23724 VSS.n83 VSS.n82 0.000501387
R23725 VSS.n1363 VSS.n1362 0.000501229
R23726 VSS.n91 VSS.n90 0.000501048
R23727 VSS.n1048 VSS.n1047 0.000501025
R23728 VSS.n1035 VSS.n1034 0.000501025
R23729 VSS.n83 VSS.n81 0.000500725
R23730 VSS.n138 VSS.n137 0.000500479
R23731 VSS.n1056 VSS.n860 0.000500181
R23732 VSS.n1032 VSS.n1031 0.000500181
R23733 VSS.n143 VSS.n142 0.000500106
R23734 VSS.n2136 VSS.n2135 0.000500075
R23735 a_1355_1794.n10 a_1355_1794.t4 60.2505
R23736 a_1355_1794.n70 a_1355_1794.t6 60.2505
R23737 a_1355_1794.n25 a_1355_1794.t9 60.2505
R23738 a_1355_1794.n47 a_1355_1794.t8 60.2505
R23739 a_1355_1794.n2 a_1355_1794.n79 9.3005
R23740 a_1355_1794.n4 a_1355_1794.n63 9.3005
R23741 a_1355_1794.n5 a_1355_1794.n56 9.3005
R23742 a_1355_1794.n7 a_1355_1794.n40 9.3005
R23743 a_1355_1794.n6 a_1355_1794.n39 9.3005
R23744 a_1355_1794.n58 a_1355_1794.n57 9.3005
R23745 a_1355_1794.n5 a_1355_1794.n55 9.3005
R23746 a_1355_1794.n55 a_1355_1794.n54 9.3005
R23747 a_1355_1794.n7 a_1355_1794.n46 9.3005
R23748 a_1355_1794.n46 a_1355_1794.n45 9.3005
R23749 a_1355_1794.n8 a_1355_1794.n33 9.3005
R23750 a_1355_1794.n35 a_1355_1794.n34 9.3005
R23751 a_1355_1794.n8 a_1355_1794.n32 9.3005
R23752 a_1355_1794.n32 a_1355_1794.n31 9.3005
R23753 a_1355_1794.n81 a_1355_1794.n80 9.3005
R23754 a_1355_1794.n2 a_1355_1794.n78 9.3005
R23755 a_1355_1794.n78 a_1355_1794.n77 9.3005
R23756 a_1355_1794.n4 a_1355_1794.n69 9.3005
R23757 a_1355_1794.n69 a_1355_1794.n68 9.3005
R23758 a_1355_1794.n3 a_1355_1794.n62 9.3005
R23759 a_1355_1794.n1 a_1355_1794.n17 9.3005
R23760 a_1355_1794.n17 a_1355_1794.n16 9.3005
R23761 a_1355_1794.n20 a_1355_1794.n19 9.3005
R23762 a_1355_1794.n1 a_1355_1794.n18 9.3005
R23763 a_1355_1794.n48 a_1355_1794.n47 8.76429
R23764 a_1355_1794.n71 a_1355_1794.n70 8.76429
R23765 a_1355_1794.n30 a_1355_1794.n29 8.21641
R23766 a_1355_1794.n53 a_1355_1794.n52 8.21641
R23767 a_1355_1794.n44 a_1355_1794.n43 8.21641
R23768 a_1355_1794.n76 a_1355_1794.n75 8.21641
R23769 a_1355_1794.n67 a_1355_1794.n66 8.21641
R23770 a_1355_1794.n15 a_1355_1794.n14 8.21641
R23771 a_1355_1794.n26 a_1355_1794.n25 6.92011
R23772 a_1355_1794.n11 a_1355_1794.n10 6.92007
R23773 a_1355_1794.n28 a_1355_1794.n27 5.64756
R23774 a_1355_1794.n51 a_1355_1794.n50 5.64756
R23775 a_1355_1794.n42 a_1355_1794.n41 5.64756
R23776 a_1355_1794.n74 a_1355_1794.n73 5.64756
R23777 a_1355_1794.n65 a_1355_1794.n64 5.64756
R23778 a_1355_1794.n13 a_1355_1794.n12 5.64756
R23779 a_1355_1794.n103 a_1355_1794.t1 5.5395
R23780 a_1355_1794.n103 a_1355_1794.t2 5.5395
R23781 a_1355_1794.t3 a_1355_1794.n129 5.5395
R23782 a_1355_1794.n129 a_1355_1794.t0 5.5395
R23783 a_1355_1794.n85 a_1355_1794.n84 5.27461
R23784 a_1355_1794.n36 a_1355_1794.n24 4.76425
R23785 a_1355_1794.n59 a_1355_1794.n23 4.76425
R23786 a_1355_1794.n38 a_1355_1794.n37 4.76425
R23787 a_1355_1794.n82 a_1355_1794.n22 4.76425
R23788 a_1355_1794.n61 a_1355_1794.n60 4.76425
R23789 a_1355_1794.n21 a_1355_1794.n9 4.76425
R23790 a_1355_1794.n49 a_1355_1794.n48 4.6505
R23791 a_1355_1794.n72 a_1355_1794.n71 4.6505
R23792 a_1355_1794.n116 a_1355_1794.n115 4.51815
R23793 a_1355_1794.n119 a_1355_1794.n118 4.51815
R23794 a_1355_1794.n86 a_1355_1794.n97 6.0005
R23795 a_1355_1794.n87 a_1355_1794.n89 4.5005
R23796 a_1355_1794.n109 a_1355_1794.n113 4.5005
R23797 a_1355_1794.n105 a_1355_1794.n108 4.5005
R23798 a_1355_1794.n98 a_1355_1794.n126 4.5005
R23799 a_1355_1794.n99 a_1355_1794.n123 4.5005
R23800 a_1355_1794.n113 a_1355_1794.n110 4.14168
R23801 a_1355_1794.n123 a_1355_1794.n120 4.14168
R23802 a_1355_1794.n1 a_1355_1794.n11 3.47842
R23803 a_1355_1794.n8 a_1355_1794.n26 3.47753
R23804 a_1355_1794.n97 a_1355_1794.n96 3.38238
R23805 a_1355_1794.n101 a_1355_1794.t5 3.3065
R23806 a_1355_1794.n101 a_1355_1794.t7 3.3065
R23807 a_1355_1794.n91 a_1355_1794.n101 3.21134
R23808 a_1355_1794.n114 a_1355_1794.n116 3.03311
R23809 a_1355_1794.n100 a_1355_1794.n119 3.03311
R23810 a_1355_1794.n129 a_1355_1794.n128 2.85325
R23811 a_1355_1794.n0 a_1355_1794.n91 2.51547
R23812 a_1355_1794.n107 a_1355_1794.n106 2.25932
R23813 a_1355_1794.n125 a_1355_1794.n124 2.25932
R23814 a_1355_1794.n113 a_1355_1794.n111 2.22452
R23815 a_1355_1794.n123 a_1355_1794.n121 2.22452
R23816 a_1355_1794.n97 a_1355_1794.n95 1.88285
R23817 a_1355_1794.n100 a_1355_1794.n0 1.68211
R23818 a_1355_1794.n104 a_1355_1794.n103 1.64453
R23819 a_1355_1794.n129 a_1355_1794.n127 1.64451
R23820 a_1355_1794.n90 a_1355_1794.n93 6.0005
R23821 a_1355_1794.n93 a_1355_1794.n92 1.12991
R23822 a_1355_1794.n31 a_1355_1794.n30 1.09595
R23823 a_1355_1794.n54 a_1355_1794.n53 1.09595
R23824 a_1355_1794.n45 a_1355_1794.n44 1.09595
R23825 a_1355_1794.n77 a_1355_1794.n76 1.09595
R23826 a_1355_1794.n68 a_1355_1794.n67 1.09595
R23827 a_1355_1794.n16 a_1355_1794.n15 1.09595
R23828 a_1355_1794.n32 a_1355_1794.n28 0.753441
R23829 a_1355_1794.n55 a_1355_1794.n51 0.753441
R23830 a_1355_1794.n46 a_1355_1794.n42 0.753441
R23831 a_1355_1794.n78 a_1355_1794.n74 0.753441
R23832 a_1355_1794.n69 a_1355_1794.n65 0.753441
R23833 a_1355_1794.n17 a_1355_1794.n13 0.753441
R23834 a_1355_1794.n95 a_1355_1794.n94 0.753441
R23835 a_1355_1794.n108 a_1355_1794.n107 0.753441
R23836 a_1355_1794.n126 a_1355_1794.n125 0.753441
R23837 a_1355_1794.n117 a_1355_1794.n102 0.571668
R23838 a_1355_1794.n61 a_1355_1794.n59 0.458354
R23839 a_1355_1794.n38 a_1355_1794.n36 0.458354
R23840 a_1355_1794.n89 a_1355_1794.n88 0.376971
R23841 a_1355_1794.n83 a_1355_1794.n21 0.229427
R23842 a_1355_1794.n83 a_1355_1794.n82 0.229427
R23843 a_1355_1794.n85 a_1355_1794.n83 0.191391
R23844 a_1355_1794.n2 a_1355_1794.n72 0.190717
R23845 a_1355_1794.n72 a_1355_1794.n4 0.190717
R23846 a_1355_1794.n5 a_1355_1794.n49 0.190717
R23847 a_1355_1794.n49 a_1355_1794.n7 0.190717
R23848 a_1355_1794.n21 a_1355_1794.n20 0.15935
R23849 a_1355_1794.n82 a_1355_1794.n81 0.15935
R23850 a_1355_1794.n3 a_1355_1794.n61 0.15935
R23851 a_1355_1794.n59 a_1355_1794.n58 0.15935
R23852 a_1355_1794.n6 a_1355_1794.n38 0.15935
R23853 a_1355_1794.n36 a_1355_1794.n35 0.15935
R23854 a_1355_1794.n90 a_1355_1794.n91 0.0960207
R23855 a_1355_1794.n98 a_1355_1794.n99 0.0905127
R23856 a_1355_1794.n109 a_1355_1794.n105 0.0900861
R23857 a_1355_1794.n86 a_1355_1794.n90 0.0765135
R23858 a_1355_1794.n87 a_1355_1794.n85 0.125375
R23859 a_1355_1794.n117 a_1355_1794.n114 0.0620415
R23860 a_1355_1794.n105 a_1355_1794.n104 0.557653
R23861 a_1355_1794.n99 a_1355_1794.n100 0.0454219
R23862 a_1355_1794.n114 a_1355_1794.n109 0.0454219
R23863 a_1355_1794.n87 a_1355_1794.n86 1.53935
R23864 a_1355_1794.n0 a_1355_1794.n117 0.709629
R23865 a_1355_1794.n35 a_1355_1794.n8 0.0466957
R23866 a_1355_1794.n7 a_1355_1794.n6 0.0466957
R23867 a_1355_1794.n58 a_1355_1794.n5 0.0466957
R23868 a_1355_1794.n4 a_1355_1794.n3 0.0466957
R23869 a_1355_1794.n81 a_1355_1794.n2 0.0466957
R23870 a_1355_1794.n20 a_1355_1794.n1 0.0466957
R23871 a_1355_1794.n111 a_1355_1794.n112 0.0303633
R23872 a_1355_1794.n121 a_1355_1794.n122 0.0303633
R23873 a_1355_1794.n127 a_1355_1794.n98 0.557387
R23874 a_1755_1820.n32 a_1755_1820.t7 60.2505
R23875 a_1755_1820.n52 a_1755_1820.t6 60.2505
R23876 a_1755_1820.n73 a_1755_1820.t2 60.2505
R23877 a_1755_1820.n85 a_1755_1820.t0 60.2505
R23878 a_1755_1820.n2 a_1755_1820.n93 9.3005
R23879 a_1755_1820.n2 a_1755_1820.n94 9.3005
R23880 a_1755_1820.n2 a_1755_1820.n92 9.3005
R23881 a_1755_1820.n92 a_1755_1820.n91 9.3005
R23882 a_1755_1820.n3 a_1755_1820.n82 9.3005
R23883 a_1755_1820.n5 a_1755_1820.n66 9.3005
R23884 a_1755_1820.n5 a_1755_1820.n65 9.3005
R23885 a_1755_1820.n5 a_1755_1820.n72 9.3005
R23886 a_1755_1820.n72 a_1755_1820.n71 9.3005
R23887 a_1755_1820.n3 a_1755_1820.n81 9.3005
R23888 a_1755_1820.n81 a_1755_1820.n80 9.3005
R23889 a_1755_1820.n3 a_1755_1820.n83 9.3005
R23890 a_1755_1820.n6 a_1755_1820.n61 9.3005
R23891 a_1755_1820.n8 a_1755_1820.n45 9.3005
R23892 a_1755_1820.n8 a_1755_1820.n44 9.3005
R23893 a_1755_1820.n8 a_1755_1820.n51 9.3005
R23894 a_1755_1820.n51 a_1755_1820.n50 9.3005
R23895 a_1755_1820.n6 a_1755_1820.n60 9.3005
R23896 a_1755_1820.n60 a_1755_1820.n59 9.3005
R23897 a_1755_1820.n6 a_1755_1820.n62 9.3005
R23898 a_1755_1820.n9 a_1755_1820.n40 9.3005
R23899 a_1755_1820.n9 a_1755_1820.n39 9.3005
R23900 a_1755_1820.n39 a_1755_1820.n38 9.3005
R23901 a_1755_1820.n9 a_1755_1820.n41 9.3005
R23902 a_1755_1820.n11 a_1755_1820.n100 9.3005
R23903 a_1755_1820.n11 a_1755_1820.n99 9.3005
R23904 a_1755_1820.n28 a_1755_1820.n101 9.3005
R23905 a_1755_1820.n27 a_1755_1820.n102 9.3005
R23906 a_1755_1820.n26 a_1755_1820.n103 9.3005
R23907 a_1755_1820.n0 a_1755_1820.n104 9.3005
R23908 a_1755_1820.n124 a_1755_1820.n111 9.909
R23909 a_1755_1820.n124 a_1755_1820.n112 11.0386
R23910 a_1755_1820.n124 a_1755_1820.n123 8.89115
R23911 a_1755_1820.n124 a_1755_1820.n120 8.88036
R23912 a_1755_1820.n124 a_1755_1820.n117 8.86963
R23913 a_1755_1820.n124 a_1755_1820.n113 8.85895
R23914 a_1755_1820.n74 a_1755_1820.n73 8.76429
R23915 a_1755_1820.n53 a_1755_1820.n52 8.76429
R23916 a_1755_1820.n37 a_1755_1820.n36 7.45411
R23917 a_1755_1820.n49 a_1755_1820.n48 7.45411
R23918 a_1755_1820.n58 a_1755_1820.n57 7.45411
R23919 a_1755_1820.n70 a_1755_1820.n69 7.45411
R23920 a_1755_1820.n79 a_1755_1820.n78 7.45411
R23921 a_1755_1820.n90 a_1755_1820.n89 7.45411
R23922 a_1755_1820.n22 a_1755_1820.n21 7.45281
R23923 a_1755_1820.n33 a_1755_1820.n32 6.80105
R23924 a_1755_1820.n86 a_1755_1820.n85 6.80105
R23925 a_1755_1820.n0 a_1755_1820.n13 6.29716
R23926 a_1755_1820.n35 a_1755_1820.n34 5.64756
R23927 a_1755_1820.n47 a_1755_1820.n46 5.64756
R23928 a_1755_1820.n56 a_1755_1820.n55 5.64756
R23929 a_1755_1820.n68 a_1755_1820.n67 5.64756
R23930 a_1755_1820.n77 a_1755_1820.n76 5.64756
R23931 a_1755_1820.n88 a_1755_1820.n87 5.64756
R23932 a_1755_1820.t3 a_1755_1820.n124 5.5395
R23933 a_1755_1820.n124 a_1755_1820.t1 5.5395
R23934 a_1755_1820.n10 a_1755_1820.n98 4.95534
R23935 a_1755_1820.n42 a_1755_1820.n31 4.73575
R23936 a_1755_1820.n7 a_1755_1820.n43 4.73575
R23937 a_1755_1820.n63 a_1755_1820.n30 4.73575
R23938 a_1755_1820.n4 a_1755_1820.n64 4.73575
R23939 a_1755_1820.n84 a_1755_1820.n29 4.73575
R23940 a_1755_1820.n96 a_1755_1820.n95 4.73575
R23941 a_1755_1820.n75 a_1755_1820.n74 4.6505
R23942 a_1755_1820.n54 a_1755_1820.n53 4.6505
R23943 a_1755_1820.n1 a_1755_1820.n23 4.5005
R23944 a_1755_1820.n1 a_1755_1820.n22 4.5005
R23945 a_1755_1820.n1 a_1755_1820.n107 4.5005
R23946 a_1755_1820.n0 a_1755_1820.n25 4.5005
R23947 a_1755_1820.n1 a_1755_1820.n109 4.5005
R23948 a_1755_1820.n9 a_1755_1820.n33 3.42768
R23949 a_1755_1820.n2 a_1755_1820.n86 3.42768
R23950 a_1755_1820.n109 a_1755_1820.n108 3.38874
R23951 a_1755_1820.n116 a_1755_1820.n115 3.38874
R23952 a_1755_1820.n19 a_1755_1820.n18 3.38238
R23953 a_1755_1820.n105 a_1755_1820.t5 3.3065
R23954 a_1755_1820.n105 a_1755_1820.t4 3.3065
R23955 a_1755_1820.n13 a_1755_1820.n105 3.21133
R23956 a_1755_1820.n22 a_1755_1820.n20 2.63579
R23957 a_1755_1820.n119 a_1755_1820.n118 2.63579
R23958 a_1755_1820.n19 a_1755_1820.n17 1.88285
R23959 a_1755_1820.n25 a_1755_1820.n24 1.88285
R23960 a_1755_1820.n122 a_1755_1820.n121 1.88285
R23961 a_1755_1820.n124 a_1755_1820.n110 1.67004
R23962 a_1755_1820.n107 a_1755_1820.n106 1.50638
R23963 a_1755_1820.n12 a_1755_1820.n15 6.0005
R23964 a_1755_1820.n15 a_1755_1820.n14 1.12991
R23965 a_1755_1820.n38 a_1755_1820.n37 0.994314
R23966 a_1755_1820.n50 a_1755_1820.n49 0.994314
R23967 a_1755_1820.n59 a_1755_1820.n58 0.994314
R23968 a_1755_1820.n71 a_1755_1820.n70 0.994314
R23969 a_1755_1820.n80 a_1755_1820.n79 0.994314
R23970 a_1755_1820.n91 a_1755_1820.n90 0.994314
R23971 a_1755_1820.n110 a_1755_1820.n1 0.944917
R23972 a_1755_1820.n17 a_1755_1820.n16 0.753441
R23973 a_1755_1820.n39 a_1755_1820.n35 0.753441
R23974 a_1755_1820.n51 a_1755_1820.n47 0.753441
R23975 a_1755_1820.n60 a_1755_1820.n56 0.753441
R23976 a_1755_1820.n72 a_1755_1820.n68 0.753441
R23977 a_1755_1820.n81 a_1755_1820.n77 0.753441
R23978 a_1755_1820.n92 a_1755_1820.n88 0.753441
R23979 a_1755_1820.n7 a_1755_1820.n42 0.458354
R23980 a_1755_1820.n4 a_1755_1820.n63 0.458354
R23981 a_1755_1820.n97 a_1755_1820.n84 0.229427
R23982 a_1755_1820.n97 a_1755_1820.n96 0.229427
R23983 a_1755_1820.n10 a_1755_1820.n97 0.215848
R23984 a_1755_1820.n27 a_1755_1820.n28 0.190717
R23985 a_1755_1820.n26 a_1755_1820.n27 0.190717
R23986 a_1755_1820.n0 a_1755_1820.n26 0.190717
R23987 a_1755_1820.n54 a_1755_1820.n8 0.190717
R23988 a_1755_1820.n6 a_1755_1820.n54 0.190717
R23989 a_1755_1820.n75 a_1755_1820.n5 0.190717
R23990 a_1755_1820.n3 a_1755_1820.n75 0.190717
R23991 a_1755_1820.n28 a_1755_1820.n11 0.174413
R23992 a_1755_1820.n113 a_1755_1820.n114 0.160869
R23993 a_1755_1820.n117 a_1755_1820.n116 0.14967
R23994 a_1755_1820.n120 a_1755_1820.n119 0.138414
R23995 a_1755_1820.n123 a_1755_1820.n122 0.127101
R23996 a_1755_1820.n12 a_1755_1820.n13 0.0960207
R23997 a_1755_1820.n19 a_1755_1820.n12 6.07651
R23998 a_1755_1820.n1 a_1755_1820.n0 0.343407
R23999 a_1755_1820.n42 a_1755_1820.n9 0.205546
R24000 a_1755_1820.n8 a_1755_1820.n7 0.205546
R24001 a_1755_1820.n63 a_1755_1820.n6 0.205546
R24002 a_1755_1820.n5 a_1755_1820.n4 0.205546
R24003 a_1755_1820.n84 a_1755_1820.n3 0.205546
R24004 a_1755_1820.n96 a_1755_1820.n2 0.205546
R24005 a_1755_1820.n11 a_1755_1820.n10 0.181081
R24006 DVDD.n11 DVDD.t39 591.327
R24007 DVDD.n16 DVDD.t22 591.327
R24008 DVDD.n121 DVDD.n112 321.882
R24009 DVDD.n134 DVDD.n112 321.882
R24010 DVDD.n134 DVDD.n109 321.882
R24011 DVDD.n138 DVDD.n109 321.882
R24012 DVDD.n139 DVDD.n138 321.882
R24013 DVDD.n139 DVDD.n108 321.882
R24014 DVDD.n55 DVDD.n46 321.882
R24015 DVDD.n68 DVDD.n46 321.882
R24016 DVDD.n68 DVDD.n43 321.882
R24017 DVDD.n72 DVDD.n43 321.882
R24018 DVDD.n73 DVDD.n72 321.882
R24019 DVDD.n73 DVDD.n42 321.882
R24020 DVDD.n135 DVDD.n111 175.386
R24021 DVDD.n137 DVDD.n136 175.386
R24022 DVDD.n69 DVDD.n45 175.386
R24023 DVDD.n71 DVDD.n70 175.386
R24024 DVDD.n121 DVDD.t10 171.452
R24025 DVDD.n55 DVDD.t35 171.452
R24026 DVDD.n252 DVDD.n251 161.37
R24027 DVDD.n227 DVDD.n226 161.37
R24028 DVDD.n207 DVDD.n206 161.37
R24029 DVDD.n180 DVDD.n179 161.37
R24030 DVDD.n1 DVDD.n0 161.37
R24031 DVDD.n143 DVDD.t21 160.743
R24032 DVDD.n77 DVDD.t26 160.743
R24033 DVDD.n125 DVDD.t11 159.81
R24034 DVDD.n59 DVDD.t36 159.81
R24035 DVDD.n19 DVDD.t40 148.294
R24036 DVDD.n140 DVDD.t2 144.327
R24037 DVDD.n74 DVDD.t14 144.327
R24038 DVDD.t20 DVDD.n140 140.673
R24039 DVDD.t25 DVDD.n74 140.673
R24040 DVDD.t18 DVDD.n247 129.546
R24041 DVDD.t0 DVDD.n222 129.546
R24042 DVDD.t31 DVDD.n202 129.546
R24043 DVDD.t33 DVDD.n175 129.546
R24044 DVDD.t37 DVDD.n4 129.546
R24045 DVDD.n148 DVDD.n141 124.013
R24046 DVDD.n82 DVDD.n75 124.013
R24047 DVDD.n248 DVDD.t18 100.874
R24048 DVDD.n223 DVDD.t0 100.874
R24049 DVDD.n203 DVDD.t31 100.874
R24050 DVDD.n176 DVDD.t33 100.874
R24051 DVDD.t6 DVDD.n135 96.8274
R24052 DVDD.t4 DVDD.n69 96.8274
R24053 DVDD.n249 DVDD.n247 92.5005
R24054 DVDD.n247 DVDD.n246 92.5005
R24055 DVDD.n224 DVDD.n222 92.5005
R24056 DVDD.n222 DVDD.n221 92.5005
R24057 DVDD.n204 DVDD.n202 92.5005
R24058 DVDD.n202 DVDD.n201 92.5005
R24059 DVDD.n177 DVDD.n175 92.5005
R24060 DVDD.n175 DVDD.n174 92.5005
R24061 DVDD.n5 DVDD.n2 92.5005
R24062 DVDD.n6 DVDD.n5 92.5005
R24063 DVDD.n136 DVDD.t6 78.5582
R24064 DVDD.n70 DVDD.t4 78.5582
R24065 DVDD.n5 DVDD.t37 67.8576
R24066 DVDD.n250 DVDD.n246 55.3934
R24067 DVDD.n225 DVDD.n221 55.3934
R24068 DVDD.n205 DVDD.n201 55.3934
R24069 DVDD.n178 DVDD.n174 55.3934
R24070 DVDD.n7 DVDD.n2 55.3934
R24071 DVDD.n19 DVDD.n15 52.9371
R24072 DVDD.n20 DVDD.n13 49.5938
R24073 DVDD.n17 DVDD.n16 47.5553
R24074 DVDD.n247 DVDD.t16 47.2949
R24075 DVDD.n222 DVDD.t8 47.2949
R24076 DVDD.n202 DVDD.t12 47.2949
R24077 DVDD.n175 DVDD.t29 47.2949
R24078 DVDD.n4 DVDD.t27 47.2949
R24079 DVDD.n250 DVDD.n249 46.2505
R24080 DVDD.n225 DVDD.n224 46.2505
R24081 DVDD.n205 DVDD.n204 46.2505
R24082 DVDD.n178 DVDD.n177 46.2505
R24083 DVDD.n19 DVDD.n18 46.2505
R24084 DVDD.n7 DVDD.n6 46.2505
R24085 DVDD.n141 DVDD.t20 37.8805
R24086 DVDD.n75 DVDD.t25 37.8805
R24087 DVDD.n122 DVDD.n113 36.1417
R24088 DVDD.n133 DVDD.n113 36.1417
R24089 DVDD.n133 DVDD.n115 36.1417
R24090 DVDD.n115 DVDD.n110 36.1417
R24091 DVDD.n110 DVDD.n107 36.1417
R24092 DVDD.n149 DVDD.n107 36.1417
R24093 DVDD.n149 DVDD.n148 36.1417
R24094 DVDD.n56 DVDD.n47 36.1417
R24095 DVDD.n67 DVDD.n47 36.1417
R24096 DVDD.n67 DVDD.n49 36.1417
R24097 DVDD.n49 DVDD.n44 36.1417
R24098 DVDD.n44 DVDD.n41 36.1417
R24099 DVDD.n83 DVDD.n41 36.1417
R24100 DVDD.n83 DVDD.n82 36.1417
R24101 DVDD.n15 DVDD.n14 34.4168
R24102 DVDD.n4 DVDD.n3 33.0167
R24103 DVDD.n251 DVDD.t19 32.8338
R24104 DVDD.n251 DVDD.t17 32.8338
R24105 DVDD.n226 DVDD.t1 32.8338
R24106 DVDD.n226 DVDD.t9 32.8338
R24107 DVDD.n206 DVDD.t32 32.8338
R24108 DVDD.n206 DVDD.t13 32.8338
R24109 DVDD.n179 DVDD.t34 32.8338
R24110 DVDD.n179 DVDD.t30 32.8338
R24111 DVDD.n0 DVDD.t28 32.8338
R24112 DVDD.n0 DVDD.t38 32.8338
R24113 DVDD.n12 DVDD.n11 32.0046
R24114 DVDD.n137 DVDD.t2 31.0582
R24115 DVDD.n71 DVDD.t14 31.0582
R24116 DVDD.n13 DVDD.n12 28.4938
R24117 DVDD.n248 DVDD.n246 26.4697
R24118 DVDD.n249 DVDD.n248 26.4697
R24119 DVDD.n223 DVDD.n221 26.4697
R24120 DVDD.n224 DVDD.n223 26.4697
R24121 DVDD.n203 DVDD.n201 26.4697
R24122 DVDD.n204 DVDD.n203 26.4697
R24123 DVDD.n176 DVDD.n174 26.4697
R24124 DVDD.n177 DVDD.n176 26.4697
R24125 DVDD.n6 DVDD.n3 26.4697
R24126 DVDD.n3 DVDD.n2 26.4697
R24127 DVDD.n25 DVDD.t23 22.8666
R24128 DVDD.n18 DVDD.n17 21.17
R24129 DVDD.n101 DVDD.t3 19.752
R24130 DVDD.n35 DVDD.t15 19.752
R24131 DVDD.n254 DVDD.n253 17.8772
R24132 DVDD.n229 DVDD.n228 17.8772
R24133 DVDD.n209 DVDD.n208 17.8772
R24134 DVDD.n182 DVDD.n181 17.8772
R24135 DVDD.n9 DVDD.n8 17.8772
R24136 DVDD.n253 DVDD.n252 17.4938
R24137 DVDD.n228 DVDD.n227 17.4938
R24138 DVDD.n208 DVDD.n207 17.4938
R24139 DVDD.n181 DVDD.n180 17.4938
R24140 DVDD.n8 DVDD.n1 17.4938
R24141 DVDD.n101 DVDD.t7 15.6579
R24142 DVDD.n35 DVDD.t5 15.6579
R24143 DVDD.n24 DVDD.n23 13.514
R24144 DVDD.t10 DVDD.n111 12.789
R24145 DVDD.t35 DVDD.n45 12.789
R24146 DVDD.n23 DVDD.t24 11.4335
R24147 DVDD.n125 DVDD.n124 9.30301
R24148 DVDD.n59 DVDD.n58 9.30301
R24149 DVDD.n157 DVDD.n98 9.3005
R24150 DVDD.n91 DVDD.n32 9.3005
R24151 DVDD.n26 DVDD.n25 9.3005
R24152 DVDD.n188 DVDD.n161 9.0245
R24153 DVDD.n122 DVDD.n121 8.85536
R24154 DVDD.n113 DVDD.n112 8.85536
R24155 DVDD.n112 DVDD.n111 8.85536
R24156 DVDD.n134 DVDD.n133 8.85536
R24157 DVDD.n135 DVDD.n134 8.85536
R24158 DVDD.n115 DVDD.n109 8.85536
R24159 DVDD.n136 DVDD.n109 8.85536
R24160 DVDD.n138 DVDD.n110 8.85536
R24161 DVDD.n138 DVDD.n137 8.85536
R24162 DVDD.n139 DVDD.n107 8.85536
R24163 DVDD.n140 DVDD.n139 8.85536
R24164 DVDD.n149 DVDD.n108 8.85536
R24165 DVDD.n56 DVDD.n55 8.85536
R24166 DVDD.n47 DVDD.n46 8.85536
R24167 DVDD.n46 DVDD.n45 8.85536
R24168 DVDD.n68 DVDD.n67 8.85536
R24169 DVDD.n69 DVDD.n68 8.85536
R24170 DVDD.n49 DVDD.n43 8.85536
R24171 DVDD.n70 DVDD.n43 8.85536
R24172 DVDD.n72 DVDD.n44 8.85536
R24173 DVDD.n72 DVDD.n71 8.85536
R24174 DVDD.n73 DVDD.n41 8.85536
R24175 DVDD.n74 DVDD.n73 8.85536
R24176 DVDD.n83 DVDD.n42 8.85536
R24177 DVDD.n157 DVDD.n101 7.96185
R24178 DVDD.n91 DVDD.n35 7.96185
R24179 DVDD.n269 DVDD.n268 5.88997
R24180 DVDD.n141 DVDD.n108 5.53567
R24181 DVDD.n75 DVDD.n42 5.53567
R24182 DVDD.n252 DVDD.n245 4.6505
R24183 DVDD.n227 DVDD.n220 4.6505
R24184 DVDD.n207 DVDD.n200 4.6505
R24185 DVDD.n180 DVDD.n173 4.6505
R24186 DVDD.n144 DVDD.n143 4.6505
R24187 DVDD.n157 DVDD.n156 4.6505
R24188 DVDD.n157 DVDD.n100 4.6505
R24189 DVDD.n126 DVDD.n125 4.6505
R24190 DVDD.n78 DVDD.n77 4.6505
R24191 DVDD.n91 DVDD.n90 4.6505
R24192 DVDD.n91 DVDD.n34 4.6505
R24193 DVDD.n60 DVDD.n59 4.6505
R24194 DVDD.n10 DVDD.n1 4.6505
R24195 DVDD.n158 DVDD.n157 4.65047
R24196 DVDD.n92 DVDD.n91 4.65047
R24197 DVDD.n125 DVDD.n120 4.65033
R24198 DVDD.n59 DVDD.n54 4.65033
R24199 DVDD.n236 DVDD.n235 4.5005
R24200 DVDD.n234 DVDD.n218 4.5005
R24201 DVDD.n233 DVDD.n232 4.5005
R24202 DVDD.n237 DVDD.n216 4.5005
R24203 DVDD.n196 DVDD.n191 4.5005
R24204 DVDD.n198 DVDD.n197 4.5005
R24205 DVDD.n199 DVDD.n190 4.5005
R24206 DVDD.n195 DVDD.n194 4.5005
R24207 DVDD.n169 DVDD.n164 4.5005
R24208 DVDD.n171 DVDD.n170 4.5005
R24209 DVDD.n172 DVDD.n163 4.5005
R24210 DVDD.n168 DVDD.n167 4.5005
R24211 DVDD.n119 DVDD.n118 4.5005
R24212 DVDD.n128 DVDD.n127 4.5005
R24213 DVDD.n129 DVDD.n116 4.5005
R24214 DVDD.n132 DVDD.n131 4.5005
R24215 DVDD.n130 DVDD.n117 4.5005
R24216 DVDD.n114 DVDD.n96 4.5005
R24217 DVDD.n99 DVDD.n97 4.5005
R24218 DVDD.n104 DVDD.n102 4.5005
R24219 DVDD.n155 DVDD.n154 4.5005
R24220 DVDD.n153 DVDD.n103 4.5005
R24221 DVDD.n152 DVDD.n151 4.5005
R24222 DVDD.n150 DVDD.n105 4.5005
R24223 DVDD.n145 DVDD.n142 4.5005
R24224 DVDD.n147 DVDD.n146 4.5005
R24225 DVDD.n53 DVDD.n52 4.5005
R24226 DVDD.n62 DVDD.n61 4.5005
R24227 DVDD.n63 DVDD.n50 4.5005
R24228 DVDD.n66 DVDD.n65 4.5005
R24229 DVDD.n64 DVDD.n51 4.5005
R24230 DVDD.n48 DVDD.n30 4.5005
R24231 DVDD.n33 DVDD.n31 4.5005
R24232 DVDD.n38 DVDD.n36 4.5005
R24233 DVDD.n89 DVDD.n88 4.5005
R24234 DVDD.n87 DVDD.n37 4.5005
R24235 DVDD.n86 DVDD.n85 4.5005
R24236 DVDD.n84 DVDD.n39 4.5005
R24237 DVDD.n79 DVDD.n76 4.5005
R24238 DVDD.n81 DVDD.n80 4.5005
R24239 DVDD.n253 DVDD.n250 4.32258
R24240 DVDD.n228 DVDD.n225 4.32258
R24241 DVDD.n208 DVDD.n205 4.32258
R24242 DVDD.n181 DVDD.n178 4.32258
R24243 DVDD.n8 DVDD.n7 4.32258
R24244 DVDD.n21 DVDD.n20 3.76521
R24245 DVDD.n185 DVDD.n184 3.4105
R24246 DVDD.n166 DVDD.n162 3.4105
R24247 DVDD.n212 DVDD.n211 3.4105
R24248 DVDD.n193 DVDD.n95 3.4105
R24249 DVDD.n231 DVDD.n219 3.4105
R24250 DVDD.n239 DVDD.n238 3.4105
R24251 DVDD.n257 DVDD.n256 3.4105
R24252 DVDD.n267 DVDD.n266 3.4105
R24253 DVDD.n20 DVDD.n19 3.34378
R24254 DVDD.n143 DVDD.n106 3.09909
R24255 DVDD.n77 DVDD.n40 3.09909
R24256 DVDD.n123 DVDD.n122 3.03311
R24257 DVDD.n127 DVDD.n113 3.03311
R24258 DVDD.n133 DVDD.n132 3.03311
R24259 DVDD.n115 DVDD.n114 3.03311
R24260 DVDD.n110 DVDD.n102 3.03311
R24261 DVDD.n107 DVDD.n103 3.03311
R24262 DVDD.n150 DVDD.n149 3.03311
R24263 DVDD.n148 DVDD.n147 3.03311
R24264 DVDD.n57 DVDD.n56 3.03311
R24265 DVDD.n61 DVDD.n47 3.03311
R24266 DVDD.n67 DVDD.n66 3.03311
R24267 DVDD.n49 DVDD.n48 3.03311
R24268 DVDD.n44 DVDD.n36 3.03311
R24269 DVDD.n41 DVDD.n37 3.03311
R24270 DVDD.n84 DVDD.n83 3.03311
R24271 DVDD.n82 DVDD.n81 3.03311
R24272 DVDD.n9 DVDD 2.87769
R24273 DVDD.n29 DVDD.n28 2.83325
R24274 DVDD.n22 DVDD.n21 2.82403
R24275 DVDD DVDD.n10 2.55963
R24276 DVDD.n27 DVDD.n26 2.54327
R24277 DVDD.n262 DVDD 2.45664
R24278 DVDD.n217 DVDD 2.45664
R24279 DVDD.n192 DVDD 2.45664
R24280 DVDD.n165 DVDD 2.45664
R24281 DVDD.n146 DVDD 2.28727
R24282 DVDD.n80 DVDD 2.28727
R24283 DVDD.n27 DVDD 1.8288
R24284 DVDD.n262 DVDD 1.67155
R24285 DVDD.n217 DVDD 1.67155
R24286 DVDD.n192 DVDD 1.67155
R24287 DVDD.n165 DVDD 1.67155
R24288 DVDD.n124 DVDD.n118 1.56265
R24289 DVDD.n58 DVDD.n52 1.56265
R24290 DVDD.n245 DVDD 1.53559
R24291 DVDD.n220 DVDD 1.53559
R24292 DVDD.n200 DVDD 1.53559
R24293 DVDD.n173 DVDD 1.53559
R24294 DVDD.n25 DVDD.n24 1.43457
R24295 DVDD DVDD.n214 1.0875
R24296 DVDD.n255 DVDD 0.966887
R24297 DVDD.n230 DVDD 0.966887
R24298 DVDD.n210 DVDD 0.966887
R24299 DVDD.n183 DVDD 0.966887
R24300 DVDD.n213 DVDD.n212 0.686051
R24301 DVDD.n214 DVDD.n95 0.686051
R24302 DVDD.n187 DVDD.n162 0.686005
R24303 DVDD.n268 DVDD.n267 0.686004
R24304 DVDD.n258 DVDD.n257 0.686004
R24305 DVDD.n240 DVDD.n239 0.686004
R24306 DVDD.n219 DVDD.n215 0.686004
R24307 DVDD.n186 DVDD.n185 0.686004
R24308 DVDD DVDD.n240 0.669357
R24309 DVDD.n188 DVDD.n187 0.669001
R24310 DVDD DVDD.n242 0.466583
R24311 DVDD DVDD.n189 0.454949
R24312 DVDD.n26 DVDD.n22 0.376971
R24313 DVDD.n255 DVDD.n254 0.325061
R24314 DVDD.n230 DVDD.n229 0.325061
R24315 DVDD.n210 DVDD.n209 0.325061
R24316 DVDD.n183 DVDD.n182 0.325061
R24317 DVDD.n241 DVDD.n94 0.280743
R24318 DVDD.n28 DVDD.n27 0.163151
R24319 DVDD.n254 DVDD.n245 0.158395
R24320 DVDD.n229 DVDD.n220 0.158395
R24321 DVDD.n209 DVDD.n200 0.158395
R24322 DVDD.n182 DVDD.n173 0.158395
R24323 DVDD.n10 DVDD.n9 0.158395
R24324 DVDD.n161 DVDD.n160 0.148924
R24325 DVDD.n189 DVDD.n161 0.139331
R24326 DVDD.n270 DVDD.n269 0.114172
R24327 DVDD.n266 DVDD.n262 0.0677269
R24328 DVDD.n238 DVDD.n217 0.0677269
R24329 DVDD.n193 DVDD.n192 0.0677269
R24330 DVDD.n166 DVDD.n165 0.0677269
R24331 DVDD.n256 DVDD 0.0425168
R24332 DVDD.n231 DVDD 0.0425168
R24333 DVDD.n211 DVDD 0.0425168
R24334 DVDD.n184 DVDD 0.0425168
R24335 DVDD.n242 DVDD 0.0408803
R24336 DVDD.n269 DVDD 0.0365511
R24337 DVDD.n187 DVDD.n186 0.0333089
R24338 DVDD.n240 DVDD.n215 0.0333089
R24339 DVDD.n268 DVDD.n258 0.0333089
R24340 DVDD.n214 DVDD.n213 0.0323971
R24341 DVDD DVDD.n270 0.0282727
R24342 DVDD DVDD.n255 0.0278109
R24343 DVDD DVDD.n230 0.0278109
R24344 DVDD DVDD.n210 0.0278109
R24345 DVDD DVDD.n183 0.0278109
R24346 DVDD.n29 DVDD 0.0269713
R24347 DVDD.n127 DVDD.n116 0.026141
R24348 DVDD.n132 DVDD.n116 0.026141
R24349 DVDD.n132 DVDD.n117 0.026141
R24350 DVDD.n102 DVDD.n99 0.026141
R24351 DVDD.n155 DVDD.n103 0.026141
R24352 DVDD.n151 DVDD.n103 0.026141
R24353 DVDD.n151 DVDD.n150 0.026141
R24354 DVDD.n147 DVDD.n142 0.026141
R24355 DVDD.n128 DVDD.n118 0.026141
R24356 DVDD.n129 DVDD.n128 0.026141
R24357 DVDD.n131 DVDD.n129 0.026141
R24358 DVDD.n131 DVDD.n130 0.026141
R24359 DVDD.n130 DVDD.n96 0.026141
R24360 DVDD.n104 DVDD.n97 0.026141
R24361 DVDD.n154 DVDD.n104 0.026141
R24362 DVDD.n154 DVDD.n153 0.026141
R24363 DVDD.n153 DVDD.n152 0.026141
R24364 DVDD.n152 DVDD.n105 0.026141
R24365 DVDD.n145 DVDD.n105 0.026141
R24366 DVDD.n146 DVDD.n145 0.026141
R24367 DVDD.n61 DVDD.n50 0.026141
R24368 DVDD.n66 DVDD.n50 0.026141
R24369 DVDD.n66 DVDD.n51 0.026141
R24370 DVDD.n36 DVDD.n33 0.026141
R24371 DVDD.n89 DVDD.n37 0.026141
R24372 DVDD.n85 DVDD.n37 0.026141
R24373 DVDD.n85 DVDD.n84 0.026141
R24374 DVDD.n81 DVDD.n76 0.026141
R24375 DVDD.n62 DVDD.n52 0.026141
R24376 DVDD.n63 DVDD.n62 0.026141
R24377 DVDD.n65 DVDD.n63 0.026141
R24378 DVDD.n65 DVDD.n64 0.026141
R24379 DVDD.n64 DVDD.n30 0.026141
R24380 DVDD.n38 DVDD.n31 0.026141
R24381 DVDD.n88 DVDD.n38 0.026141
R24382 DVDD.n88 DVDD.n87 0.026141
R24383 DVDD.n87 DVDD.n86 0.026141
R24384 DVDD.n86 DVDD.n39 0.026141
R24385 DVDD.n79 DVDD.n39 0.026141
R24386 DVDD.n80 DVDD.n79 0.026141
R24387 DVDD.n261 DVDD.n260 0.0248644
R24388 DVDD.n235 DVDD.n216 0.0248644
R24389 DVDD.n234 DVDD.n233 0.0248644
R24390 DVDD.n196 DVDD.n195 0.0248644
R24391 DVDD.n197 DVDD.n190 0.0248644
R24392 DVDD.n169 DVDD.n168 0.0248644
R24393 DVDD.n170 DVDD.n163 0.0248644
R24394 DVDD.n120 DVDD.n119 0.0247712
R24395 DVDD.n54 DVDD.n53 0.0247712
R24396 DVDD.n265 DVDD.n264 0.0246597
R24397 DVDD.n237 DVDD.n236 0.0246597
R24398 DVDD.n232 DVDD.n218 0.0246597
R24399 DVDD.n194 DVDD.n191 0.0246597
R24400 DVDD.n199 DVDD.n198 0.0246597
R24401 DVDD.n167 DVDD.n164 0.0246597
R24402 DVDD.n172 DVDD.n171 0.0246597
R24403 DVDD.n114 DVDD.n100 0.0245385
R24404 DVDD.n156 DVDD.n155 0.0245385
R24405 DVDD.n48 DVDD.n34 0.0245385
R24406 DVDD.n90 DVDD.n89 0.0245385
R24407 DVDD.n241 DVDD 0.0232879
R24408 DVDD.n189 DVDD 0.0229632
R24409 DVDD DVDD.n144 0.0224017
R24410 DVDD DVDD.n78 0.0224017
R24411 DVDD.n186 DVDD 0.0220387
R24412 DVDD.n215 DVDD 0.0220387
R24413 DVDD.n258 DVDD 0.0220387
R24414 DVDD.n213 DVDD 0.0214379
R24415 DVDD.n150 DVDD.n106 0.0198496
R24416 DVDD.n84 DVDD.n40 0.0198496
R24417 DVDD.n260 DVDD.n259 0.0195678
R24418 DVDD.n235 DVDD.n234 0.0195678
R24419 DVDD.n197 DVDD.n196 0.0195678
R24420 DVDD.n170 DVDD.n169 0.0195678
R24421 DVDD.n264 DVDD.n263 0.0194076
R24422 DVDD.n236 DVDD.n218 0.0194076
R24423 DVDD.n198 DVDD.n191 0.0194076
R24424 DVDD.n171 DVDD.n164 0.0194076
R24425 DVDD.n160 DVDD.n96 0.0143889
R24426 DVDD.n94 DVDD.n30 0.0143889
R24427 DVDD.n126 DVDD.n119 0.0138547
R24428 DVDD.n60 DVDD.n53 0.0138547
R24429 DVDD.n127 DVDD.n126 0.0127863
R24430 DVDD.n61 DVDD.n60 0.0127863
R24431 DVDD.n160 DVDD.n97 0.0122521
R24432 DVDD.n94 DVDD.n31 0.0122521
R24433 DVDD.n158 DVDD.n99 0.0111495
R24434 DVDD.n92 DVDD.n33 0.0111495
R24435 DVDD.n142 DVDD.n106 0.00878597
R24436 DVDD.n76 DVDD.n40 0.00878597
R24437 DVDD.n114 DVDD.n98 0.00797863
R24438 DVDD.n48 DVDD.n32 0.00797863
R24439 DVDD.n159 DVDD.n98 0.00691026
R24440 DVDD.n93 DVDD.n32 0.00691026
R24441 DVDD.n124 DVDD.n123 0.00486531
R24442 DVDD.n58 DVDD.n57 0.00486531
R24443 DVDD.n147 DVDD.n144 0.00423932
R24444 DVDD.n81 DVDD.n78 0.00423932
R24445 DVDD.n267 DVDD.n261 0.00367797
R24446 DVDD.n257 DVDD.n243 0.00367797
R24447 DVDD.n239 DVDD.n216 0.00367797
R24448 DVDD.n233 DVDD.n219 0.00367797
R24449 DVDD.n195 DVDD.n95 0.00367797
R24450 DVDD.n212 DVDD.n190 0.00367797
R24451 DVDD.n168 DVDD.n162 0.00367797
R24452 DVDD.n185 DVDD.n163 0.00367797
R24453 DVDD.n266 DVDD.n265 0.00365126
R24454 DVDD.n256 DVDD.n244 0.00365126
R24455 DVDD.n238 DVDD.n237 0.00365126
R24456 DVDD.n232 DVDD.n231 0.00365126
R24457 DVDD.n194 DVDD.n193 0.00365126
R24458 DVDD.n211 DVDD.n199 0.00365126
R24459 DVDD.n167 DVDD.n166 0.00365126
R24460 DVDD.n184 DVDD.n172 0.00365126
R24461 DVDD.n242 DVDD.n241 0.00299242
R24462 DVDD.n123 DVDD.n120 0.00286947
R24463 DVDD.n57 DVDD.n54 0.00286947
R24464 DVDD.n159 DVDD.n158 0.00260244
R24465 DVDD.n93 DVDD.n92 0.00260244
R24466 DVDD.n270 DVDD.n29 0.00212069
R24467 DVDD.n117 DVDD.n100 0.00210256
R24468 DVDD.n156 DVDD.n102 0.00210256
R24469 DVDD.n51 DVDD.n34 0.00210256
R24470 DVDD.n90 DVDD.n36 0.00210256
R24471 DVDD DVDD.n188 0.000856061
R24472 DVDD.n160 DVDD.n159 0.000500107
R24473 DVDD.n94 DVDD.n93 0.000500107
R24474 DVSS.n3344 DVSS.n3342 22998.7
R24475 DVSS.n4939 DVSS.n4938 19002.1
R24476 DVSS.n1726 DVSS.n1725 17372
R24477 DVSS.n1346 DVSS.n1345 11671.2
R24478 DVSS.n3 DVSS.t163 10257.4
R24479 DVSS.n6407 DVSS.n6406 9711.48
R24480 DVSS.n1741 DVSS.n1740 4670.27
R24481 DVSS.n1061 DVSS.t2 4455
R24482 DVSS.n6549 DVSS.n6548 3233.9
R24483 DVSS.n1345 DVSS.n963 2811.93
R24484 DVSS.n5059 DVSS.n5058 2240.16
R24485 DVSS.n1847 DVSS.n1846 2240.16
R24486 DVSS.t245 DVSS.t53 2192.97
R24487 DVSS.t163 DVSS.t165 2165.3
R24488 DVSS.n3463 DVSS.n3462 1972.41
R24489 DVSS.n5058 DVSS.n5057 1972.41
R24490 DVSS.n1846 DVSS.n1845 1972.41
R24491 DVSS.n1117 DVSS.n1054 1892.22
R24492 DVSS.n1124 DVSS.n969 1711.76
R24493 DVSS.n1345 DVSS.n1344 1573.68
R24494 DVSS.n1344 DVSS.n1343 1461.05
R24495 DVSS.n1230 DVSS.n1229 1372.22
R24496 DVSS.n3464 DVSS.n3463 1338.74
R24497 DVSS.n1157 DVSS.t5 1265
R24498 DVSS.n6650 DVSS.t131 1193.69
R24499 DVSS.n1892 DVSS.t114 1193.69
R24500 DVSS.n4 DVSS.n3 1170.69
R24501 DVSS.n6699 DVSS.t55 1108.71
R24502 DVSS.n6734 DVSS.t93 1108.71
R24503 DVSS.n6548 DVSS.n6547 1053.42
R24504 DVSS.n1321 DVSS.t247 1034.58
R24505 DVSS.n3917 DVSS.n3780 1013.97
R24506 DVSS.n3915 DVSS.n3781 1013.97
R24507 DVSS.n3907 DVSS.n3906 1013.97
R24508 DVSS.n3909 DVSS.n3901 1013.97
R24509 DVSS.n4382 DVSS.n4245 1013.97
R24510 DVSS.n4380 DVSS.n4246 1013.97
R24511 DVSS.n4372 DVSS.n4371 1013.97
R24512 DVSS.n4374 DVSS.n4366 1013.97
R24513 DVSS.n2321 DVSS.n2184 1013.97
R24514 DVSS.n2319 DVSS.n2185 1013.97
R24515 DVSS.n2311 DVSS.n2310 1013.97
R24516 DVSS.n2313 DVSS.n2305 1013.97
R24517 DVSS.n2786 DVSS.n2649 1013.97
R24518 DVSS.n2784 DVSS.n2650 1013.97
R24519 DVSS.n2776 DVSS.n2775 1013.97
R24520 DVSS.n2778 DVSS.n2770 1013.97
R24521 DVSS.n5385 DVSS.n5248 1013.97
R24522 DVSS.n5383 DVSS.n5249 1013.97
R24523 DVSS.n5375 DVSS.n5374 1013.97
R24524 DVSS.n5377 DVSS.n5369 1013.97
R24525 DVSS.n5850 DVSS.n5713 1013.97
R24526 DVSS.n5848 DVSS.n5714 1013.97
R24527 DVSS.n5840 DVSS.n5839 1013.97
R24528 DVSS.n5842 DVSS.n5834 1013.97
R24529 DVSS.n320 DVSS.n183 1013.97
R24530 DVSS.n318 DVSS.n184 1013.97
R24531 DVSS.n310 DVSS.n309 1013.97
R24532 DVSS.n312 DVSS.n304 1013.97
R24533 DVSS.n785 DVSS.n648 1013.97
R24534 DVSS.n783 DVSS.n649 1013.97
R24535 DVSS.n775 DVSS.n774 1013.97
R24536 DVSS.n777 DVSS.n769 1013.97
R24537 DVSS.n3478 DVSS.n3476 968.973
R24538 DVSS.n1227 DVSS.t0 868.74
R24539 DVSS.n1347 DVSS.n1346 863.648
R24540 DVSS.n1343 DVSS.n1342 755.345
R24541 DVSS.n6408 DVSS.n6407 751.22
R24542 DVSS.n4940 DVSS.n4939 751.22
R24543 DVSS.n3345 DVSS.n3344 751.22
R24544 DVSS.n1727 DVSS.n1726 751.22
R24545 DVSS.n1229 DVSS.n1228 738.889
R24546 DVSS.n3796 DVSS.n3788 728.663
R24547 DVSS.n3937 DVSS.n3762 728.663
R24548 DVSS.n4261 DVSS.n4253 728.663
R24549 DVSS.n4402 DVSS.n4227 728.663
R24550 DVSS.n2200 DVSS.n2192 728.663
R24551 DVSS.n2341 DVSS.n2166 728.663
R24552 DVSS.n2665 DVSS.n2657 728.663
R24553 DVSS.n2806 DVSS.n2631 728.663
R24554 DVSS.n5264 DVSS.n5256 728.663
R24555 DVSS.n5405 DVSS.n5230 728.663
R24556 DVSS.n5729 DVSS.n5721 728.663
R24557 DVSS.n5870 DVSS.n5695 728.663
R24558 DVSS.n199 DVSS.n191 728.663
R24559 DVSS.n340 DVSS.n165 728.663
R24560 DVSS.n664 DVSS.n656 728.663
R24561 DVSS.n805 DVSS.n630 728.663
R24562 DVSS.n1156 DVSS.t262 693.934
R24563 DVSS.n3892 DVSS.n3787 668.5
R24564 DVSS.n3890 DVSS.n3790 668.5
R24565 DVSS.n3939 DVSS.n3759 668.5
R24566 DVSS.n3899 DVSS.n3763 668.5
R24567 DVSS.n3867 DVSS.n3846 668.5
R24568 DVSS.n3871 DVSS.n3848 668.5
R24569 DVSS.n3882 DVSS.n3844 668.5
R24570 DVSS.n3885 DVSS.n3884 668.5
R24571 DVSS.n3712 DVSS.n3684 668.5
R24572 DVSS.n3697 DVSS.n3682 668.5
R24573 DVSS.n4054 DVSS.n4053 668.5
R24574 DVSS.n4070 DVSS.n4069 668.5
R24575 DVSS.n4357 DVSS.n4252 668.5
R24576 DVSS.n4355 DVSS.n4255 668.5
R24577 DVSS.n4404 DVSS.n4224 668.5
R24578 DVSS.n4364 DVSS.n4228 668.5
R24579 DVSS.n4332 DVSS.n4311 668.5
R24580 DVSS.n4336 DVSS.n4313 668.5
R24581 DVSS.n4347 DVSS.n4309 668.5
R24582 DVSS.n4350 DVSS.n4349 668.5
R24583 DVSS.n4177 DVSS.n4149 668.5
R24584 DVSS.n4162 DVSS.n4147 668.5
R24585 DVSS.n4519 DVSS.n4518 668.5
R24586 DVSS.n4534 DVSS.n4533 668.5
R24587 DVSS.n2296 DVSS.n2191 668.5
R24588 DVSS.n2294 DVSS.n2194 668.5
R24589 DVSS.n2343 DVSS.n2163 668.5
R24590 DVSS.n2303 DVSS.n2167 668.5
R24591 DVSS.n2271 DVSS.n2250 668.5
R24592 DVSS.n2275 DVSS.n2252 668.5
R24593 DVSS.n2286 DVSS.n2248 668.5
R24594 DVSS.n2289 DVSS.n2288 668.5
R24595 DVSS.n2116 DVSS.n2088 668.5
R24596 DVSS.n2101 DVSS.n2086 668.5
R24597 DVSS.n2458 DVSS.n2457 668.5
R24598 DVSS.n2474 DVSS.n2473 668.5
R24599 DVSS.n2761 DVSS.n2656 668.5
R24600 DVSS.n2759 DVSS.n2659 668.5
R24601 DVSS.n2808 DVSS.n2628 668.5
R24602 DVSS.n2768 DVSS.n2632 668.5
R24603 DVSS.n2736 DVSS.n2715 668.5
R24604 DVSS.n2740 DVSS.n2717 668.5
R24605 DVSS.n2751 DVSS.n2713 668.5
R24606 DVSS.n2754 DVSS.n2753 668.5
R24607 DVSS.n2581 DVSS.n2553 668.5
R24608 DVSS.n2566 DVSS.n2551 668.5
R24609 DVSS.n2923 DVSS.n2922 668.5
R24610 DVSS.n2938 DVSS.n2937 668.5
R24611 DVSS.n5360 DVSS.n5255 668.5
R24612 DVSS.n5358 DVSS.n5258 668.5
R24613 DVSS.n5407 DVSS.n5227 668.5
R24614 DVSS.n5367 DVSS.n5231 668.5
R24615 DVSS.n5335 DVSS.n5314 668.5
R24616 DVSS.n5339 DVSS.n5316 668.5
R24617 DVSS.n5350 DVSS.n5312 668.5
R24618 DVSS.n5353 DVSS.n5352 668.5
R24619 DVSS.n5180 DVSS.n5152 668.5
R24620 DVSS.n5165 DVSS.n5150 668.5
R24621 DVSS.n5522 DVSS.n5521 668.5
R24622 DVSS.n5538 DVSS.n5537 668.5
R24623 DVSS.n5825 DVSS.n5720 668.5
R24624 DVSS.n5823 DVSS.n5723 668.5
R24625 DVSS.n5872 DVSS.n5692 668.5
R24626 DVSS.n5832 DVSS.n5696 668.5
R24627 DVSS.n5800 DVSS.n5779 668.5
R24628 DVSS.n5804 DVSS.n5781 668.5
R24629 DVSS.n5815 DVSS.n5777 668.5
R24630 DVSS.n5818 DVSS.n5817 668.5
R24631 DVSS.n5645 DVSS.n5617 668.5
R24632 DVSS.n5630 DVSS.n5615 668.5
R24633 DVSS.n5987 DVSS.n5986 668.5
R24634 DVSS.n6002 DVSS.n6001 668.5
R24635 DVSS.n295 DVSS.n190 668.5
R24636 DVSS.n293 DVSS.n193 668.5
R24637 DVSS.n342 DVSS.n162 668.5
R24638 DVSS.n302 DVSS.n166 668.5
R24639 DVSS.n270 DVSS.n249 668.5
R24640 DVSS.n274 DVSS.n251 668.5
R24641 DVSS.n285 DVSS.n247 668.5
R24642 DVSS.n288 DVSS.n287 668.5
R24643 DVSS.n115 DVSS.n87 668.5
R24644 DVSS.n100 DVSS.n85 668.5
R24645 DVSS.n457 DVSS.n456 668.5
R24646 DVSS.n473 DVSS.n472 668.5
R24647 DVSS.n760 DVSS.n655 668.5
R24648 DVSS.n758 DVSS.n658 668.5
R24649 DVSS.n807 DVSS.n627 668.5
R24650 DVSS.n767 DVSS.n631 668.5
R24651 DVSS.n735 DVSS.n714 668.5
R24652 DVSS.n739 DVSS.n716 668.5
R24653 DVSS.n750 DVSS.n712 668.5
R24654 DVSS.n753 DVSS.n752 668.5
R24655 DVSS.n580 DVSS.n552 668.5
R24656 DVSS.n565 DVSS.n550 668.5
R24657 DVSS.n922 DVSS.n921 668.5
R24658 DVSS.n937 DVSS.n936 668.5
R24659 DVSS.t172 DVSS.n1157 643.51
R24660 DVSS.n1054 DVSS.n1053 590.426
R24661 DVSS.n3981 DVSS.n3646 562.173
R24662 DVSS.n4029 DVSS.n3630 562.173
R24663 DVSS.n4446 DVSS.n4111 562.173
R24664 DVSS.n4494 DVSS.n4095 562.173
R24665 DVSS.n2385 DVSS.n2050 562.173
R24666 DVSS.n2433 DVSS.n2034 562.173
R24667 DVSS.n2850 DVSS.n2515 562.173
R24668 DVSS.n2898 DVSS.n2499 562.173
R24669 DVSS.n5449 DVSS.n5114 562.173
R24670 DVSS.n5497 DVSS.n5098 562.173
R24671 DVSS.n5914 DVSS.n5579 562.173
R24672 DVSS.n5962 DVSS.n5563 562.173
R24673 DVSS.n384 DVSS.n49 562.173
R24674 DVSS.n432 DVSS.n33 562.173
R24675 DVSS.n849 DVSS.n514 562.173
R24676 DVSS.n897 DVSS.n498 562.173
R24677 DVSS.n3908 DVSS.n3904 535.801
R24678 DVSS.n4373 DVSS.n4369 535.801
R24679 DVSS.n2312 DVSS.n2308 535.801
R24680 DVSS.n2777 DVSS.n2773 535.801
R24681 DVSS.n5376 DVSS.n5372 535.801
R24682 DVSS.n5841 DVSS.n5837 535.801
R24683 DVSS.n311 DVSS.n307 535.801
R24684 DVSS.n776 DVSS.n772 535.801
R24685 DVSS.n3869 DVSS.n3847 518.471
R24686 DVSS.n3883 DVSS.n3796 518.471
R24687 DVSS.n3891 DVSS.n3788 518.471
R24688 DVSS.n3937 DVSS.n3761 518.471
R24689 DVSS.n4334 DVSS.n4312 518.471
R24690 DVSS.n4348 DVSS.n4261 518.471
R24691 DVSS.n4356 DVSS.n4253 518.471
R24692 DVSS.n4402 DVSS.n4226 518.471
R24693 DVSS.n2273 DVSS.n2251 518.471
R24694 DVSS.n2287 DVSS.n2200 518.471
R24695 DVSS.n2295 DVSS.n2192 518.471
R24696 DVSS.n2341 DVSS.n2165 518.471
R24697 DVSS.n2738 DVSS.n2716 518.471
R24698 DVSS.n2752 DVSS.n2665 518.471
R24699 DVSS.n2760 DVSS.n2657 518.471
R24700 DVSS.n2806 DVSS.n2630 518.471
R24701 DVSS.n5337 DVSS.n5315 518.471
R24702 DVSS.n5351 DVSS.n5264 518.471
R24703 DVSS.n5359 DVSS.n5256 518.471
R24704 DVSS.n5405 DVSS.n5229 518.471
R24705 DVSS.n5802 DVSS.n5780 518.471
R24706 DVSS.n5816 DVSS.n5729 518.471
R24707 DVSS.n5824 DVSS.n5721 518.471
R24708 DVSS.n5870 DVSS.n5694 518.471
R24709 DVSS.n272 DVSS.n250 518.471
R24710 DVSS.n286 DVSS.n199 518.471
R24711 DVSS.n294 DVSS.n191 518.471
R24712 DVSS.n340 DVSS.n164 518.471
R24713 DVSS.n737 DVSS.n715 518.471
R24714 DVSS.n751 DVSS.n664 518.471
R24715 DVSS.n759 DVSS.n656 518.471
R24716 DVSS.n805 DVSS.n629 518.471
R24717 DVSS.n3477 DVSS.t245 506.07
R24718 DVSS.n3711 DVSS.n3683 491.349
R24719 DVSS.n3967 DVSS.n3646 491.349
R24720 DVSS.n3630 DVSS.n3621 491.349
R24721 DVSS.n4051 DVSS.n3615 491.349
R24722 DVSS.n4176 DVSS.n4148 491.349
R24723 DVSS.n4432 DVSS.n4111 491.349
R24724 DVSS.n4095 DVSS.n4086 491.349
R24725 DVSS.n4516 DVSS.n4080 491.349
R24726 DVSS.n2115 DVSS.n2087 491.349
R24727 DVSS.n2371 DVSS.n2050 491.349
R24728 DVSS.n2034 DVSS.n2025 491.349
R24729 DVSS.n2455 DVSS.n2019 491.349
R24730 DVSS.n2580 DVSS.n2552 491.349
R24731 DVSS.n2836 DVSS.n2515 491.349
R24732 DVSS.n2499 DVSS.n2490 491.349
R24733 DVSS.n2920 DVSS.n2484 491.349
R24734 DVSS.n5179 DVSS.n5151 491.349
R24735 DVSS.n5435 DVSS.n5114 491.349
R24736 DVSS.n5098 DVSS.n5089 491.349
R24737 DVSS.n5519 DVSS.n5083 491.349
R24738 DVSS.n5644 DVSS.n5616 491.349
R24739 DVSS.n5900 DVSS.n5579 491.349
R24740 DVSS.n5563 DVSS.n5554 491.349
R24741 DVSS.n5984 DVSS.n5548 491.349
R24742 DVSS.n114 DVSS.n86 491.349
R24743 DVSS.n370 DVSS.n49 491.349
R24744 DVSS.n33 DVSS.n24 491.349
R24745 DVSS.n454 DVSS.n18 491.349
R24746 DVSS.n579 DVSS.n551 491.349
R24747 DVSS.n835 DVSS.n514 491.349
R24748 DVSS.n498 DVSS.n489 491.349
R24749 DVSS.n919 DVSS.n483 491.349
R24750 DVSS.n6645 DVSS.n6644 469.046
R24751 DVSS.n3506 DVSS.n3505 468.613
R24752 DVSS.n1904 DVSS.n1903 468.277
R24753 DVSS.n6859 DVSS.n6858 468.277
R24754 DVSS.n1117 DVSS.t154 468.178
R24755 DVSS.n3903 DVSS.n3762 448.409
R24756 DVSS.n4368 DVSS.n4227 448.409
R24757 DVSS.n2307 DVSS.n2166 448.409
R24758 DVSS.n2772 DVSS.n2631 448.409
R24759 DVSS.n5371 DVSS.n5230 448.409
R24760 DVSS.n5836 DVSS.n5695 448.409
R24761 DVSS.n306 DVSS.n165 448.409
R24762 DVSS.n771 DVSS.n630 448.409
R24763 DVSS.n3901 DVSS.n3781 394
R24764 DVSS.n4366 DVSS.n4246 394
R24765 DVSS.n2305 DVSS.n2185 394
R24766 DVSS.n2770 DVSS.n2650 394
R24767 DVSS.n5369 DVSS.n5249 394
R24768 DVSS.n5834 DVSS.n5714 394
R24769 DVSS.n304 DVSS.n184 394
R24770 DVSS.n769 DVSS.n649 394
R24771 DVSS.n6718 DVSS.n6717 390.654
R24772 DVSS.n6693 DVSS.n6692 390.654
R24773 DVSS.t0 DVSS.t157 390.324
R24774 DVSS.n6753 DVSS.n6752 389.442
R24775 DVSS.n6728 DVSS.n6727 389.442
R24776 DVSS.n4005 DVSS.n3628 366.841
R24777 DVSS.n4020 DVSS.n3632 366.841
R24778 DVSS.n3659 DVSS.n3645 366.841
R24779 DVSS.n3675 DVSS.n3648 366.841
R24780 DVSS.n4470 DVSS.n4093 366.841
R24781 DVSS.n4485 DVSS.n4097 366.841
R24782 DVSS.n4124 DVSS.n4110 366.841
R24783 DVSS.n4140 DVSS.n4113 366.841
R24784 DVSS.n2409 DVSS.n2032 366.841
R24785 DVSS.n2424 DVSS.n2036 366.841
R24786 DVSS.n2063 DVSS.n2049 366.841
R24787 DVSS.n2079 DVSS.n2052 366.841
R24788 DVSS.n2874 DVSS.n2497 366.841
R24789 DVSS.n2889 DVSS.n2501 366.841
R24790 DVSS.n2528 DVSS.n2514 366.841
R24791 DVSS.n2544 DVSS.n2517 366.841
R24792 DVSS.n5473 DVSS.n5096 366.841
R24793 DVSS.n5488 DVSS.n5100 366.841
R24794 DVSS.n5127 DVSS.n5113 366.841
R24795 DVSS.n5143 DVSS.n5116 366.841
R24796 DVSS.n5938 DVSS.n5561 366.841
R24797 DVSS.n5953 DVSS.n5565 366.841
R24798 DVSS.n5592 DVSS.n5578 366.841
R24799 DVSS.n5608 DVSS.n5581 366.841
R24800 DVSS.n408 DVSS.n31 366.841
R24801 DVSS.n423 DVSS.n35 366.841
R24802 DVSS.n62 DVSS.n48 366.841
R24803 DVSS.n78 DVSS.n51 366.841
R24804 DVSS.n873 DVSS.n496 366.841
R24805 DVSS.n888 DVSS.n500 366.841
R24806 DVSS.n527 DVSS.n513 366.841
R24807 DVSS.n543 DVSS.n516 366.841
R24808 DVSS.n1124 DVSS.t145 356.863
R24809 DVSS.t160 DVSS.n1061 349.909
R24810 DVSS.n1755 DVSS.t232 339.149
R24811 DVSS.n4967 DVSS.t170 339.149
R24812 DVSS.n3372 DVSS.t69 339.149
R24813 DVSS.n6435 DVSS.t258 339.149
R24814 DVSS.n3877 DVSS.n3847 317.623
R24815 DVSS.n3883 DVSS.n3795 317.623
R24816 DVSS.n3891 DVSS.n3789 317.623
R24817 DVSS.n3897 DVSS.n3761 317.623
R24818 DVSS.n4342 DVSS.n4312 317.623
R24819 DVSS.n4348 DVSS.n4260 317.623
R24820 DVSS.n4356 DVSS.n4254 317.623
R24821 DVSS.n4362 DVSS.n4226 317.623
R24822 DVSS.n2281 DVSS.n2251 317.623
R24823 DVSS.n2287 DVSS.n2199 317.623
R24824 DVSS.n2295 DVSS.n2193 317.623
R24825 DVSS.n2301 DVSS.n2165 317.623
R24826 DVSS.n2746 DVSS.n2716 317.623
R24827 DVSS.n2752 DVSS.n2664 317.623
R24828 DVSS.n2760 DVSS.n2658 317.623
R24829 DVSS.n2766 DVSS.n2630 317.623
R24830 DVSS.n5345 DVSS.n5315 317.623
R24831 DVSS.n5351 DVSS.n5263 317.623
R24832 DVSS.n5359 DVSS.n5257 317.623
R24833 DVSS.n5365 DVSS.n5229 317.623
R24834 DVSS.n5810 DVSS.n5780 317.623
R24835 DVSS.n5816 DVSS.n5728 317.623
R24836 DVSS.n5824 DVSS.n5722 317.623
R24837 DVSS.n5830 DVSS.n5694 317.623
R24838 DVSS.n280 DVSS.n250 317.623
R24839 DVSS.n286 DVSS.n198 317.623
R24840 DVSS.n294 DVSS.n192 317.623
R24841 DVSS.n300 DVSS.n164 317.623
R24842 DVSS.n745 DVSS.n715 317.623
R24843 DVSS.n751 DVSS.n663 317.623
R24844 DVSS.n759 DVSS.n657 317.623
R24845 DVSS.n765 DVSS.n629 317.623
R24846 DVSS.n3980 DVSS.n3648 306.26
R24847 DVSS.n4028 DVSS.n3632 306.26
R24848 DVSS.n3982 DVSS.n3645 306.26
R24849 DVSS.n4030 DVSS.n3628 306.26
R24850 DVSS.n4445 DVSS.n4113 306.26
R24851 DVSS.n4493 DVSS.n4097 306.26
R24852 DVSS.n4447 DVSS.n4110 306.26
R24853 DVSS.n4495 DVSS.n4093 306.26
R24854 DVSS.n2384 DVSS.n2052 306.26
R24855 DVSS.n2432 DVSS.n2036 306.26
R24856 DVSS.n2386 DVSS.n2049 306.26
R24857 DVSS.n2434 DVSS.n2032 306.26
R24858 DVSS.n2849 DVSS.n2517 306.26
R24859 DVSS.n2897 DVSS.n2501 306.26
R24860 DVSS.n2851 DVSS.n2514 306.26
R24861 DVSS.n2899 DVSS.n2497 306.26
R24862 DVSS.n5448 DVSS.n5116 306.26
R24863 DVSS.n5496 DVSS.n5100 306.26
R24864 DVSS.n5450 DVSS.n5113 306.26
R24865 DVSS.n5498 DVSS.n5096 306.26
R24866 DVSS.n5913 DVSS.n5581 306.26
R24867 DVSS.n5961 DVSS.n5565 306.26
R24868 DVSS.n5915 DVSS.n5578 306.26
R24869 DVSS.n5963 DVSS.n5561 306.26
R24870 DVSS.n383 DVSS.n51 306.26
R24871 DVSS.n431 DVSS.n35 306.26
R24872 DVSS.n385 DVSS.n48 306.26
R24873 DVSS.n433 DVSS.n31 306.26
R24874 DVSS.n848 DVSS.n516 306.26
R24875 DVSS.n896 DVSS.n500 306.26
R24876 DVSS.n850 DVSS.n513 306.26
R24877 DVSS.n898 DVSS.n496 306.26
R24878 DVSS.n3961 DVSS.n3683 301.007
R24879 DVSS.n3967 DVSS.n3679 301.007
R24880 DVSS.n3981 DVSS.n3647 301.007
R24881 DVSS.n3988 DVSS.n3641 301.007
R24882 DVSS.n4029 DVSS.n3629 301.007
R24883 DVSS.n4059 DVSS.n3621 301.007
R24884 DVSS.n3623 DVSS.n3615 301.007
R24885 DVSS.n4426 DVSS.n4148 301.007
R24886 DVSS.n4432 DVSS.n4144 301.007
R24887 DVSS.n4446 DVSS.n4112 301.007
R24888 DVSS.n4453 DVSS.n4106 301.007
R24889 DVSS.n4494 DVSS.n4094 301.007
R24890 DVSS.n4524 DVSS.n4086 301.007
R24891 DVSS.n4088 DVSS.n4080 301.007
R24892 DVSS.n2365 DVSS.n2087 301.007
R24893 DVSS.n2371 DVSS.n2083 301.007
R24894 DVSS.n2385 DVSS.n2051 301.007
R24895 DVSS.n2392 DVSS.n2045 301.007
R24896 DVSS.n2433 DVSS.n2033 301.007
R24897 DVSS.n2463 DVSS.n2025 301.007
R24898 DVSS.n2027 DVSS.n2019 301.007
R24899 DVSS.n2830 DVSS.n2552 301.007
R24900 DVSS.n2836 DVSS.n2548 301.007
R24901 DVSS.n2850 DVSS.n2516 301.007
R24902 DVSS.n2857 DVSS.n2510 301.007
R24903 DVSS.n2898 DVSS.n2498 301.007
R24904 DVSS.n2928 DVSS.n2490 301.007
R24905 DVSS.n2492 DVSS.n2484 301.007
R24906 DVSS.n5429 DVSS.n5151 301.007
R24907 DVSS.n5435 DVSS.n5147 301.007
R24908 DVSS.n5449 DVSS.n5115 301.007
R24909 DVSS.n5456 DVSS.n5109 301.007
R24910 DVSS.n5497 DVSS.n5097 301.007
R24911 DVSS.n5527 DVSS.n5089 301.007
R24912 DVSS.n5091 DVSS.n5083 301.007
R24913 DVSS.n5894 DVSS.n5616 301.007
R24914 DVSS.n5900 DVSS.n5612 301.007
R24915 DVSS.n5914 DVSS.n5580 301.007
R24916 DVSS.n5921 DVSS.n5574 301.007
R24917 DVSS.n5962 DVSS.n5562 301.007
R24918 DVSS.n5992 DVSS.n5554 301.007
R24919 DVSS.n5556 DVSS.n5548 301.007
R24920 DVSS.n364 DVSS.n86 301.007
R24921 DVSS.n370 DVSS.n82 301.007
R24922 DVSS.n384 DVSS.n50 301.007
R24923 DVSS.n391 DVSS.n44 301.007
R24924 DVSS.n432 DVSS.n32 301.007
R24925 DVSS.n462 DVSS.n24 301.007
R24926 DVSS.n26 DVSS.n18 301.007
R24927 DVSS.n829 DVSS.n551 301.007
R24928 DVSS.n835 DVSS.n547 301.007
R24929 DVSS.n849 DVSS.n515 301.007
R24930 DVSS.n856 DVSS.n509 301.007
R24931 DVSS.n897 DVSS.n497 301.007
R24932 DVSS.n927 DVSS.n489 301.007
R24933 DVSS.n491 DVSS.n483 301.007
R24934 DVSS.n3884 DVSS.n3791 292.5
R24935 DVSS.n3884 DVSS.n3883 292.5
R24936 DVSS.n3900 DVSS.n3899 292.5
R24937 DVSS.n3899 DVSS.n3761 292.5
R24938 DVSS.n3867 DVSS.n3866 292.5
R24939 DVSS.n3865 DVSS.n3854 292.5
R24940 DVSS.n3864 DVSS.n3863 292.5
R24941 DVSS.n3862 DVSS.n3861 292.5
R24942 DVSS.n3860 DVSS.n3859 292.5
R24943 DVSS.n3858 DVSS.n3857 292.5
R24944 DVSS.n3856 DVSS.n3855 292.5
R24945 DVSS.n3850 DVSS.n3849 292.5
R24946 DVSS.n3898 DVSS.n3783 292.5
R24947 DVSS.n3898 DVSS.n3897 292.5
R24948 DVSS.n3888 DVSS.n3784 292.5
R24949 DVSS.n3789 DVSS.n3784 292.5
R24950 DVSS.n3876 DVSS.n3875 292.5
R24951 DVSS.n3877 DVSS.n3876 292.5
R24952 DVSS.n3874 DVSS.n3794 292.5
R24953 DVSS.n3795 DVSS.n3794 292.5
R24954 DVSS.n3890 DVSS.n3889 292.5
R24955 DVSS.n3891 DVSS.n3890 292.5
R24956 DVSS.n3872 DVSS.n3871 292.5
R24957 DVSS.n3873 DVSS.n3848 292.5
R24958 DVSS.n3848 DVSS.n3847 292.5
R24959 DVSS.n3911 DVSS.n3901 292.5
R24960 DVSS.n3904 DVSS.n3901 292.5
R24961 DVSS.n3912 DVSS.n3781 292.5
R24962 DVSS.n3903 DVSS.n3781 292.5
R24963 DVSS.n3910 DVSS.n3909 292.5
R24964 DVSS.n3907 DVSS.n3902 292.5
R24965 DVSS.n3918 DVSS.n3917 292.5
R24966 DVSS.n3920 DVSS.n3919 292.5
R24967 DVSS.n3782 DVSS.n3763 292.5
R24968 DVSS.n3937 DVSS.n3763 292.5
R24969 DVSS.n3915 DVSS.n3914 292.5
R24970 DVSS.n3906 DVSS.n3904 292.5
R24971 DVSS.n3903 DVSS.n3780 292.5
R24972 DVSS.n3778 DVSS.n3777 292.5
R24973 DVSS.n3926 DVSS.n3925 292.5
R24974 DVSS.n3929 DVSS.n3928 292.5
R24975 DVSS.n3772 DVSS.n3771 292.5
R24976 DVSS.n3935 DVSS.n3934 292.5
R24977 DVSS.n3769 DVSS.n3760 292.5
R24978 DVSS.n3940 DVSS.n3939 292.5
R24979 DVSS.n3759 DVSS.n3757 292.5
R24980 DVSS.n3761 DVSS.n3759 292.5
R24981 DVSS.n3896 DVSS.n3895 292.5
R24982 DVSS.n3897 DVSS.n3896 292.5
R24983 DVSS.n3894 DVSS.n3785 292.5
R24984 DVSS.n3789 DVSS.n3785 292.5
R24985 DVSS.n3893 DVSS.n3892 292.5
R24986 DVSS.n3892 DVSS.n3891 292.5
R24987 DVSS.n3846 DVSS.n3845 292.5
R24988 DVSS.n3847 DVSS.n3846 292.5
R24989 DVSS.n3879 DVSS.n3878 292.5
R24990 DVSS.n3878 DVSS.n3877 292.5
R24991 DVSS.n3880 DVSS.n3797 292.5
R24992 DVSS.n3797 DVSS.n3795 292.5
R24993 DVSS.n3882 DVSS.n3881 292.5
R24994 DVSS.n3883 DVSS.n3882 292.5
R24995 DVSS.n3886 DVSS.n3790 292.5
R24996 DVSS.n3844 DVSS.n3843 292.5
R24997 DVSS.n3843 DVSS.n3787 292.5
R24998 DVSS.n3802 DVSS.n3800 292.5
R24999 DVSS.n3807 DVSS.n3800 292.5
R25000 DVSS.n3838 DVSS.n3804 292.5
R25001 DVSS.n3838 DVSS.n3837 292.5
R25002 DVSS.n3812 DVSS.n3809 292.5
R25003 DVSS.n3836 DVSS.n3809 292.5
R25004 DVSS.n3833 DVSS.n3814 292.5
R25005 DVSS.n3834 DVSS.n3833 292.5
R25006 DVSS.n3819 DVSS.n3815 292.5
R25007 DVSS.n3815 DVSS.n3810 292.5
R25008 DVSS.n3828 DVSS.n3821 292.5
R25009 DVSS.n3828 DVSS.n3827 292.5
R25010 DVSS.n3826 DVSS.n3824 292.5
R25011 DVSS.n3824 DVSS.n3823 292.5
R25012 DVSS.n3886 DVSS.n3885 292.5
R25013 DVSS.n3698 DVSS.n3697 292.5
R25014 DVSS.n3689 DVSS.n3688 292.5
R25015 DVSS.n3701 DVSS.n3700 292.5
R25016 DVSS.n3703 DVSS.n3702 292.5
R25017 DVSS.n3705 DVSS.n3704 292.5
R25018 DVSS.n3707 DVSS.n3706 292.5
R25019 DVSS.n3709 DVSS.n3708 292.5
R25020 DVSS.n3699 DVSS.n3696 292.5
R25021 DVSS.n3713 DVSS.n3712 292.5
R25022 DVSS.n3712 DVSS.n3711 292.5
R25023 DVSS.n4005 DVSS.n3625 292.5
R25024 DVSS.n4005 DVSS.n3630 292.5
R25025 DVSS.n4018 DVSS.n4001 292.5
R25026 DVSS.n4017 DVSS.n4016 292.5
R25027 DVSS.n4015 DVSS.n4014 292.5
R25028 DVSS.n4013 DVSS.n4003 292.5
R25029 DVSS.n4011 DVSS.n4010 292.5
R25030 DVSS.n4009 DVSS.n4004 292.5
R25031 DVSS.n4008 DVSS.n4007 292.5
R25032 DVSS.n4021 DVSS.n4020 292.5
R25033 DVSS.n3661 DVSS.n3657 292.5
R25034 DVSS.n3674 DVSS.n3653 292.5
R25035 DVSS.n3672 DVSS.n3671 292.5
R25036 DVSS.n3670 DVSS.n3669 292.5
R25037 DVSS.n3667 DVSS.n3655 292.5
R25038 DVSS.n3665 DVSS.n3664 292.5
R25039 DVSS.n3663 DVSS.n3662 292.5
R25040 DVSS.n3676 DVSS.n3675 292.5
R25041 DVSS.n3675 DVSS.n3646 292.5
R25042 DVSS.n3659 DVSS.n3658 292.5
R25043 DVSS.n4055 DVSS.n4054 292.5
R25044 DVSS.n4054 DVSS.n3615 292.5
R25045 DVSS.n4056 DVSS.n3624 292.5
R25046 DVSS.n3624 DVSS.n3623 292.5
R25047 DVSS.n4058 DVSS.n4057 292.5
R25048 DVSS.n4059 DVSS.n4058 292.5
R25049 DVSS.n4033 DVSS.n3622 292.5
R25050 DVSS.n3622 DVSS.n3621 292.5
R25051 DVSS.n4031 DVSS.n4030 292.5
R25052 DVSS.n4030 DVSS.n4029 292.5
R25053 DVSS.n3627 DVSS.n3626 292.5
R25054 DVSS.n3629 DVSS.n3627 292.5
R25055 DVSS.n3985 DVSS.n3643 292.5
R25056 DVSS.n3643 DVSS.n3641 292.5
R25057 DVSS.n3987 DVSS.n3986 292.5
R25058 DVSS.n3988 DVSS.n3987 292.5
R25059 DVSS.n3984 DVSS.n3642 292.5
R25060 DVSS.n3647 DVSS.n3642 292.5
R25061 DVSS.n3983 DVSS.n3982 292.5
R25062 DVSS.n3982 DVSS.n3981 292.5
R25063 DVSS.n3966 DVSS.n3965 292.5
R25064 DVSS.n3967 DVSS.n3966 292.5
R25065 DVSS.n3964 DVSS.n3680 292.5
R25066 DVSS.n3680 DVSS.n3679 292.5
R25067 DVSS.n3963 DVSS.n3962 292.5
R25068 DVSS.n3962 DVSS.n3961 292.5
R25069 DVSS.n3682 DVSS.n3681 292.5
R25070 DVSS.n3683 DVSS.n3682 292.5
R25071 DVSS.n4053 DVSS.n4034 292.5
R25072 DVSS.n4039 DVSS.n4035 292.5
R25073 DVSS.n4049 DVSS.n4048 292.5
R25074 DVSS.n4047 DVSS.n4038 292.5
R25075 DVSS.n4046 DVSS.n4045 292.5
R25076 DVSS.n4044 DVSS.n4043 292.5
R25077 DVSS.n4042 DVSS.n4041 292.5
R25078 DVSS.n4040 DVSS.n3612 292.5
R25079 DVSS.n4071 DVSS.n4070 292.5
R25080 DVSS.n4349 DVSS.n4256 292.5
R25081 DVSS.n4349 DVSS.n4348 292.5
R25082 DVSS.n4365 DVSS.n4364 292.5
R25083 DVSS.n4364 DVSS.n4226 292.5
R25084 DVSS.n4332 DVSS.n4331 292.5
R25085 DVSS.n4330 DVSS.n4319 292.5
R25086 DVSS.n4329 DVSS.n4328 292.5
R25087 DVSS.n4327 DVSS.n4326 292.5
R25088 DVSS.n4325 DVSS.n4324 292.5
R25089 DVSS.n4323 DVSS.n4322 292.5
R25090 DVSS.n4321 DVSS.n4320 292.5
R25091 DVSS.n4315 DVSS.n4314 292.5
R25092 DVSS.n4363 DVSS.n4248 292.5
R25093 DVSS.n4363 DVSS.n4362 292.5
R25094 DVSS.n4353 DVSS.n4249 292.5
R25095 DVSS.n4254 DVSS.n4249 292.5
R25096 DVSS.n4341 DVSS.n4340 292.5
R25097 DVSS.n4342 DVSS.n4341 292.5
R25098 DVSS.n4339 DVSS.n4259 292.5
R25099 DVSS.n4260 DVSS.n4259 292.5
R25100 DVSS.n4355 DVSS.n4354 292.5
R25101 DVSS.n4356 DVSS.n4355 292.5
R25102 DVSS.n4337 DVSS.n4336 292.5
R25103 DVSS.n4338 DVSS.n4313 292.5
R25104 DVSS.n4313 DVSS.n4312 292.5
R25105 DVSS.n4376 DVSS.n4366 292.5
R25106 DVSS.n4369 DVSS.n4366 292.5
R25107 DVSS.n4377 DVSS.n4246 292.5
R25108 DVSS.n4368 DVSS.n4246 292.5
R25109 DVSS.n4375 DVSS.n4374 292.5
R25110 DVSS.n4372 DVSS.n4367 292.5
R25111 DVSS.n4383 DVSS.n4382 292.5
R25112 DVSS.n4385 DVSS.n4384 292.5
R25113 DVSS.n4247 DVSS.n4228 292.5
R25114 DVSS.n4402 DVSS.n4228 292.5
R25115 DVSS.n4380 DVSS.n4379 292.5
R25116 DVSS.n4371 DVSS.n4369 292.5
R25117 DVSS.n4368 DVSS.n4245 292.5
R25118 DVSS.n4243 DVSS.n4242 292.5
R25119 DVSS.n4391 DVSS.n4390 292.5
R25120 DVSS.n4394 DVSS.n4393 292.5
R25121 DVSS.n4237 DVSS.n4236 292.5
R25122 DVSS.n4400 DVSS.n4399 292.5
R25123 DVSS.n4234 DVSS.n4225 292.5
R25124 DVSS.n4405 DVSS.n4404 292.5
R25125 DVSS.n4224 DVSS.n4222 292.5
R25126 DVSS.n4226 DVSS.n4224 292.5
R25127 DVSS.n4361 DVSS.n4360 292.5
R25128 DVSS.n4362 DVSS.n4361 292.5
R25129 DVSS.n4359 DVSS.n4250 292.5
R25130 DVSS.n4254 DVSS.n4250 292.5
R25131 DVSS.n4358 DVSS.n4357 292.5
R25132 DVSS.n4357 DVSS.n4356 292.5
R25133 DVSS.n4311 DVSS.n4310 292.5
R25134 DVSS.n4312 DVSS.n4311 292.5
R25135 DVSS.n4344 DVSS.n4343 292.5
R25136 DVSS.n4343 DVSS.n4342 292.5
R25137 DVSS.n4345 DVSS.n4262 292.5
R25138 DVSS.n4262 DVSS.n4260 292.5
R25139 DVSS.n4347 DVSS.n4346 292.5
R25140 DVSS.n4348 DVSS.n4347 292.5
R25141 DVSS.n4351 DVSS.n4255 292.5
R25142 DVSS.n4309 DVSS.n4308 292.5
R25143 DVSS.n4308 DVSS.n4252 292.5
R25144 DVSS.n4267 DVSS.n4265 292.5
R25145 DVSS.n4272 DVSS.n4265 292.5
R25146 DVSS.n4303 DVSS.n4269 292.5
R25147 DVSS.n4303 DVSS.n4302 292.5
R25148 DVSS.n4277 DVSS.n4274 292.5
R25149 DVSS.n4301 DVSS.n4274 292.5
R25150 DVSS.n4298 DVSS.n4279 292.5
R25151 DVSS.n4299 DVSS.n4298 292.5
R25152 DVSS.n4284 DVSS.n4280 292.5
R25153 DVSS.n4280 DVSS.n4275 292.5
R25154 DVSS.n4293 DVSS.n4286 292.5
R25155 DVSS.n4293 DVSS.n4292 292.5
R25156 DVSS.n4291 DVSS.n4289 292.5
R25157 DVSS.n4289 DVSS.n4288 292.5
R25158 DVSS.n4351 DVSS.n4350 292.5
R25159 DVSS.n4163 DVSS.n4162 292.5
R25160 DVSS.n4154 DVSS.n4153 292.5
R25161 DVSS.n4166 DVSS.n4165 292.5
R25162 DVSS.n4168 DVSS.n4167 292.5
R25163 DVSS.n4170 DVSS.n4169 292.5
R25164 DVSS.n4172 DVSS.n4171 292.5
R25165 DVSS.n4174 DVSS.n4173 292.5
R25166 DVSS.n4164 DVSS.n4161 292.5
R25167 DVSS.n4178 DVSS.n4177 292.5
R25168 DVSS.n4177 DVSS.n4176 292.5
R25169 DVSS.n4470 DVSS.n4090 292.5
R25170 DVSS.n4470 DVSS.n4095 292.5
R25171 DVSS.n4483 DVSS.n4466 292.5
R25172 DVSS.n4482 DVSS.n4481 292.5
R25173 DVSS.n4480 DVSS.n4479 292.5
R25174 DVSS.n4478 DVSS.n4468 292.5
R25175 DVSS.n4476 DVSS.n4475 292.5
R25176 DVSS.n4474 DVSS.n4469 292.5
R25177 DVSS.n4473 DVSS.n4472 292.5
R25178 DVSS.n4486 DVSS.n4485 292.5
R25179 DVSS.n4126 DVSS.n4122 292.5
R25180 DVSS.n4139 DVSS.n4118 292.5
R25181 DVSS.n4137 DVSS.n4136 292.5
R25182 DVSS.n4135 DVSS.n4134 292.5
R25183 DVSS.n4132 DVSS.n4120 292.5
R25184 DVSS.n4130 DVSS.n4129 292.5
R25185 DVSS.n4128 DVSS.n4127 292.5
R25186 DVSS.n4141 DVSS.n4140 292.5
R25187 DVSS.n4140 DVSS.n4111 292.5
R25188 DVSS.n4124 DVSS.n4123 292.5
R25189 DVSS.n4520 DVSS.n4519 292.5
R25190 DVSS.n4519 DVSS.n4080 292.5
R25191 DVSS.n4521 DVSS.n4089 292.5
R25192 DVSS.n4089 DVSS.n4088 292.5
R25193 DVSS.n4523 DVSS.n4522 292.5
R25194 DVSS.n4524 DVSS.n4523 292.5
R25195 DVSS.n4498 DVSS.n4087 292.5
R25196 DVSS.n4087 DVSS.n4086 292.5
R25197 DVSS.n4496 DVSS.n4495 292.5
R25198 DVSS.n4495 DVSS.n4494 292.5
R25199 DVSS.n4092 DVSS.n4091 292.5
R25200 DVSS.n4094 DVSS.n4092 292.5
R25201 DVSS.n4450 DVSS.n4108 292.5
R25202 DVSS.n4108 DVSS.n4106 292.5
R25203 DVSS.n4452 DVSS.n4451 292.5
R25204 DVSS.n4453 DVSS.n4452 292.5
R25205 DVSS.n4449 DVSS.n4107 292.5
R25206 DVSS.n4112 DVSS.n4107 292.5
R25207 DVSS.n4448 DVSS.n4447 292.5
R25208 DVSS.n4447 DVSS.n4446 292.5
R25209 DVSS.n4431 DVSS.n4430 292.5
R25210 DVSS.n4432 DVSS.n4431 292.5
R25211 DVSS.n4429 DVSS.n4145 292.5
R25212 DVSS.n4145 DVSS.n4144 292.5
R25213 DVSS.n4428 DVSS.n4427 292.5
R25214 DVSS.n4427 DVSS.n4426 292.5
R25215 DVSS.n4147 DVSS.n4146 292.5
R25216 DVSS.n4148 DVSS.n4147 292.5
R25217 DVSS.n4518 DVSS.n4499 292.5
R25218 DVSS.n4504 DVSS.n4500 292.5
R25219 DVSS.n4514 DVSS.n4513 292.5
R25220 DVSS.n4512 DVSS.n4503 292.5
R25221 DVSS.n4511 DVSS.n4510 292.5
R25222 DVSS.n4509 DVSS.n4508 292.5
R25223 DVSS.n4507 DVSS.n4506 292.5
R25224 DVSS.n4505 DVSS.n4077 292.5
R25225 DVSS.n4535 DVSS.n4534 292.5
R25226 DVSS.n6400 DVSS.n6399 292.5
R25227 DVSS.n6402 DVSS.n6401 292.5
R25228 DVSS.n6405 DVSS.n6404 292.5
R25229 DVSS.n6411 DVSS.n6410 292.5
R25230 DVSS.n6397 DVSS.n6396 292.5
R25231 DVSS.n6378 DVSS.n6376 292.5
R25232 DVSS.n6363 DVSS.n6361 292.5
R25233 DVSS.n6348 DVSS.n6346 292.5
R25234 DVSS.n6345 DVSS.n6344 292.5
R25235 DVSS.n6322 DVSS.n6321 292.5
R25236 DVSS.n6320 DVSS.n6319 292.5
R25237 DVSS.n6304 DVSS.n6303 292.5
R25238 DVSS.n6289 DVSS.n6288 292.5
R25239 DVSS.n6274 DVSS.n6273 292.5
R25240 DVSS.n6259 DVSS.n6258 292.5
R25241 DVSS.n6244 DVSS.n6243 292.5
R25242 DVSS.n6229 DVSS.n6228 292.5
R25243 DVSS.n6214 DVSS.n6213 292.5
R25244 DVSS.n6203 DVSS.n6201 292.5
R25245 DVSS.n6188 DVSS.n6186 292.5
R25246 DVSS.n6173 DVSS.n6171 292.5
R25247 DVSS.n6158 DVSS.n6156 292.5
R25248 DVSS.n6143 DVSS.n6141 292.5
R25249 DVSS.n6128 DVSS.n6126 292.5
R25250 DVSS.n6113 DVSS.n6111 292.5
R25251 DVSS.n6098 DVSS.n6096 292.5
R25252 DVSS.n6095 DVSS.n6094 292.5
R25253 DVSS.n6072 DVSS.n6071 292.5
R25254 DVSS.n6070 DVSS.n6069 292.5
R25255 DVSS.n6054 DVSS.n6053 292.5
R25256 DVSS.n6027 DVSS.n6026 292.5
R25257 DVSS.n6025 DVSS.n6024 292.5
R25258 DVSS.n6022 DVSS.n6021 292.5
R25259 DVSS.n6020 DVSS.n6019 292.5
R25260 DVSS.n6039 DVSS.n6038 292.5
R25261 DVSS.n6031 DVSS.n6030 292.5
R25262 DVSS.n4932 DVSS.n4931 292.5
R25263 DVSS.n4934 DVSS.n4933 292.5
R25264 DVSS.n4937 DVSS.n4936 292.5
R25265 DVSS.n4943 DVSS.n4942 292.5
R25266 DVSS.n4929 DVSS.n4928 292.5
R25267 DVSS.n4910 DVSS.n4908 292.5
R25268 DVSS.n4895 DVSS.n4893 292.5
R25269 DVSS.n4880 DVSS.n4878 292.5
R25270 DVSS.n4877 DVSS.n4876 292.5
R25271 DVSS.n4854 DVSS.n4853 292.5
R25272 DVSS.n4852 DVSS.n4851 292.5
R25273 DVSS.n4836 DVSS.n4835 292.5
R25274 DVSS.n4821 DVSS.n4820 292.5
R25275 DVSS.n4806 DVSS.n4805 292.5
R25276 DVSS.n4791 DVSS.n4790 292.5
R25277 DVSS.n4776 DVSS.n4775 292.5
R25278 DVSS.n4761 DVSS.n4760 292.5
R25279 DVSS.n4746 DVSS.n4745 292.5
R25280 DVSS.n4735 DVSS.n4733 292.5
R25281 DVSS.n4720 DVSS.n4718 292.5
R25282 DVSS.n4705 DVSS.n4703 292.5
R25283 DVSS.n4690 DVSS.n4688 292.5
R25284 DVSS.n4675 DVSS.n4673 292.5
R25285 DVSS.n4660 DVSS.n4658 292.5
R25286 DVSS.n4645 DVSS.n4643 292.5
R25287 DVSS.n4630 DVSS.n4628 292.5
R25288 DVSS.n4627 DVSS.n4626 292.5
R25289 DVSS.n4604 DVSS.n4603 292.5
R25290 DVSS.n4602 DVSS.n4601 292.5
R25291 DVSS.n4586 DVSS.n4585 292.5
R25292 DVSS.n4559 DVSS.n4558 292.5
R25293 DVSS.n4557 DVSS.n4556 292.5
R25294 DVSS.n4554 DVSS.n4553 292.5
R25295 DVSS.n4552 DVSS.n4551 292.5
R25296 DVSS.n4571 DVSS.n4570 292.5
R25297 DVSS.n4563 DVSS.n4562 292.5
R25298 DVSS.n2288 DVSS.n2195 292.5
R25299 DVSS.n2288 DVSS.n2287 292.5
R25300 DVSS.n2304 DVSS.n2303 292.5
R25301 DVSS.n2303 DVSS.n2165 292.5
R25302 DVSS.n2271 DVSS.n2270 292.5
R25303 DVSS.n2269 DVSS.n2258 292.5
R25304 DVSS.n2268 DVSS.n2267 292.5
R25305 DVSS.n2266 DVSS.n2265 292.5
R25306 DVSS.n2264 DVSS.n2263 292.5
R25307 DVSS.n2262 DVSS.n2261 292.5
R25308 DVSS.n2260 DVSS.n2259 292.5
R25309 DVSS.n2254 DVSS.n2253 292.5
R25310 DVSS.n2302 DVSS.n2187 292.5
R25311 DVSS.n2302 DVSS.n2301 292.5
R25312 DVSS.n2292 DVSS.n2188 292.5
R25313 DVSS.n2193 DVSS.n2188 292.5
R25314 DVSS.n2280 DVSS.n2279 292.5
R25315 DVSS.n2281 DVSS.n2280 292.5
R25316 DVSS.n2278 DVSS.n2198 292.5
R25317 DVSS.n2199 DVSS.n2198 292.5
R25318 DVSS.n2294 DVSS.n2293 292.5
R25319 DVSS.n2295 DVSS.n2294 292.5
R25320 DVSS.n2276 DVSS.n2275 292.5
R25321 DVSS.n2277 DVSS.n2252 292.5
R25322 DVSS.n2252 DVSS.n2251 292.5
R25323 DVSS.n2315 DVSS.n2305 292.5
R25324 DVSS.n2308 DVSS.n2305 292.5
R25325 DVSS.n2316 DVSS.n2185 292.5
R25326 DVSS.n2307 DVSS.n2185 292.5
R25327 DVSS.n2314 DVSS.n2313 292.5
R25328 DVSS.n2311 DVSS.n2306 292.5
R25329 DVSS.n2322 DVSS.n2321 292.5
R25330 DVSS.n2324 DVSS.n2323 292.5
R25331 DVSS.n2186 DVSS.n2167 292.5
R25332 DVSS.n2341 DVSS.n2167 292.5
R25333 DVSS.n2319 DVSS.n2318 292.5
R25334 DVSS.n2310 DVSS.n2308 292.5
R25335 DVSS.n2307 DVSS.n2184 292.5
R25336 DVSS.n2182 DVSS.n2181 292.5
R25337 DVSS.n2330 DVSS.n2329 292.5
R25338 DVSS.n2333 DVSS.n2332 292.5
R25339 DVSS.n2176 DVSS.n2175 292.5
R25340 DVSS.n2339 DVSS.n2338 292.5
R25341 DVSS.n2173 DVSS.n2164 292.5
R25342 DVSS.n2344 DVSS.n2343 292.5
R25343 DVSS.n2163 DVSS.n2161 292.5
R25344 DVSS.n2165 DVSS.n2163 292.5
R25345 DVSS.n2300 DVSS.n2299 292.5
R25346 DVSS.n2301 DVSS.n2300 292.5
R25347 DVSS.n2298 DVSS.n2189 292.5
R25348 DVSS.n2193 DVSS.n2189 292.5
R25349 DVSS.n2297 DVSS.n2296 292.5
R25350 DVSS.n2296 DVSS.n2295 292.5
R25351 DVSS.n2250 DVSS.n2249 292.5
R25352 DVSS.n2251 DVSS.n2250 292.5
R25353 DVSS.n2283 DVSS.n2282 292.5
R25354 DVSS.n2282 DVSS.n2281 292.5
R25355 DVSS.n2284 DVSS.n2201 292.5
R25356 DVSS.n2201 DVSS.n2199 292.5
R25357 DVSS.n2286 DVSS.n2285 292.5
R25358 DVSS.n2287 DVSS.n2286 292.5
R25359 DVSS.n2290 DVSS.n2194 292.5
R25360 DVSS.n2248 DVSS.n2247 292.5
R25361 DVSS.n2247 DVSS.n2191 292.5
R25362 DVSS.n2206 DVSS.n2204 292.5
R25363 DVSS.n2211 DVSS.n2204 292.5
R25364 DVSS.n2242 DVSS.n2208 292.5
R25365 DVSS.n2242 DVSS.n2241 292.5
R25366 DVSS.n2216 DVSS.n2213 292.5
R25367 DVSS.n2240 DVSS.n2213 292.5
R25368 DVSS.n2237 DVSS.n2218 292.5
R25369 DVSS.n2238 DVSS.n2237 292.5
R25370 DVSS.n2223 DVSS.n2219 292.5
R25371 DVSS.n2219 DVSS.n2214 292.5
R25372 DVSS.n2232 DVSS.n2225 292.5
R25373 DVSS.n2232 DVSS.n2231 292.5
R25374 DVSS.n2230 DVSS.n2228 292.5
R25375 DVSS.n2228 DVSS.n2227 292.5
R25376 DVSS.n2290 DVSS.n2289 292.5
R25377 DVSS.n2102 DVSS.n2101 292.5
R25378 DVSS.n2093 DVSS.n2092 292.5
R25379 DVSS.n2105 DVSS.n2104 292.5
R25380 DVSS.n2107 DVSS.n2106 292.5
R25381 DVSS.n2109 DVSS.n2108 292.5
R25382 DVSS.n2111 DVSS.n2110 292.5
R25383 DVSS.n2113 DVSS.n2112 292.5
R25384 DVSS.n2103 DVSS.n2100 292.5
R25385 DVSS.n2117 DVSS.n2116 292.5
R25386 DVSS.n2116 DVSS.n2115 292.5
R25387 DVSS.n2409 DVSS.n2029 292.5
R25388 DVSS.n2409 DVSS.n2034 292.5
R25389 DVSS.n2422 DVSS.n2405 292.5
R25390 DVSS.n2421 DVSS.n2420 292.5
R25391 DVSS.n2419 DVSS.n2418 292.5
R25392 DVSS.n2417 DVSS.n2407 292.5
R25393 DVSS.n2415 DVSS.n2414 292.5
R25394 DVSS.n2413 DVSS.n2408 292.5
R25395 DVSS.n2412 DVSS.n2411 292.5
R25396 DVSS.n2425 DVSS.n2424 292.5
R25397 DVSS.n2065 DVSS.n2061 292.5
R25398 DVSS.n2078 DVSS.n2057 292.5
R25399 DVSS.n2076 DVSS.n2075 292.5
R25400 DVSS.n2074 DVSS.n2073 292.5
R25401 DVSS.n2071 DVSS.n2059 292.5
R25402 DVSS.n2069 DVSS.n2068 292.5
R25403 DVSS.n2067 DVSS.n2066 292.5
R25404 DVSS.n2080 DVSS.n2079 292.5
R25405 DVSS.n2079 DVSS.n2050 292.5
R25406 DVSS.n2063 DVSS.n2062 292.5
R25407 DVSS.n2459 DVSS.n2458 292.5
R25408 DVSS.n2458 DVSS.n2019 292.5
R25409 DVSS.n2460 DVSS.n2028 292.5
R25410 DVSS.n2028 DVSS.n2027 292.5
R25411 DVSS.n2462 DVSS.n2461 292.5
R25412 DVSS.n2463 DVSS.n2462 292.5
R25413 DVSS.n2437 DVSS.n2026 292.5
R25414 DVSS.n2026 DVSS.n2025 292.5
R25415 DVSS.n2435 DVSS.n2434 292.5
R25416 DVSS.n2434 DVSS.n2433 292.5
R25417 DVSS.n2031 DVSS.n2030 292.5
R25418 DVSS.n2033 DVSS.n2031 292.5
R25419 DVSS.n2389 DVSS.n2047 292.5
R25420 DVSS.n2047 DVSS.n2045 292.5
R25421 DVSS.n2391 DVSS.n2390 292.5
R25422 DVSS.n2392 DVSS.n2391 292.5
R25423 DVSS.n2388 DVSS.n2046 292.5
R25424 DVSS.n2051 DVSS.n2046 292.5
R25425 DVSS.n2387 DVSS.n2386 292.5
R25426 DVSS.n2386 DVSS.n2385 292.5
R25427 DVSS.n2370 DVSS.n2369 292.5
R25428 DVSS.n2371 DVSS.n2370 292.5
R25429 DVSS.n2368 DVSS.n2084 292.5
R25430 DVSS.n2084 DVSS.n2083 292.5
R25431 DVSS.n2367 DVSS.n2366 292.5
R25432 DVSS.n2366 DVSS.n2365 292.5
R25433 DVSS.n2086 DVSS.n2085 292.5
R25434 DVSS.n2087 DVSS.n2086 292.5
R25435 DVSS.n2457 DVSS.n2438 292.5
R25436 DVSS.n2443 DVSS.n2439 292.5
R25437 DVSS.n2453 DVSS.n2452 292.5
R25438 DVSS.n2451 DVSS.n2442 292.5
R25439 DVSS.n2450 DVSS.n2449 292.5
R25440 DVSS.n2448 DVSS.n2447 292.5
R25441 DVSS.n2446 DVSS.n2445 292.5
R25442 DVSS.n2444 DVSS.n2016 292.5
R25443 DVSS.n2475 DVSS.n2474 292.5
R25444 DVSS.n2753 DVSS.n2660 292.5
R25445 DVSS.n2753 DVSS.n2752 292.5
R25446 DVSS.n2769 DVSS.n2768 292.5
R25447 DVSS.n2768 DVSS.n2630 292.5
R25448 DVSS.n2736 DVSS.n2735 292.5
R25449 DVSS.n2734 DVSS.n2723 292.5
R25450 DVSS.n2733 DVSS.n2732 292.5
R25451 DVSS.n2731 DVSS.n2730 292.5
R25452 DVSS.n2729 DVSS.n2728 292.5
R25453 DVSS.n2727 DVSS.n2726 292.5
R25454 DVSS.n2725 DVSS.n2724 292.5
R25455 DVSS.n2719 DVSS.n2718 292.5
R25456 DVSS.n2767 DVSS.n2652 292.5
R25457 DVSS.n2767 DVSS.n2766 292.5
R25458 DVSS.n2757 DVSS.n2653 292.5
R25459 DVSS.n2658 DVSS.n2653 292.5
R25460 DVSS.n2745 DVSS.n2744 292.5
R25461 DVSS.n2746 DVSS.n2745 292.5
R25462 DVSS.n2743 DVSS.n2663 292.5
R25463 DVSS.n2664 DVSS.n2663 292.5
R25464 DVSS.n2759 DVSS.n2758 292.5
R25465 DVSS.n2760 DVSS.n2759 292.5
R25466 DVSS.n2741 DVSS.n2740 292.5
R25467 DVSS.n2742 DVSS.n2717 292.5
R25468 DVSS.n2717 DVSS.n2716 292.5
R25469 DVSS.n2780 DVSS.n2770 292.5
R25470 DVSS.n2773 DVSS.n2770 292.5
R25471 DVSS.n2781 DVSS.n2650 292.5
R25472 DVSS.n2772 DVSS.n2650 292.5
R25473 DVSS.n2779 DVSS.n2778 292.5
R25474 DVSS.n2776 DVSS.n2771 292.5
R25475 DVSS.n2787 DVSS.n2786 292.5
R25476 DVSS.n2789 DVSS.n2788 292.5
R25477 DVSS.n2651 DVSS.n2632 292.5
R25478 DVSS.n2806 DVSS.n2632 292.5
R25479 DVSS.n2784 DVSS.n2783 292.5
R25480 DVSS.n2775 DVSS.n2773 292.5
R25481 DVSS.n2772 DVSS.n2649 292.5
R25482 DVSS.n2647 DVSS.n2646 292.5
R25483 DVSS.n2795 DVSS.n2794 292.5
R25484 DVSS.n2798 DVSS.n2797 292.5
R25485 DVSS.n2641 DVSS.n2640 292.5
R25486 DVSS.n2804 DVSS.n2803 292.5
R25487 DVSS.n2638 DVSS.n2629 292.5
R25488 DVSS.n2809 DVSS.n2808 292.5
R25489 DVSS.n2628 DVSS.n2626 292.5
R25490 DVSS.n2630 DVSS.n2628 292.5
R25491 DVSS.n2765 DVSS.n2764 292.5
R25492 DVSS.n2766 DVSS.n2765 292.5
R25493 DVSS.n2763 DVSS.n2654 292.5
R25494 DVSS.n2658 DVSS.n2654 292.5
R25495 DVSS.n2762 DVSS.n2761 292.5
R25496 DVSS.n2761 DVSS.n2760 292.5
R25497 DVSS.n2715 DVSS.n2714 292.5
R25498 DVSS.n2716 DVSS.n2715 292.5
R25499 DVSS.n2748 DVSS.n2747 292.5
R25500 DVSS.n2747 DVSS.n2746 292.5
R25501 DVSS.n2749 DVSS.n2666 292.5
R25502 DVSS.n2666 DVSS.n2664 292.5
R25503 DVSS.n2751 DVSS.n2750 292.5
R25504 DVSS.n2752 DVSS.n2751 292.5
R25505 DVSS.n2755 DVSS.n2659 292.5
R25506 DVSS.n2713 DVSS.n2712 292.5
R25507 DVSS.n2712 DVSS.n2656 292.5
R25508 DVSS.n2671 DVSS.n2669 292.5
R25509 DVSS.n2676 DVSS.n2669 292.5
R25510 DVSS.n2707 DVSS.n2673 292.5
R25511 DVSS.n2707 DVSS.n2706 292.5
R25512 DVSS.n2681 DVSS.n2678 292.5
R25513 DVSS.n2705 DVSS.n2678 292.5
R25514 DVSS.n2702 DVSS.n2683 292.5
R25515 DVSS.n2703 DVSS.n2702 292.5
R25516 DVSS.n2688 DVSS.n2684 292.5
R25517 DVSS.n2684 DVSS.n2679 292.5
R25518 DVSS.n2697 DVSS.n2690 292.5
R25519 DVSS.n2697 DVSS.n2696 292.5
R25520 DVSS.n2695 DVSS.n2693 292.5
R25521 DVSS.n2693 DVSS.n2692 292.5
R25522 DVSS.n2755 DVSS.n2754 292.5
R25523 DVSS.n2567 DVSS.n2566 292.5
R25524 DVSS.n2558 DVSS.n2557 292.5
R25525 DVSS.n2570 DVSS.n2569 292.5
R25526 DVSS.n2572 DVSS.n2571 292.5
R25527 DVSS.n2574 DVSS.n2573 292.5
R25528 DVSS.n2576 DVSS.n2575 292.5
R25529 DVSS.n2578 DVSS.n2577 292.5
R25530 DVSS.n2568 DVSS.n2565 292.5
R25531 DVSS.n2582 DVSS.n2581 292.5
R25532 DVSS.n2581 DVSS.n2580 292.5
R25533 DVSS.n2874 DVSS.n2494 292.5
R25534 DVSS.n2874 DVSS.n2499 292.5
R25535 DVSS.n2887 DVSS.n2870 292.5
R25536 DVSS.n2886 DVSS.n2885 292.5
R25537 DVSS.n2884 DVSS.n2883 292.5
R25538 DVSS.n2882 DVSS.n2872 292.5
R25539 DVSS.n2880 DVSS.n2879 292.5
R25540 DVSS.n2878 DVSS.n2873 292.5
R25541 DVSS.n2877 DVSS.n2876 292.5
R25542 DVSS.n2890 DVSS.n2889 292.5
R25543 DVSS.n2530 DVSS.n2526 292.5
R25544 DVSS.n2543 DVSS.n2522 292.5
R25545 DVSS.n2541 DVSS.n2540 292.5
R25546 DVSS.n2539 DVSS.n2538 292.5
R25547 DVSS.n2536 DVSS.n2524 292.5
R25548 DVSS.n2534 DVSS.n2533 292.5
R25549 DVSS.n2532 DVSS.n2531 292.5
R25550 DVSS.n2545 DVSS.n2544 292.5
R25551 DVSS.n2544 DVSS.n2515 292.5
R25552 DVSS.n2528 DVSS.n2527 292.5
R25553 DVSS.n2924 DVSS.n2923 292.5
R25554 DVSS.n2923 DVSS.n2484 292.5
R25555 DVSS.n2925 DVSS.n2493 292.5
R25556 DVSS.n2493 DVSS.n2492 292.5
R25557 DVSS.n2927 DVSS.n2926 292.5
R25558 DVSS.n2928 DVSS.n2927 292.5
R25559 DVSS.n2902 DVSS.n2491 292.5
R25560 DVSS.n2491 DVSS.n2490 292.5
R25561 DVSS.n2900 DVSS.n2899 292.5
R25562 DVSS.n2899 DVSS.n2898 292.5
R25563 DVSS.n2496 DVSS.n2495 292.5
R25564 DVSS.n2498 DVSS.n2496 292.5
R25565 DVSS.n2854 DVSS.n2512 292.5
R25566 DVSS.n2512 DVSS.n2510 292.5
R25567 DVSS.n2856 DVSS.n2855 292.5
R25568 DVSS.n2857 DVSS.n2856 292.5
R25569 DVSS.n2853 DVSS.n2511 292.5
R25570 DVSS.n2516 DVSS.n2511 292.5
R25571 DVSS.n2852 DVSS.n2851 292.5
R25572 DVSS.n2851 DVSS.n2850 292.5
R25573 DVSS.n2835 DVSS.n2834 292.5
R25574 DVSS.n2836 DVSS.n2835 292.5
R25575 DVSS.n2833 DVSS.n2549 292.5
R25576 DVSS.n2549 DVSS.n2548 292.5
R25577 DVSS.n2832 DVSS.n2831 292.5
R25578 DVSS.n2831 DVSS.n2830 292.5
R25579 DVSS.n2551 DVSS.n2550 292.5
R25580 DVSS.n2552 DVSS.n2551 292.5
R25581 DVSS.n2922 DVSS.n2903 292.5
R25582 DVSS.n2908 DVSS.n2904 292.5
R25583 DVSS.n2918 DVSS.n2917 292.5
R25584 DVSS.n2916 DVSS.n2907 292.5
R25585 DVSS.n2915 DVSS.n2914 292.5
R25586 DVSS.n2913 DVSS.n2912 292.5
R25587 DVSS.n2911 DVSS.n2910 292.5
R25588 DVSS.n2909 DVSS.n2481 292.5
R25589 DVSS.n2939 DVSS.n2938 292.5
R25590 DVSS.n3336 DVSS.n3335 292.5
R25591 DVSS.n3338 DVSS.n3337 292.5
R25592 DVSS.n3341 DVSS.n3340 292.5
R25593 DVSS.n3348 DVSS.n3347 292.5
R25594 DVSS.n3333 DVSS.n3332 292.5
R25595 DVSS.n3314 DVSS.n3312 292.5
R25596 DVSS.n3299 DVSS.n3297 292.5
R25597 DVSS.n3284 DVSS.n3282 292.5
R25598 DVSS.n3281 DVSS.n3280 292.5
R25599 DVSS.n3258 DVSS.n3257 292.5
R25600 DVSS.n3256 DVSS.n3255 292.5
R25601 DVSS.n3240 DVSS.n3239 292.5
R25602 DVSS.n3225 DVSS.n3224 292.5
R25603 DVSS.n3210 DVSS.n3209 292.5
R25604 DVSS.n3195 DVSS.n3194 292.5
R25605 DVSS.n3180 DVSS.n3179 292.5
R25606 DVSS.n3165 DVSS.n3164 292.5
R25607 DVSS.n3150 DVSS.n3149 292.5
R25608 DVSS.n3139 DVSS.n3137 292.5
R25609 DVSS.n3124 DVSS.n3122 292.5
R25610 DVSS.n3109 DVSS.n3107 292.5
R25611 DVSS.n3094 DVSS.n3092 292.5
R25612 DVSS.n3079 DVSS.n3077 292.5
R25613 DVSS.n3064 DVSS.n3062 292.5
R25614 DVSS.n3049 DVSS.n3047 292.5
R25615 DVSS.n3034 DVSS.n3032 292.5
R25616 DVSS.n3031 DVSS.n3030 292.5
R25617 DVSS.n3008 DVSS.n3007 292.5
R25618 DVSS.n3006 DVSS.n3005 292.5
R25619 DVSS.n2990 DVSS.n2989 292.5
R25620 DVSS.n2963 DVSS.n2962 292.5
R25621 DVSS.n2961 DVSS.n2960 292.5
R25622 DVSS.n2958 DVSS.n2957 292.5
R25623 DVSS.n2956 DVSS.n2955 292.5
R25624 DVSS.n2975 DVSS.n2974 292.5
R25625 DVSS.n2967 DVSS.n2966 292.5
R25626 DVSS.n5352 DVSS.n5259 292.5
R25627 DVSS.n5352 DVSS.n5351 292.5
R25628 DVSS.n5368 DVSS.n5367 292.5
R25629 DVSS.n5367 DVSS.n5229 292.5
R25630 DVSS.n5335 DVSS.n5334 292.5
R25631 DVSS.n5333 DVSS.n5322 292.5
R25632 DVSS.n5332 DVSS.n5331 292.5
R25633 DVSS.n5330 DVSS.n5329 292.5
R25634 DVSS.n5328 DVSS.n5327 292.5
R25635 DVSS.n5326 DVSS.n5325 292.5
R25636 DVSS.n5324 DVSS.n5323 292.5
R25637 DVSS.n5318 DVSS.n5317 292.5
R25638 DVSS.n5366 DVSS.n5251 292.5
R25639 DVSS.n5366 DVSS.n5365 292.5
R25640 DVSS.n5356 DVSS.n5252 292.5
R25641 DVSS.n5257 DVSS.n5252 292.5
R25642 DVSS.n5344 DVSS.n5343 292.5
R25643 DVSS.n5345 DVSS.n5344 292.5
R25644 DVSS.n5342 DVSS.n5262 292.5
R25645 DVSS.n5263 DVSS.n5262 292.5
R25646 DVSS.n5358 DVSS.n5357 292.5
R25647 DVSS.n5359 DVSS.n5358 292.5
R25648 DVSS.n5340 DVSS.n5339 292.5
R25649 DVSS.n5341 DVSS.n5316 292.5
R25650 DVSS.n5316 DVSS.n5315 292.5
R25651 DVSS.n5379 DVSS.n5369 292.5
R25652 DVSS.n5372 DVSS.n5369 292.5
R25653 DVSS.n5380 DVSS.n5249 292.5
R25654 DVSS.n5371 DVSS.n5249 292.5
R25655 DVSS.n5378 DVSS.n5377 292.5
R25656 DVSS.n5375 DVSS.n5370 292.5
R25657 DVSS.n5386 DVSS.n5385 292.5
R25658 DVSS.n5388 DVSS.n5387 292.5
R25659 DVSS.n5250 DVSS.n5231 292.5
R25660 DVSS.n5405 DVSS.n5231 292.5
R25661 DVSS.n5383 DVSS.n5382 292.5
R25662 DVSS.n5374 DVSS.n5372 292.5
R25663 DVSS.n5371 DVSS.n5248 292.5
R25664 DVSS.n5246 DVSS.n5245 292.5
R25665 DVSS.n5394 DVSS.n5393 292.5
R25666 DVSS.n5397 DVSS.n5396 292.5
R25667 DVSS.n5240 DVSS.n5239 292.5
R25668 DVSS.n5403 DVSS.n5402 292.5
R25669 DVSS.n5237 DVSS.n5228 292.5
R25670 DVSS.n5408 DVSS.n5407 292.5
R25671 DVSS.n5227 DVSS.n5225 292.5
R25672 DVSS.n5229 DVSS.n5227 292.5
R25673 DVSS.n5364 DVSS.n5363 292.5
R25674 DVSS.n5365 DVSS.n5364 292.5
R25675 DVSS.n5362 DVSS.n5253 292.5
R25676 DVSS.n5257 DVSS.n5253 292.5
R25677 DVSS.n5361 DVSS.n5360 292.5
R25678 DVSS.n5360 DVSS.n5359 292.5
R25679 DVSS.n5314 DVSS.n5313 292.5
R25680 DVSS.n5315 DVSS.n5314 292.5
R25681 DVSS.n5347 DVSS.n5346 292.5
R25682 DVSS.n5346 DVSS.n5345 292.5
R25683 DVSS.n5348 DVSS.n5265 292.5
R25684 DVSS.n5265 DVSS.n5263 292.5
R25685 DVSS.n5350 DVSS.n5349 292.5
R25686 DVSS.n5351 DVSS.n5350 292.5
R25687 DVSS.n5354 DVSS.n5258 292.5
R25688 DVSS.n5312 DVSS.n5311 292.5
R25689 DVSS.n5311 DVSS.n5255 292.5
R25690 DVSS.n5270 DVSS.n5268 292.5
R25691 DVSS.n5275 DVSS.n5268 292.5
R25692 DVSS.n5306 DVSS.n5272 292.5
R25693 DVSS.n5306 DVSS.n5305 292.5
R25694 DVSS.n5280 DVSS.n5277 292.5
R25695 DVSS.n5304 DVSS.n5277 292.5
R25696 DVSS.n5301 DVSS.n5282 292.5
R25697 DVSS.n5302 DVSS.n5301 292.5
R25698 DVSS.n5287 DVSS.n5283 292.5
R25699 DVSS.n5283 DVSS.n5278 292.5
R25700 DVSS.n5296 DVSS.n5289 292.5
R25701 DVSS.n5296 DVSS.n5295 292.5
R25702 DVSS.n5294 DVSS.n5292 292.5
R25703 DVSS.n5292 DVSS.n5291 292.5
R25704 DVSS.n5354 DVSS.n5353 292.5
R25705 DVSS.n5166 DVSS.n5165 292.5
R25706 DVSS.n5157 DVSS.n5156 292.5
R25707 DVSS.n5169 DVSS.n5168 292.5
R25708 DVSS.n5171 DVSS.n5170 292.5
R25709 DVSS.n5173 DVSS.n5172 292.5
R25710 DVSS.n5175 DVSS.n5174 292.5
R25711 DVSS.n5177 DVSS.n5176 292.5
R25712 DVSS.n5167 DVSS.n5164 292.5
R25713 DVSS.n5181 DVSS.n5180 292.5
R25714 DVSS.n5180 DVSS.n5179 292.5
R25715 DVSS.n5473 DVSS.n5093 292.5
R25716 DVSS.n5473 DVSS.n5098 292.5
R25717 DVSS.n5486 DVSS.n5469 292.5
R25718 DVSS.n5485 DVSS.n5484 292.5
R25719 DVSS.n5483 DVSS.n5482 292.5
R25720 DVSS.n5481 DVSS.n5471 292.5
R25721 DVSS.n5479 DVSS.n5478 292.5
R25722 DVSS.n5477 DVSS.n5472 292.5
R25723 DVSS.n5476 DVSS.n5475 292.5
R25724 DVSS.n5489 DVSS.n5488 292.5
R25725 DVSS.n5129 DVSS.n5125 292.5
R25726 DVSS.n5142 DVSS.n5121 292.5
R25727 DVSS.n5140 DVSS.n5139 292.5
R25728 DVSS.n5138 DVSS.n5137 292.5
R25729 DVSS.n5135 DVSS.n5123 292.5
R25730 DVSS.n5133 DVSS.n5132 292.5
R25731 DVSS.n5131 DVSS.n5130 292.5
R25732 DVSS.n5144 DVSS.n5143 292.5
R25733 DVSS.n5143 DVSS.n5114 292.5
R25734 DVSS.n5127 DVSS.n5126 292.5
R25735 DVSS.n5523 DVSS.n5522 292.5
R25736 DVSS.n5522 DVSS.n5083 292.5
R25737 DVSS.n5524 DVSS.n5092 292.5
R25738 DVSS.n5092 DVSS.n5091 292.5
R25739 DVSS.n5526 DVSS.n5525 292.5
R25740 DVSS.n5527 DVSS.n5526 292.5
R25741 DVSS.n5501 DVSS.n5090 292.5
R25742 DVSS.n5090 DVSS.n5089 292.5
R25743 DVSS.n5499 DVSS.n5498 292.5
R25744 DVSS.n5498 DVSS.n5497 292.5
R25745 DVSS.n5095 DVSS.n5094 292.5
R25746 DVSS.n5097 DVSS.n5095 292.5
R25747 DVSS.n5453 DVSS.n5111 292.5
R25748 DVSS.n5111 DVSS.n5109 292.5
R25749 DVSS.n5455 DVSS.n5454 292.5
R25750 DVSS.n5456 DVSS.n5455 292.5
R25751 DVSS.n5452 DVSS.n5110 292.5
R25752 DVSS.n5115 DVSS.n5110 292.5
R25753 DVSS.n5451 DVSS.n5450 292.5
R25754 DVSS.n5450 DVSS.n5449 292.5
R25755 DVSS.n5434 DVSS.n5433 292.5
R25756 DVSS.n5435 DVSS.n5434 292.5
R25757 DVSS.n5432 DVSS.n5148 292.5
R25758 DVSS.n5148 DVSS.n5147 292.5
R25759 DVSS.n5431 DVSS.n5430 292.5
R25760 DVSS.n5430 DVSS.n5429 292.5
R25761 DVSS.n5150 DVSS.n5149 292.5
R25762 DVSS.n5151 DVSS.n5150 292.5
R25763 DVSS.n5521 DVSS.n5502 292.5
R25764 DVSS.n5507 DVSS.n5503 292.5
R25765 DVSS.n5517 DVSS.n5516 292.5
R25766 DVSS.n5515 DVSS.n5506 292.5
R25767 DVSS.n5514 DVSS.n5513 292.5
R25768 DVSS.n5512 DVSS.n5511 292.5
R25769 DVSS.n5510 DVSS.n5509 292.5
R25770 DVSS.n5508 DVSS.n5080 292.5
R25771 DVSS.n5539 DVSS.n5538 292.5
R25772 DVSS.n5817 DVSS.n5724 292.5
R25773 DVSS.n5817 DVSS.n5816 292.5
R25774 DVSS.n5833 DVSS.n5832 292.5
R25775 DVSS.n5832 DVSS.n5694 292.5
R25776 DVSS.n5800 DVSS.n5799 292.5
R25777 DVSS.n5798 DVSS.n5787 292.5
R25778 DVSS.n5797 DVSS.n5796 292.5
R25779 DVSS.n5795 DVSS.n5794 292.5
R25780 DVSS.n5793 DVSS.n5792 292.5
R25781 DVSS.n5791 DVSS.n5790 292.5
R25782 DVSS.n5789 DVSS.n5788 292.5
R25783 DVSS.n5783 DVSS.n5782 292.5
R25784 DVSS.n5831 DVSS.n5716 292.5
R25785 DVSS.n5831 DVSS.n5830 292.5
R25786 DVSS.n5821 DVSS.n5717 292.5
R25787 DVSS.n5722 DVSS.n5717 292.5
R25788 DVSS.n5809 DVSS.n5808 292.5
R25789 DVSS.n5810 DVSS.n5809 292.5
R25790 DVSS.n5807 DVSS.n5727 292.5
R25791 DVSS.n5728 DVSS.n5727 292.5
R25792 DVSS.n5823 DVSS.n5822 292.5
R25793 DVSS.n5824 DVSS.n5823 292.5
R25794 DVSS.n5805 DVSS.n5804 292.5
R25795 DVSS.n5806 DVSS.n5781 292.5
R25796 DVSS.n5781 DVSS.n5780 292.5
R25797 DVSS.n5844 DVSS.n5834 292.5
R25798 DVSS.n5837 DVSS.n5834 292.5
R25799 DVSS.n5845 DVSS.n5714 292.5
R25800 DVSS.n5836 DVSS.n5714 292.5
R25801 DVSS.n5843 DVSS.n5842 292.5
R25802 DVSS.n5840 DVSS.n5835 292.5
R25803 DVSS.n5851 DVSS.n5850 292.5
R25804 DVSS.n5853 DVSS.n5852 292.5
R25805 DVSS.n5715 DVSS.n5696 292.5
R25806 DVSS.n5870 DVSS.n5696 292.5
R25807 DVSS.n5848 DVSS.n5847 292.5
R25808 DVSS.n5839 DVSS.n5837 292.5
R25809 DVSS.n5836 DVSS.n5713 292.5
R25810 DVSS.n5711 DVSS.n5710 292.5
R25811 DVSS.n5859 DVSS.n5858 292.5
R25812 DVSS.n5862 DVSS.n5861 292.5
R25813 DVSS.n5705 DVSS.n5704 292.5
R25814 DVSS.n5868 DVSS.n5867 292.5
R25815 DVSS.n5702 DVSS.n5693 292.5
R25816 DVSS.n5873 DVSS.n5872 292.5
R25817 DVSS.n5692 DVSS.n5690 292.5
R25818 DVSS.n5694 DVSS.n5692 292.5
R25819 DVSS.n5829 DVSS.n5828 292.5
R25820 DVSS.n5830 DVSS.n5829 292.5
R25821 DVSS.n5827 DVSS.n5718 292.5
R25822 DVSS.n5722 DVSS.n5718 292.5
R25823 DVSS.n5826 DVSS.n5825 292.5
R25824 DVSS.n5825 DVSS.n5824 292.5
R25825 DVSS.n5779 DVSS.n5778 292.5
R25826 DVSS.n5780 DVSS.n5779 292.5
R25827 DVSS.n5812 DVSS.n5811 292.5
R25828 DVSS.n5811 DVSS.n5810 292.5
R25829 DVSS.n5813 DVSS.n5730 292.5
R25830 DVSS.n5730 DVSS.n5728 292.5
R25831 DVSS.n5815 DVSS.n5814 292.5
R25832 DVSS.n5816 DVSS.n5815 292.5
R25833 DVSS.n5819 DVSS.n5723 292.5
R25834 DVSS.n5777 DVSS.n5776 292.5
R25835 DVSS.n5776 DVSS.n5720 292.5
R25836 DVSS.n5735 DVSS.n5733 292.5
R25837 DVSS.n5740 DVSS.n5733 292.5
R25838 DVSS.n5771 DVSS.n5737 292.5
R25839 DVSS.n5771 DVSS.n5770 292.5
R25840 DVSS.n5745 DVSS.n5742 292.5
R25841 DVSS.n5769 DVSS.n5742 292.5
R25842 DVSS.n5766 DVSS.n5747 292.5
R25843 DVSS.n5767 DVSS.n5766 292.5
R25844 DVSS.n5752 DVSS.n5748 292.5
R25845 DVSS.n5748 DVSS.n5743 292.5
R25846 DVSS.n5761 DVSS.n5754 292.5
R25847 DVSS.n5761 DVSS.n5760 292.5
R25848 DVSS.n5759 DVSS.n5757 292.5
R25849 DVSS.n5757 DVSS.n5756 292.5
R25850 DVSS.n5819 DVSS.n5818 292.5
R25851 DVSS.n5631 DVSS.n5630 292.5
R25852 DVSS.n5622 DVSS.n5621 292.5
R25853 DVSS.n5634 DVSS.n5633 292.5
R25854 DVSS.n5636 DVSS.n5635 292.5
R25855 DVSS.n5638 DVSS.n5637 292.5
R25856 DVSS.n5640 DVSS.n5639 292.5
R25857 DVSS.n5642 DVSS.n5641 292.5
R25858 DVSS.n5632 DVSS.n5629 292.5
R25859 DVSS.n5646 DVSS.n5645 292.5
R25860 DVSS.n5645 DVSS.n5644 292.5
R25861 DVSS.n5938 DVSS.n5558 292.5
R25862 DVSS.n5938 DVSS.n5563 292.5
R25863 DVSS.n5951 DVSS.n5934 292.5
R25864 DVSS.n5950 DVSS.n5949 292.5
R25865 DVSS.n5948 DVSS.n5947 292.5
R25866 DVSS.n5946 DVSS.n5936 292.5
R25867 DVSS.n5944 DVSS.n5943 292.5
R25868 DVSS.n5942 DVSS.n5937 292.5
R25869 DVSS.n5941 DVSS.n5940 292.5
R25870 DVSS.n5954 DVSS.n5953 292.5
R25871 DVSS.n5594 DVSS.n5590 292.5
R25872 DVSS.n5607 DVSS.n5586 292.5
R25873 DVSS.n5605 DVSS.n5604 292.5
R25874 DVSS.n5603 DVSS.n5602 292.5
R25875 DVSS.n5600 DVSS.n5588 292.5
R25876 DVSS.n5598 DVSS.n5597 292.5
R25877 DVSS.n5596 DVSS.n5595 292.5
R25878 DVSS.n5609 DVSS.n5608 292.5
R25879 DVSS.n5608 DVSS.n5579 292.5
R25880 DVSS.n5592 DVSS.n5591 292.5
R25881 DVSS.n5988 DVSS.n5987 292.5
R25882 DVSS.n5987 DVSS.n5548 292.5
R25883 DVSS.n5989 DVSS.n5557 292.5
R25884 DVSS.n5557 DVSS.n5556 292.5
R25885 DVSS.n5991 DVSS.n5990 292.5
R25886 DVSS.n5992 DVSS.n5991 292.5
R25887 DVSS.n5966 DVSS.n5555 292.5
R25888 DVSS.n5555 DVSS.n5554 292.5
R25889 DVSS.n5964 DVSS.n5963 292.5
R25890 DVSS.n5963 DVSS.n5962 292.5
R25891 DVSS.n5560 DVSS.n5559 292.5
R25892 DVSS.n5562 DVSS.n5560 292.5
R25893 DVSS.n5918 DVSS.n5576 292.5
R25894 DVSS.n5576 DVSS.n5574 292.5
R25895 DVSS.n5920 DVSS.n5919 292.5
R25896 DVSS.n5921 DVSS.n5920 292.5
R25897 DVSS.n5917 DVSS.n5575 292.5
R25898 DVSS.n5580 DVSS.n5575 292.5
R25899 DVSS.n5916 DVSS.n5915 292.5
R25900 DVSS.n5915 DVSS.n5914 292.5
R25901 DVSS.n5899 DVSS.n5898 292.5
R25902 DVSS.n5900 DVSS.n5899 292.5
R25903 DVSS.n5897 DVSS.n5613 292.5
R25904 DVSS.n5613 DVSS.n5612 292.5
R25905 DVSS.n5896 DVSS.n5895 292.5
R25906 DVSS.n5895 DVSS.n5894 292.5
R25907 DVSS.n5615 DVSS.n5614 292.5
R25908 DVSS.n5616 DVSS.n5615 292.5
R25909 DVSS.n5986 DVSS.n5967 292.5
R25910 DVSS.n5972 DVSS.n5968 292.5
R25911 DVSS.n5982 DVSS.n5981 292.5
R25912 DVSS.n5980 DVSS.n5971 292.5
R25913 DVSS.n5979 DVSS.n5978 292.5
R25914 DVSS.n5977 DVSS.n5976 292.5
R25915 DVSS.n5975 DVSS.n5974 292.5
R25916 DVSS.n5973 DVSS.n5545 292.5
R25917 DVSS.n6003 DVSS.n6002 292.5
R25918 DVSS.n287 DVSS.n194 292.5
R25919 DVSS.n287 DVSS.n286 292.5
R25920 DVSS.n303 DVSS.n302 292.5
R25921 DVSS.n302 DVSS.n164 292.5
R25922 DVSS.n270 DVSS.n269 292.5
R25923 DVSS.n268 DVSS.n257 292.5
R25924 DVSS.n267 DVSS.n266 292.5
R25925 DVSS.n265 DVSS.n264 292.5
R25926 DVSS.n263 DVSS.n262 292.5
R25927 DVSS.n261 DVSS.n260 292.5
R25928 DVSS.n259 DVSS.n258 292.5
R25929 DVSS.n253 DVSS.n252 292.5
R25930 DVSS.n301 DVSS.n186 292.5
R25931 DVSS.n301 DVSS.n300 292.5
R25932 DVSS.n291 DVSS.n187 292.5
R25933 DVSS.n192 DVSS.n187 292.5
R25934 DVSS.n279 DVSS.n278 292.5
R25935 DVSS.n280 DVSS.n279 292.5
R25936 DVSS.n277 DVSS.n197 292.5
R25937 DVSS.n198 DVSS.n197 292.5
R25938 DVSS.n293 DVSS.n292 292.5
R25939 DVSS.n294 DVSS.n293 292.5
R25940 DVSS.n275 DVSS.n274 292.5
R25941 DVSS.n276 DVSS.n251 292.5
R25942 DVSS.n251 DVSS.n250 292.5
R25943 DVSS.n314 DVSS.n304 292.5
R25944 DVSS.n307 DVSS.n304 292.5
R25945 DVSS.n315 DVSS.n184 292.5
R25946 DVSS.n306 DVSS.n184 292.5
R25947 DVSS.n313 DVSS.n312 292.5
R25948 DVSS.n310 DVSS.n305 292.5
R25949 DVSS.n321 DVSS.n320 292.5
R25950 DVSS.n323 DVSS.n322 292.5
R25951 DVSS.n185 DVSS.n166 292.5
R25952 DVSS.n340 DVSS.n166 292.5
R25953 DVSS.n318 DVSS.n317 292.5
R25954 DVSS.n309 DVSS.n307 292.5
R25955 DVSS.n306 DVSS.n183 292.5
R25956 DVSS.n181 DVSS.n180 292.5
R25957 DVSS.n329 DVSS.n328 292.5
R25958 DVSS.n332 DVSS.n331 292.5
R25959 DVSS.n175 DVSS.n174 292.5
R25960 DVSS.n338 DVSS.n337 292.5
R25961 DVSS.n172 DVSS.n163 292.5
R25962 DVSS.n343 DVSS.n342 292.5
R25963 DVSS.n162 DVSS.n160 292.5
R25964 DVSS.n164 DVSS.n162 292.5
R25965 DVSS.n299 DVSS.n298 292.5
R25966 DVSS.n300 DVSS.n299 292.5
R25967 DVSS.n297 DVSS.n188 292.5
R25968 DVSS.n192 DVSS.n188 292.5
R25969 DVSS.n296 DVSS.n295 292.5
R25970 DVSS.n295 DVSS.n294 292.5
R25971 DVSS.n249 DVSS.n248 292.5
R25972 DVSS.n250 DVSS.n249 292.5
R25973 DVSS.n282 DVSS.n281 292.5
R25974 DVSS.n281 DVSS.n280 292.5
R25975 DVSS.n283 DVSS.n200 292.5
R25976 DVSS.n200 DVSS.n198 292.5
R25977 DVSS.n285 DVSS.n284 292.5
R25978 DVSS.n286 DVSS.n285 292.5
R25979 DVSS.n289 DVSS.n193 292.5
R25980 DVSS.n247 DVSS.n246 292.5
R25981 DVSS.n246 DVSS.n190 292.5
R25982 DVSS.n205 DVSS.n203 292.5
R25983 DVSS.n210 DVSS.n203 292.5
R25984 DVSS.n241 DVSS.n207 292.5
R25985 DVSS.n241 DVSS.n240 292.5
R25986 DVSS.n215 DVSS.n212 292.5
R25987 DVSS.n239 DVSS.n212 292.5
R25988 DVSS.n236 DVSS.n217 292.5
R25989 DVSS.n237 DVSS.n236 292.5
R25990 DVSS.n222 DVSS.n218 292.5
R25991 DVSS.n218 DVSS.n213 292.5
R25992 DVSS.n231 DVSS.n224 292.5
R25993 DVSS.n231 DVSS.n230 292.5
R25994 DVSS.n229 DVSS.n227 292.5
R25995 DVSS.n227 DVSS.n226 292.5
R25996 DVSS.n289 DVSS.n288 292.5
R25997 DVSS.n101 DVSS.n100 292.5
R25998 DVSS.n92 DVSS.n91 292.5
R25999 DVSS.n104 DVSS.n103 292.5
R26000 DVSS.n106 DVSS.n105 292.5
R26001 DVSS.n108 DVSS.n107 292.5
R26002 DVSS.n110 DVSS.n109 292.5
R26003 DVSS.n112 DVSS.n111 292.5
R26004 DVSS.n102 DVSS.n99 292.5
R26005 DVSS.n116 DVSS.n115 292.5
R26006 DVSS.n115 DVSS.n114 292.5
R26007 DVSS.n408 DVSS.n28 292.5
R26008 DVSS.n408 DVSS.n33 292.5
R26009 DVSS.n421 DVSS.n404 292.5
R26010 DVSS.n420 DVSS.n419 292.5
R26011 DVSS.n418 DVSS.n417 292.5
R26012 DVSS.n416 DVSS.n406 292.5
R26013 DVSS.n414 DVSS.n413 292.5
R26014 DVSS.n412 DVSS.n407 292.5
R26015 DVSS.n411 DVSS.n410 292.5
R26016 DVSS.n424 DVSS.n423 292.5
R26017 DVSS.n64 DVSS.n60 292.5
R26018 DVSS.n77 DVSS.n56 292.5
R26019 DVSS.n75 DVSS.n74 292.5
R26020 DVSS.n73 DVSS.n72 292.5
R26021 DVSS.n70 DVSS.n58 292.5
R26022 DVSS.n68 DVSS.n67 292.5
R26023 DVSS.n66 DVSS.n65 292.5
R26024 DVSS.n79 DVSS.n78 292.5
R26025 DVSS.n78 DVSS.n49 292.5
R26026 DVSS.n62 DVSS.n61 292.5
R26027 DVSS.n458 DVSS.n457 292.5
R26028 DVSS.n457 DVSS.n18 292.5
R26029 DVSS.n459 DVSS.n27 292.5
R26030 DVSS.n27 DVSS.n26 292.5
R26031 DVSS.n461 DVSS.n460 292.5
R26032 DVSS.n462 DVSS.n461 292.5
R26033 DVSS.n436 DVSS.n25 292.5
R26034 DVSS.n25 DVSS.n24 292.5
R26035 DVSS.n434 DVSS.n433 292.5
R26036 DVSS.n433 DVSS.n432 292.5
R26037 DVSS.n30 DVSS.n29 292.5
R26038 DVSS.n32 DVSS.n30 292.5
R26039 DVSS.n388 DVSS.n46 292.5
R26040 DVSS.n46 DVSS.n44 292.5
R26041 DVSS.n390 DVSS.n389 292.5
R26042 DVSS.n391 DVSS.n390 292.5
R26043 DVSS.n387 DVSS.n45 292.5
R26044 DVSS.n50 DVSS.n45 292.5
R26045 DVSS.n386 DVSS.n385 292.5
R26046 DVSS.n385 DVSS.n384 292.5
R26047 DVSS.n369 DVSS.n368 292.5
R26048 DVSS.n370 DVSS.n369 292.5
R26049 DVSS.n367 DVSS.n83 292.5
R26050 DVSS.n83 DVSS.n82 292.5
R26051 DVSS.n366 DVSS.n365 292.5
R26052 DVSS.n365 DVSS.n364 292.5
R26053 DVSS.n85 DVSS.n84 292.5
R26054 DVSS.n86 DVSS.n85 292.5
R26055 DVSS.n456 DVSS.n437 292.5
R26056 DVSS.n442 DVSS.n438 292.5
R26057 DVSS.n452 DVSS.n451 292.5
R26058 DVSS.n450 DVSS.n441 292.5
R26059 DVSS.n449 DVSS.n448 292.5
R26060 DVSS.n447 DVSS.n446 292.5
R26061 DVSS.n445 DVSS.n444 292.5
R26062 DVSS.n443 DVSS.n15 292.5
R26063 DVSS.n474 DVSS.n473 292.5
R26064 DVSS.n752 DVSS.n659 292.5
R26065 DVSS.n752 DVSS.n751 292.5
R26066 DVSS.n768 DVSS.n767 292.5
R26067 DVSS.n767 DVSS.n629 292.5
R26068 DVSS.n735 DVSS.n734 292.5
R26069 DVSS.n733 DVSS.n722 292.5
R26070 DVSS.n732 DVSS.n731 292.5
R26071 DVSS.n730 DVSS.n729 292.5
R26072 DVSS.n728 DVSS.n727 292.5
R26073 DVSS.n726 DVSS.n725 292.5
R26074 DVSS.n724 DVSS.n723 292.5
R26075 DVSS.n718 DVSS.n717 292.5
R26076 DVSS.n766 DVSS.n651 292.5
R26077 DVSS.n766 DVSS.n765 292.5
R26078 DVSS.n756 DVSS.n652 292.5
R26079 DVSS.n657 DVSS.n652 292.5
R26080 DVSS.n744 DVSS.n743 292.5
R26081 DVSS.n745 DVSS.n744 292.5
R26082 DVSS.n742 DVSS.n662 292.5
R26083 DVSS.n663 DVSS.n662 292.5
R26084 DVSS.n758 DVSS.n757 292.5
R26085 DVSS.n759 DVSS.n758 292.5
R26086 DVSS.n740 DVSS.n739 292.5
R26087 DVSS.n741 DVSS.n716 292.5
R26088 DVSS.n716 DVSS.n715 292.5
R26089 DVSS.n779 DVSS.n769 292.5
R26090 DVSS.n772 DVSS.n769 292.5
R26091 DVSS.n780 DVSS.n649 292.5
R26092 DVSS.n771 DVSS.n649 292.5
R26093 DVSS.n778 DVSS.n777 292.5
R26094 DVSS.n775 DVSS.n770 292.5
R26095 DVSS.n786 DVSS.n785 292.5
R26096 DVSS.n788 DVSS.n787 292.5
R26097 DVSS.n650 DVSS.n631 292.5
R26098 DVSS.n805 DVSS.n631 292.5
R26099 DVSS.n783 DVSS.n782 292.5
R26100 DVSS.n774 DVSS.n772 292.5
R26101 DVSS.n771 DVSS.n648 292.5
R26102 DVSS.n646 DVSS.n645 292.5
R26103 DVSS.n794 DVSS.n793 292.5
R26104 DVSS.n797 DVSS.n796 292.5
R26105 DVSS.n640 DVSS.n639 292.5
R26106 DVSS.n803 DVSS.n802 292.5
R26107 DVSS.n637 DVSS.n628 292.5
R26108 DVSS.n808 DVSS.n807 292.5
R26109 DVSS.n627 DVSS.n625 292.5
R26110 DVSS.n629 DVSS.n627 292.5
R26111 DVSS.n764 DVSS.n763 292.5
R26112 DVSS.n765 DVSS.n764 292.5
R26113 DVSS.n762 DVSS.n653 292.5
R26114 DVSS.n657 DVSS.n653 292.5
R26115 DVSS.n761 DVSS.n760 292.5
R26116 DVSS.n760 DVSS.n759 292.5
R26117 DVSS.n714 DVSS.n713 292.5
R26118 DVSS.n715 DVSS.n714 292.5
R26119 DVSS.n747 DVSS.n746 292.5
R26120 DVSS.n746 DVSS.n745 292.5
R26121 DVSS.n748 DVSS.n665 292.5
R26122 DVSS.n665 DVSS.n663 292.5
R26123 DVSS.n750 DVSS.n749 292.5
R26124 DVSS.n751 DVSS.n750 292.5
R26125 DVSS.n754 DVSS.n658 292.5
R26126 DVSS.n712 DVSS.n711 292.5
R26127 DVSS.n711 DVSS.n655 292.5
R26128 DVSS.n670 DVSS.n668 292.5
R26129 DVSS.n675 DVSS.n668 292.5
R26130 DVSS.n706 DVSS.n672 292.5
R26131 DVSS.n706 DVSS.n705 292.5
R26132 DVSS.n680 DVSS.n677 292.5
R26133 DVSS.n704 DVSS.n677 292.5
R26134 DVSS.n701 DVSS.n682 292.5
R26135 DVSS.n702 DVSS.n701 292.5
R26136 DVSS.n687 DVSS.n683 292.5
R26137 DVSS.n683 DVSS.n678 292.5
R26138 DVSS.n696 DVSS.n689 292.5
R26139 DVSS.n696 DVSS.n695 292.5
R26140 DVSS.n694 DVSS.n692 292.5
R26141 DVSS.n692 DVSS.n691 292.5
R26142 DVSS.n754 DVSS.n753 292.5
R26143 DVSS.n566 DVSS.n565 292.5
R26144 DVSS.n557 DVSS.n556 292.5
R26145 DVSS.n569 DVSS.n568 292.5
R26146 DVSS.n571 DVSS.n570 292.5
R26147 DVSS.n573 DVSS.n572 292.5
R26148 DVSS.n575 DVSS.n574 292.5
R26149 DVSS.n577 DVSS.n576 292.5
R26150 DVSS.n567 DVSS.n564 292.5
R26151 DVSS.n581 DVSS.n580 292.5
R26152 DVSS.n580 DVSS.n579 292.5
R26153 DVSS.n873 DVSS.n493 292.5
R26154 DVSS.n873 DVSS.n498 292.5
R26155 DVSS.n886 DVSS.n869 292.5
R26156 DVSS.n885 DVSS.n884 292.5
R26157 DVSS.n883 DVSS.n882 292.5
R26158 DVSS.n881 DVSS.n871 292.5
R26159 DVSS.n879 DVSS.n878 292.5
R26160 DVSS.n877 DVSS.n872 292.5
R26161 DVSS.n876 DVSS.n875 292.5
R26162 DVSS.n889 DVSS.n888 292.5
R26163 DVSS.n529 DVSS.n525 292.5
R26164 DVSS.n542 DVSS.n521 292.5
R26165 DVSS.n540 DVSS.n539 292.5
R26166 DVSS.n538 DVSS.n537 292.5
R26167 DVSS.n535 DVSS.n523 292.5
R26168 DVSS.n533 DVSS.n532 292.5
R26169 DVSS.n531 DVSS.n530 292.5
R26170 DVSS.n544 DVSS.n543 292.5
R26171 DVSS.n543 DVSS.n514 292.5
R26172 DVSS.n527 DVSS.n526 292.5
R26173 DVSS.n923 DVSS.n922 292.5
R26174 DVSS.n922 DVSS.n483 292.5
R26175 DVSS.n924 DVSS.n492 292.5
R26176 DVSS.n492 DVSS.n491 292.5
R26177 DVSS.n926 DVSS.n925 292.5
R26178 DVSS.n927 DVSS.n926 292.5
R26179 DVSS.n901 DVSS.n490 292.5
R26180 DVSS.n490 DVSS.n489 292.5
R26181 DVSS.n899 DVSS.n898 292.5
R26182 DVSS.n898 DVSS.n897 292.5
R26183 DVSS.n495 DVSS.n494 292.5
R26184 DVSS.n497 DVSS.n495 292.5
R26185 DVSS.n853 DVSS.n511 292.5
R26186 DVSS.n511 DVSS.n509 292.5
R26187 DVSS.n855 DVSS.n854 292.5
R26188 DVSS.n856 DVSS.n855 292.5
R26189 DVSS.n852 DVSS.n510 292.5
R26190 DVSS.n515 DVSS.n510 292.5
R26191 DVSS.n851 DVSS.n850 292.5
R26192 DVSS.n850 DVSS.n849 292.5
R26193 DVSS.n834 DVSS.n833 292.5
R26194 DVSS.n835 DVSS.n834 292.5
R26195 DVSS.n832 DVSS.n548 292.5
R26196 DVSS.n548 DVSS.n547 292.5
R26197 DVSS.n831 DVSS.n830 292.5
R26198 DVSS.n830 DVSS.n829 292.5
R26199 DVSS.n550 DVSS.n549 292.5
R26200 DVSS.n551 DVSS.n550 292.5
R26201 DVSS.n921 DVSS.n902 292.5
R26202 DVSS.n907 DVSS.n903 292.5
R26203 DVSS.n917 DVSS.n916 292.5
R26204 DVSS.n915 DVSS.n906 292.5
R26205 DVSS.n914 DVSS.n913 292.5
R26206 DVSS.n912 DVSS.n911 292.5
R26207 DVSS.n910 DVSS.n909 292.5
R26208 DVSS.n908 DVSS.n480 292.5
R26209 DVSS.n938 DVSS.n937 292.5
R26210 DVSS.n1719 DVSS.n1718 292.5
R26211 DVSS.n1721 DVSS.n1720 292.5
R26212 DVSS.n1724 DVSS.n1723 292.5
R26213 DVSS.n1730 DVSS.n1729 292.5
R26214 DVSS.n1716 DVSS.n1715 292.5
R26215 DVSS.n1697 DVSS.n1695 292.5
R26216 DVSS.n1682 DVSS.n1680 292.5
R26217 DVSS.n1667 DVSS.n1665 292.5
R26218 DVSS.n1664 DVSS.n1663 292.5
R26219 DVSS.n1641 DVSS.n1640 292.5
R26220 DVSS.n1639 DVSS.n1638 292.5
R26221 DVSS.n1623 DVSS.n1622 292.5
R26222 DVSS.n1608 DVSS.n1607 292.5
R26223 DVSS.n1593 DVSS.n1592 292.5
R26224 DVSS.n1578 DVSS.n1577 292.5
R26225 DVSS.n1563 DVSS.n1562 292.5
R26226 DVSS.n1548 DVSS.n1547 292.5
R26227 DVSS.n1533 DVSS.n1532 292.5
R26228 DVSS.n1522 DVSS.n1520 292.5
R26229 DVSS.n1507 DVSS.n1505 292.5
R26230 DVSS.n1492 DVSS.n1490 292.5
R26231 DVSS.n1477 DVSS.n1475 292.5
R26232 DVSS.n1462 DVSS.n1460 292.5
R26233 DVSS.n1447 DVSS.n1445 292.5
R26234 DVSS.n1432 DVSS.n1430 292.5
R26235 DVSS.n1417 DVSS.n1415 292.5
R26236 DVSS.n1414 DVSS.n1413 292.5
R26237 DVSS.n1391 DVSS.n1390 292.5
R26238 DVSS.n1389 DVSS.n1388 292.5
R26239 DVSS.n1373 DVSS.n1372 292.5
R26240 DVSS.n962 DVSS.n961 292.5
R26241 DVSS.n960 DVSS.n959 292.5
R26242 DVSS.n957 DVSS.n956 292.5
R26243 DVSS.n955 DVSS.n954 292.5
R26244 DVSS.n1358 DVSS.n1357 292.5
R26245 DVSS.n1350 DVSS.n1349 292.5
R26246 DVSS.t260 DVSS.n1062 277.438
R26247 DVSS.n6073 DVSS.n6072 270.849
R26248 DVSS.n6099 DVSS.n6095 270.849
R26249 DVSS.n6323 DVSS.n6322 270.849
R26250 DVSS.n6349 DVSS.n6345 270.849
R26251 DVSS.n4605 DVSS.n4604 270.849
R26252 DVSS.n4631 DVSS.n4627 270.849
R26253 DVSS.n4855 DVSS.n4854 270.849
R26254 DVSS.n4881 DVSS.n4877 270.849
R26255 DVSS.n3009 DVSS.n3008 270.849
R26256 DVSS.n3035 DVSS.n3031 270.849
R26257 DVSS.n3259 DVSS.n3258 270.849
R26258 DVSS.n3285 DVSS.n3281 270.849
R26259 DVSS.n1392 DVSS.n1391 270.849
R26260 DVSS.n1418 DVSS.n1414 270.849
R26261 DVSS.n1642 DVSS.n1641 270.849
R26262 DVSS.n1668 DVSS.n1664 270.849
R26263 DVSS.n3968 DVSS.n3648 270.034
R26264 DVSS.n3628 DVSS.n3622 270.034
R26265 DVSS.n3632 DVSS.n3620 270.034
R26266 DVSS.n3966 DVSS.n3645 270.034
R26267 DVSS.n4433 DVSS.n4113 270.034
R26268 DVSS.n4093 DVSS.n4087 270.034
R26269 DVSS.n4097 DVSS.n4085 270.034
R26270 DVSS.n4431 DVSS.n4110 270.034
R26271 DVSS.n2372 DVSS.n2052 270.034
R26272 DVSS.n2032 DVSS.n2026 270.034
R26273 DVSS.n2036 DVSS.n2024 270.034
R26274 DVSS.n2370 DVSS.n2049 270.034
R26275 DVSS.n2837 DVSS.n2517 270.034
R26276 DVSS.n2497 DVSS.n2491 270.034
R26277 DVSS.n2501 DVSS.n2489 270.034
R26278 DVSS.n2835 DVSS.n2514 270.034
R26279 DVSS.n5436 DVSS.n5116 270.034
R26280 DVSS.n5096 DVSS.n5090 270.034
R26281 DVSS.n5100 DVSS.n5088 270.034
R26282 DVSS.n5434 DVSS.n5113 270.034
R26283 DVSS.n5901 DVSS.n5581 270.034
R26284 DVSS.n5561 DVSS.n5555 270.034
R26285 DVSS.n5565 DVSS.n5553 270.034
R26286 DVSS.n5899 DVSS.n5578 270.034
R26287 DVSS.n371 DVSS.n51 270.034
R26288 DVSS.n31 DVSS.n25 270.034
R26289 DVSS.n35 DVSS.n23 270.034
R26290 DVSS.n369 DVSS.n48 270.034
R26291 DVSS.n836 DVSS.n516 270.034
R26292 DVSS.n496 DVSS.n490 270.034
R26293 DVSS.n500 DVSS.n488 270.034
R26294 DVSS.n834 DVSS.n513 270.034
R26295 DVSS.n6525 DVSS.n6524 255.838
R26296 DVSS.n1255 DVSS.t149 252.812
R26297 DVSS.n3654 DVSS.n3646 248.683
R26298 DVSS.n3668 DVSS.n3646 248.683
R26299 DVSS.n3666 DVSS.n3646 248.683
R26300 DVSS.n4119 DVSS.n4111 248.683
R26301 DVSS.n4133 DVSS.n4111 248.683
R26302 DVSS.n4131 DVSS.n4111 248.683
R26303 DVSS.n2058 DVSS.n2050 248.683
R26304 DVSS.n2072 DVSS.n2050 248.683
R26305 DVSS.n2070 DVSS.n2050 248.683
R26306 DVSS.n2523 DVSS.n2515 248.683
R26307 DVSS.n2537 DVSS.n2515 248.683
R26308 DVSS.n2535 DVSS.n2515 248.683
R26309 DVSS.n5122 DVSS.n5114 248.683
R26310 DVSS.n5136 DVSS.n5114 248.683
R26311 DVSS.n5134 DVSS.n5114 248.683
R26312 DVSS.n5587 DVSS.n5579 248.683
R26313 DVSS.n5601 DVSS.n5579 248.683
R26314 DVSS.n5599 DVSS.n5579 248.683
R26315 DVSS.n57 DVSS.n49 248.683
R26316 DVSS.n71 DVSS.n49 248.683
R26317 DVSS.n69 DVSS.n49 248.683
R26318 DVSS.n522 DVSS.n514 248.683
R26319 DVSS.n536 DVSS.n514 248.683
R26320 DVSS.n534 DVSS.n514 248.683
R26321 DVSS.n3937 DVSS.n3765 245.512
R26322 DVSS.n3937 DVSS.n3766 245.512
R26323 DVSS.n3937 DVSS.n3767 245.512
R26324 DVSS.n3937 DVSS.n3768 245.512
R26325 DVSS.n3937 DVSS.n3936 245.512
R26326 DVSS.n3711 DVSS.n3692 245.512
R26327 DVSS.n3711 DVSS.n3693 245.512
R26328 DVSS.n3711 DVSS.n3694 245.512
R26329 DVSS.n3711 DVSS.n3695 245.512
R26330 DVSS.n3711 DVSS.n3710 245.512
R26331 DVSS.n4402 DVSS.n4230 245.512
R26332 DVSS.n4402 DVSS.n4231 245.512
R26333 DVSS.n4402 DVSS.n4232 245.512
R26334 DVSS.n4402 DVSS.n4233 245.512
R26335 DVSS.n4402 DVSS.n4401 245.512
R26336 DVSS.n4176 DVSS.n4157 245.512
R26337 DVSS.n4176 DVSS.n4158 245.512
R26338 DVSS.n4176 DVSS.n4159 245.512
R26339 DVSS.n4176 DVSS.n4160 245.512
R26340 DVSS.n4176 DVSS.n4175 245.512
R26341 DVSS.n2341 DVSS.n2169 245.512
R26342 DVSS.n2341 DVSS.n2170 245.512
R26343 DVSS.n2341 DVSS.n2171 245.512
R26344 DVSS.n2341 DVSS.n2172 245.512
R26345 DVSS.n2341 DVSS.n2340 245.512
R26346 DVSS.n2115 DVSS.n2096 245.512
R26347 DVSS.n2115 DVSS.n2097 245.512
R26348 DVSS.n2115 DVSS.n2098 245.512
R26349 DVSS.n2115 DVSS.n2099 245.512
R26350 DVSS.n2115 DVSS.n2114 245.512
R26351 DVSS.n2806 DVSS.n2634 245.512
R26352 DVSS.n2806 DVSS.n2635 245.512
R26353 DVSS.n2806 DVSS.n2636 245.512
R26354 DVSS.n2806 DVSS.n2637 245.512
R26355 DVSS.n2806 DVSS.n2805 245.512
R26356 DVSS.n2580 DVSS.n2561 245.512
R26357 DVSS.n2580 DVSS.n2562 245.512
R26358 DVSS.n2580 DVSS.n2563 245.512
R26359 DVSS.n2580 DVSS.n2564 245.512
R26360 DVSS.n2580 DVSS.n2579 245.512
R26361 DVSS.n5405 DVSS.n5233 245.512
R26362 DVSS.n5405 DVSS.n5234 245.512
R26363 DVSS.n5405 DVSS.n5235 245.512
R26364 DVSS.n5405 DVSS.n5236 245.512
R26365 DVSS.n5405 DVSS.n5404 245.512
R26366 DVSS.n5179 DVSS.n5160 245.512
R26367 DVSS.n5179 DVSS.n5161 245.512
R26368 DVSS.n5179 DVSS.n5162 245.512
R26369 DVSS.n5179 DVSS.n5163 245.512
R26370 DVSS.n5179 DVSS.n5178 245.512
R26371 DVSS.n5870 DVSS.n5698 245.512
R26372 DVSS.n5870 DVSS.n5699 245.512
R26373 DVSS.n5870 DVSS.n5700 245.512
R26374 DVSS.n5870 DVSS.n5701 245.512
R26375 DVSS.n5870 DVSS.n5869 245.512
R26376 DVSS.n5644 DVSS.n5625 245.512
R26377 DVSS.n5644 DVSS.n5626 245.512
R26378 DVSS.n5644 DVSS.n5627 245.512
R26379 DVSS.n5644 DVSS.n5628 245.512
R26380 DVSS.n5644 DVSS.n5643 245.512
R26381 DVSS.n340 DVSS.n168 245.512
R26382 DVSS.n340 DVSS.n169 245.512
R26383 DVSS.n340 DVSS.n170 245.512
R26384 DVSS.n340 DVSS.n171 245.512
R26385 DVSS.n340 DVSS.n339 245.512
R26386 DVSS.n114 DVSS.n95 245.512
R26387 DVSS.n114 DVSS.n96 245.512
R26388 DVSS.n114 DVSS.n97 245.512
R26389 DVSS.n114 DVSS.n98 245.512
R26390 DVSS.n114 DVSS.n113 245.512
R26391 DVSS.n805 DVSS.n633 245.512
R26392 DVSS.n805 DVSS.n634 245.512
R26393 DVSS.n805 DVSS.n635 245.512
R26394 DVSS.n805 DVSS.n636 245.512
R26395 DVSS.n805 DVSS.n804 245.512
R26396 DVSS.n579 DVSS.n560 245.512
R26397 DVSS.n579 DVSS.n561 245.512
R26398 DVSS.n579 DVSS.n562 245.512
R26399 DVSS.n579 DVSS.n563 245.512
R26400 DVSS.n579 DVSS.n578 245.512
R26401 DVSS.n3401 DVSS.t15 232.049
R26402 DVSS.n4996 DVSS.t204 232.049
R26403 DVSS.n1784 DVSS.t141 232.049
R26404 DVSS.n3422 DVSS.t7 230.262
R26405 DVSS.n5017 DVSS.t208 230.262
R26406 DVSS.n1805 DVSS.t137 230.262
R26407 DVSS.n6485 DVSS.t210 230.262
R26408 DVSS.n3837 DVSS.n3836 223.931
R26409 DVSS.n3834 DVSS.n3810 223.931
R26410 DVSS.n3827 DVSS.n3826 223.931
R26411 DVSS.n3892 DVSS.n3785 223.931
R26412 DVSS.n3896 DVSS.n3785 223.931
R26413 DVSS.n3896 DVSS.n3759 223.931
R26414 DVSS.n3919 DVSS.n3763 223.931
R26415 DVSS.n3890 DVSS.n3784 223.931
R26416 DVSS.n3898 DVSS.n3784 223.931
R26417 DVSS.n3899 DVSS.n3898 223.931
R26418 DVSS.n3863 DVSS.n3862 223.931
R26419 DVSS.n3859 DVSS.n3858 223.931
R26420 DVSS.n3855 DVSS.n3850 223.931
R26421 DVSS.n3878 DVSS.n3846 223.931
R26422 DVSS.n3878 DVSS.n3797 223.931
R26423 DVSS.n3882 DVSS.n3797 223.931
R26424 DVSS.n3812 DVSS.n3804 223.931
R26425 DVSS.n3819 DVSS.n3814 223.931
R26426 DVSS.n3823 DVSS.n3821 223.931
R26427 DVSS.n3876 DVSS.n3848 223.931
R26428 DVSS.n3876 DVSS.n3794 223.931
R26429 DVSS.n3884 DVSS.n3794 223.931
R26430 DVSS.n3960 DVSS.n3684 223.931
R26431 DVSS.n3960 DVSS.n3678 223.931
R26432 DVSS.n3968 DVSS.n3678 223.931
R26433 DVSS.n3712 DVSS.n3689 223.931
R26434 DVSS.n4058 DVSS.n3622 223.931
R26435 DVSS.n4058 DVSS.n3624 223.931
R26436 DVSS.n4054 DVSS.n3624 223.931
R26437 DVSS.n4049 DVSS.n4038 223.931
R26438 DVSS.n4045 DVSS.n4044 223.931
R26439 DVSS.n4041 DVSS.n4040 223.931
R26440 DVSS.n4060 DVSS.n3620 223.931
R26441 DVSS.n4060 DVSS.n3614 223.931
R26442 DVSS.n4069 DVSS.n3614 223.931
R26443 DVSS.n3980 DVSS.n3639 223.931
R26444 DVSS.n3989 DVSS.n3639 223.931
R26445 DVSS.n3989 DVSS.n3640 223.931
R26446 DVSS.n3640 DVSS.n3631 223.931
R26447 DVSS.n4028 DVSS.n3631 223.931
R26448 DVSS.n3982 DVSS.n3642 223.931
R26449 DVSS.n3987 DVSS.n3642 223.931
R26450 DVSS.n3987 DVSS.n3643 223.931
R26451 DVSS.n3643 DVSS.n3627 223.931
R26452 DVSS.n4030 DVSS.n3627 223.931
R26453 DVSS.n3962 DVSS.n3682 223.931
R26454 DVSS.n3962 DVSS.n3680 223.931
R26455 DVSS.n3966 DVSS.n3680 223.931
R26456 DVSS.n4302 DVSS.n4301 223.931
R26457 DVSS.n4299 DVSS.n4275 223.931
R26458 DVSS.n4292 DVSS.n4291 223.931
R26459 DVSS.n4357 DVSS.n4250 223.931
R26460 DVSS.n4361 DVSS.n4250 223.931
R26461 DVSS.n4361 DVSS.n4224 223.931
R26462 DVSS.n4384 DVSS.n4228 223.931
R26463 DVSS.n4355 DVSS.n4249 223.931
R26464 DVSS.n4363 DVSS.n4249 223.931
R26465 DVSS.n4364 DVSS.n4363 223.931
R26466 DVSS.n4328 DVSS.n4327 223.931
R26467 DVSS.n4324 DVSS.n4323 223.931
R26468 DVSS.n4320 DVSS.n4315 223.931
R26469 DVSS.n4343 DVSS.n4311 223.931
R26470 DVSS.n4343 DVSS.n4262 223.931
R26471 DVSS.n4347 DVSS.n4262 223.931
R26472 DVSS.n4277 DVSS.n4269 223.931
R26473 DVSS.n4284 DVSS.n4279 223.931
R26474 DVSS.n4288 DVSS.n4286 223.931
R26475 DVSS.n4341 DVSS.n4313 223.931
R26476 DVSS.n4341 DVSS.n4259 223.931
R26477 DVSS.n4349 DVSS.n4259 223.931
R26478 DVSS.n4425 DVSS.n4149 223.931
R26479 DVSS.n4425 DVSS.n4143 223.931
R26480 DVSS.n4433 DVSS.n4143 223.931
R26481 DVSS.n4177 DVSS.n4154 223.931
R26482 DVSS.n4523 DVSS.n4087 223.931
R26483 DVSS.n4523 DVSS.n4089 223.931
R26484 DVSS.n4519 DVSS.n4089 223.931
R26485 DVSS.n4514 DVSS.n4503 223.931
R26486 DVSS.n4510 DVSS.n4509 223.931
R26487 DVSS.n4506 DVSS.n4505 223.931
R26488 DVSS.n4525 DVSS.n4085 223.931
R26489 DVSS.n4525 DVSS.n4079 223.931
R26490 DVSS.n4533 DVSS.n4079 223.931
R26491 DVSS.n4445 DVSS.n4104 223.931
R26492 DVSS.n4454 DVSS.n4104 223.931
R26493 DVSS.n4454 DVSS.n4105 223.931
R26494 DVSS.n4105 DVSS.n4096 223.931
R26495 DVSS.n4493 DVSS.n4096 223.931
R26496 DVSS.n4447 DVSS.n4107 223.931
R26497 DVSS.n4452 DVSS.n4107 223.931
R26498 DVSS.n4452 DVSS.n4108 223.931
R26499 DVSS.n4108 DVSS.n4092 223.931
R26500 DVSS.n4495 DVSS.n4092 223.931
R26501 DVSS.n4427 DVSS.n4147 223.931
R26502 DVSS.n4427 DVSS.n4145 223.931
R26503 DVSS.n4431 DVSS.n4145 223.931
R26504 DVSS.n2241 DVSS.n2240 223.931
R26505 DVSS.n2238 DVSS.n2214 223.931
R26506 DVSS.n2231 DVSS.n2230 223.931
R26507 DVSS.n2296 DVSS.n2189 223.931
R26508 DVSS.n2300 DVSS.n2189 223.931
R26509 DVSS.n2300 DVSS.n2163 223.931
R26510 DVSS.n2323 DVSS.n2167 223.931
R26511 DVSS.n2294 DVSS.n2188 223.931
R26512 DVSS.n2302 DVSS.n2188 223.931
R26513 DVSS.n2303 DVSS.n2302 223.931
R26514 DVSS.n2267 DVSS.n2266 223.931
R26515 DVSS.n2263 DVSS.n2262 223.931
R26516 DVSS.n2259 DVSS.n2254 223.931
R26517 DVSS.n2282 DVSS.n2250 223.931
R26518 DVSS.n2282 DVSS.n2201 223.931
R26519 DVSS.n2286 DVSS.n2201 223.931
R26520 DVSS.n2216 DVSS.n2208 223.931
R26521 DVSS.n2223 DVSS.n2218 223.931
R26522 DVSS.n2227 DVSS.n2225 223.931
R26523 DVSS.n2280 DVSS.n2252 223.931
R26524 DVSS.n2280 DVSS.n2198 223.931
R26525 DVSS.n2288 DVSS.n2198 223.931
R26526 DVSS.n2364 DVSS.n2088 223.931
R26527 DVSS.n2364 DVSS.n2082 223.931
R26528 DVSS.n2372 DVSS.n2082 223.931
R26529 DVSS.n2116 DVSS.n2093 223.931
R26530 DVSS.n2462 DVSS.n2026 223.931
R26531 DVSS.n2462 DVSS.n2028 223.931
R26532 DVSS.n2458 DVSS.n2028 223.931
R26533 DVSS.n2453 DVSS.n2442 223.931
R26534 DVSS.n2449 DVSS.n2448 223.931
R26535 DVSS.n2445 DVSS.n2444 223.931
R26536 DVSS.n2464 DVSS.n2024 223.931
R26537 DVSS.n2464 DVSS.n2018 223.931
R26538 DVSS.n2473 DVSS.n2018 223.931
R26539 DVSS.n2384 DVSS.n2043 223.931
R26540 DVSS.n2393 DVSS.n2043 223.931
R26541 DVSS.n2393 DVSS.n2044 223.931
R26542 DVSS.n2044 DVSS.n2035 223.931
R26543 DVSS.n2432 DVSS.n2035 223.931
R26544 DVSS.n2386 DVSS.n2046 223.931
R26545 DVSS.n2391 DVSS.n2046 223.931
R26546 DVSS.n2391 DVSS.n2047 223.931
R26547 DVSS.n2047 DVSS.n2031 223.931
R26548 DVSS.n2434 DVSS.n2031 223.931
R26549 DVSS.n2366 DVSS.n2086 223.931
R26550 DVSS.n2366 DVSS.n2084 223.931
R26551 DVSS.n2370 DVSS.n2084 223.931
R26552 DVSS.n2706 DVSS.n2705 223.931
R26553 DVSS.n2703 DVSS.n2679 223.931
R26554 DVSS.n2696 DVSS.n2695 223.931
R26555 DVSS.n2761 DVSS.n2654 223.931
R26556 DVSS.n2765 DVSS.n2654 223.931
R26557 DVSS.n2765 DVSS.n2628 223.931
R26558 DVSS.n2788 DVSS.n2632 223.931
R26559 DVSS.n2759 DVSS.n2653 223.931
R26560 DVSS.n2767 DVSS.n2653 223.931
R26561 DVSS.n2768 DVSS.n2767 223.931
R26562 DVSS.n2732 DVSS.n2731 223.931
R26563 DVSS.n2728 DVSS.n2727 223.931
R26564 DVSS.n2724 DVSS.n2719 223.931
R26565 DVSS.n2747 DVSS.n2715 223.931
R26566 DVSS.n2747 DVSS.n2666 223.931
R26567 DVSS.n2751 DVSS.n2666 223.931
R26568 DVSS.n2681 DVSS.n2673 223.931
R26569 DVSS.n2688 DVSS.n2683 223.931
R26570 DVSS.n2692 DVSS.n2690 223.931
R26571 DVSS.n2745 DVSS.n2717 223.931
R26572 DVSS.n2745 DVSS.n2663 223.931
R26573 DVSS.n2753 DVSS.n2663 223.931
R26574 DVSS.n2829 DVSS.n2553 223.931
R26575 DVSS.n2829 DVSS.n2547 223.931
R26576 DVSS.n2837 DVSS.n2547 223.931
R26577 DVSS.n2581 DVSS.n2558 223.931
R26578 DVSS.n2927 DVSS.n2491 223.931
R26579 DVSS.n2927 DVSS.n2493 223.931
R26580 DVSS.n2923 DVSS.n2493 223.931
R26581 DVSS.n2918 DVSS.n2907 223.931
R26582 DVSS.n2914 DVSS.n2913 223.931
R26583 DVSS.n2910 DVSS.n2909 223.931
R26584 DVSS.n2929 DVSS.n2489 223.931
R26585 DVSS.n2929 DVSS.n2483 223.931
R26586 DVSS.n2937 DVSS.n2483 223.931
R26587 DVSS.n2849 DVSS.n2508 223.931
R26588 DVSS.n2858 DVSS.n2508 223.931
R26589 DVSS.n2858 DVSS.n2509 223.931
R26590 DVSS.n2509 DVSS.n2500 223.931
R26591 DVSS.n2897 DVSS.n2500 223.931
R26592 DVSS.n2851 DVSS.n2511 223.931
R26593 DVSS.n2856 DVSS.n2511 223.931
R26594 DVSS.n2856 DVSS.n2512 223.931
R26595 DVSS.n2512 DVSS.n2496 223.931
R26596 DVSS.n2899 DVSS.n2496 223.931
R26597 DVSS.n2831 DVSS.n2551 223.931
R26598 DVSS.n2831 DVSS.n2549 223.931
R26599 DVSS.n2835 DVSS.n2549 223.931
R26600 DVSS.n5305 DVSS.n5304 223.931
R26601 DVSS.n5302 DVSS.n5278 223.931
R26602 DVSS.n5295 DVSS.n5294 223.931
R26603 DVSS.n5360 DVSS.n5253 223.931
R26604 DVSS.n5364 DVSS.n5253 223.931
R26605 DVSS.n5364 DVSS.n5227 223.931
R26606 DVSS.n5387 DVSS.n5231 223.931
R26607 DVSS.n5358 DVSS.n5252 223.931
R26608 DVSS.n5366 DVSS.n5252 223.931
R26609 DVSS.n5367 DVSS.n5366 223.931
R26610 DVSS.n5331 DVSS.n5330 223.931
R26611 DVSS.n5327 DVSS.n5326 223.931
R26612 DVSS.n5323 DVSS.n5318 223.931
R26613 DVSS.n5346 DVSS.n5314 223.931
R26614 DVSS.n5346 DVSS.n5265 223.931
R26615 DVSS.n5350 DVSS.n5265 223.931
R26616 DVSS.n5280 DVSS.n5272 223.931
R26617 DVSS.n5287 DVSS.n5282 223.931
R26618 DVSS.n5291 DVSS.n5289 223.931
R26619 DVSS.n5344 DVSS.n5316 223.931
R26620 DVSS.n5344 DVSS.n5262 223.931
R26621 DVSS.n5352 DVSS.n5262 223.931
R26622 DVSS.n5428 DVSS.n5152 223.931
R26623 DVSS.n5428 DVSS.n5146 223.931
R26624 DVSS.n5436 DVSS.n5146 223.931
R26625 DVSS.n5180 DVSS.n5157 223.931
R26626 DVSS.n5526 DVSS.n5090 223.931
R26627 DVSS.n5526 DVSS.n5092 223.931
R26628 DVSS.n5522 DVSS.n5092 223.931
R26629 DVSS.n5517 DVSS.n5506 223.931
R26630 DVSS.n5513 DVSS.n5512 223.931
R26631 DVSS.n5509 DVSS.n5508 223.931
R26632 DVSS.n5528 DVSS.n5088 223.931
R26633 DVSS.n5528 DVSS.n5082 223.931
R26634 DVSS.n5537 DVSS.n5082 223.931
R26635 DVSS.n5448 DVSS.n5107 223.931
R26636 DVSS.n5457 DVSS.n5107 223.931
R26637 DVSS.n5457 DVSS.n5108 223.931
R26638 DVSS.n5108 DVSS.n5099 223.931
R26639 DVSS.n5496 DVSS.n5099 223.931
R26640 DVSS.n5450 DVSS.n5110 223.931
R26641 DVSS.n5455 DVSS.n5110 223.931
R26642 DVSS.n5455 DVSS.n5111 223.931
R26643 DVSS.n5111 DVSS.n5095 223.931
R26644 DVSS.n5498 DVSS.n5095 223.931
R26645 DVSS.n5430 DVSS.n5150 223.931
R26646 DVSS.n5430 DVSS.n5148 223.931
R26647 DVSS.n5434 DVSS.n5148 223.931
R26648 DVSS.n5770 DVSS.n5769 223.931
R26649 DVSS.n5767 DVSS.n5743 223.931
R26650 DVSS.n5760 DVSS.n5759 223.931
R26651 DVSS.n5825 DVSS.n5718 223.931
R26652 DVSS.n5829 DVSS.n5718 223.931
R26653 DVSS.n5829 DVSS.n5692 223.931
R26654 DVSS.n5852 DVSS.n5696 223.931
R26655 DVSS.n5823 DVSS.n5717 223.931
R26656 DVSS.n5831 DVSS.n5717 223.931
R26657 DVSS.n5832 DVSS.n5831 223.931
R26658 DVSS.n5796 DVSS.n5795 223.931
R26659 DVSS.n5792 DVSS.n5791 223.931
R26660 DVSS.n5788 DVSS.n5783 223.931
R26661 DVSS.n5811 DVSS.n5779 223.931
R26662 DVSS.n5811 DVSS.n5730 223.931
R26663 DVSS.n5815 DVSS.n5730 223.931
R26664 DVSS.n5745 DVSS.n5737 223.931
R26665 DVSS.n5752 DVSS.n5747 223.931
R26666 DVSS.n5756 DVSS.n5754 223.931
R26667 DVSS.n5809 DVSS.n5781 223.931
R26668 DVSS.n5809 DVSS.n5727 223.931
R26669 DVSS.n5817 DVSS.n5727 223.931
R26670 DVSS.n5893 DVSS.n5617 223.931
R26671 DVSS.n5893 DVSS.n5611 223.931
R26672 DVSS.n5901 DVSS.n5611 223.931
R26673 DVSS.n5645 DVSS.n5622 223.931
R26674 DVSS.n5991 DVSS.n5555 223.931
R26675 DVSS.n5991 DVSS.n5557 223.931
R26676 DVSS.n5987 DVSS.n5557 223.931
R26677 DVSS.n5982 DVSS.n5971 223.931
R26678 DVSS.n5978 DVSS.n5977 223.931
R26679 DVSS.n5974 DVSS.n5973 223.931
R26680 DVSS.n5993 DVSS.n5553 223.931
R26681 DVSS.n5993 DVSS.n5547 223.931
R26682 DVSS.n6001 DVSS.n5547 223.931
R26683 DVSS.n5913 DVSS.n5572 223.931
R26684 DVSS.n5922 DVSS.n5572 223.931
R26685 DVSS.n5922 DVSS.n5573 223.931
R26686 DVSS.n5573 DVSS.n5564 223.931
R26687 DVSS.n5961 DVSS.n5564 223.931
R26688 DVSS.n5915 DVSS.n5575 223.931
R26689 DVSS.n5920 DVSS.n5575 223.931
R26690 DVSS.n5920 DVSS.n5576 223.931
R26691 DVSS.n5576 DVSS.n5560 223.931
R26692 DVSS.n5963 DVSS.n5560 223.931
R26693 DVSS.n5895 DVSS.n5615 223.931
R26694 DVSS.n5895 DVSS.n5613 223.931
R26695 DVSS.n5899 DVSS.n5613 223.931
R26696 DVSS.n240 DVSS.n239 223.931
R26697 DVSS.n237 DVSS.n213 223.931
R26698 DVSS.n230 DVSS.n229 223.931
R26699 DVSS.n295 DVSS.n188 223.931
R26700 DVSS.n299 DVSS.n188 223.931
R26701 DVSS.n299 DVSS.n162 223.931
R26702 DVSS.n322 DVSS.n166 223.931
R26703 DVSS.n293 DVSS.n187 223.931
R26704 DVSS.n301 DVSS.n187 223.931
R26705 DVSS.n302 DVSS.n301 223.931
R26706 DVSS.n266 DVSS.n265 223.931
R26707 DVSS.n262 DVSS.n261 223.931
R26708 DVSS.n258 DVSS.n253 223.931
R26709 DVSS.n281 DVSS.n249 223.931
R26710 DVSS.n281 DVSS.n200 223.931
R26711 DVSS.n285 DVSS.n200 223.931
R26712 DVSS.n215 DVSS.n207 223.931
R26713 DVSS.n222 DVSS.n217 223.931
R26714 DVSS.n226 DVSS.n224 223.931
R26715 DVSS.n279 DVSS.n251 223.931
R26716 DVSS.n279 DVSS.n197 223.931
R26717 DVSS.n287 DVSS.n197 223.931
R26718 DVSS.n363 DVSS.n87 223.931
R26719 DVSS.n363 DVSS.n81 223.931
R26720 DVSS.n371 DVSS.n81 223.931
R26721 DVSS.n115 DVSS.n92 223.931
R26722 DVSS.n461 DVSS.n25 223.931
R26723 DVSS.n461 DVSS.n27 223.931
R26724 DVSS.n457 DVSS.n27 223.931
R26725 DVSS.n452 DVSS.n441 223.931
R26726 DVSS.n448 DVSS.n447 223.931
R26727 DVSS.n444 DVSS.n443 223.931
R26728 DVSS.n463 DVSS.n23 223.931
R26729 DVSS.n463 DVSS.n17 223.931
R26730 DVSS.n472 DVSS.n17 223.931
R26731 DVSS.n383 DVSS.n42 223.931
R26732 DVSS.n392 DVSS.n42 223.931
R26733 DVSS.n392 DVSS.n43 223.931
R26734 DVSS.n43 DVSS.n34 223.931
R26735 DVSS.n431 DVSS.n34 223.931
R26736 DVSS.n385 DVSS.n45 223.931
R26737 DVSS.n390 DVSS.n45 223.931
R26738 DVSS.n390 DVSS.n46 223.931
R26739 DVSS.n46 DVSS.n30 223.931
R26740 DVSS.n433 DVSS.n30 223.931
R26741 DVSS.n365 DVSS.n85 223.931
R26742 DVSS.n365 DVSS.n83 223.931
R26743 DVSS.n369 DVSS.n83 223.931
R26744 DVSS.n705 DVSS.n704 223.931
R26745 DVSS.n702 DVSS.n678 223.931
R26746 DVSS.n695 DVSS.n694 223.931
R26747 DVSS.n760 DVSS.n653 223.931
R26748 DVSS.n764 DVSS.n653 223.931
R26749 DVSS.n764 DVSS.n627 223.931
R26750 DVSS.n787 DVSS.n631 223.931
R26751 DVSS.n758 DVSS.n652 223.931
R26752 DVSS.n766 DVSS.n652 223.931
R26753 DVSS.n767 DVSS.n766 223.931
R26754 DVSS.n731 DVSS.n730 223.931
R26755 DVSS.n727 DVSS.n726 223.931
R26756 DVSS.n723 DVSS.n718 223.931
R26757 DVSS.n746 DVSS.n714 223.931
R26758 DVSS.n746 DVSS.n665 223.931
R26759 DVSS.n750 DVSS.n665 223.931
R26760 DVSS.n680 DVSS.n672 223.931
R26761 DVSS.n687 DVSS.n682 223.931
R26762 DVSS.n691 DVSS.n689 223.931
R26763 DVSS.n744 DVSS.n716 223.931
R26764 DVSS.n744 DVSS.n662 223.931
R26765 DVSS.n752 DVSS.n662 223.931
R26766 DVSS.n828 DVSS.n552 223.931
R26767 DVSS.n828 DVSS.n546 223.931
R26768 DVSS.n836 DVSS.n546 223.931
R26769 DVSS.n580 DVSS.n557 223.931
R26770 DVSS.n926 DVSS.n490 223.931
R26771 DVSS.n926 DVSS.n492 223.931
R26772 DVSS.n922 DVSS.n492 223.931
R26773 DVSS.n917 DVSS.n906 223.931
R26774 DVSS.n913 DVSS.n912 223.931
R26775 DVSS.n909 DVSS.n908 223.931
R26776 DVSS.n928 DVSS.n488 223.931
R26777 DVSS.n928 DVSS.n482 223.931
R26778 DVSS.n936 DVSS.n482 223.931
R26779 DVSS.n848 DVSS.n507 223.931
R26780 DVSS.n857 DVSS.n507 223.931
R26781 DVSS.n857 DVSS.n508 223.931
R26782 DVSS.n508 DVSS.n499 223.931
R26783 DVSS.n896 DVSS.n499 223.931
R26784 DVSS.n850 DVSS.n510 223.931
R26785 DVSS.n855 DVSS.n510 223.931
R26786 DVSS.n855 DVSS.n511 223.931
R26787 DVSS.n511 DVSS.n495 223.931
R26788 DVSS.n898 DVSS.n495 223.931
R26789 DVSS.n830 DVSS.n550 223.931
R26790 DVSS.n830 DVSS.n548 223.931
R26791 DVSS.n834 DVSS.n548 223.931
R26792 DVSS.n4007 DVSS.n4005 206.16
R26793 DVSS.n4011 DVSS.n4004 206.16
R26794 DVSS.n4014 DVSS.n4013 206.16
R26795 DVSS.n4018 DVSS.n4017 206.16
R26796 DVSS.n3662 DVSS.n3661 206.16
R26797 DVSS.n3675 DVSS.n3674 206.16
R26798 DVSS.n4472 DVSS.n4470 206.16
R26799 DVSS.n4476 DVSS.n4469 206.16
R26800 DVSS.n4479 DVSS.n4478 206.16
R26801 DVSS.n4483 DVSS.n4482 206.16
R26802 DVSS.n4127 DVSS.n4126 206.16
R26803 DVSS.n4140 DVSS.n4139 206.16
R26804 DVSS.n2411 DVSS.n2409 206.16
R26805 DVSS.n2415 DVSS.n2408 206.16
R26806 DVSS.n2418 DVSS.n2417 206.16
R26807 DVSS.n2422 DVSS.n2421 206.16
R26808 DVSS.n2066 DVSS.n2065 206.16
R26809 DVSS.n2079 DVSS.n2078 206.16
R26810 DVSS.n2876 DVSS.n2874 206.16
R26811 DVSS.n2880 DVSS.n2873 206.16
R26812 DVSS.n2883 DVSS.n2882 206.16
R26813 DVSS.n2887 DVSS.n2886 206.16
R26814 DVSS.n2531 DVSS.n2530 206.16
R26815 DVSS.n2544 DVSS.n2543 206.16
R26816 DVSS.n5475 DVSS.n5473 206.16
R26817 DVSS.n5479 DVSS.n5472 206.16
R26818 DVSS.n5482 DVSS.n5481 206.16
R26819 DVSS.n5486 DVSS.n5485 206.16
R26820 DVSS.n5130 DVSS.n5129 206.16
R26821 DVSS.n5143 DVSS.n5142 206.16
R26822 DVSS.n5940 DVSS.n5938 206.16
R26823 DVSS.n5944 DVSS.n5937 206.16
R26824 DVSS.n5947 DVSS.n5946 206.16
R26825 DVSS.n5951 DVSS.n5950 206.16
R26826 DVSS.n5595 DVSS.n5594 206.16
R26827 DVSS.n5608 DVSS.n5607 206.16
R26828 DVSS.n410 DVSS.n408 206.16
R26829 DVSS.n414 DVSS.n407 206.16
R26830 DVSS.n417 DVSS.n416 206.16
R26831 DVSS.n421 DVSS.n420 206.16
R26832 DVSS.n65 DVSS.n64 206.16
R26833 DVSS.n78 DVSS.n77 206.16
R26834 DVSS.n875 DVSS.n873 206.16
R26835 DVSS.n879 DVSS.n872 206.16
R26836 DVSS.n882 DVSS.n881 206.16
R26837 DVSS.n886 DVSS.n885 206.16
R26838 DVSS.n530 DVSS.n529 206.16
R26839 DVSS.n543 DVSS.n542 206.16
R26840 DVSS.n969 DVSS.n963 200.287
R26841 DVSS.n3988 DVSS.t66 199.196
R26842 DVSS.n3641 DVSS.t222 199.196
R26843 DVSS.n4453 DVSS.t96 199.196
R26844 DVSS.n4106 DVSS.t38 199.196
R26845 DVSS.n2392 DVSS.t74 199.196
R26846 DVSS.n2045 DVSS.t73 199.196
R26847 DVSS.n2857 DVSS.t22 199.196
R26848 DVSS.n2510 DVSS.t21 199.196
R26849 DVSS.n5456 DVSS.t20 199.196
R26850 DVSS.n5109 DVSS.t162 199.196
R26851 DVSS.n5921 DVSS.t107 199.196
R26852 DVSS.n5574 DVSS.t153 199.196
R26853 DVSS.n391 DVSS.t68 199.196
R26854 DVSS.n44 DVSS.t67 199.196
R26855 DVSS.n856 DVSS.t174 199.196
R26856 DVSS.n509 DVSS.t37 199.196
R26857 DVSS.n1264 DVSS.t238 199.023
R26858 DVSS.n3438 DVSS.t11 196.35
R26859 DVSS.n5033 DVSS.t198 196.35
R26860 DVSS.n1821 DVSS.t139 196.35
R26861 DVSS.n1343 DVSS.n1156 194.454
R26862 DVSS.n3751 DVSS.n3738 185
R26863 DVSS.n3753 DVSS.n3752 185
R26864 DVSS.n3730 DVSS.n3717 185
R26865 DVSS.n3732 DVSS.n3731 185
R26866 DVSS.n4216 DVSS.n4203 185
R26867 DVSS.n4218 DVSS.n4217 185
R26868 DVSS.n4195 DVSS.n4182 185
R26869 DVSS.n4197 DVSS.n4196 185
R26870 DVSS.n2155 DVSS.n2142 185
R26871 DVSS.n2157 DVSS.n2156 185
R26872 DVSS.n2134 DVSS.n2121 185
R26873 DVSS.n2136 DVSS.n2135 185
R26874 DVSS.n2620 DVSS.n2607 185
R26875 DVSS.n2622 DVSS.n2621 185
R26876 DVSS.n2599 DVSS.n2586 185
R26877 DVSS.n2601 DVSS.n2600 185
R26878 DVSS.n5219 DVSS.n5206 185
R26879 DVSS.n5221 DVSS.n5220 185
R26880 DVSS.n5198 DVSS.n5185 185
R26881 DVSS.n5200 DVSS.n5199 185
R26882 DVSS.n5684 DVSS.n5671 185
R26883 DVSS.n5686 DVSS.n5685 185
R26884 DVSS.n5663 DVSS.n5650 185
R26885 DVSS.n5665 DVSS.n5664 185
R26886 DVSS.n154 DVSS.n141 185
R26887 DVSS.n156 DVSS.n155 185
R26888 DVSS.n133 DVSS.n120 185
R26889 DVSS.n135 DVSS.n134 185
R26890 DVSS.n619 DVSS.n606 185
R26891 DVSS.n621 DVSS.n620 185
R26892 DVSS.n598 DVSS.n585 185
R26893 DVSS.n600 DVSS.n599 185
R26894 DVSS.n1057 DVSS.n1055 184.572
R26895 DVSS.n1100 DVSS.n1098 184.572
R26896 DVSS.n1106 DVSS.n1104 184.572
R26897 DVSS.n1393 DVSS.n1386 174.535
R26898 DVSS.n1419 DVSS.n1410 174.535
R26899 DVSS.n1643 DVSS.n1636 174.535
R26900 DVSS.n1669 DVSS.n1660 174.535
R26901 DVSS.n4606 DVSS.n4599 174.535
R26902 DVSS.n4632 DVSS.n4623 174.535
R26903 DVSS.n4856 DVSS.n4849 174.535
R26904 DVSS.n4882 DVSS.n4873 174.535
R26905 DVSS.n6074 DVSS.n6067 174.535
R26906 DVSS.n6100 DVSS.n6091 174.535
R26907 DVSS.n6324 DVSS.n6317 174.535
R26908 DVSS.n6350 DVSS.n6341 174.535
R26909 DVSS.n3010 DVSS.n3003 174.535
R26910 DVSS.n3036 DVSS.n3027 174.535
R26911 DVSS.n3260 DVSS.n3253 174.535
R26912 DVSS.n3286 DVSS.n3277 174.535
R26913 DVSS.n3435 DVSS.n3434 161.605
R26914 DVSS.n5030 DVSS.n5029 161.605
R26915 DVSS.n1818 DVSS.n1817 161.605
R26916 DVSS.n3877 DVSS.t81 158.811
R26917 DVSS.t81 DVSS.n3795 158.811
R26918 DVSS.n3789 DVSS.t185 158.811
R26919 DVSS.n3897 DVSS.t185 158.811
R26920 DVSS.t83 DVSS.n3903 158.811
R26921 DVSS.n3904 DVSS.t83 158.811
R26922 DVSS.n4342 DVSS.t84 158.811
R26923 DVSS.t84 DVSS.n4260 158.811
R26924 DVSS.n4254 DVSS.t118 158.811
R26925 DVSS.n4362 DVSS.t118 158.811
R26926 DVSS.t86 DVSS.n4368 158.811
R26927 DVSS.n4369 DVSS.t86 158.811
R26928 DVSS.n2281 DVSS.t124 158.811
R26929 DVSS.t124 DVSS.n2199 158.811
R26930 DVSS.n2193 DVSS.t223 158.811
R26931 DVSS.n2301 DVSS.t223 158.811
R26932 DVSS.t123 DVSS.n2307 158.811
R26933 DVSS.n2308 DVSS.t123 158.811
R26934 DVSS.n2746 DVSS.t120 158.811
R26935 DVSS.t120 DVSS.n2664 158.811
R26936 DVSS.n2658 DVSS.t61 158.811
R26937 DVSS.n2766 DVSS.t61 158.811
R26938 DVSS.t122 DVSS.n2772 158.811
R26939 DVSS.n2773 DVSS.t122 158.811
R26940 DVSS.n5345 DVSS.t79 158.811
R26941 DVSS.t79 DVSS.n5263 158.811
R26942 DVSS.n5257 DVSS.t91 158.811
R26943 DVSS.n5365 DVSS.t91 158.811
R26944 DVSS.t78 DVSS.n5371 158.811
R26945 DVSS.n5372 DVSS.t78 158.811
R26946 DVSS.n5810 DVSS.t76 158.811
R26947 DVSS.t76 DVSS.n5728 158.811
R26948 DVSS.n5722 DVSS.t151 158.811
R26949 DVSS.n5830 DVSS.t151 158.811
R26950 DVSS.t75 DVSS.n5836 158.811
R26951 DVSS.n5837 DVSS.t75 158.811
R26952 DVSS.n280 DVSS.t112 158.811
R26953 DVSS.t112 DVSS.n198 158.811
R26954 DVSS.n192 DVSS.t187 158.811
R26955 DVSS.n300 DVSS.t187 158.811
R26956 DVSS.t108 DVSS.n306 158.811
R26957 DVSS.n307 DVSS.t108 158.811
R26958 DVSS.n745 DVSS.t109 158.811
R26959 DVSS.t109 DVSS.n663 158.811
R26960 DVSS.n657 DVSS.t230 158.811
R26961 DVSS.n765 DVSS.t230 158.811
R26962 DVSS.t111 DVSS.n771 158.811
R26963 DVSS.n772 DVSS.t111 158.811
R26964 DVSS.n3656 DVSS.n3646 157.904
R26965 DVSS.n4121 DVSS.n4111 157.904
R26966 DVSS.n2060 DVSS.n2050 157.904
R26967 DVSS.n2525 DVSS.n2515 157.904
R26968 DVSS.n5124 DVSS.n5114 157.904
R26969 DVSS.n5589 DVSS.n5579 157.904
R26970 DVSS.n59 DVSS.n49 157.904
R26971 DVSS.n524 DVSS.n514 157.904
R26972 DVSS.n3673 DVSS.n3646 157.904
R26973 DVSS.n4138 DVSS.n4111 157.904
R26974 DVSS.n2077 DVSS.n2050 157.904
R26975 DVSS.n2542 DVSS.n2515 157.904
R26976 DVSS.n5141 DVSS.n5114 157.904
R26977 DVSS.n5606 DVSS.n5579 157.904
R26978 DVSS.n76 DVSS.n49 157.904
R26979 DVSS.n541 DVSS.n514 157.904
R26980 DVSS.n3938 DVSS.n3937 155.356
R26981 DVSS.n4403 DVSS.n4402 155.356
R26982 DVSS.n6409 DVSS.n6408 155.356
R26983 DVSS.n4941 DVSS.n4940 155.356
R26984 DVSS.n2342 DVSS.n2341 155.356
R26985 DVSS.n2807 DVSS.n2806 155.356
R26986 DVSS.n3346 DVSS.n3345 155.356
R26987 DVSS.n5406 DVSS.n5405 155.356
R26988 DVSS.n5871 DVSS.n5870 155.356
R26989 DVSS.n341 DVSS.n340 155.356
R26990 DVSS.n806 DVSS.n805 155.356
R26991 DVSS.n1728 DVSS.n1727 155.356
R26992 DVSS.n3869 DVSS.n3868 155.356
R26993 DVSS.n3869 DVSS.n3853 155.356
R26994 DVSS.n3937 DVSS.n3764 155.356
R26995 DVSS.n3798 DVSS.n3796 155.356
R26996 DVSS.n3806 DVSS.n3788 155.356
R26997 DVSS.n3803 DVSS.n3796 155.356
R26998 DVSS.n3808 DVSS.n3788 155.356
R26999 DVSS.n3711 DVSS.n3690 155.356
R27000 DVSS.n3711 DVSS.n3691 155.356
R27001 DVSS.n4052 DVSS.n4051 155.356
R27002 DVSS.n4051 DVSS.n4050 155.356
R27003 DVSS.n4334 DVSS.n4333 155.356
R27004 DVSS.n4334 DVSS.n4318 155.356
R27005 DVSS.n4402 DVSS.n4229 155.356
R27006 DVSS.n4263 DVSS.n4261 155.356
R27007 DVSS.n4271 DVSS.n4253 155.356
R27008 DVSS.n4268 DVSS.n4261 155.356
R27009 DVSS.n4273 DVSS.n4253 155.356
R27010 DVSS.n4176 DVSS.n4155 155.356
R27011 DVSS.n4176 DVSS.n4156 155.356
R27012 DVSS.n4517 DVSS.n4516 155.356
R27013 DVSS.n4516 DVSS.n4515 155.356
R27014 DVSS.n2273 DVSS.n2272 155.356
R27015 DVSS.n2273 DVSS.n2257 155.356
R27016 DVSS.n2341 DVSS.n2168 155.356
R27017 DVSS.n2202 DVSS.n2200 155.356
R27018 DVSS.n2210 DVSS.n2192 155.356
R27019 DVSS.n2207 DVSS.n2200 155.356
R27020 DVSS.n2212 DVSS.n2192 155.356
R27021 DVSS.n2115 DVSS.n2094 155.356
R27022 DVSS.n2115 DVSS.n2095 155.356
R27023 DVSS.n2456 DVSS.n2455 155.356
R27024 DVSS.n2455 DVSS.n2454 155.356
R27025 DVSS.n2738 DVSS.n2737 155.356
R27026 DVSS.n2738 DVSS.n2722 155.356
R27027 DVSS.n2806 DVSS.n2633 155.356
R27028 DVSS.n2667 DVSS.n2665 155.356
R27029 DVSS.n2675 DVSS.n2657 155.356
R27030 DVSS.n2672 DVSS.n2665 155.356
R27031 DVSS.n2677 DVSS.n2657 155.356
R27032 DVSS.n2580 DVSS.n2559 155.356
R27033 DVSS.n2580 DVSS.n2560 155.356
R27034 DVSS.n2921 DVSS.n2920 155.356
R27035 DVSS.n2920 DVSS.n2919 155.356
R27036 DVSS.n5337 DVSS.n5336 155.356
R27037 DVSS.n5337 DVSS.n5321 155.356
R27038 DVSS.n5405 DVSS.n5232 155.356
R27039 DVSS.n5266 DVSS.n5264 155.356
R27040 DVSS.n5274 DVSS.n5256 155.356
R27041 DVSS.n5271 DVSS.n5264 155.356
R27042 DVSS.n5276 DVSS.n5256 155.356
R27043 DVSS.n5179 DVSS.n5158 155.356
R27044 DVSS.n5179 DVSS.n5159 155.356
R27045 DVSS.n5520 DVSS.n5519 155.356
R27046 DVSS.n5519 DVSS.n5518 155.356
R27047 DVSS.n5802 DVSS.n5801 155.356
R27048 DVSS.n5802 DVSS.n5786 155.356
R27049 DVSS.n5870 DVSS.n5697 155.356
R27050 DVSS.n5731 DVSS.n5729 155.356
R27051 DVSS.n5739 DVSS.n5721 155.356
R27052 DVSS.n5736 DVSS.n5729 155.356
R27053 DVSS.n5741 DVSS.n5721 155.356
R27054 DVSS.n5644 DVSS.n5623 155.356
R27055 DVSS.n5644 DVSS.n5624 155.356
R27056 DVSS.n5985 DVSS.n5984 155.356
R27057 DVSS.n5984 DVSS.n5983 155.356
R27058 DVSS.n272 DVSS.n271 155.356
R27059 DVSS.n272 DVSS.n256 155.356
R27060 DVSS.n340 DVSS.n167 155.356
R27061 DVSS.n201 DVSS.n199 155.356
R27062 DVSS.n209 DVSS.n191 155.356
R27063 DVSS.n206 DVSS.n199 155.356
R27064 DVSS.n211 DVSS.n191 155.356
R27065 DVSS.n114 DVSS.n93 155.356
R27066 DVSS.n114 DVSS.n94 155.356
R27067 DVSS.n455 DVSS.n454 155.356
R27068 DVSS.n454 DVSS.n453 155.356
R27069 DVSS.n737 DVSS.n736 155.356
R27070 DVSS.n737 DVSS.n721 155.356
R27071 DVSS.n805 DVSS.n632 155.356
R27072 DVSS.n666 DVSS.n664 155.356
R27073 DVSS.n674 DVSS.n656 155.356
R27074 DVSS.n671 DVSS.n664 155.356
R27075 DVSS.n676 DVSS.n656 155.356
R27076 DVSS.n579 DVSS.n558 155.356
R27077 DVSS.n579 DVSS.n559 155.356
R27078 DVSS.n920 DVSS.n919 155.356
R27079 DVSS.n919 DVSS.n918 155.356
R27080 DVSS.n3961 DVSS.t65 150.504
R27081 DVSS.t65 DVSS.n3679 150.504
R27082 DVSS.n4059 DVSS.t19 150.504
R27083 DVSS.n3623 DVSS.t19 150.504
R27084 DVSS.n4426 DVSS.t52 150.504
R27085 DVSS.t52 DVSS.n4144 150.504
R27086 DVSS.n4524 DVSS.t51 150.504
R27087 DVSS.n4088 DVSS.t51 150.504
R27088 DVSS.n2365 DVSS.t225 150.504
R27089 DVSS.t225 DVSS.n2083 150.504
R27090 DVSS.n2463 DVSS.t193 150.504
R27091 DVSS.n2027 DVSS.t193 150.504
R27092 DVSS.n2830 DVSS.t130 150.504
R27093 DVSS.t130 DVSS.n2548 150.504
R27094 DVSS.n2928 DVSS.t129 150.504
R27095 DVSS.n2492 DVSS.t129 150.504
R27096 DVSS.n5429 DVSS.t169 150.504
R27097 DVSS.t169 DVSS.n5147 150.504
R27098 DVSS.n5527 DVSS.t234 150.504
R27099 DVSS.n5091 DVSS.t234 150.504
R27100 DVSS.n5894 DVSS.t147 150.504
R27101 DVSS.t147 DVSS.n5612 150.504
R27102 DVSS.n5992 DVSS.t148 150.504
R27103 DVSS.n5556 DVSS.t148 150.504
R27104 DVSS.n364 DVSS.t95 150.504
R27105 DVSS.t95 DVSS.n82 150.504
R27106 DVSS.n462 DVSS.t126 150.504
R27107 DVSS.n26 DVSS.t126 150.504
R27108 DVSS.n829 DVSS.t167 150.504
R27109 DVSS.t167 DVSS.n547 150.504
R27110 DVSS.n927 DVSS.t168 150.504
R27111 DVSS.n491 DVSS.t168 150.504
R27112 DVSS.n6665 DVSS.t254 147.352
R27113 DVSS.t145 DVSS.t235 147.06
R27114 DVSS.n1869 DVSS.t59 146.894
R27115 DVSS.n6464 DVSS.t218 130.149
R27116 DVSS.n1243 DVSS.n1242 129.095
R27117 DVSS.t15 DVSS.n3400 125.389
R27118 DVSS.t204 DVSS.n4995 125.389
R27119 DVSS.t141 DVSS.n1783 125.389
R27120 DVSS.t55 DVSS.n6698 124.132
R27121 DVSS.t93 DVSS.n6733 124.132
R27122 DVSS.n6717 DVSS.n6716 122.674
R27123 DVSS.n6754 DVSS.n6753 122.472
R27124 DVSS.n3746 DVSS.t186 119.998
R27125 DVSS.n3725 DVSS.t82 119.998
R27126 DVSS.n4211 DVSS.t119 119.998
R27127 DVSS.n4190 DVSS.t85 119.998
R27128 DVSS.n2150 DVSS.t224 119.998
R27129 DVSS.n2129 DVSS.t125 119.998
R27130 DVSS.n2615 DVSS.t62 119.998
R27131 DVSS.n2594 DVSS.t121 119.998
R27132 DVSS.n5214 DVSS.t92 119.998
R27133 DVSS.n5193 DVSS.t80 119.998
R27134 DVSS.n5679 DVSS.t152 119.998
R27135 DVSS.n5658 DVSS.t77 119.998
R27136 DVSS.n149 DVSS.t188 119.998
R27137 DVSS.n128 DVSS.t113 119.998
R27138 DVSS.n614 DVSS.t231 119.998
R27139 DVSS.n593 DVSS.t110 119.998
R27140 DVSS.n3938 DVSS.n3760 118.938
R27141 DVSS.n4403 DVSS.n4225 118.938
R27142 DVSS.n2342 DVSS.n2164 118.938
R27143 DVSS.n2807 DVSS.n2629 118.938
R27144 DVSS.n5406 DVSS.n5228 118.938
R27145 DVSS.n5871 DVSS.n5693 118.938
R27146 DVSS.n341 DVSS.n163 118.938
R27147 DVSS.n806 DVSS.n628 118.938
R27148 DVSS.n3868 DVSS.n3854 118.936
R27149 DVSS.n3854 DVSS.n3853 118.936
R27150 DVSS.n3777 DVSS.n3764 118.936
R27151 DVSS.n3802 DVSS.n3798 118.936
R27152 DVSS.n3807 DVSS.n3806 118.936
R27153 DVSS.n3803 DVSS.n3802 118.936
R27154 DVSS.n3808 DVSS.n3807 118.936
R27155 DVSS.n3696 DVSS.n3690 118.936
R27156 DVSS.n3700 DVSS.n3691 118.936
R27157 DVSS.n4052 DVSS.n4035 118.936
R27158 DVSS.n4050 DVSS.n4035 118.936
R27159 DVSS.n4333 DVSS.n4319 118.936
R27160 DVSS.n4319 DVSS.n4318 118.936
R27161 DVSS.n4242 DVSS.n4229 118.936
R27162 DVSS.n4267 DVSS.n4263 118.936
R27163 DVSS.n4272 DVSS.n4271 118.936
R27164 DVSS.n4268 DVSS.n4267 118.936
R27165 DVSS.n4273 DVSS.n4272 118.936
R27166 DVSS.n4161 DVSS.n4155 118.936
R27167 DVSS.n4165 DVSS.n4156 118.936
R27168 DVSS.n4517 DVSS.n4500 118.936
R27169 DVSS.n4515 DVSS.n4500 118.936
R27170 DVSS.n2272 DVSS.n2258 118.936
R27171 DVSS.n2258 DVSS.n2257 118.936
R27172 DVSS.n2181 DVSS.n2168 118.936
R27173 DVSS.n2206 DVSS.n2202 118.936
R27174 DVSS.n2211 DVSS.n2210 118.936
R27175 DVSS.n2207 DVSS.n2206 118.936
R27176 DVSS.n2212 DVSS.n2211 118.936
R27177 DVSS.n2100 DVSS.n2094 118.936
R27178 DVSS.n2104 DVSS.n2095 118.936
R27179 DVSS.n2456 DVSS.n2439 118.936
R27180 DVSS.n2454 DVSS.n2439 118.936
R27181 DVSS.n2737 DVSS.n2723 118.936
R27182 DVSS.n2723 DVSS.n2722 118.936
R27183 DVSS.n2646 DVSS.n2633 118.936
R27184 DVSS.n2671 DVSS.n2667 118.936
R27185 DVSS.n2676 DVSS.n2675 118.936
R27186 DVSS.n2672 DVSS.n2671 118.936
R27187 DVSS.n2677 DVSS.n2676 118.936
R27188 DVSS.n2565 DVSS.n2559 118.936
R27189 DVSS.n2569 DVSS.n2560 118.936
R27190 DVSS.n2921 DVSS.n2904 118.936
R27191 DVSS.n2919 DVSS.n2904 118.936
R27192 DVSS.n5336 DVSS.n5322 118.936
R27193 DVSS.n5322 DVSS.n5321 118.936
R27194 DVSS.n5245 DVSS.n5232 118.936
R27195 DVSS.n5270 DVSS.n5266 118.936
R27196 DVSS.n5275 DVSS.n5274 118.936
R27197 DVSS.n5271 DVSS.n5270 118.936
R27198 DVSS.n5276 DVSS.n5275 118.936
R27199 DVSS.n5164 DVSS.n5158 118.936
R27200 DVSS.n5168 DVSS.n5159 118.936
R27201 DVSS.n5520 DVSS.n5503 118.936
R27202 DVSS.n5518 DVSS.n5503 118.936
R27203 DVSS.n5801 DVSS.n5787 118.936
R27204 DVSS.n5787 DVSS.n5786 118.936
R27205 DVSS.n5710 DVSS.n5697 118.936
R27206 DVSS.n5735 DVSS.n5731 118.936
R27207 DVSS.n5740 DVSS.n5739 118.936
R27208 DVSS.n5736 DVSS.n5735 118.936
R27209 DVSS.n5741 DVSS.n5740 118.936
R27210 DVSS.n5629 DVSS.n5623 118.936
R27211 DVSS.n5633 DVSS.n5624 118.936
R27212 DVSS.n5985 DVSS.n5968 118.936
R27213 DVSS.n5983 DVSS.n5968 118.936
R27214 DVSS.n271 DVSS.n257 118.936
R27215 DVSS.n257 DVSS.n256 118.936
R27216 DVSS.n180 DVSS.n167 118.936
R27217 DVSS.n205 DVSS.n201 118.936
R27218 DVSS.n210 DVSS.n209 118.936
R27219 DVSS.n206 DVSS.n205 118.936
R27220 DVSS.n211 DVSS.n210 118.936
R27221 DVSS.n99 DVSS.n93 118.936
R27222 DVSS.n103 DVSS.n94 118.936
R27223 DVSS.n455 DVSS.n438 118.936
R27224 DVSS.n453 DVSS.n438 118.936
R27225 DVSS.n736 DVSS.n722 118.936
R27226 DVSS.n722 DVSS.n721 118.936
R27227 DVSS.n645 DVSS.n632 118.936
R27228 DVSS.n670 DVSS.n666 118.936
R27229 DVSS.n675 DVSS.n674 118.936
R27230 DVSS.n671 DVSS.n670 118.936
R27231 DVSS.n676 DVSS.n675 118.936
R27232 DVSS.n564 DVSS.n558 118.936
R27233 DVSS.n568 DVSS.n559 118.936
R27234 DVSS.n920 DVSS.n903 118.936
R27235 DVSS.n918 DVSS.n903 118.936
R27236 DVSS.n3909 DVSS.n3908 117.719
R27237 DVSS.n3917 DVSS.n3916 117.719
R27238 DVSS.n3906 DVSS.n3905 117.719
R27239 DVSS.n4374 DVSS.n4373 117.719
R27240 DVSS.n4382 DVSS.n4381 117.719
R27241 DVSS.n4371 DVSS.n4370 117.719
R27242 DVSS.n2313 DVSS.n2312 117.719
R27243 DVSS.n2321 DVSS.n2320 117.719
R27244 DVSS.n2310 DVSS.n2309 117.719
R27245 DVSS.n2778 DVSS.n2777 117.719
R27246 DVSS.n2786 DVSS.n2785 117.719
R27247 DVSS.n2775 DVSS.n2774 117.719
R27248 DVSS.n5377 DVSS.n5376 117.719
R27249 DVSS.n5385 DVSS.n5384 117.719
R27250 DVSS.n5374 DVSS.n5373 117.719
R27251 DVSS.n5842 DVSS.n5841 117.719
R27252 DVSS.n5850 DVSS.n5849 117.719
R27253 DVSS.n5839 DVSS.n5838 117.719
R27254 DVSS.n312 DVSS.n311 117.719
R27255 DVSS.n320 DVSS.n319 117.719
R27256 DVSS.n309 DVSS.n308 117.719
R27257 DVSS.n777 DVSS.n776 117.719
R27258 DVSS.n785 DVSS.n784 117.719
R27259 DVSS.n774 DVSS.n773 117.719
R27260 DVSS.n3916 DVSS.n3915 117.719
R27261 DVSS.n3905 DVSS.n3780 117.719
R27262 DVSS.n4381 DVSS.n4380 117.719
R27263 DVSS.n4370 DVSS.n4245 117.719
R27264 DVSS.n2320 DVSS.n2319 117.719
R27265 DVSS.n2309 DVSS.n2184 117.719
R27266 DVSS.n2785 DVSS.n2784 117.719
R27267 DVSS.n2774 DVSS.n2649 117.719
R27268 DVSS.n5384 DVSS.n5383 117.719
R27269 DVSS.n5373 DVSS.n5248 117.719
R27270 DVSS.n5849 DVSS.n5848 117.719
R27271 DVSS.n5838 DVSS.n5713 117.719
R27272 DVSS.n319 DVSS.n318 117.719
R27273 DVSS.n308 DVSS.n183 117.719
R27274 DVSS.n784 DVSS.n783 117.719
R27275 DVSS.n773 DVSS.n648 117.719
R27276 DVSS.n3908 DVSS.n3907 117.719
R27277 DVSS.n4373 DVSS.n4372 117.719
R27278 DVSS.n2312 DVSS.n2311 117.719
R27279 DVSS.n2777 DVSS.n2776 117.719
R27280 DVSS.n5376 DVSS.n5375 117.719
R27281 DVSS.n5841 DVSS.n5840 117.719
R27282 DVSS.n311 DVSS.n310 117.719
R27283 DVSS.n776 DVSS.n775 117.719
R27284 DVSS.n1078 DVSS.t161 115.689
R27285 DVSS.n7 DVSS.t164 114.245
R27286 DVSS.n3481 DVSS.t246 114.245
R27287 DVSS.n6705 DVSS.t56 114.245
R27288 DVSS.n6740 DVSS.t94 114.245
R27289 DVSS.n1180 DVSS.t3 113.74
R27290 DVSS.n3754 DVSS.n3753 112.831
R27291 DVSS.n3733 DVSS.n3732 112.831
R27292 DVSS.n4219 DVSS.n4218 112.831
R27293 DVSS.n4198 DVSS.n4197 112.831
R27294 DVSS.n2158 DVSS.n2157 112.831
R27295 DVSS.n2137 DVSS.n2136 112.831
R27296 DVSS.n2623 DVSS.n2622 112.831
R27297 DVSS.n2602 DVSS.n2601 112.831
R27298 DVSS.n5222 DVSS.n5221 112.831
R27299 DVSS.n5201 DVSS.n5200 112.831
R27300 DVSS.n5687 DVSS.n5686 112.831
R27301 DVSS.n5666 DVSS.n5665 112.831
R27302 DVSS.n157 DVSS.n156 112.831
R27303 DVSS.n136 DVSS.n135 112.831
R27304 DVSS.n622 DVSS.n621 112.831
R27305 DVSS.n601 DVSS.n600 112.831
R27306 DVSS.n964 DVSS.t266 112.501
R27307 DVSS.n1859 DVSS.t40 112.499
R27308 DVSS.n3483 DVSS.t88 112.499
R27309 DVSS.n3665 DVSS.n3656 111.293
R27310 DVSS.n4130 DVSS.n4121 111.293
R27311 DVSS.n2069 DVSS.n2060 111.293
R27312 DVSS.n2534 DVSS.n2525 111.293
R27313 DVSS.n5133 DVSS.n5124 111.293
R27314 DVSS.n5598 DVSS.n5589 111.293
R27315 DVSS.n68 DVSS.n59 111.293
R27316 DVSS.n533 DVSS.n524 111.293
R27317 DVSS.n3673 DVSS.n3672 111.293
R27318 DVSS.n4138 DVSS.n4137 111.293
R27319 DVSS.n2077 DVSS.n2076 111.293
R27320 DVSS.n2542 DVSS.n2541 111.293
R27321 DVSS.n5141 DVSS.n5140 111.293
R27322 DVSS.n5606 DVSS.n5605 111.293
R27323 DVSS.n76 DVSS.n75 111.293
R27324 DVSS.n541 DVSS.n540 111.293
R27325 DVSS.n6502 DVSS.t216 110.126
R27326 DVSS.n6694 DVSS.n6693 108.242
R27327 DVSS.n3660 DVSS.n3646 108.141
R27328 DVSS.n4125 DVSS.n4111 108.141
R27329 DVSS.n2064 DVSS.n2050 108.141
R27330 DVSS.n2529 DVSS.n2515 108.141
R27331 DVSS.n5128 DVSS.n5114 108.141
R27332 DVSS.n5593 DVSS.n5579 108.141
R27333 DVSS.n63 DVSS.n49 108.141
R27334 DVSS.n528 DVSS.n514 108.141
R27335 DVSS.n4006 DVSS.n3630 108.141
R27336 DVSS.n4012 DVSS.n3630 108.141
R27337 DVSS.n4002 DVSS.n3630 108.141
R27338 DVSS.n4019 DVSS.n3630 108.141
R27339 DVSS.n4471 DVSS.n4095 108.141
R27340 DVSS.n4477 DVSS.n4095 108.141
R27341 DVSS.n4467 DVSS.n4095 108.141
R27342 DVSS.n4484 DVSS.n4095 108.141
R27343 DVSS.n2410 DVSS.n2034 108.141
R27344 DVSS.n2416 DVSS.n2034 108.141
R27345 DVSS.n2406 DVSS.n2034 108.141
R27346 DVSS.n2423 DVSS.n2034 108.141
R27347 DVSS.n2875 DVSS.n2499 108.141
R27348 DVSS.n2881 DVSS.n2499 108.141
R27349 DVSS.n2871 DVSS.n2499 108.141
R27350 DVSS.n2888 DVSS.n2499 108.141
R27351 DVSS.n5474 DVSS.n5098 108.141
R27352 DVSS.n5480 DVSS.n5098 108.141
R27353 DVSS.n5470 DVSS.n5098 108.141
R27354 DVSS.n5487 DVSS.n5098 108.141
R27355 DVSS.n5939 DVSS.n5563 108.141
R27356 DVSS.n5945 DVSS.n5563 108.141
R27357 DVSS.n5935 DVSS.n5563 108.141
R27358 DVSS.n5952 DVSS.n5563 108.141
R27359 DVSS.n409 DVSS.n33 108.141
R27360 DVSS.n415 DVSS.n33 108.141
R27361 DVSS.n405 DVSS.n33 108.141
R27362 DVSS.n422 DVSS.n33 108.141
R27363 DVSS.n874 DVSS.n498 108.141
R27364 DVSS.n880 DVSS.n498 108.141
R27365 DVSS.n870 DVSS.n498 108.141
R27366 DVSS.n887 DVSS.n498 108.141
R27367 DVSS.n6729 DVSS.n6728 108.064
R27368 DVSS.n1198 DVSS.t173 108.037
R27369 DVSS.n3825 DVSS.n3788 105.766
R27370 DVSS.n4290 DVSS.n4253 105.766
R27371 DVSS.n6029 DVSS.n6028 105.766
R27372 DVSS.n4561 DVSS.n4560 105.766
R27373 DVSS.n2229 DVSS.n2192 105.766
R27374 DVSS.n2694 DVSS.n2657 105.766
R27375 DVSS.n2965 DVSS.n2964 105.766
R27376 DVSS.n5293 DVSS.n5256 105.766
R27377 DVSS.n5758 DVSS.n5721 105.766
R27378 DVSS.n228 DVSS.n191 105.766
R27379 DVSS.n693 DVSS.n656 105.766
R27380 DVSS.n1348 DVSS.n1347 105.766
R27381 DVSS.n3869 DVSS.n3852 105.766
R27382 DVSS.n3869 DVSS.n3851 105.766
R27383 DVSS.n3870 DVSS.n3869 105.766
R27384 DVSS.n3813 DVSS.n3796 105.766
R27385 DVSS.n3835 DVSS.n3788 105.766
R27386 DVSS.n3820 DVSS.n3796 105.766
R27387 DVSS.n3822 DVSS.n3788 105.766
R27388 DVSS.n3796 DVSS.n3793 105.766
R27389 DVSS.n4051 DVSS.n4037 105.766
R27390 DVSS.n4051 DVSS.n4036 105.766
R27391 DVSS.n4051 DVSS.n3613 105.766
R27392 DVSS.n4334 DVSS.n4317 105.766
R27393 DVSS.n4334 DVSS.n4316 105.766
R27394 DVSS.n4335 DVSS.n4334 105.766
R27395 DVSS.n4278 DVSS.n4261 105.766
R27396 DVSS.n4300 DVSS.n4253 105.766
R27397 DVSS.n4285 DVSS.n4261 105.766
R27398 DVSS.n4287 DVSS.n4253 105.766
R27399 DVSS.n4261 DVSS.n4258 105.766
R27400 DVSS.n4516 DVSS.n4502 105.766
R27401 DVSS.n4516 DVSS.n4501 105.766
R27402 DVSS.n4516 DVSS.n4078 105.766
R27403 DVSS.n2273 DVSS.n2256 105.766
R27404 DVSS.n2273 DVSS.n2255 105.766
R27405 DVSS.n2274 DVSS.n2273 105.766
R27406 DVSS.n2217 DVSS.n2200 105.766
R27407 DVSS.n2239 DVSS.n2192 105.766
R27408 DVSS.n2224 DVSS.n2200 105.766
R27409 DVSS.n2226 DVSS.n2192 105.766
R27410 DVSS.n2200 DVSS.n2197 105.766
R27411 DVSS.n2455 DVSS.n2441 105.766
R27412 DVSS.n2455 DVSS.n2440 105.766
R27413 DVSS.n2455 DVSS.n2017 105.766
R27414 DVSS.n2738 DVSS.n2721 105.766
R27415 DVSS.n2738 DVSS.n2720 105.766
R27416 DVSS.n2739 DVSS.n2738 105.766
R27417 DVSS.n2682 DVSS.n2665 105.766
R27418 DVSS.n2704 DVSS.n2657 105.766
R27419 DVSS.n2689 DVSS.n2665 105.766
R27420 DVSS.n2691 DVSS.n2657 105.766
R27421 DVSS.n2665 DVSS.n2662 105.766
R27422 DVSS.n2920 DVSS.n2906 105.766
R27423 DVSS.n2920 DVSS.n2905 105.766
R27424 DVSS.n2920 DVSS.n2482 105.766
R27425 DVSS.n5337 DVSS.n5320 105.766
R27426 DVSS.n5337 DVSS.n5319 105.766
R27427 DVSS.n5338 DVSS.n5337 105.766
R27428 DVSS.n5281 DVSS.n5264 105.766
R27429 DVSS.n5303 DVSS.n5256 105.766
R27430 DVSS.n5288 DVSS.n5264 105.766
R27431 DVSS.n5290 DVSS.n5256 105.766
R27432 DVSS.n5264 DVSS.n5261 105.766
R27433 DVSS.n5519 DVSS.n5505 105.766
R27434 DVSS.n5519 DVSS.n5504 105.766
R27435 DVSS.n5519 DVSS.n5081 105.766
R27436 DVSS.n5802 DVSS.n5785 105.766
R27437 DVSS.n5802 DVSS.n5784 105.766
R27438 DVSS.n5803 DVSS.n5802 105.766
R27439 DVSS.n5746 DVSS.n5729 105.766
R27440 DVSS.n5768 DVSS.n5721 105.766
R27441 DVSS.n5753 DVSS.n5729 105.766
R27442 DVSS.n5755 DVSS.n5721 105.766
R27443 DVSS.n5729 DVSS.n5726 105.766
R27444 DVSS.n5984 DVSS.n5970 105.766
R27445 DVSS.n5984 DVSS.n5969 105.766
R27446 DVSS.n5984 DVSS.n5546 105.766
R27447 DVSS.n272 DVSS.n255 105.766
R27448 DVSS.n272 DVSS.n254 105.766
R27449 DVSS.n273 DVSS.n272 105.766
R27450 DVSS.n216 DVSS.n199 105.766
R27451 DVSS.n238 DVSS.n191 105.766
R27452 DVSS.n223 DVSS.n199 105.766
R27453 DVSS.n225 DVSS.n191 105.766
R27454 DVSS.n199 DVSS.n196 105.766
R27455 DVSS.n454 DVSS.n440 105.766
R27456 DVSS.n454 DVSS.n439 105.766
R27457 DVSS.n454 DVSS.n16 105.766
R27458 DVSS.n737 DVSS.n720 105.766
R27459 DVSS.n737 DVSS.n719 105.766
R27460 DVSS.n738 DVSS.n737 105.766
R27461 DVSS.n681 DVSS.n664 105.766
R27462 DVSS.n703 DVSS.n656 105.766
R27463 DVSS.n688 DVSS.n664 105.766
R27464 DVSS.n690 DVSS.n656 105.766
R27465 DVSS.n664 DVSS.n661 105.766
R27466 DVSS.n919 DVSS.n905 105.766
R27467 DVSS.n919 DVSS.n904 105.766
R27468 DVSS.n919 DVSS.n481 105.766
R27469 DVSS.n3749 DVSS.n3748 104.172
R27470 DVSS.n3728 DVSS.n3727 104.172
R27471 DVSS.n4214 DVSS.n4213 104.172
R27472 DVSS.n4193 DVSS.n4192 104.172
R27473 DVSS.n2153 DVSS.n2152 104.172
R27474 DVSS.n2132 DVSS.n2131 104.172
R27475 DVSS.n2618 DVSS.n2617 104.172
R27476 DVSS.n2597 DVSS.n2596 104.172
R27477 DVSS.n5217 DVSS.n5216 104.172
R27478 DVSS.n5196 DVSS.n5195 104.172
R27479 DVSS.n5682 DVSS.n5681 104.172
R27480 DVSS.n5661 DVSS.n5660 104.172
R27481 DVSS.n152 DVSS.n151 104.172
R27482 DVSS.n131 DVSS.n130 104.172
R27483 DVSS.n617 DVSS.n616 104.172
R27484 DVSS.n596 DVSS.n595 104.172
R27485 DVSS.n1330 DVSS.t263 102.794
R27486 DVSS.n1890 DVSS.t90 102.794
R27487 DVSS.n6686 DVSS.t128 102.794
R27488 DVSS.n3647 DVSS.t66 101.811
R27489 DVSS.t222 DVSS.n3629 101.811
R27490 DVSS.n4112 DVSS.t96 101.811
R27491 DVSS.t38 DVSS.n4094 101.811
R27492 DVSS.n2051 DVSS.t74 101.811
R27493 DVSS.t73 DVSS.n2033 101.811
R27494 DVSS.n2516 DVSS.t22 101.811
R27495 DVSS.t21 DVSS.n2498 101.811
R27496 DVSS.n5115 DVSS.t20 101.811
R27497 DVSS.t162 DVSS.n5097 101.811
R27498 DVSS.n5580 DVSS.t107 101.811
R27499 DVSS.t153 DVSS.n5562 101.811
R27500 DVSS.n50 DVSS.t68 101.811
R27501 DVSS.t67 DVSS.n32 101.811
R27502 DVSS.n515 DVSS.t174 101.811
R27503 DVSS.t37 DVSS.n497 101.811
R27504 DVSS.n8 DVSS.t166 101.038
R27505 DVSS.n3500 DVSS.t54 101.038
R27506 DVSS.n5070 DVSS.t132 101.038
R27507 DVSS.n1898 DVSS.t115 101.038
R27508 DVSS.n1743 DVSS.t25 98.1749
R27509 DVSS.n4955 DVSS.t256 98.1749
R27510 DVSS.n3358 DVSS.t23 98.1749
R27511 DVSS.n6423 DVSS.t63 98.1749
R27512 DVSS.n3478 DVSS.n3477 95.4569
R27513 DVSS.n3936 DVSS.n3935 93.9796
R27514 DVSS.n3771 DVSS.n3768 93.9796
R27515 DVSS.n3928 DVSS.n3767 93.9796
R27516 DVSS.n3925 DVSS.n3766 93.9796
R27517 DVSS.n3777 DVSS.n3765 93.9796
R27518 DVSS.n3925 DVSS.n3765 93.9796
R27519 DVSS.n3928 DVSS.n3766 93.9796
R27520 DVSS.n3771 DVSS.n3767 93.9796
R27521 DVSS.n3935 DVSS.n3768 93.9796
R27522 DVSS.n3936 DVSS.n3760 93.9796
R27523 DVSS.n3710 DVSS.n3709 93.9796
R27524 DVSS.n3706 DVSS.n3695 93.9796
R27525 DVSS.n3704 DVSS.n3694 93.9796
R27526 DVSS.n3702 DVSS.n3693 93.9796
R27527 DVSS.n3700 DVSS.n3692 93.9796
R27528 DVSS.n3709 DVSS.n3695 93.9796
R27529 DVSS.n3706 DVSS.n3694 93.9796
R27530 DVSS.n3704 DVSS.n3693 93.9796
R27531 DVSS.n3702 DVSS.n3692 93.9796
R27532 DVSS.n3710 DVSS.n3696 93.9796
R27533 DVSS.n4401 DVSS.n4400 93.9796
R27534 DVSS.n4236 DVSS.n4233 93.9796
R27535 DVSS.n4393 DVSS.n4232 93.9796
R27536 DVSS.n4390 DVSS.n4231 93.9796
R27537 DVSS.n4242 DVSS.n4230 93.9796
R27538 DVSS.n4390 DVSS.n4230 93.9796
R27539 DVSS.n4393 DVSS.n4231 93.9796
R27540 DVSS.n4236 DVSS.n4232 93.9796
R27541 DVSS.n4400 DVSS.n4233 93.9796
R27542 DVSS.n4401 DVSS.n4225 93.9796
R27543 DVSS.n4175 DVSS.n4174 93.9796
R27544 DVSS.n4171 DVSS.n4160 93.9796
R27545 DVSS.n4169 DVSS.n4159 93.9796
R27546 DVSS.n4167 DVSS.n4158 93.9796
R27547 DVSS.n4165 DVSS.n4157 93.9796
R27548 DVSS.n4174 DVSS.n4160 93.9796
R27549 DVSS.n4171 DVSS.n4159 93.9796
R27550 DVSS.n4169 DVSS.n4158 93.9796
R27551 DVSS.n4167 DVSS.n4157 93.9796
R27552 DVSS.n4175 DVSS.n4161 93.9796
R27553 DVSS.n6404 DVSS.n6403 93.9796
R27554 DVSS.n4936 DVSS.n4935 93.9796
R27555 DVSS.n2340 DVSS.n2339 93.9796
R27556 DVSS.n2175 DVSS.n2172 93.9796
R27557 DVSS.n2332 DVSS.n2171 93.9796
R27558 DVSS.n2329 DVSS.n2170 93.9796
R27559 DVSS.n2181 DVSS.n2169 93.9796
R27560 DVSS.n2329 DVSS.n2169 93.9796
R27561 DVSS.n2332 DVSS.n2170 93.9796
R27562 DVSS.n2175 DVSS.n2171 93.9796
R27563 DVSS.n2339 DVSS.n2172 93.9796
R27564 DVSS.n2340 DVSS.n2164 93.9796
R27565 DVSS.n2114 DVSS.n2113 93.9796
R27566 DVSS.n2110 DVSS.n2099 93.9796
R27567 DVSS.n2108 DVSS.n2098 93.9796
R27568 DVSS.n2106 DVSS.n2097 93.9796
R27569 DVSS.n2104 DVSS.n2096 93.9796
R27570 DVSS.n2113 DVSS.n2099 93.9796
R27571 DVSS.n2110 DVSS.n2098 93.9796
R27572 DVSS.n2108 DVSS.n2097 93.9796
R27573 DVSS.n2106 DVSS.n2096 93.9796
R27574 DVSS.n2114 DVSS.n2100 93.9796
R27575 DVSS.n2805 DVSS.n2804 93.9796
R27576 DVSS.n2640 DVSS.n2637 93.9796
R27577 DVSS.n2797 DVSS.n2636 93.9796
R27578 DVSS.n2794 DVSS.n2635 93.9796
R27579 DVSS.n2646 DVSS.n2634 93.9796
R27580 DVSS.n2794 DVSS.n2634 93.9796
R27581 DVSS.n2797 DVSS.n2635 93.9796
R27582 DVSS.n2640 DVSS.n2636 93.9796
R27583 DVSS.n2804 DVSS.n2637 93.9796
R27584 DVSS.n2805 DVSS.n2629 93.9796
R27585 DVSS.n2579 DVSS.n2578 93.9796
R27586 DVSS.n2575 DVSS.n2564 93.9796
R27587 DVSS.n2573 DVSS.n2563 93.9796
R27588 DVSS.n2571 DVSS.n2562 93.9796
R27589 DVSS.n2569 DVSS.n2561 93.9796
R27590 DVSS.n2578 DVSS.n2564 93.9796
R27591 DVSS.n2575 DVSS.n2563 93.9796
R27592 DVSS.n2573 DVSS.n2562 93.9796
R27593 DVSS.n2571 DVSS.n2561 93.9796
R27594 DVSS.n2579 DVSS.n2565 93.9796
R27595 DVSS.n3340 DVSS.n3339 93.9796
R27596 DVSS.n5404 DVSS.n5403 93.9796
R27597 DVSS.n5239 DVSS.n5236 93.9796
R27598 DVSS.n5396 DVSS.n5235 93.9796
R27599 DVSS.n5393 DVSS.n5234 93.9796
R27600 DVSS.n5245 DVSS.n5233 93.9796
R27601 DVSS.n5393 DVSS.n5233 93.9796
R27602 DVSS.n5396 DVSS.n5234 93.9796
R27603 DVSS.n5239 DVSS.n5235 93.9796
R27604 DVSS.n5403 DVSS.n5236 93.9796
R27605 DVSS.n5404 DVSS.n5228 93.9796
R27606 DVSS.n5178 DVSS.n5177 93.9796
R27607 DVSS.n5174 DVSS.n5163 93.9796
R27608 DVSS.n5172 DVSS.n5162 93.9796
R27609 DVSS.n5170 DVSS.n5161 93.9796
R27610 DVSS.n5168 DVSS.n5160 93.9796
R27611 DVSS.n5177 DVSS.n5163 93.9796
R27612 DVSS.n5174 DVSS.n5162 93.9796
R27613 DVSS.n5172 DVSS.n5161 93.9796
R27614 DVSS.n5170 DVSS.n5160 93.9796
R27615 DVSS.n5178 DVSS.n5164 93.9796
R27616 DVSS.n5869 DVSS.n5868 93.9796
R27617 DVSS.n5704 DVSS.n5701 93.9796
R27618 DVSS.n5861 DVSS.n5700 93.9796
R27619 DVSS.n5858 DVSS.n5699 93.9796
R27620 DVSS.n5710 DVSS.n5698 93.9796
R27621 DVSS.n5858 DVSS.n5698 93.9796
R27622 DVSS.n5861 DVSS.n5699 93.9796
R27623 DVSS.n5704 DVSS.n5700 93.9796
R27624 DVSS.n5868 DVSS.n5701 93.9796
R27625 DVSS.n5869 DVSS.n5693 93.9796
R27626 DVSS.n5643 DVSS.n5642 93.9796
R27627 DVSS.n5639 DVSS.n5628 93.9796
R27628 DVSS.n5637 DVSS.n5627 93.9796
R27629 DVSS.n5635 DVSS.n5626 93.9796
R27630 DVSS.n5633 DVSS.n5625 93.9796
R27631 DVSS.n5642 DVSS.n5628 93.9796
R27632 DVSS.n5639 DVSS.n5627 93.9796
R27633 DVSS.n5637 DVSS.n5626 93.9796
R27634 DVSS.n5635 DVSS.n5625 93.9796
R27635 DVSS.n5643 DVSS.n5629 93.9796
R27636 DVSS.n339 DVSS.n338 93.9796
R27637 DVSS.n174 DVSS.n171 93.9796
R27638 DVSS.n331 DVSS.n170 93.9796
R27639 DVSS.n328 DVSS.n169 93.9796
R27640 DVSS.n180 DVSS.n168 93.9796
R27641 DVSS.n328 DVSS.n168 93.9796
R27642 DVSS.n331 DVSS.n169 93.9796
R27643 DVSS.n174 DVSS.n170 93.9796
R27644 DVSS.n338 DVSS.n171 93.9796
R27645 DVSS.n339 DVSS.n163 93.9796
R27646 DVSS.n113 DVSS.n112 93.9796
R27647 DVSS.n109 DVSS.n98 93.9796
R27648 DVSS.n107 DVSS.n97 93.9796
R27649 DVSS.n105 DVSS.n96 93.9796
R27650 DVSS.n103 DVSS.n95 93.9796
R27651 DVSS.n112 DVSS.n98 93.9796
R27652 DVSS.n109 DVSS.n97 93.9796
R27653 DVSS.n107 DVSS.n96 93.9796
R27654 DVSS.n105 DVSS.n95 93.9796
R27655 DVSS.n113 DVSS.n99 93.9796
R27656 DVSS.n804 DVSS.n803 93.9796
R27657 DVSS.n639 DVSS.n636 93.9796
R27658 DVSS.n796 DVSS.n635 93.9796
R27659 DVSS.n793 DVSS.n634 93.9796
R27660 DVSS.n645 DVSS.n633 93.9796
R27661 DVSS.n793 DVSS.n633 93.9796
R27662 DVSS.n796 DVSS.n634 93.9796
R27663 DVSS.n639 DVSS.n635 93.9796
R27664 DVSS.n803 DVSS.n636 93.9796
R27665 DVSS.n804 DVSS.n628 93.9796
R27666 DVSS.n578 DVSS.n577 93.9796
R27667 DVSS.n574 DVSS.n563 93.9796
R27668 DVSS.n572 DVSS.n562 93.9796
R27669 DVSS.n570 DVSS.n561 93.9796
R27670 DVSS.n568 DVSS.n560 93.9796
R27671 DVSS.n577 DVSS.n563 93.9796
R27672 DVSS.n574 DVSS.n562 93.9796
R27673 DVSS.n572 DVSS.n561 93.9796
R27674 DVSS.n570 DVSS.n560 93.9796
R27675 DVSS.n578 DVSS.n564 93.9796
R27676 DVSS.n1723 DVSS.n1722 93.9796
R27677 DVSS.n1140 DVSS.n1139 92.5005
R27678 DVSS.n1874 DVSS.n1873 92.5005
R27679 DVSS.n6670 DVSS.n6669 92.5005
R27680 DVSS.n3748 DVSS.n3747 92.5005
R27681 DVSS.n3727 DVSS.n3726 92.5005
R27682 DVSS.n4213 DVSS.n4212 92.5005
R27683 DVSS.n4192 DVSS.n4191 92.5005
R27684 DVSS.n2152 DVSS.n2151 92.5005
R27685 DVSS.n2131 DVSS.n2130 92.5005
R27686 DVSS.n2617 DVSS.n2616 92.5005
R27687 DVSS.n2596 DVSS.n2595 92.5005
R27688 DVSS.n5216 DVSS.n5215 92.5005
R27689 DVSS.n5195 DVSS.n5194 92.5005
R27690 DVSS.n5681 DVSS.n5680 92.5005
R27691 DVSS.n5660 DVSS.n5659 92.5005
R27692 DVSS.n151 DVSS.n150 92.5005
R27693 DVSS.n130 DVSS.n129 92.5005
R27694 DVSS.n616 DVSS.n615 92.5005
R27695 DVSS.n595 DVSS.n594 92.5005
R27696 DVSS.n6212 DVSS.t57 91.9866
R27697 DVSS.n4744 DVSS.t243 91.9866
R27698 DVSS.n3148 DVSS.t189 91.9866
R27699 DVSS.n1531 DVSS.t196 91.9866
R27700 DVSS.n1181 DVSS.t4 91.1965
R27701 DVSS.n1180 DVSS.t6 91.1965
R27702 DVSS.n10 DVSS.t34 90.704
R27703 DVSS.n3556 DVSS.t44 90.704
R27704 DVSS.n6595 DVSS.t104 90.704
R27705 DVSS.n1953 DVSS.t180 90.704
R27706 DVSS.n1038 DVSS.t237 90.7037
R27707 DVSS.n1284 DVSS.t252 90.7036
R27708 DVSS.n1825 DVSS.t140 90.703
R27709 DVSS.n5037 DVSS.t199 90.703
R27710 DVSS.n3442 DVSS.t12 90.703
R27711 DVSS.n6506 DVSS.t217 90.703
R27712 DVSS.n3413 DVSS.t9 89.25
R27713 DVSS.n5008 DVSS.t206 89.25
R27714 DVSS.n1796 DVSS.t135 89.25
R27715 DVSS.n3667 DVSS.n3666 87.6383
R27716 DVSS.n3669 DVSS.n3668 87.6383
R27717 DVSS.n3672 DVSS.n3654 87.6383
R27718 DVSS.n3666 DVSS.n3665 87.6383
R27719 DVSS.n3668 DVSS.n3667 87.6383
R27720 DVSS.n3669 DVSS.n3654 87.6383
R27721 DVSS.n4132 DVSS.n4131 87.6383
R27722 DVSS.n4134 DVSS.n4133 87.6383
R27723 DVSS.n4137 DVSS.n4119 87.6383
R27724 DVSS.n4131 DVSS.n4130 87.6383
R27725 DVSS.n4133 DVSS.n4132 87.6383
R27726 DVSS.n4134 DVSS.n4119 87.6383
R27727 DVSS.n2071 DVSS.n2070 87.6383
R27728 DVSS.n2073 DVSS.n2072 87.6383
R27729 DVSS.n2076 DVSS.n2058 87.6383
R27730 DVSS.n2070 DVSS.n2069 87.6383
R27731 DVSS.n2072 DVSS.n2071 87.6383
R27732 DVSS.n2073 DVSS.n2058 87.6383
R27733 DVSS.n2536 DVSS.n2535 87.6383
R27734 DVSS.n2538 DVSS.n2537 87.6383
R27735 DVSS.n2541 DVSS.n2523 87.6383
R27736 DVSS.n2535 DVSS.n2534 87.6383
R27737 DVSS.n2537 DVSS.n2536 87.6383
R27738 DVSS.n2538 DVSS.n2523 87.6383
R27739 DVSS.n5135 DVSS.n5134 87.6383
R27740 DVSS.n5137 DVSS.n5136 87.6383
R27741 DVSS.n5140 DVSS.n5122 87.6383
R27742 DVSS.n5134 DVSS.n5133 87.6383
R27743 DVSS.n5136 DVSS.n5135 87.6383
R27744 DVSS.n5137 DVSS.n5122 87.6383
R27745 DVSS.n5600 DVSS.n5599 87.6383
R27746 DVSS.n5602 DVSS.n5601 87.6383
R27747 DVSS.n5605 DVSS.n5587 87.6383
R27748 DVSS.n5599 DVSS.n5598 87.6383
R27749 DVSS.n5601 DVSS.n5600 87.6383
R27750 DVSS.n5602 DVSS.n5587 87.6383
R27751 DVSS.n70 DVSS.n69 87.6383
R27752 DVSS.n72 DVSS.n71 87.6383
R27753 DVSS.n75 DVSS.n57 87.6383
R27754 DVSS.n69 DVSS.n68 87.6383
R27755 DVSS.n71 DVSS.n70 87.6383
R27756 DVSS.n72 DVSS.n57 87.6383
R27757 DVSS.n535 DVSS.n534 87.6383
R27758 DVSS.n537 DVSS.n536 87.6383
R27759 DVSS.n540 DVSS.n522 87.6383
R27760 DVSS.n534 DVSS.n533 87.6383
R27761 DVSS.n536 DVSS.n535 87.6383
R27762 DVSS.n537 DVSS.n522 87.6383
R27763 DVSS.n3916 DVSS.n3762 87.3927
R27764 DVSS.n3905 DVSS.n3775 87.3927
R27765 DVSS.n4381 DVSS.n4227 87.3927
R27766 DVSS.n4370 DVSS.n4240 87.3927
R27767 DVSS.n2320 DVSS.n2166 87.3927
R27768 DVSS.n2309 DVSS.n2179 87.3927
R27769 DVSS.n2785 DVSS.n2631 87.3927
R27770 DVSS.n2774 DVSS.n2644 87.3927
R27771 DVSS.n5384 DVSS.n5230 87.3927
R27772 DVSS.n5373 DVSS.n5243 87.3927
R27773 DVSS.n5849 DVSS.n5695 87.3927
R27774 DVSS.n5838 DVSS.n5708 87.3927
R27775 DVSS.n319 DVSS.n165 87.3927
R27776 DVSS.n308 DVSS.n178 87.3927
R27777 DVSS.n784 DVSS.n630 87.3927
R27778 DVSS.n773 DVSS.n643 87.3927
R27779 DVSS.n6598 DVSS.n6597 85.7982
R27780 DVSS.n3586 DVSS.t71 84.7893
R27781 DVSS.n6564 DVSS.t228 84.7893
R27782 DVSS.n1983 DVSS.t191 84.6505
R27783 DVSS.n6776 DVSS.t116 84.6505
R27784 DVSS.n6203 DVSS.n6202 81.7659
R27785 DVSS.n6214 DVSS.n6212 81.7659
R27786 DVSS.n4735 DVSS.n4734 81.7659
R27787 DVSS.n4746 DVSS.n4744 81.7659
R27788 DVSS.n3139 DVSS.n3138 81.7659
R27789 DVSS.n3150 DVSS.n3148 81.7659
R27790 DVSS.n1522 DVSS.n1521 81.7659
R27791 DVSS.n1533 DVSS.n1531 81.7659
R27792 DVSS.n3825 DVSS.n3790 80.9725
R27793 DVSS.n4290 DVSS.n4255 80.9725
R27794 DVSS.n6024 DVSS.n6023 80.9725
R27795 DVSS.n4556 DVSS.n4555 80.9725
R27796 DVSS.n2229 DVSS.n2194 80.9725
R27797 DVSS.n2694 DVSS.n2659 80.9725
R27798 DVSS.n2960 DVSS.n2959 80.9725
R27799 DVSS.n5293 DVSS.n5258 80.9725
R27800 DVSS.n5758 DVSS.n5723 80.9725
R27801 DVSS.n228 DVSS.n193 80.9725
R27802 DVSS.n693 DVSS.n658 80.9725
R27803 DVSS.n959 DVSS.n958 80.9725
R27804 DVSS.n3826 DVSS.n3825 80.9721
R27805 DVSS.n4291 DVSS.n4290 80.9721
R27806 DVSS.n6030 DVSS.n6029 80.9721
R27807 DVSS.n4562 DVSS.n4561 80.9721
R27808 DVSS.n2230 DVSS.n2229 80.9721
R27809 DVSS.n2695 DVSS.n2694 80.9721
R27810 DVSS.n2966 DVSS.n2965 80.9721
R27811 DVSS.n5294 DVSS.n5293 80.9721
R27812 DVSS.n5759 DVSS.n5758 80.9721
R27813 DVSS.n229 DVSS.n228 80.9721
R27814 DVSS.n694 DVSS.n693 80.9721
R27815 DVSS.n1349 DVSS.n1348 80.9721
R27816 DVSS.n3835 DVSS.n3834 80.9719
R27817 DVSS.n3827 DVSS.n3822 80.9719
R27818 DVSS.n3859 DVSS.n3852 80.9719
R27819 DVSS.n3855 DVSS.n3851 80.9719
R27820 DVSS.n3871 DVSS.n3870 80.9719
R27821 DVSS.n3814 DVSS.n3813 80.9719
R27822 DVSS.n3821 DVSS.n3820 80.9719
R27823 DVSS.n3885 DVSS.n3793 80.9719
R27824 DVSS.n3862 DVSS.n3852 80.9719
R27825 DVSS.n3858 DVSS.n3851 80.9719
R27826 DVSS.n3870 DVSS.n3850 80.9719
R27827 DVSS.n3813 DVSS.n3812 80.9719
R27828 DVSS.n3836 DVSS.n3835 80.9719
R27829 DVSS.n3820 DVSS.n3819 80.9719
R27830 DVSS.n3822 DVSS.n3810 80.9719
R27831 DVSS.n3823 DVSS.n3793 80.9719
R27832 DVSS.n4045 DVSS.n4037 80.9719
R27833 DVSS.n4041 DVSS.n4036 80.9719
R27834 DVSS.n4070 DVSS.n3613 80.9719
R27835 DVSS.n4038 DVSS.n4037 80.9719
R27836 DVSS.n4044 DVSS.n4036 80.9719
R27837 DVSS.n4040 DVSS.n3613 80.9719
R27838 DVSS.n4300 DVSS.n4299 80.9719
R27839 DVSS.n4292 DVSS.n4287 80.9719
R27840 DVSS.n4324 DVSS.n4317 80.9719
R27841 DVSS.n4320 DVSS.n4316 80.9719
R27842 DVSS.n4336 DVSS.n4335 80.9719
R27843 DVSS.n4279 DVSS.n4278 80.9719
R27844 DVSS.n4286 DVSS.n4285 80.9719
R27845 DVSS.n4350 DVSS.n4258 80.9719
R27846 DVSS.n4327 DVSS.n4317 80.9719
R27847 DVSS.n4323 DVSS.n4316 80.9719
R27848 DVSS.n4335 DVSS.n4315 80.9719
R27849 DVSS.n4278 DVSS.n4277 80.9719
R27850 DVSS.n4301 DVSS.n4300 80.9719
R27851 DVSS.n4285 DVSS.n4284 80.9719
R27852 DVSS.n4287 DVSS.n4275 80.9719
R27853 DVSS.n4288 DVSS.n4258 80.9719
R27854 DVSS.n4510 DVSS.n4502 80.9719
R27855 DVSS.n4506 DVSS.n4501 80.9719
R27856 DVSS.n4534 DVSS.n4078 80.9719
R27857 DVSS.n4503 DVSS.n4502 80.9719
R27858 DVSS.n4509 DVSS.n4501 80.9719
R27859 DVSS.n4505 DVSS.n4078 80.9719
R27860 DVSS.n2239 DVSS.n2238 80.9719
R27861 DVSS.n2231 DVSS.n2226 80.9719
R27862 DVSS.n2263 DVSS.n2256 80.9719
R27863 DVSS.n2259 DVSS.n2255 80.9719
R27864 DVSS.n2275 DVSS.n2274 80.9719
R27865 DVSS.n2218 DVSS.n2217 80.9719
R27866 DVSS.n2225 DVSS.n2224 80.9719
R27867 DVSS.n2289 DVSS.n2197 80.9719
R27868 DVSS.n2266 DVSS.n2256 80.9719
R27869 DVSS.n2262 DVSS.n2255 80.9719
R27870 DVSS.n2274 DVSS.n2254 80.9719
R27871 DVSS.n2217 DVSS.n2216 80.9719
R27872 DVSS.n2240 DVSS.n2239 80.9719
R27873 DVSS.n2224 DVSS.n2223 80.9719
R27874 DVSS.n2226 DVSS.n2214 80.9719
R27875 DVSS.n2227 DVSS.n2197 80.9719
R27876 DVSS.n2449 DVSS.n2441 80.9719
R27877 DVSS.n2445 DVSS.n2440 80.9719
R27878 DVSS.n2474 DVSS.n2017 80.9719
R27879 DVSS.n2442 DVSS.n2441 80.9719
R27880 DVSS.n2448 DVSS.n2440 80.9719
R27881 DVSS.n2444 DVSS.n2017 80.9719
R27882 DVSS.n2704 DVSS.n2703 80.9719
R27883 DVSS.n2696 DVSS.n2691 80.9719
R27884 DVSS.n2728 DVSS.n2721 80.9719
R27885 DVSS.n2724 DVSS.n2720 80.9719
R27886 DVSS.n2740 DVSS.n2739 80.9719
R27887 DVSS.n2683 DVSS.n2682 80.9719
R27888 DVSS.n2690 DVSS.n2689 80.9719
R27889 DVSS.n2754 DVSS.n2662 80.9719
R27890 DVSS.n2731 DVSS.n2721 80.9719
R27891 DVSS.n2727 DVSS.n2720 80.9719
R27892 DVSS.n2739 DVSS.n2719 80.9719
R27893 DVSS.n2682 DVSS.n2681 80.9719
R27894 DVSS.n2705 DVSS.n2704 80.9719
R27895 DVSS.n2689 DVSS.n2688 80.9719
R27896 DVSS.n2691 DVSS.n2679 80.9719
R27897 DVSS.n2692 DVSS.n2662 80.9719
R27898 DVSS.n2914 DVSS.n2906 80.9719
R27899 DVSS.n2910 DVSS.n2905 80.9719
R27900 DVSS.n2938 DVSS.n2482 80.9719
R27901 DVSS.n2907 DVSS.n2906 80.9719
R27902 DVSS.n2913 DVSS.n2905 80.9719
R27903 DVSS.n2909 DVSS.n2482 80.9719
R27904 DVSS.n5303 DVSS.n5302 80.9719
R27905 DVSS.n5295 DVSS.n5290 80.9719
R27906 DVSS.n5327 DVSS.n5320 80.9719
R27907 DVSS.n5323 DVSS.n5319 80.9719
R27908 DVSS.n5339 DVSS.n5338 80.9719
R27909 DVSS.n5282 DVSS.n5281 80.9719
R27910 DVSS.n5289 DVSS.n5288 80.9719
R27911 DVSS.n5353 DVSS.n5261 80.9719
R27912 DVSS.n5330 DVSS.n5320 80.9719
R27913 DVSS.n5326 DVSS.n5319 80.9719
R27914 DVSS.n5338 DVSS.n5318 80.9719
R27915 DVSS.n5281 DVSS.n5280 80.9719
R27916 DVSS.n5304 DVSS.n5303 80.9719
R27917 DVSS.n5288 DVSS.n5287 80.9719
R27918 DVSS.n5290 DVSS.n5278 80.9719
R27919 DVSS.n5291 DVSS.n5261 80.9719
R27920 DVSS.n5513 DVSS.n5505 80.9719
R27921 DVSS.n5509 DVSS.n5504 80.9719
R27922 DVSS.n5538 DVSS.n5081 80.9719
R27923 DVSS.n5506 DVSS.n5505 80.9719
R27924 DVSS.n5512 DVSS.n5504 80.9719
R27925 DVSS.n5508 DVSS.n5081 80.9719
R27926 DVSS.n5768 DVSS.n5767 80.9719
R27927 DVSS.n5760 DVSS.n5755 80.9719
R27928 DVSS.n5792 DVSS.n5785 80.9719
R27929 DVSS.n5788 DVSS.n5784 80.9719
R27930 DVSS.n5804 DVSS.n5803 80.9719
R27931 DVSS.n5747 DVSS.n5746 80.9719
R27932 DVSS.n5754 DVSS.n5753 80.9719
R27933 DVSS.n5818 DVSS.n5726 80.9719
R27934 DVSS.n5795 DVSS.n5785 80.9719
R27935 DVSS.n5791 DVSS.n5784 80.9719
R27936 DVSS.n5803 DVSS.n5783 80.9719
R27937 DVSS.n5746 DVSS.n5745 80.9719
R27938 DVSS.n5769 DVSS.n5768 80.9719
R27939 DVSS.n5753 DVSS.n5752 80.9719
R27940 DVSS.n5755 DVSS.n5743 80.9719
R27941 DVSS.n5756 DVSS.n5726 80.9719
R27942 DVSS.n5978 DVSS.n5970 80.9719
R27943 DVSS.n5974 DVSS.n5969 80.9719
R27944 DVSS.n6002 DVSS.n5546 80.9719
R27945 DVSS.n5971 DVSS.n5970 80.9719
R27946 DVSS.n5977 DVSS.n5969 80.9719
R27947 DVSS.n5973 DVSS.n5546 80.9719
R27948 DVSS.n238 DVSS.n237 80.9719
R27949 DVSS.n230 DVSS.n225 80.9719
R27950 DVSS.n262 DVSS.n255 80.9719
R27951 DVSS.n258 DVSS.n254 80.9719
R27952 DVSS.n274 DVSS.n273 80.9719
R27953 DVSS.n217 DVSS.n216 80.9719
R27954 DVSS.n224 DVSS.n223 80.9719
R27955 DVSS.n288 DVSS.n196 80.9719
R27956 DVSS.n265 DVSS.n255 80.9719
R27957 DVSS.n261 DVSS.n254 80.9719
R27958 DVSS.n273 DVSS.n253 80.9719
R27959 DVSS.n216 DVSS.n215 80.9719
R27960 DVSS.n239 DVSS.n238 80.9719
R27961 DVSS.n223 DVSS.n222 80.9719
R27962 DVSS.n225 DVSS.n213 80.9719
R27963 DVSS.n226 DVSS.n196 80.9719
R27964 DVSS.n448 DVSS.n440 80.9719
R27965 DVSS.n444 DVSS.n439 80.9719
R27966 DVSS.n473 DVSS.n16 80.9719
R27967 DVSS.n441 DVSS.n440 80.9719
R27968 DVSS.n447 DVSS.n439 80.9719
R27969 DVSS.n443 DVSS.n16 80.9719
R27970 DVSS.n703 DVSS.n702 80.9719
R27971 DVSS.n695 DVSS.n690 80.9719
R27972 DVSS.n727 DVSS.n720 80.9719
R27973 DVSS.n723 DVSS.n719 80.9719
R27974 DVSS.n739 DVSS.n738 80.9719
R27975 DVSS.n682 DVSS.n681 80.9719
R27976 DVSS.n689 DVSS.n688 80.9719
R27977 DVSS.n753 DVSS.n661 80.9719
R27978 DVSS.n730 DVSS.n720 80.9719
R27979 DVSS.n726 DVSS.n719 80.9719
R27980 DVSS.n738 DVSS.n718 80.9719
R27981 DVSS.n681 DVSS.n680 80.9719
R27982 DVSS.n704 DVSS.n703 80.9719
R27983 DVSS.n688 DVSS.n687 80.9719
R27984 DVSS.n690 DVSS.n678 80.9719
R27985 DVSS.n691 DVSS.n661 80.9719
R27986 DVSS.n913 DVSS.n905 80.9719
R27987 DVSS.n909 DVSS.n904 80.9719
R27988 DVSS.n937 DVSS.n481 80.9719
R27989 DVSS.n906 DVSS.n905 80.9719
R27990 DVSS.n912 DVSS.n904 80.9719
R27991 DVSS.n908 DVSS.n481 80.9719
R27992 DVSS.n3559 DVSS.n3558 78.5406
R27993 DVSS.n1956 DVSS.n1955 78.4133
R27994 DVSS.n6804 DVSS.n6803 78.4133
R27995 DVSS.n6651 DVSS.n6650 77.5733
R27996 DVSS.n6591 DVSS.t103 77.5733
R27997 DVSS.n1893 DVSS.n1892 77.4463
R27998 DVSS.n3559 DVSS.t43 76.7556
R27999 DVSS.n6073 DVSS.n6070 76.6556
R28000 DVSS.n6099 DVSS.n6098 76.6556
R28001 DVSS.n6323 DVSS.n6320 76.6556
R28002 DVSS.n6349 DVSS.n6348 76.6556
R28003 DVSS.n4605 DVSS.n4602 76.6556
R28004 DVSS.n4631 DVSS.n4630 76.6556
R28005 DVSS.n4855 DVSS.n4852 76.6556
R28006 DVSS.n4881 DVSS.n4880 76.6556
R28007 DVSS.n3009 DVSS.n3006 76.6556
R28008 DVSS.n3035 DVSS.n3034 76.6556
R28009 DVSS.n3259 DVSS.n3256 76.6556
R28010 DVSS.n3285 DVSS.n3284 76.6556
R28011 DVSS.n1392 DVSS.n1389 76.6556
R28012 DVSS.n1418 DVSS.n1417 76.6556
R28013 DVSS.n1642 DVSS.n1639 76.6556
R28014 DVSS.n1668 DVSS.n1667 76.6556
R28015 DVSS.n1956 DVSS.t179 76.6312
R28016 DVSS.n6804 DVSS.t33 76.6312
R28017 DVSS.n1716 DVSS.n1714 76.424
R28018 DVSS.n955 DVSS.n953 76.424
R28019 DVSS.n4929 DVSS.n4927 76.424
R28020 DVSS.n4552 DVSS.n4550 76.424
R28021 DVSS.n6397 DVSS.n6395 76.424
R28022 DVSS.n6020 DVSS.n6018 76.424
R28023 DVSS.n3333 DVSS.n3331 76.424
R28024 DVSS.n2956 DVSS.n2954 76.424
R28025 DVSS.n1228 DVSS.n1227 76.4173
R28026 DVSS.n3661 DVSS.n3660 76.2208
R28027 DVSS.n4126 DVSS.n4125 76.2208
R28028 DVSS.n2065 DVSS.n2064 76.2208
R28029 DVSS.n2530 DVSS.n2529 76.2208
R28030 DVSS.n5129 DVSS.n5128 76.2208
R28031 DVSS.n5594 DVSS.n5593 76.2208
R28032 DVSS.n64 DVSS.n63 76.2208
R28033 DVSS.n529 DVSS.n528 76.2208
R28034 DVSS.n3660 DVSS.n3659 76.2204
R28035 DVSS.n4125 DVSS.n4124 76.2204
R28036 DVSS.n2064 DVSS.n2063 76.2204
R28037 DVSS.n2529 DVSS.n2528 76.2204
R28038 DVSS.n5128 DVSS.n5127 76.2204
R28039 DVSS.n5593 DVSS.n5592 76.2204
R28040 DVSS.n63 DVSS.n62 76.2204
R28041 DVSS.n528 DVSS.n527 76.2204
R28042 DVSS.n4006 DVSS.n4004 76.2201
R28043 DVSS.n4013 DVSS.n4012 76.2201
R28044 DVSS.n4017 DVSS.n4002 76.2201
R28045 DVSS.n4020 DVSS.n4019 76.2201
R28046 DVSS.n4007 DVSS.n4006 76.2201
R28047 DVSS.n4012 DVSS.n4011 76.2201
R28048 DVSS.n4014 DVSS.n4002 76.2201
R28049 DVSS.n4019 DVSS.n4018 76.2201
R28050 DVSS.n4471 DVSS.n4469 76.2201
R28051 DVSS.n4478 DVSS.n4477 76.2201
R28052 DVSS.n4482 DVSS.n4467 76.2201
R28053 DVSS.n4485 DVSS.n4484 76.2201
R28054 DVSS.n4472 DVSS.n4471 76.2201
R28055 DVSS.n4477 DVSS.n4476 76.2201
R28056 DVSS.n4479 DVSS.n4467 76.2201
R28057 DVSS.n4484 DVSS.n4483 76.2201
R28058 DVSS.n2410 DVSS.n2408 76.2201
R28059 DVSS.n2417 DVSS.n2416 76.2201
R28060 DVSS.n2421 DVSS.n2406 76.2201
R28061 DVSS.n2424 DVSS.n2423 76.2201
R28062 DVSS.n2411 DVSS.n2410 76.2201
R28063 DVSS.n2416 DVSS.n2415 76.2201
R28064 DVSS.n2418 DVSS.n2406 76.2201
R28065 DVSS.n2423 DVSS.n2422 76.2201
R28066 DVSS.n2875 DVSS.n2873 76.2201
R28067 DVSS.n2882 DVSS.n2881 76.2201
R28068 DVSS.n2886 DVSS.n2871 76.2201
R28069 DVSS.n2889 DVSS.n2888 76.2201
R28070 DVSS.n2876 DVSS.n2875 76.2201
R28071 DVSS.n2881 DVSS.n2880 76.2201
R28072 DVSS.n2883 DVSS.n2871 76.2201
R28073 DVSS.n2888 DVSS.n2887 76.2201
R28074 DVSS.n5474 DVSS.n5472 76.2201
R28075 DVSS.n5481 DVSS.n5480 76.2201
R28076 DVSS.n5485 DVSS.n5470 76.2201
R28077 DVSS.n5488 DVSS.n5487 76.2201
R28078 DVSS.n5475 DVSS.n5474 76.2201
R28079 DVSS.n5480 DVSS.n5479 76.2201
R28080 DVSS.n5482 DVSS.n5470 76.2201
R28081 DVSS.n5487 DVSS.n5486 76.2201
R28082 DVSS.n5939 DVSS.n5937 76.2201
R28083 DVSS.n5946 DVSS.n5945 76.2201
R28084 DVSS.n5950 DVSS.n5935 76.2201
R28085 DVSS.n5953 DVSS.n5952 76.2201
R28086 DVSS.n5940 DVSS.n5939 76.2201
R28087 DVSS.n5945 DVSS.n5944 76.2201
R28088 DVSS.n5947 DVSS.n5935 76.2201
R28089 DVSS.n5952 DVSS.n5951 76.2201
R28090 DVSS.n409 DVSS.n407 76.2201
R28091 DVSS.n416 DVSS.n415 76.2201
R28092 DVSS.n420 DVSS.n405 76.2201
R28093 DVSS.n423 DVSS.n422 76.2201
R28094 DVSS.n410 DVSS.n409 76.2201
R28095 DVSS.n415 DVSS.n414 76.2201
R28096 DVSS.n417 DVSS.n405 76.2201
R28097 DVSS.n422 DVSS.n421 76.2201
R28098 DVSS.n874 DVSS.n872 76.2201
R28099 DVSS.n881 DVSS.n880 76.2201
R28100 DVSS.n885 DVSS.n870 76.2201
R28101 DVSS.n888 DVSS.n887 76.2201
R28102 DVSS.n875 DVSS.n874 76.2201
R28103 DVSS.n880 DVSS.n879 76.2201
R28104 DVSS.n882 DVSS.n870 76.2201
R28105 DVSS.n887 DVSS.n886 76.2201
R28106 DVSS.n6188 DVSS.n6187 71.5452
R28107 DVSS.n6229 DVSS.n6227 71.5452
R28108 DVSS.n4720 DVSS.n4719 71.5452
R28109 DVSS.n4761 DVSS.n4759 71.5452
R28110 DVSS.n3124 DVSS.n3123 71.5452
R28111 DVSS.n3165 DVSS.n3163 71.5452
R28112 DVSS.n1507 DVSS.n1506 71.5452
R28113 DVSS.n1548 DVSS.n1546 71.5452
R28114 DVSS.t154 DVSS.t260 71.5276
R28115 DVSS.n3430 DVSS.t13 70.0806
R28116 DVSS.n5025 DVSS.t200 70.0806
R28117 DVSS.n1813 DVSS.t143 70.0806
R28118 DVSS.n6493 DVSS.t214 70.0801
R28119 DVSS.t216 DVSS.n6501 70.0801
R28120 DVSS.n1262 DVSS.n1260 69.3226
R28121 DVSS.n6783 DVSS.n6781 69.3226
R28122 DVSS.n3583 DVSS.n3581 69.3226
R28123 DVSS.n6571 DVSS.n6569 69.3226
R28124 DVSS.n1980 DVSS.n1978 69.3226
R28125 DVSS.n1062 DVSS.t160 69.0146
R28126 DVSS.n3748 DVSS.t186 66.8281
R28127 DVSS.n3727 DVSS.t82 66.8281
R28128 DVSS.n4213 DVSS.t119 66.8281
R28129 DVSS.n4192 DVSS.t85 66.8281
R28130 DVSS.n2152 DVSS.t224 66.8281
R28131 DVSS.n2131 DVSS.t125 66.8281
R28132 DVSS.n2617 DVSS.t62 66.8281
R28133 DVSS.n2596 DVSS.t121 66.8281
R28134 DVSS.n5216 DVSS.t92 66.8281
R28135 DVSS.n5195 DVSS.t80 66.8281
R28136 DVSS.n5681 DVSS.t152 66.8281
R28137 DVSS.n5660 DVSS.t77 66.8281
R28138 DVSS.n151 DVSS.t188 66.8281
R28139 DVSS.n130 DVSS.t113 66.8281
R28140 DVSS.n616 DVSS.t231 66.8281
R28141 DVSS.n595 DVSS.t110 66.8281
R28142 DVSS.n3577 DVSS.t202 66.7492
R28143 DVSS.n6573 DVSS.t212 66.7492
R28144 DVSS.n1974 DVSS.t17 66.6399
R28145 DVSS.n6785 DVSS.t133 66.6399
R28146 DVSS.n6055 DVSS.n6054 66.4349
R28147 DVSS.n6114 DVSS.n6113 66.4349
R28148 DVSS.n6305 DVSS.n6304 66.4349
R28149 DVSS.n6364 DVSS.n6363 66.4349
R28150 DVSS.n4587 DVSS.n4586 66.4349
R28151 DVSS.n4646 DVSS.n4645 66.4349
R28152 DVSS.n4837 DVSS.n4836 66.4349
R28153 DVSS.n4896 DVSS.n4895 66.4349
R28154 DVSS.n2991 DVSS.n2990 66.4349
R28155 DVSS.n3050 DVSS.n3049 66.4349
R28156 DVSS.n3241 DVSS.n3240 66.4349
R28157 DVSS.n3300 DVSS.n3299 66.4349
R28158 DVSS.n1374 DVSS.n1373 66.4349
R28159 DVSS.n1433 DVSS.n1432 66.4349
R28160 DVSS.n1624 DVSS.n1623 66.4349
R28161 DVSS.n1683 DVSS.n1682 66.4349
R28162 DVSS.n6682 DVSS.t127 65.1095
R28163 DVSS.n1886 DVSS.t89 64.9073
R28164 DVSS.n6173 DVSS.n6172 61.3245
R28165 DVSS.n6244 DVSS.n6242 61.3245
R28166 DVSS.n4705 DVSS.n4704 61.3245
R28167 DVSS.n4776 DVSS.n4774 61.3245
R28168 DVSS.n3109 DVSS.n3108 61.3245
R28169 DVSS.n3180 DVSS.n3178 61.3245
R28170 DVSS.n1492 DVSS.n1491 61.3245
R28171 DVSS.n1563 DVSS.n1561 61.3245
R28172 DVSS.n3939 DVSS.n3938 59.4692
R28173 DVSS.n4404 DVSS.n4403 59.4692
R28174 DVSS.n6410 DVSS.n6409 59.4692
R28175 DVSS.n4942 DVSS.n4941 59.4692
R28176 DVSS.n2343 DVSS.n2342 59.4692
R28177 DVSS.n2808 DVSS.n2807 59.4692
R28178 DVSS.n3347 DVSS.n3346 59.4692
R28179 DVSS.n5407 DVSS.n5406 59.4692
R28180 DVSS.n5872 DVSS.n5871 59.4692
R28181 DVSS.n342 DVSS.n341 59.4692
R28182 DVSS.n807 DVSS.n806 59.4692
R28183 DVSS.n1729 DVSS.n1728 59.4692
R28184 DVSS.n1718 DVSS.n1717 59.4689
R28185 DVSS.n4931 DVSS.n4930 59.4689
R28186 DVSS.n3806 DVSS.n3787 59.4689
R28187 DVSS.n3837 DVSS.n3808 59.4689
R28188 DVSS.n3919 DVSS.n3764 59.4689
R28189 DVSS.n3868 DVSS.n3867 59.4689
R28190 DVSS.n3863 DVSS.n3853 59.4689
R28191 DVSS.n3844 DVSS.n3798 59.4689
R28192 DVSS.n3804 DVSS.n3803 59.4689
R28193 DVSS.n3697 DVSS.n3690 59.4689
R28194 DVSS.n3691 DVSS.n3689 59.4689
R28195 DVSS.n4053 DVSS.n4052 59.4689
R28196 DVSS.n4050 DVSS.n4049 59.4689
R28197 DVSS.n4271 DVSS.n4252 59.4689
R28198 DVSS.n4302 DVSS.n4273 59.4689
R28199 DVSS.n4384 DVSS.n4229 59.4689
R28200 DVSS.n4333 DVSS.n4332 59.4689
R28201 DVSS.n4328 DVSS.n4318 59.4689
R28202 DVSS.n4309 DVSS.n4263 59.4689
R28203 DVSS.n4269 DVSS.n4268 59.4689
R28204 DVSS.n4162 DVSS.n4155 59.4689
R28205 DVSS.n4156 DVSS.n4154 59.4689
R28206 DVSS.n4518 DVSS.n4517 59.4689
R28207 DVSS.n4515 DVSS.n4514 59.4689
R28208 DVSS.n6399 DVSS.n6398 59.4689
R28209 DVSS.n3335 DVSS.n3334 59.4689
R28210 DVSS.n2210 DVSS.n2191 59.4689
R28211 DVSS.n2241 DVSS.n2212 59.4689
R28212 DVSS.n2323 DVSS.n2168 59.4689
R28213 DVSS.n2272 DVSS.n2271 59.4689
R28214 DVSS.n2267 DVSS.n2257 59.4689
R28215 DVSS.n2248 DVSS.n2202 59.4689
R28216 DVSS.n2208 DVSS.n2207 59.4689
R28217 DVSS.n2101 DVSS.n2094 59.4689
R28218 DVSS.n2095 DVSS.n2093 59.4689
R28219 DVSS.n2457 DVSS.n2456 59.4689
R28220 DVSS.n2454 DVSS.n2453 59.4689
R28221 DVSS.n2675 DVSS.n2656 59.4689
R28222 DVSS.n2706 DVSS.n2677 59.4689
R28223 DVSS.n2788 DVSS.n2633 59.4689
R28224 DVSS.n2737 DVSS.n2736 59.4689
R28225 DVSS.n2732 DVSS.n2722 59.4689
R28226 DVSS.n2713 DVSS.n2667 59.4689
R28227 DVSS.n2673 DVSS.n2672 59.4689
R28228 DVSS.n2566 DVSS.n2559 59.4689
R28229 DVSS.n2560 DVSS.n2558 59.4689
R28230 DVSS.n2922 DVSS.n2921 59.4689
R28231 DVSS.n2919 DVSS.n2918 59.4689
R28232 DVSS.n5274 DVSS.n5255 59.4689
R28233 DVSS.n5305 DVSS.n5276 59.4689
R28234 DVSS.n5387 DVSS.n5232 59.4689
R28235 DVSS.n5336 DVSS.n5335 59.4689
R28236 DVSS.n5331 DVSS.n5321 59.4689
R28237 DVSS.n5312 DVSS.n5266 59.4689
R28238 DVSS.n5272 DVSS.n5271 59.4689
R28239 DVSS.n5165 DVSS.n5158 59.4689
R28240 DVSS.n5159 DVSS.n5157 59.4689
R28241 DVSS.n5521 DVSS.n5520 59.4689
R28242 DVSS.n5518 DVSS.n5517 59.4689
R28243 DVSS.n5739 DVSS.n5720 59.4689
R28244 DVSS.n5770 DVSS.n5741 59.4689
R28245 DVSS.n5852 DVSS.n5697 59.4689
R28246 DVSS.n5801 DVSS.n5800 59.4689
R28247 DVSS.n5796 DVSS.n5786 59.4689
R28248 DVSS.n5777 DVSS.n5731 59.4689
R28249 DVSS.n5737 DVSS.n5736 59.4689
R28250 DVSS.n5630 DVSS.n5623 59.4689
R28251 DVSS.n5624 DVSS.n5622 59.4689
R28252 DVSS.n5986 DVSS.n5985 59.4689
R28253 DVSS.n5983 DVSS.n5982 59.4689
R28254 DVSS.n209 DVSS.n190 59.4689
R28255 DVSS.n240 DVSS.n211 59.4689
R28256 DVSS.n322 DVSS.n167 59.4689
R28257 DVSS.n271 DVSS.n270 59.4689
R28258 DVSS.n266 DVSS.n256 59.4689
R28259 DVSS.n247 DVSS.n201 59.4689
R28260 DVSS.n207 DVSS.n206 59.4689
R28261 DVSS.n100 DVSS.n93 59.4689
R28262 DVSS.n94 DVSS.n92 59.4689
R28263 DVSS.n456 DVSS.n455 59.4689
R28264 DVSS.n453 DVSS.n452 59.4689
R28265 DVSS.n674 DVSS.n655 59.4689
R28266 DVSS.n705 DVSS.n676 59.4689
R28267 DVSS.n787 DVSS.n632 59.4689
R28268 DVSS.n736 DVSS.n735 59.4689
R28269 DVSS.n731 DVSS.n721 59.4689
R28270 DVSS.n712 DVSS.n666 59.4689
R28271 DVSS.n672 DVSS.n671 59.4689
R28272 DVSS.n565 DVSS.n558 59.4689
R28273 DVSS.n559 DVSS.n557 59.4689
R28274 DVSS.n921 DVSS.n920 59.4689
R28275 DVSS.n918 DVSS.n917 59.4689
R28276 DVSS.n1159 DVSS.n1158 59.3519
R28277 DVSS.n1064 DVSS.n1063 59.3519
R28278 DVSS.n6673 DVSS.t194 58.256
R28279 DVSS.n1877 DVSS.t226 58.075
R28280 DVSS.n1731 DVSS.n1730 57.6005
R28281 DVSS.n1351 DVSS.n1350 57.6005
R28282 DVSS.n4944 DVSS.n4943 57.6005
R28283 DVSS.n4564 DVSS.n4563 57.6005
R28284 DVSS.n6412 DVSS.n6411 57.6005
R28285 DVSS.n6032 DVSS.n6031 57.6005
R28286 DVSS.n3349 DVSS.n3348 57.6005
R28287 DVSS.n2968 DVSS.n2967 57.6005
R28288 DVSS.n3431 DVSS.n3430 56.5671
R28289 DVSS.n5026 DVSS.n5025 56.5671
R28290 DVSS.n1814 DVSS.n1813 56.5671
R28291 DVSS.n6040 DVSS.n6039 56.2142
R28292 DVSS.n6129 DVSS.n6128 56.2142
R28293 DVSS.n6290 DVSS.n6289 56.2142
R28294 DVSS.n6379 DVSS.n6378 56.2142
R28295 DVSS.n4572 DVSS.n4571 56.2142
R28296 DVSS.n4661 DVSS.n4660 56.2142
R28297 DVSS.n4822 DVSS.n4821 56.2142
R28298 DVSS.n4911 DVSS.n4910 56.2142
R28299 DVSS.n2976 DVSS.n2975 56.2142
R28300 DVSS.n3065 DVSS.n3064 56.2142
R28301 DVSS.n3226 DVSS.n3225 56.2142
R28302 DVSS.n3315 DVSS.n3314 56.2142
R28303 DVSS.n1359 DVSS.n1358 56.2142
R28304 DVSS.n1448 DVSS.n1447 56.2142
R28305 DVSS.n1609 DVSS.n1608 56.2142
R28306 DVSS.n1698 DVSS.n1697 56.2142
R28307 DVSS.n3531 DVSS.t41 55.9251
R28308 DVSS.n6619 DVSS.t105 55.9251
R28309 DVSS.n1928 DVSS.t177 55.8335
R28310 DVSS.n6830 DVSS.t27 55.8335
R28311 DVSS.n3662 DVSS.n3656 55.6474
R28312 DVSS.n4127 DVSS.n4121 55.6474
R28313 DVSS.n2066 DVSS.n2060 55.6474
R28314 DVSS.n2531 DVSS.n2525 55.6474
R28315 DVSS.n5130 DVSS.n5124 55.6474
R28316 DVSS.n5595 DVSS.n5589 55.6474
R28317 DVSS.n65 DVSS.n59 55.6474
R28318 DVSS.n530 DVSS.n524 55.6474
R28319 DVSS.n3674 DVSS.n3673 55.6471
R28320 DVSS.n4139 DVSS.n4138 55.6471
R28321 DVSS.n2078 DVSS.n2077 55.6471
R28322 DVSS.n2543 DVSS.n2542 55.6471
R28323 DVSS.n5142 DVSS.n5141 55.6471
R28324 DVSS.n5607 DVSS.n5606 55.6471
R28325 DVSS.n77 DVSS.n76 55.6471
R28326 DVSS.n542 DVSS.n541 55.6471
R28327 DVSS.t218 DVSS.n6463 55.0631
R28328 DVSS.n1519 DVSS.n1518 52.6902
R28329 DVSS.n1530 DVSS.n1529 52.6902
R28330 DVSS.n4732 DVSS.n4731 52.6902
R28331 DVSS.n4743 DVSS.n4742 52.6902
R28332 DVSS.n6200 DVSS.n6199 52.6902
R28333 DVSS.n6211 DVSS.n6210 52.6902
R28334 DVSS.n3136 DVSS.n3135 52.6902
R28335 DVSS.n3147 DVSS.n3146 52.6902
R28336 DVSS.n3535 DVSS.t45 52.317
R28337 DVSS.n6615 DVSS.t97 52.317
R28338 DVSS.n971 DVSS.n970 52.3069
R28339 DVSS.n1753 DVSS.n1752 52.3069
R28340 DVSS.n4965 DVSS.n4964 52.3069
R28341 DVSS.n3370 DVSS.n3369 52.3069
R28342 DVSS.n6433 DVSS.n6432 52.3069
R28343 DVSS.n1932 DVSS.t181 52.2314
R28344 DVSS.n6826 DVSS.t29 52.2314
R28345 DVSS.n6158 DVSS.n6157 51.1039
R28346 DVSS.n6259 DVSS.n6257 51.1039
R28347 DVSS.n4690 DVSS.n4689 51.1039
R28348 DVSS.n4791 DVSS.n4789 51.1039
R28349 DVSS.n3094 DVSS.n3093 51.1039
R28350 DVSS.n3195 DVSS.n3193 51.1039
R28351 DVSS.n1477 DVSS.n1476 51.1039
R28352 DVSS.n1578 DVSS.n1576 51.1039
R28353 DVSS.n6550 DVSS.n6549 50.513
R28354 DVSS.n6476 DVSS.t220 50.0574
R28355 DVSS.n1393 DVSS.n1385 49.397
R28356 DVSS.n1419 DVSS.n1412 49.397
R28357 DVSS.n1643 DVSS.n1635 49.397
R28358 DVSS.n1669 DVSS.n1662 49.397
R28359 DVSS.n4606 DVSS.n4598 49.397
R28360 DVSS.n4632 DVSS.n4625 49.397
R28361 DVSS.n4856 DVSS.n4848 49.397
R28362 DVSS.n4882 DVSS.n4875 49.397
R28363 DVSS.n6074 DVSS.n6066 49.397
R28364 DVSS.n6100 DVSS.n6093 49.397
R28365 DVSS.n6324 DVSS.n6316 49.397
R28366 DVSS.n6350 DVSS.n6343 49.397
R28367 DVSS.n3010 DVSS.n3002 49.397
R28368 DVSS.n3036 DVSS.n3029 49.397
R28369 DVSS.n3260 DVSS.n3252 49.397
R28370 DVSS.n3286 DVSS.n3279 49.397
R28371 DVSS.n4946 DVSS.t244 47.1806
R28372 DVSS.n6414 DVSS.t58 47.1806
R28373 DVSS.n3351 DVSS.t190 47.1806
R28374 DVSS.n1733 DVSS.t197 47.1519
R28375 DVSS.n1504 DVSS.n1503 46.104
R28376 DVSS.n1545 DVSS.n1544 46.104
R28377 DVSS.n4717 DVSS.n4716 46.104
R28378 DVSS.n4758 DVSS.n4757 46.104
R28379 DVSS.n6185 DVSS.n6184 46.104
R28380 DVSS.n6226 DVSS.n6225 46.104
R28381 DVSS.n3121 DVSS.n3120 46.104
R28382 DVSS.n3162 DVSS.n3161 46.104
R28383 DVSS.n6144 DVSS.n6143 45.9935
R28384 DVSS.n6275 DVSS.n6274 45.9935
R28385 DVSS.n4676 DVSS.n4675 45.9935
R28386 DVSS.n4807 DVSS.n4806 45.9935
R28387 DVSS.n3080 DVSS.n3079 45.9935
R28388 DVSS.n3211 DVSS.n3210 45.9935
R28389 DVSS.n1463 DVSS.n1462 45.9935
R28390 DVSS.n1594 DVSS.n1593 45.9935
R28391 DVSS.n3866 DVSS.n3845 45.5782
R28392 DVSS.n3873 DVSS.n3872 45.5782
R28393 DVSS.n4331 DVSS.n4310 45.5782
R28394 DVSS.n4338 DVSS.n4337 45.5782
R28395 DVSS.n2270 DVSS.n2249 45.5782
R28396 DVSS.n2277 DVSS.n2276 45.5782
R28397 DVSS.n2735 DVSS.n2714 45.5782
R28398 DVSS.n2742 DVSS.n2741 45.5782
R28399 DVSS.n5334 DVSS.n5313 45.5782
R28400 DVSS.n5341 DVSS.n5340 45.5782
R28401 DVSS.n5799 DVSS.n5778 45.5782
R28402 DVSS.n5806 DVSS.n5805 45.5782
R28403 DVSS.n269 DVSS.n248 45.5782
R28404 DVSS.n276 DVSS.n275 45.5782
R28405 DVSS.n734 DVSS.n713 45.5782
R28406 DVSS.n741 DVSS.n740 45.5782
R28407 DVSS.n1078 DVSS.n1077 43.8838
R28408 DVSS.n1375 DVSS.n1370 42.8108
R28409 DVSS.n1434 DVSS.n1429 42.8108
R28410 DVSS.n1625 DVSS.n1620 42.8108
R28411 DVSS.n1684 DVSS.n1679 42.8108
R28412 DVSS.n4588 DVSS.n4583 42.8108
R28413 DVSS.n4647 DVSS.n4642 42.8108
R28414 DVSS.n4838 DVSS.n4833 42.8108
R28415 DVSS.n4897 DVSS.n4892 42.8108
R28416 DVSS.n6056 DVSS.n6051 42.8108
R28417 DVSS.n6115 DVSS.n6110 42.8108
R28418 DVSS.n6306 DVSS.n6301 42.8108
R28419 DVSS.n6365 DVSS.n6360 42.8108
R28420 DVSS.n2992 DVSS.n2987 42.8108
R28421 DVSS.n3051 DVSS.n3046 42.8108
R28422 DVSS.n3242 DVSS.n3237 42.8108
R28423 DVSS.n3301 DVSS.n3296 42.8108
R28424 DVSS.n3911 DVSS.n3910 42.4097
R28425 DVSS.n4376 DVSS.n4375 42.4097
R28426 DVSS.n2315 DVSS.n2314 42.4097
R28427 DVSS.n2780 DVSS.n2779 42.4097
R28428 DVSS.n5379 DVSS.n5378 42.4097
R28429 DVSS.n5844 DVSS.n5843 42.4097
R28430 DVSS.n314 DVSS.n313 42.4097
R28431 DVSS.n779 DVSS.n778 42.4097
R28432 DVSS.n6143 DVSS.n6142 40.8832
R28433 DVSS.n6274 DVSS.n6272 40.8832
R28434 DVSS.n4675 DVSS.n4674 40.8832
R28435 DVSS.n4806 DVSS.n4804 40.8832
R28436 DVSS.n3079 DVSS.n3078 40.8832
R28437 DVSS.n3210 DVSS.n3208 40.8832
R28438 DVSS.n1462 DVSS.n1461 40.8832
R28439 DVSS.n1593 DVSS.n1591 40.8832
R28440 DVSS.n1489 DVSS.n1488 39.5177
R28441 DVSS.n1560 DVSS.n1559 39.5177
R28442 DVSS.n4702 DVSS.n4701 39.5177
R28443 DVSS.n4773 DVSS.n4772 39.5177
R28444 DVSS.n6170 DVSS.n6169 39.5177
R28445 DVSS.n6241 DVSS.n6240 39.5177
R28446 DVSS.n3106 DVSS.n3105 39.5177
R28447 DVSS.n3177 DVSS.n3176 39.5177
R28448 DVSS.n3941 DVSS.n3757 36.7611
R28449 DVSS.n4406 DVSS.n4222 36.7611
R28450 DVSS.n2345 DVSS.n2161 36.7611
R28451 DVSS.n2810 DVSS.n2626 36.7611
R28452 DVSS.n5409 DVSS.n5225 36.7611
R28453 DVSS.n5874 DVSS.n5690 36.7611
R28454 DVSS.n344 DVSS.n160 36.7611
R28455 DVSS.n809 DVSS.n625 36.7611
R28456 DVSS.n1360 DVSS.n1355 36.2246
R28457 DVSS.n1449 DVSS.n1444 36.2246
R28458 DVSS.n1610 DVSS.n1605 36.2246
R28459 DVSS.n1699 DVSS.n1694 36.2246
R28460 DVSS.n4573 DVSS.n4568 36.2246
R28461 DVSS.n4662 DVSS.n4657 36.2246
R28462 DVSS.n4823 DVSS.n4818 36.2246
R28463 DVSS.n4912 DVSS.n4907 36.2246
R28464 DVSS.n6041 DVSS.n6036 36.2246
R28465 DVSS.n6130 DVSS.n6125 36.2246
R28466 DVSS.n6291 DVSS.n6286 36.2246
R28467 DVSS.n6380 DVSS.n6375 36.2246
R28468 DVSS.n2977 DVSS.n2972 36.2246
R28469 DVSS.n3066 DVSS.n3061 36.2246
R28470 DVSS.n3227 DVSS.n3222 36.2246
R28471 DVSS.n3316 DVSS.n3311 36.2246
R28472 DVSS.t0 DVSS.t172 36.1979
R28473 DVSS.n6558 DVSS.n6557 36.1417
R28474 DVSS.n3599 DVSS.n3598 36.1417
R28475 DVSS.n1997 DVSS.n1994 36.1417
R28476 DVSS.n6770 DVSS.n6767 36.1417
R28477 DVSS.n6159 DVSS.n6158 35.7729
R28478 DVSS.n6260 DVSS.n6259 35.7729
R28479 DVSS.n4691 DVSS.n4690 35.7729
R28480 DVSS.n4792 DVSS.n4791 35.7729
R28481 DVSS.n3095 DVSS.n3094 35.7729
R28482 DVSS.n3196 DVSS.n3195 35.7729
R28483 DVSS.n1478 DVSS.n1477 35.7729
R28484 DVSS.n1579 DVSS.n1578 35.7729
R28485 DVSS.n3889 DVSS.n3887 35.3887
R28486 DVSS.n3913 DVSS.n3900 35.3887
R28487 DVSS.n3887 DVSS.n3791 35.3887
R28488 DVSS.n3893 DVSS.n3786 35.3887
R28489 DVSS.n3881 DVSS.n3786 35.3887
R28490 DVSS.n4354 DVSS.n4352 35.3887
R28491 DVSS.n4378 DVSS.n4365 35.3887
R28492 DVSS.n4352 DVSS.n4256 35.3887
R28493 DVSS.n4358 DVSS.n4251 35.3887
R28494 DVSS.n4346 DVSS.n4251 35.3887
R28495 DVSS.n2293 DVSS.n2291 35.3887
R28496 DVSS.n2317 DVSS.n2304 35.3887
R28497 DVSS.n2291 DVSS.n2195 35.3887
R28498 DVSS.n2297 DVSS.n2190 35.3887
R28499 DVSS.n2285 DVSS.n2190 35.3887
R28500 DVSS.n2758 DVSS.n2756 35.3887
R28501 DVSS.n2782 DVSS.n2769 35.3887
R28502 DVSS.n2756 DVSS.n2660 35.3887
R28503 DVSS.n2762 DVSS.n2655 35.3887
R28504 DVSS.n2750 DVSS.n2655 35.3887
R28505 DVSS.n5357 DVSS.n5355 35.3887
R28506 DVSS.n5381 DVSS.n5368 35.3887
R28507 DVSS.n5355 DVSS.n5259 35.3887
R28508 DVSS.n5361 DVSS.n5254 35.3887
R28509 DVSS.n5349 DVSS.n5254 35.3887
R28510 DVSS.n5822 DVSS.n5820 35.3887
R28511 DVSS.n5846 DVSS.n5833 35.3887
R28512 DVSS.n5820 DVSS.n5724 35.3887
R28513 DVSS.n5826 DVSS.n5719 35.3887
R28514 DVSS.n5814 DVSS.n5719 35.3887
R28515 DVSS.n292 DVSS.n290 35.3887
R28516 DVSS.n316 DVSS.n303 35.3887
R28517 DVSS.n290 DVSS.n194 35.3887
R28518 DVSS.n296 DVSS.n189 35.3887
R28519 DVSS.n284 DVSS.n189 35.3887
R28520 DVSS.n757 DVSS.n755 35.3887
R28521 DVSS.n781 DVSS.n768 35.3887
R28522 DVSS.n755 DVSS.n659 35.3887
R28523 DVSS.n761 DVSS.n654 35.3887
R28524 DVSS.n749 DVSS.n654 35.3887
R28525 DVSS.n1158 DVSS.t158 35.0689
R28526 DVSS.n1063 DVSS.t261 35.0689
R28527 DVSS.n4032 DVSS.n3625 34.1338
R28528 DVSS.n3658 DVSS.n3644 34.1338
R28529 DVSS.n4497 DVSS.n4090 34.1338
R28530 DVSS.n4123 DVSS.n4109 34.1338
R28531 DVSS.n2436 DVSS.n2029 34.1338
R28532 DVSS.n2062 DVSS.n2048 34.1338
R28533 DVSS.n2901 DVSS.n2494 34.1338
R28534 DVSS.n2527 DVSS.n2513 34.1338
R28535 DVSS.n5500 DVSS.n5093 34.1338
R28536 DVSS.n5126 DVSS.n5112 34.1338
R28537 DVSS.n5965 DVSS.n5558 34.1338
R28538 DVSS.n5591 DVSS.n5577 34.1338
R28539 DVSS.n435 DVSS.n28 34.1338
R28540 DVSS.n61 DVSS.n47 34.1338
R28541 DVSS.n900 DVSS.n493 34.1338
R28542 DVSS.n526 DVSS.n512 34.1338
R28543 DVSS.n1314 DVSS.n1313 33.5205
R28544 DVSS.n1299 DVSS.n1297 33.5205
R28545 DVSS.n1021 DVSS.n1020 33.5205
R28546 DVSS.n1006 DVSS.n1005 33.5205
R28547 DVSS.n1794 DVSS.n1793 33.5205
R28548 DVSS.n1811 DVSS.n1810 33.5205
R28549 DVSS.n6840 DVSS.n6839 33.5205
R28550 DVSS.n6824 DVSS.n6822 33.5205
R28551 DVSS.n3524 DVSS.n3523 33.5205
R28552 DVSS.n3541 DVSS.n3539 33.5205
R28553 DVSS.n6613 DVSS.n6611 33.5205
R28554 DVSS.n5073 DVSS.n5072 33.5205
R28555 DVSS.n5006 DVSS.n5005 33.5205
R28556 DVSS.n5023 DVSS.n5022 33.5205
R28557 DVSS.n1938 DVSS.n1936 33.5205
R28558 DVSS.n1921 DVSS.n1920 33.5205
R28559 DVSS.n3411 DVSS.n3410 33.5205
R28560 DVSS.n3428 DVSS.n3427 33.5205
R28561 DVSS.n6474 DVSS.n6473 33.5205
R28562 DVSS.n6491 DVSS.n6490 33.5205
R28563 DVSS.n3423 DVSS.n3422 32.9668
R28564 DVSS.n5018 DVSS.n5017 32.9668
R28565 DVSS.n1806 DVSS.n1805 32.9668
R28566 DVSS.n1474 DVSS.n1473 32.9315
R28567 DVSS.n1575 DVSS.n1574 32.9315
R28568 DVSS.n4687 DVSS.n4686 32.9315
R28569 DVSS.n4788 DVSS.n4787 32.9315
R28570 DVSS.n6155 DVSS.n6154 32.9315
R28571 DVSS.n6256 DVSS.n6255 32.9315
R28572 DVSS.n3091 DVSS.n3090 32.9315
R28573 DVSS.n3192 DVSS.n3191 32.9315
R28574 DVSS.n6039 DVSS.n6037 30.6625
R28575 DVSS.n6128 DVSS.n6127 30.6625
R28576 DVSS.n6289 DVSS.n6287 30.6625
R28577 DVSS.n6378 DVSS.n6377 30.6625
R28578 DVSS.n4571 DVSS.n4569 30.6625
R28579 DVSS.n4660 DVSS.n4659 30.6625
R28580 DVSS.n4821 DVSS.n4819 30.6625
R28581 DVSS.n4910 DVSS.n4909 30.6625
R28582 DVSS.n2975 DVSS.n2973 30.6625
R28583 DVSS.n3064 DVSS.n3063 30.6625
R28584 DVSS.n3225 DVSS.n3223 30.6625
R28585 DVSS.n3314 DVSS.n3313 30.6625
R28586 DVSS.n1358 DVSS.n1356 30.6625
R28587 DVSS.n1447 DVSS.n1446 30.6625
R28588 DVSS.n1608 DVSS.n1606 30.6625
R28589 DVSS.n1697 DVSS.n1696 30.6625
R28590 DVSS.n1181 DVSS.n1180 30.5709
R28591 DVSS.n3913 DVSS.n3912 29.7417
R28592 DVSS.n4378 DVSS.n4377 29.7417
R28593 DVSS.n2317 DVSS.n2316 29.7417
R28594 DVSS.n2782 DVSS.n2781 29.7417
R28595 DVSS.n5381 DVSS.n5380 29.7417
R28596 DVSS.n5846 DVSS.n5845 29.7417
R28597 DVSS.n316 DVSS.n315 29.7417
R28598 DVSS.n781 DVSS.n780 29.7417
R28599 DVSS.n1464 DVSS.n1459 29.6384
R28600 DVSS.n1595 DVSS.n1590 29.6384
R28601 DVSS.n4677 DVSS.n4672 29.6384
R28602 DVSS.n4808 DVSS.n4803 29.6384
R28603 DVSS.n6145 DVSS.n6140 29.6384
R28604 DVSS.n6276 DVSS.n6271 29.6384
R28605 DVSS.n3081 DVSS.n3076 29.6384
R28606 DVSS.n3212 DVSS.n3207 29.6384
R28607 DVSS.n3749 DVSS.n3738 29.4833
R28608 DVSS.n3728 DVSS.n3717 29.4833
R28609 DVSS.n4214 DVSS.n4203 29.4833
R28610 DVSS.n4193 DVSS.n4182 29.4833
R28611 DVSS.n2153 DVSS.n2142 29.4833
R28612 DVSS.n2132 DVSS.n2121 29.4833
R28613 DVSS.n2618 DVSS.n2607 29.4833
R28614 DVSS.n2597 DVSS.n2586 29.4833
R28615 DVSS.n5217 DVSS.n5206 29.4833
R28616 DVSS.n5196 DVSS.n5185 29.4833
R28617 DVSS.n5682 DVSS.n5671 29.4833
R28618 DVSS.n5661 DVSS.n5650 29.4833
R28619 DVSS.n152 DVSS.n141 29.4833
R28620 DVSS.n131 DVSS.n120 29.4833
R28621 DVSS.n617 DVSS.n606 29.4833
R28622 DVSS.n596 DVSS.n585 29.4833
R28623 DVSS.n3698 DVSS.n3681 29.1989
R28624 DVSS.n4055 DVSS.n4034 29.1989
R28625 DVSS.n4163 DVSS.n4146 29.1989
R28626 DVSS.n4520 DVSS.n4499 29.1989
R28627 DVSS.n2102 DVSS.n2085 29.1989
R28628 DVSS.n2459 DVSS.n2438 29.1989
R28629 DVSS.n2567 DVSS.n2550 29.1989
R28630 DVSS.n2924 DVSS.n2903 29.1989
R28631 DVSS.n5166 DVSS.n5149 29.1989
R28632 DVSS.n5523 DVSS.n5502 29.1989
R28633 DVSS.n5631 DVSS.n5614 29.1989
R28634 DVSS.n5988 DVSS.n5967 29.1989
R28635 DVSS.n101 DVSS.n84 29.1989
R28636 DVSS.n458 DVSS.n437 29.1989
R28637 DVSS.n566 DVSS.n549 29.1989
R28638 DVSS.n923 DVSS.n902 29.1989
R28639 DVSS.n970 DVSS.t253 28.1205
R28640 DVSS.n1752 DVSS.t233 28.1205
R28641 DVSS.n4964 DVSS.t171 28.1205
R28642 DVSS.n3369 DVSS.t70 28.1205
R28643 DVSS.n6432 DVSS.t259 28.1205
R28644 DVSS.n1459 DVSS.n1458 26.3453
R28645 DVSS.n1590 DVSS.n1589 26.3453
R28646 DVSS.n4672 DVSS.n4671 26.3453
R28647 DVSS.n4803 DVSS.n4802 26.3453
R28648 DVSS.n6140 DVSS.n6139 26.3453
R28649 DVSS.n6271 DVSS.n6270 26.3453
R28650 DVSS.n3076 DVSS.n3075 26.3453
R28651 DVSS.n3207 DVSS.n3206 26.3453
R28652 DVSS.n1730 DVSS.n1724 25.6005
R28653 DVSS.n1724 DVSS.n1721 25.6005
R28654 DVSS.n1721 DVSS.n1719 25.6005
R28655 DVSS.n1719 DVSS.n1716 25.6005
R28656 DVSS.n953 DVSS.n952 25.6005
R28657 DVSS.n952 DVSS.n951 25.6005
R28658 DVSS.n951 DVSS.n950 25.6005
R28659 DVSS.n950 DVSS.n949 25.6005
R28660 DVSS.n949 DVSS.n948 25.6005
R28661 DVSS.n948 DVSS.n947 25.6005
R28662 DVSS.n947 DVSS.n946 25.6005
R28663 DVSS.n946 DVSS.n945 25.6005
R28664 DVSS.n945 DVSS.n944 25.6005
R28665 DVSS.n944 DVSS.n943 25.6005
R28666 DVSS.n943 DVSS.n942 25.6005
R28667 DVSS.n942 DVSS.n941 25.6005
R28668 DVSS.n1703 DVSS.n1702 25.6005
R28669 DVSS.n1704 DVSS.n1703 25.6005
R28670 DVSS.n1705 DVSS.n1704 25.6005
R28671 DVSS.n1706 DVSS.n1705 25.6005
R28672 DVSS.n1707 DVSS.n1706 25.6005
R28673 DVSS.n1708 DVSS.n1707 25.6005
R28674 DVSS.n1709 DVSS.n1708 25.6005
R28675 DVSS.n1710 DVSS.n1709 25.6005
R28676 DVSS.n1711 DVSS.n1710 25.6005
R28677 DVSS.n1712 DVSS.n1711 25.6005
R28678 DVSS.n1713 DVSS.n1712 25.6005
R28679 DVSS.n1714 DVSS.n1713 25.6005
R28680 DVSS.n1350 DVSS.n962 25.6005
R28681 DVSS.n962 DVSS.n960 25.6005
R28682 DVSS.n960 DVSS.n957 25.6005
R28683 DVSS.n957 DVSS.n955 25.6005
R28684 DVSS.n4943 DVSS.n4937 25.6005
R28685 DVSS.n4937 DVSS.n4934 25.6005
R28686 DVSS.n4934 DVSS.n4932 25.6005
R28687 DVSS.n4932 DVSS.n4929 25.6005
R28688 DVSS.n4550 DVSS.n4549 25.6005
R28689 DVSS.n4549 DVSS.n4548 25.6005
R28690 DVSS.n4548 DVSS.n4547 25.6005
R28691 DVSS.n4547 DVSS.n4546 25.6005
R28692 DVSS.n4546 DVSS.n4545 25.6005
R28693 DVSS.n4545 DVSS.n4544 25.6005
R28694 DVSS.n4544 DVSS.n4543 25.6005
R28695 DVSS.n4543 DVSS.n4542 25.6005
R28696 DVSS.n4542 DVSS.n4541 25.6005
R28697 DVSS.n4541 DVSS.n4540 25.6005
R28698 DVSS.n4540 DVSS.n4539 25.6005
R28699 DVSS.n4539 DVSS.n4538 25.6005
R28700 DVSS.n4916 DVSS.n4915 25.6005
R28701 DVSS.n4917 DVSS.n4916 25.6005
R28702 DVSS.n4918 DVSS.n4917 25.6005
R28703 DVSS.n4919 DVSS.n4918 25.6005
R28704 DVSS.n4920 DVSS.n4919 25.6005
R28705 DVSS.n4921 DVSS.n4920 25.6005
R28706 DVSS.n4922 DVSS.n4921 25.6005
R28707 DVSS.n4923 DVSS.n4922 25.6005
R28708 DVSS.n4924 DVSS.n4923 25.6005
R28709 DVSS.n4925 DVSS.n4924 25.6005
R28710 DVSS.n4926 DVSS.n4925 25.6005
R28711 DVSS.n4927 DVSS.n4926 25.6005
R28712 DVSS.n4563 DVSS.n4559 25.6005
R28713 DVSS.n4559 DVSS.n4557 25.6005
R28714 DVSS.n4557 DVSS.n4554 25.6005
R28715 DVSS.n4554 DVSS.n4552 25.6005
R28716 DVSS.n3889 DVSS.n3888 25.6005
R28717 DVSS.n3888 DVSS.n3783 25.6005
R28718 DVSS.n3900 DVSS.n3783 25.6005
R28719 DVSS.n3875 DVSS.n3873 25.6005
R28720 DVSS.n3875 DVSS.n3874 25.6005
R28721 DVSS.n3874 DVSS.n3791 25.6005
R28722 DVSS.n3912 DVSS.n3911 25.6005
R28723 DVSS.n3894 DVSS.n3893 25.6005
R28724 DVSS.n3895 DVSS.n3894 25.6005
R28725 DVSS.n3895 DVSS.n3757 25.6005
R28726 DVSS.n3879 DVSS.n3845 25.6005
R28727 DVSS.n3880 DVSS.n3879 25.6005
R28728 DVSS.n3881 DVSS.n3880 25.6005
R28729 DVSS.n4354 DVSS.n4353 25.6005
R28730 DVSS.n4353 DVSS.n4248 25.6005
R28731 DVSS.n4365 DVSS.n4248 25.6005
R28732 DVSS.n4340 DVSS.n4338 25.6005
R28733 DVSS.n4340 DVSS.n4339 25.6005
R28734 DVSS.n4339 DVSS.n4256 25.6005
R28735 DVSS.n4377 DVSS.n4376 25.6005
R28736 DVSS.n4359 DVSS.n4358 25.6005
R28737 DVSS.n4360 DVSS.n4359 25.6005
R28738 DVSS.n4360 DVSS.n4222 25.6005
R28739 DVSS.n4344 DVSS.n4310 25.6005
R28740 DVSS.n4345 DVSS.n4344 25.6005
R28741 DVSS.n4346 DVSS.n4345 25.6005
R28742 DVSS.n6411 DVSS.n6405 25.6005
R28743 DVSS.n6405 DVSS.n6402 25.6005
R28744 DVSS.n6402 DVSS.n6400 25.6005
R28745 DVSS.n6400 DVSS.n6397 25.6005
R28746 DVSS.n6018 DVSS.n6017 25.6005
R28747 DVSS.n6017 DVSS.n6016 25.6005
R28748 DVSS.n6016 DVSS.n6015 25.6005
R28749 DVSS.n6015 DVSS.n6014 25.6005
R28750 DVSS.n6014 DVSS.n6013 25.6005
R28751 DVSS.n6013 DVSS.n6012 25.6005
R28752 DVSS.n6012 DVSS.n6011 25.6005
R28753 DVSS.n6011 DVSS.n6010 25.6005
R28754 DVSS.n6010 DVSS.n6009 25.6005
R28755 DVSS.n6009 DVSS.n6008 25.6005
R28756 DVSS.n6008 DVSS.n6007 25.6005
R28757 DVSS.n6007 DVSS.n6006 25.6005
R28758 DVSS.n6384 DVSS.n6383 25.6005
R28759 DVSS.n6385 DVSS.n6384 25.6005
R28760 DVSS.n6386 DVSS.n6385 25.6005
R28761 DVSS.n6387 DVSS.n6386 25.6005
R28762 DVSS.n6388 DVSS.n6387 25.6005
R28763 DVSS.n6389 DVSS.n6388 25.6005
R28764 DVSS.n6390 DVSS.n6389 25.6005
R28765 DVSS.n6391 DVSS.n6390 25.6005
R28766 DVSS.n6392 DVSS.n6391 25.6005
R28767 DVSS.n6393 DVSS.n6392 25.6005
R28768 DVSS.n6394 DVSS.n6393 25.6005
R28769 DVSS.n6395 DVSS.n6394 25.6005
R28770 DVSS.n6031 DVSS.n6027 25.6005
R28771 DVSS.n6027 DVSS.n6025 25.6005
R28772 DVSS.n6025 DVSS.n6022 25.6005
R28773 DVSS.n6022 DVSS.n6020 25.6005
R28774 DVSS.n3348 DVSS.n3341 25.6005
R28775 DVSS.n3341 DVSS.n3338 25.6005
R28776 DVSS.n3338 DVSS.n3336 25.6005
R28777 DVSS.n3336 DVSS.n3333 25.6005
R28778 DVSS.n2954 DVSS.n2953 25.6005
R28779 DVSS.n2953 DVSS.n2952 25.6005
R28780 DVSS.n2952 DVSS.n2951 25.6005
R28781 DVSS.n2951 DVSS.n2950 25.6005
R28782 DVSS.n2950 DVSS.n2949 25.6005
R28783 DVSS.n2949 DVSS.n2948 25.6005
R28784 DVSS.n2948 DVSS.n2947 25.6005
R28785 DVSS.n2947 DVSS.n2946 25.6005
R28786 DVSS.n2946 DVSS.n2945 25.6005
R28787 DVSS.n2945 DVSS.n2944 25.6005
R28788 DVSS.n2944 DVSS.n2943 25.6005
R28789 DVSS.n2943 DVSS.n2942 25.6005
R28790 DVSS.n3320 DVSS.n3319 25.6005
R28791 DVSS.n3321 DVSS.n3320 25.6005
R28792 DVSS.n3322 DVSS.n3321 25.6005
R28793 DVSS.n3323 DVSS.n3322 25.6005
R28794 DVSS.n3324 DVSS.n3323 25.6005
R28795 DVSS.n3325 DVSS.n3324 25.6005
R28796 DVSS.n3326 DVSS.n3325 25.6005
R28797 DVSS.n3327 DVSS.n3326 25.6005
R28798 DVSS.n3328 DVSS.n3327 25.6005
R28799 DVSS.n3329 DVSS.n3328 25.6005
R28800 DVSS.n3330 DVSS.n3329 25.6005
R28801 DVSS.n3331 DVSS.n3330 25.6005
R28802 DVSS.n2967 DVSS.n2963 25.6005
R28803 DVSS.n2963 DVSS.n2961 25.6005
R28804 DVSS.n2961 DVSS.n2958 25.6005
R28805 DVSS.n2958 DVSS.n2956 25.6005
R28806 DVSS.n2293 DVSS.n2292 25.6005
R28807 DVSS.n2292 DVSS.n2187 25.6005
R28808 DVSS.n2304 DVSS.n2187 25.6005
R28809 DVSS.n2279 DVSS.n2277 25.6005
R28810 DVSS.n2279 DVSS.n2278 25.6005
R28811 DVSS.n2278 DVSS.n2195 25.6005
R28812 DVSS.n2316 DVSS.n2315 25.6005
R28813 DVSS.n2298 DVSS.n2297 25.6005
R28814 DVSS.n2299 DVSS.n2298 25.6005
R28815 DVSS.n2299 DVSS.n2161 25.6005
R28816 DVSS.n2283 DVSS.n2249 25.6005
R28817 DVSS.n2284 DVSS.n2283 25.6005
R28818 DVSS.n2285 DVSS.n2284 25.6005
R28819 DVSS.n2758 DVSS.n2757 25.6005
R28820 DVSS.n2757 DVSS.n2652 25.6005
R28821 DVSS.n2769 DVSS.n2652 25.6005
R28822 DVSS.n2744 DVSS.n2742 25.6005
R28823 DVSS.n2744 DVSS.n2743 25.6005
R28824 DVSS.n2743 DVSS.n2660 25.6005
R28825 DVSS.n2781 DVSS.n2780 25.6005
R28826 DVSS.n2763 DVSS.n2762 25.6005
R28827 DVSS.n2764 DVSS.n2763 25.6005
R28828 DVSS.n2764 DVSS.n2626 25.6005
R28829 DVSS.n2748 DVSS.n2714 25.6005
R28830 DVSS.n2749 DVSS.n2748 25.6005
R28831 DVSS.n2750 DVSS.n2749 25.6005
R28832 DVSS.n5357 DVSS.n5356 25.6005
R28833 DVSS.n5356 DVSS.n5251 25.6005
R28834 DVSS.n5368 DVSS.n5251 25.6005
R28835 DVSS.n5343 DVSS.n5341 25.6005
R28836 DVSS.n5343 DVSS.n5342 25.6005
R28837 DVSS.n5342 DVSS.n5259 25.6005
R28838 DVSS.n5380 DVSS.n5379 25.6005
R28839 DVSS.n5362 DVSS.n5361 25.6005
R28840 DVSS.n5363 DVSS.n5362 25.6005
R28841 DVSS.n5363 DVSS.n5225 25.6005
R28842 DVSS.n5347 DVSS.n5313 25.6005
R28843 DVSS.n5348 DVSS.n5347 25.6005
R28844 DVSS.n5349 DVSS.n5348 25.6005
R28845 DVSS.n5822 DVSS.n5821 25.6005
R28846 DVSS.n5821 DVSS.n5716 25.6005
R28847 DVSS.n5833 DVSS.n5716 25.6005
R28848 DVSS.n5808 DVSS.n5806 25.6005
R28849 DVSS.n5808 DVSS.n5807 25.6005
R28850 DVSS.n5807 DVSS.n5724 25.6005
R28851 DVSS.n5845 DVSS.n5844 25.6005
R28852 DVSS.n5827 DVSS.n5826 25.6005
R28853 DVSS.n5828 DVSS.n5827 25.6005
R28854 DVSS.n5828 DVSS.n5690 25.6005
R28855 DVSS.n5812 DVSS.n5778 25.6005
R28856 DVSS.n5813 DVSS.n5812 25.6005
R28857 DVSS.n5814 DVSS.n5813 25.6005
R28858 DVSS.n292 DVSS.n291 25.6005
R28859 DVSS.n291 DVSS.n186 25.6005
R28860 DVSS.n303 DVSS.n186 25.6005
R28861 DVSS.n278 DVSS.n276 25.6005
R28862 DVSS.n278 DVSS.n277 25.6005
R28863 DVSS.n277 DVSS.n194 25.6005
R28864 DVSS.n315 DVSS.n314 25.6005
R28865 DVSS.n297 DVSS.n296 25.6005
R28866 DVSS.n298 DVSS.n297 25.6005
R28867 DVSS.n298 DVSS.n160 25.6005
R28868 DVSS.n282 DVSS.n248 25.6005
R28869 DVSS.n283 DVSS.n282 25.6005
R28870 DVSS.n284 DVSS.n283 25.6005
R28871 DVSS.n757 DVSS.n756 25.6005
R28872 DVSS.n756 DVSS.n651 25.6005
R28873 DVSS.n768 DVSS.n651 25.6005
R28874 DVSS.n743 DVSS.n741 25.6005
R28875 DVSS.n743 DVSS.n742 25.6005
R28876 DVSS.n742 DVSS.n659 25.6005
R28877 DVSS.n780 DVSS.n779 25.6005
R28878 DVSS.n762 DVSS.n761 25.6005
R28879 DVSS.n763 DVSS.n762 25.6005
R28880 DVSS.n763 DVSS.n625 25.6005
R28881 DVSS.n747 DVSS.n713 25.6005
R28882 DVSS.n748 DVSS.n747 25.6005
R28883 DVSS.n749 DVSS.n748 25.6005
R28884 DVSS.n6174 DVSS.n6173 25.5522
R28885 DVSS.n6245 DVSS.n6244 25.5522
R28886 DVSS.n4706 DVSS.n4705 25.5522
R28887 DVSS.n4777 DVSS.n4776 25.5522
R28888 DVSS.n3110 DVSS.n3109 25.5522
R28889 DVSS.n3181 DVSS.n3180 25.5522
R28890 DVSS.n1493 DVSS.n1492 25.5522
R28891 DVSS.n1564 DVSS.n1563 25.5522
R28892 DVSS.n1321 DVSS.n1319 24.1542
R28893 DVSS.n6656 DVSS.t87 23.988
R28894 DVSS.n1860 DVSS.t39 23.9135
R28895 DVSS.n1479 DVSS.n1474 23.0522
R28896 DVSS.n1580 DVSS.n1575 23.0522
R28897 DVSS.n4692 DVSS.n4687 23.0522
R28898 DVSS.n4793 DVSS.n4788 23.0522
R28899 DVSS.n6160 DVSS.n6155 23.0522
R28900 DVSS.n6261 DVSS.n6256 23.0522
R28901 DVSS.n3096 DVSS.n3091 23.0522
R28902 DVSS.n3197 DVSS.n3192 23.0522
R28903 DVSS.n4008 DVSS.n3625 22.3184
R28904 DVSS.n4009 DVSS.n4008 22.3184
R28905 DVSS.n4010 DVSS.n4009 22.3184
R28906 DVSS.n4010 DVSS.n4003 22.3184
R28907 DVSS.n4015 DVSS.n4003 22.3184
R28908 DVSS.n4016 DVSS.n4015 22.3184
R28909 DVSS.n4016 DVSS.n4001 22.3184
R28910 DVSS.n4021 DVSS.n4001 22.3184
R28911 DVSS.n3658 DVSS.n3657 22.3184
R28912 DVSS.n3663 DVSS.n3657 22.3184
R28913 DVSS.n3664 DVSS.n3663 22.3184
R28914 DVSS.n3664 DVSS.n3655 22.3184
R28915 DVSS.n3670 DVSS.n3655 22.3184
R28916 DVSS.n3671 DVSS.n3670 22.3184
R28917 DVSS.n3671 DVSS.n3653 22.3184
R28918 DVSS.n3676 DVSS.n3653 22.3184
R28919 DVSS.n4473 DVSS.n4090 22.3184
R28920 DVSS.n4474 DVSS.n4473 22.3184
R28921 DVSS.n4475 DVSS.n4474 22.3184
R28922 DVSS.n4475 DVSS.n4468 22.3184
R28923 DVSS.n4480 DVSS.n4468 22.3184
R28924 DVSS.n4481 DVSS.n4480 22.3184
R28925 DVSS.n4481 DVSS.n4466 22.3184
R28926 DVSS.n4486 DVSS.n4466 22.3184
R28927 DVSS.n4123 DVSS.n4122 22.3184
R28928 DVSS.n4128 DVSS.n4122 22.3184
R28929 DVSS.n4129 DVSS.n4128 22.3184
R28930 DVSS.n4129 DVSS.n4120 22.3184
R28931 DVSS.n4135 DVSS.n4120 22.3184
R28932 DVSS.n4136 DVSS.n4135 22.3184
R28933 DVSS.n4136 DVSS.n4118 22.3184
R28934 DVSS.n4141 DVSS.n4118 22.3184
R28935 DVSS.n2412 DVSS.n2029 22.3184
R28936 DVSS.n2413 DVSS.n2412 22.3184
R28937 DVSS.n2414 DVSS.n2413 22.3184
R28938 DVSS.n2414 DVSS.n2407 22.3184
R28939 DVSS.n2419 DVSS.n2407 22.3184
R28940 DVSS.n2420 DVSS.n2419 22.3184
R28941 DVSS.n2420 DVSS.n2405 22.3184
R28942 DVSS.n2425 DVSS.n2405 22.3184
R28943 DVSS.n2062 DVSS.n2061 22.3184
R28944 DVSS.n2067 DVSS.n2061 22.3184
R28945 DVSS.n2068 DVSS.n2067 22.3184
R28946 DVSS.n2068 DVSS.n2059 22.3184
R28947 DVSS.n2074 DVSS.n2059 22.3184
R28948 DVSS.n2075 DVSS.n2074 22.3184
R28949 DVSS.n2075 DVSS.n2057 22.3184
R28950 DVSS.n2080 DVSS.n2057 22.3184
R28951 DVSS.n2877 DVSS.n2494 22.3184
R28952 DVSS.n2878 DVSS.n2877 22.3184
R28953 DVSS.n2879 DVSS.n2878 22.3184
R28954 DVSS.n2879 DVSS.n2872 22.3184
R28955 DVSS.n2884 DVSS.n2872 22.3184
R28956 DVSS.n2885 DVSS.n2884 22.3184
R28957 DVSS.n2885 DVSS.n2870 22.3184
R28958 DVSS.n2890 DVSS.n2870 22.3184
R28959 DVSS.n2527 DVSS.n2526 22.3184
R28960 DVSS.n2532 DVSS.n2526 22.3184
R28961 DVSS.n2533 DVSS.n2532 22.3184
R28962 DVSS.n2533 DVSS.n2524 22.3184
R28963 DVSS.n2539 DVSS.n2524 22.3184
R28964 DVSS.n2540 DVSS.n2539 22.3184
R28965 DVSS.n2540 DVSS.n2522 22.3184
R28966 DVSS.n2545 DVSS.n2522 22.3184
R28967 DVSS.n5476 DVSS.n5093 22.3184
R28968 DVSS.n5477 DVSS.n5476 22.3184
R28969 DVSS.n5478 DVSS.n5477 22.3184
R28970 DVSS.n5478 DVSS.n5471 22.3184
R28971 DVSS.n5483 DVSS.n5471 22.3184
R28972 DVSS.n5484 DVSS.n5483 22.3184
R28973 DVSS.n5484 DVSS.n5469 22.3184
R28974 DVSS.n5489 DVSS.n5469 22.3184
R28975 DVSS.n5126 DVSS.n5125 22.3184
R28976 DVSS.n5131 DVSS.n5125 22.3184
R28977 DVSS.n5132 DVSS.n5131 22.3184
R28978 DVSS.n5132 DVSS.n5123 22.3184
R28979 DVSS.n5138 DVSS.n5123 22.3184
R28980 DVSS.n5139 DVSS.n5138 22.3184
R28981 DVSS.n5139 DVSS.n5121 22.3184
R28982 DVSS.n5144 DVSS.n5121 22.3184
R28983 DVSS.n5941 DVSS.n5558 22.3184
R28984 DVSS.n5942 DVSS.n5941 22.3184
R28985 DVSS.n5943 DVSS.n5942 22.3184
R28986 DVSS.n5943 DVSS.n5936 22.3184
R28987 DVSS.n5948 DVSS.n5936 22.3184
R28988 DVSS.n5949 DVSS.n5948 22.3184
R28989 DVSS.n5949 DVSS.n5934 22.3184
R28990 DVSS.n5954 DVSS.n5934 22.3184
R28991 DVSS.n5591 DVSS.n5590 22.3184
R28992 DVSS.n5596 DVSS.n5590 22.3184
R28993 DVSS.n5597 DVSS.n5596 22.3184
R28994 DVSS.n5597 DVSS.n5588 22.3184
R28995 DVSS.n5603 DVSS.n5588 22.3184
R28996 DVSS.n5604 DVSS.n5603 22.3184
R28997 DVSS.n5604 DVSS.n5586 22.3184
R28998 DVSS.n5609 DVSS.n5586 22.3184
R28999 DVSS.n411 DVSS.n28 22.3184
R29000 DVSS.n412 DVSS.n411 22.3184
R29001 DVSS.n413 DVSS.n412 22.3184
R29002 DVSS.n413 DVSS.n406 22.3184
R29003 DVSS.n418 DVSS.n406 22.3184
R29004 DVSS.n419 DVSS.n418 22.3184
R29005 DVSS.n419 DVSS.n404 22.3184
R29006 DVSS.n424 DVSS.n404 22.3184
R29007 DVSS.n61 DVSS.n60 22.3184
R29008 DVSS.n66 DVSS.n60 22.3184
R29009 DVSS.n67 DVSS.n66 22.3184
R29010 DVSS.n67 DVSS.n58 22.3184
R29011 DVSS.n73 DVSS.n58 22.3184
R29012 DVSS.n74 DVSS.n73 22.3184
R29013 DVSS.n74 DVSS.n56 22.3184
R29014 DVSS.n79 DVSS.n56 22.3184
R29015 DVSS.n876 DVSS.n493 22.3184
R29016 DVSS.n877 DVSS.n876 22.3184
R29017 DVSS.n878 DVSS.n877 22.3184
R29018 DVSS.n878 DVSS.n871 22.3184
R29019 DVSS.n883 DVSS.n871 22.3184
R29020 DVSS.n884 DVSS.n883 22.3184
R29021 DVSS.n884 DVSS.n869 22.3184
R29022 DVSS.n889 DVSS.n869 22.3184
R29023 DVSS.n526 DVSS.n525 22.3184
R29024 DVSS.n531 DVSS.n525 22.3184
R29025 DVSS.n532 DVSS.n531 22.3184
R29026 DVSS.n532 DVSS.n523 22.3184
R29027 DVSS.n538 DVSS.n523 22.3184
R29028 DVSS.n539 DVSS.n538 22.3184
R29029 DVSS.n539 DVSS.n521 22.3184
R29030 DVSS.n544 DVSS.n521 22.3184
R29031 DVSS.n1158 DVSS.t1 22.2377
R29032 DVSS.n1063 DVSS.t159 22.2377
R29033 DVSS.n1139 DVSS.t265 21.2805
R29034 DVSS.n1139 DVSS.t264 21.2805
R29035 DVSS.n970 DVSS.t146 21.2805
R29036 DVSS.n1077 DVSS.t155 21.2805
R29037 DVSS.n1077 DVSS.t156 21.2805
R29038 DVSS.n1752 DVSS.t26 21.2805
R29039 DVSS.n1873 DVSS.t60 21.2805
R29040 DVSS.n1873 DVSS.t227 21.2805
R29041 DVSS.n6669 DVSS.t255 21.2805
R29042 DVSS.n6669 DVSS.t195 21.2805
R29043 DVSS.n4964 DVSS.t257 21.2805
R29044 DVSS.n3369 DVSS.t24 21.2805
R29045 DVSS.n6432 DVSS.t64 21.2805
R29046 DVSS.n6054 DVSS.n6052 20.4418
R29047 DVSS.n6113 DVSS.n6112 20.4418
R29048 DVSS.n6304 DVSS.n6302 20.4418
R29049 DVSS.n6363 DVSS.n6362 20.4418
R29050 DVSS.n4586 DVSS.n4584 20.4418
R29051 DVSS.n4645 DVSS.n4644 20.4418
R29052 DVSS.n4836 DVSS.n4834 20.4418
R29053 DVSS.n4895 DVSS.n4894 20.4418
R29054 DVSS.n2990 DVSS.n2988 20.4418
R29055 DVSS.n3049 DVSS.n3048 20.4418
R29056 DVSS.n3240 DVSS.n3238 20.4418
R29057 DVSS.n3299 DVSS.n3298 20.4418
R29058 DVSS.n1373 DVSS.n1371 20.4418
R29059 DVSS.n1432 DVSS.n1431 20.4418
R29060 DVSS.n1623 DVSS.n1621 20.4418
R29061 DVSS.n1682 DVSS.n1681 20.4418
R29062 DVSS.n4022 DVSS.n4021 20.3492
R29063 DVSS.n3677 DVSS.n3676 20.3492
R29064 DVSS.n4487 DVSS.n4486 20.3492
R29065 DVSS.n4142 DVSS.n4141 20.3492
R29066 DVSS.n2426 DVSS.n2425 20.3492
R29067 DVSS.n2081 DVSS.n2080 20.3492
R29068 DVSS.n2891 DVSS.n2890 20.3492
R29069 DVSS.n2546 DVSS.n2545 20.3492
R29070 DVSS.n5490 DVSS.n5489 20.3492
R29071 DVSS.n5145 DVSS.n5144 20.3492
R29072 DVSS.n5955 DVSS.n5954 20.3492
R29073 DVSS.n5610 DVSS.n5609 20.3492
R29074 DVSS.n425 DVSS.n424 20.3492
R29075 DVSS.n80 DVSS.n79 20.3492
R29076 DVSS.n890 DVSS.n889 20.3492
R29077 DVSS.n545 DVSS.n544 20.3492
R29078 DVSS.n1260 DVSS.t150 20.0005
R29079 DVSS.n1260 DVSS.t239 20.0005
R29080 DVSS.n6781 DVSS.t134 20.0005
R29081 DVSS.n6781 DVSS.t117 20.0005
R29082 DVSS.n3581 DVSS.t203 20.0005
R29083 DVSS.n3581 DVSS.t72 20.0005
R29084 DVSS.n6569 DVSS.t213 20.0005
R29085 DVSS.n6569 DVSS.t229 20.0005
R29086 DVSS.n1978 DVSS.t18 20.0005
R29087 DVSS.n1978 DVSS.t192 20.0005
R29088 DVSS.n1355 DVSS.n1354 19.7591
R29089 DVSS.n1444 DVSS.n1443 19.7591
R29090 DVSS.n1605 DVSS.n1604 19.7591
R29091 DVSS.n1694 DVSS.n1693 19.7591
R29092 DVSS.n4568 DVSS.n4567 19.7591
R29093 DVSS.n4657 DVSS.n4656 19.7591
R29094 DVSS.n4818 DVSS.n4817 19.7591
R29095 DVSS.n4907 DVSS.n4906 19.7591
R29096 DVSS.n6036 DVSS.n6035 19.7591
R29097 DVSS.n6125 DVSS.n6124 19.7591
R29098 DVSS.n6286 DVSS.n6285 19.7591
R29099 DVSS.n6375 DVSS.n6374 19.7591
R29100 DVSS.n2972 DVSS.n2971 19.7591
R29101 DVSS.n3061 DVSS.n3060 19.7591
R29102 DVSS.n3222 DVSS.n3221 19.7591
R29103 DVSS.n3311 DVSS.n3310 19.7591
R29104 DVSS.n3344 DVSS.n3343 18.4105
R29105 DVSS.n1336 DVSS.n1335 18.0103
R29106 DVSS.n1119 DVSS.n1118 18.0093
R29107 DVSS.n1126 DVSS.n1125 18.0093
R29108 DVSS.n1135 DVSS.n1131 18.0093
R29109 DVSS.n1123 DVSS.n1122 18.0093
R29110 DVSS.n1161 DVSS.n1160 18.007
R29111 DVSS.n1116 DVSS.n1115 17.2422
R29112 DVSS.n4032 DVSS.n4031 17.0218
R29113 DVSS.n4497 DVSS.n4496 17.0218
R29114 DVSS.n2436 DVSS.n2435 17.0218
R29115 DVSS.n2901 DVSS.n2900 17.0218
R29116 DVSS.n5500 DVSS.n5499 17.0218
R29117 DVSS.n5965 DVSS.n5964 17.0218
R29118 DVSS.n435 DVSS.n434 17.0218
R29119 DVSS.n900 DVSS.n899 17.0218
R29120 DVSS.n3983 DVSS.n3644 16.8856
R29121 DVSS.n4448 DVSS.n4109 16.8856
R29122 DVSS.n2387 DVSS.n2048 16.8856
R29123 DVSS.n2852 DVSS.n2513 16.8856
R29124 DVSS.n5451 DVSS.n5112 16.8856
R29125 DVSS.n5916 DVSS.n5577 16.8856
R29126 DVSS.n386 DVSS.n47 16.8856
R29127 DVSS.n851 DVSS.n512 16.8856
R29128 DVSS.n1494 DVSS.n1489 16.466
R29129 DVSS.n1565 DVSS.n1560 16.466
R29130 DVSS.n4707 DVSS.n4702 16.466
R29131 DVSS.n4778 DVSS.n4773 16.466
R29132 DVSS.n6175 DVSS.n6170 16.466
R29133 DVSS.n6246 DVSS.n6241 16.466
R29134 DVSS.n3111 DVSS.n3106 16.466
R29135 DVSS.n3182 DVSS.n3177 16.466
R29136 DVSS.n3965 DVSS.n3644 15.5239
R29137 DVSS.n4430 DVSS.n4109 15.5239
R29138 DVSS.n2369 DVSS.n2048 15.5239
R29139 DVSS.n2834 DVSS.n2513 15.5239
R29140 DVSS.n5433 DVSS.n5112 15.5239
R29141 DVSS.n5898 DVSS.n5577 15.5239
R29142 DVSS.n368 DVSS.n47 15.5239
R29143 DVSS.n833 DVSS.n512 15.5239
R29144 DVSS.n3747 DVSS.n3746 15.463
R29145 DVSS.n3726 DVSS.n3725 15.463
R29146 DVSS.n4212 DVSS.n4211 15.463
R29147 DVSS.n4191 DVSS.n4190 15.463
R29148 DVSS.n2151 DVSS.n2150 15.463
R29149 DVSS.n2130 DVSS.n2129 15.463
R29150 DVSS.n2616 DVSS.n2615 15.463
R29151 DVSS.n2595 DVSS.n2594 15.463
R29152 DVSS.n5215 DVSS.n5214 15.463
R29153 DVSS.n5194 DVSS.n5193 15.463
R29154 DVSS.n5680 DVSS.n5679 15.463
R29155 DVSS.n5659 DVSS.n5658 15.463
R29156 DVSS.n150 DVSS.n149 15.463
R29157 DVSS.n129 DVSS.n128 15.463
R29158 DVSS.n615 DVSS.n614 15.463
R29159 DVSS.n594 DVSS.n593 15.463
R29160 DVSS.n4033 DVSS.n4032 15.3877
R29161 DVSS.n4498 DVSS.n4497 15.3877
R29162 DVSS.n2437 DVSS.n2436 15.3877
R29163 DVSS.n2902 DVSS.n2901 15.3877
R29164 DVSS.n5501 DVSS.n5500 15.3877
R29165 DVSS.n5966 DVSS.n5965 15.3877
R29166 DVSS.n436 DVSS.n435 15.3877
R29167 DVSS.n901 DVSS.n900 15.3877
R29168 DVSS.n6189 DVSS.n6188 15.3315
R29169 DVSS.n6230 DVSS.n6229 15.3315
R29170 DVSS.n4721 DVSS.n4720 15.3315
R29171 DVSS.n4762 DVSS.n4761 15.3315
R29172 DVSS.n3125 DVSS.n3124 15.3315
R29173 DVSS.n3166 DVSS.n3165 15.3315
R29174 DVSS.n1508 DVSS.n1507 15.3315
R29175 DVSS.n1549 DVSS.n1548 15.3315
R29176 DVSS.n1182 DVSS.n1181 14.4554
R29177 DVSS.n1079 DVSS.n1078 14.4288
R29178 DVSS.n3752 DVSS.n3739 13.5534
R29179 DVSS.n3747 DVSS.n3743 13.5534
R29180 DVSS.n3731 DVSS.n3718 13.5534
R29181 DVSS.n3726 DVSS.n3722 13.5534
R29182 DVSS.n4217 DVSS.n4204 13.5534
R29183 DVSS.n4212 DVSS.n4208 13.5534
R29184 DVSS.n4196 DVSS.n4183 13.5534
R29185 DVSS.n4191 DVSS.n4187 13.5534
R29186 DVSS.n2156 DVSS.n2143 13.5534
R29187 DVSS.n2151 DVSS.n2147 13.5534
R29188 DVSS.n2135 DVSS.n2122 13.5534
R29189 DVSS.n2130 DVSS.n2126 13.5534
R29190 DVSS.n2621 DVSS.n2608 13.5534
R29191 DVSS.n2616 DVSS.n2612 13.5534
R29192 DVSS.n2600 DVSS.n2587 13.5534
R29193 DVSS.n2595 DVSS.n2591 13.5534
R29194 DVSS.n5220 DVSS.n5207 13.5534
R29195 DVSS.n5215 DVSS.n5211 13.5534
R29196 DVSS.n5199 DVSS.n5186 13.5534
R29197 DVSS.n5194 DVSS.n5190 13.5534
R29198 DVSS.n5685 DVSS.n5672 13.5534
R29199 DVSS.n5680 DVSS.n5676 13.5534
R29200 DVSS.n5664 DVSS.n5651 13.5534
R29201 DVSS.n5659 DVSS.n5655 13.5534
R29202 DVSS.n155 DVSS.n142 13.5534
R29203 DVSS.n150 DVSS.n146 13.5534
R29204 DVSS.n134 DVSS.n121 13.5534
R29205 DVSS.n129 DVSS.n125 13.5534
R29206 DVSS.n620 DVSS.n607 13.5534
R29207 DVSS.n615 DVSS.n611 13.5534
R29208 DVSS.n599 DVSS.n586 13.5534
R29209 DVSS.n594 DVSS.n590 13.5534
R29210 DVSS.n1370 DVSS.n1369 13.1729
R29211 DVSS.n1429 DVSS.n1428 13.1729
R29212 DVSS.n1620 DVSS.n1619 13.1729
R29213 DVSS.n1679 DVSS.n1678 13.1729
R29214 DVSS.n4583 DVSS.n4582 13.1729
R29215 DVSS.n4642 DVSS.n4641 13.1729
R29216 DVSS.n4833 DVSS.n4832 13.1729
R29217 DVSS.n4892 DVSS.n4891 13.1729
R29218 DVSS.n6051 DVSS.n6050 13.1729
R29219 DVSS.n6110 DVSS.n6109 13.1729
R29220 DVSS.n6301 DVSS.n6300 13.1729
R29221 DVSS.n6360 DVSS.n6359 13.1729
R29222 DVSS.n2987 DVSS.n2986 13.1729
R29223 DVSS.n3046 DVSS.n3045 13.1729
R29224 DVSS.n3237 DVSS.n3236 13.1729
R29225 DVSS.n3296 DVSS.n3295 13.1729
R29226 DVSS.n1746 DVSS.n1742 12.8977
R29227 DVSS.n4958 DVSS.n4954 12.8977
R29228 DVSS.n3363 DVSS.n3362 12.8977
R29229 DVSS.n6426 DVSS.n6422 12.8977
R29230 DVSS.n1222 DVSS.n1218 12.8862
R29231 DVSS.n1402 DVSS.n1400 12.8005
R29232 DVSS.n1402 DVSS.n1401 12.8005
R29233 DVSS.n1652 DVSS.n1650 12.8005
R29234 DVSS.n1652 DVSS.n1651 12.8005
R29235 DVSS.n4615 DVSS.n4613 12.8005
R29236 DVSS.n4615 DVSS.n4614 12.8005
R29237 DVSS.n4865 DVSS.n4863 12.8005
R29238 DVSS.n4865 DVSS.n4864 12.8005
R29239 DVSS.n6083 DVSS.n6081 12.8005
R29240 DVSS.n6083 DVSS.n6082 12.8005
R29241 DVSS.n6333 DVSS.n6331 12.8005
R29242 DVSS.n6333 DVSS.n6332 12.8005
R29243 DVSS.n3019 DVSS.n3017 12.8005
R29244 DVSS.n3019 DVSS.n3018 12.8005
R29245 DVSS.n3269 DVSS.n3267 12.8005
R29246 DVSS.n3269 DVSS.n3268 12.8005
R29247 DVSS.n3548 DVSS.t49 12.6286
R29248 DVSS.n6602 DVSS.t99 12.6286
R29249 DVSS.n1945 DVSS.t183 12.608
R29250 DVSS.n6813 DVSS.t31 12.608
R29251 DVSS.n3544 DVSS.n3543 12.2862
R29252 DVSS.n6608 DVSS.n6607 12.2862
R29253 DVSS.n1941 DVSS.n1940 12.2762
R29254 DVSS.n6819 DVSS.n6818 12.2762
R29255 DVSS.n6625 DVSS.n6624 12.261
R29256 DVSS.n3527 DVSS.n3526 12.261
R29257 DVSS.n1924 DVSS.n1923 12.2511
R29258 DVSS.n6836 DVSS.n6835 12.2511
R29259 DVSS.n1313 DVSS.t248 10.6405
R29260 DVSS.n1313 DVSS.t250 10.6405
R29261 DVSS.n1297 DVSS.t251 10.6405
R29262 DVSS.n1297 DVSS.t249 10.6405
R29263 DVSS.n1005 DVSS.t242 10.6405
R29264 DVSS.n1005 DVSS.t236 10.6405
R29265 DVSS.n1020 DVSS.t240 10.6405
R29266 DVSS.n1020 DVSS.t241 10.6405
R29267 DVSS.n1793 DVSS.t142 10.6405
R29268 DVSS.n1793 DVSS.t136 10.6405
R29269 DVSS.n1810 DVSS.t138 10.6405
R29270 DVSS.n1810 DVSS.t144 10.6405
R29271 DVSS.n6839 DVSS.t36 10.6405
R29272 DVSS.n6839 DVSS.t28 10.6405
R29273 DVSS.n6822 DVSS.t30 10.6405
R29274 DVSS.n6822 DVSS.t32 10.6405
R29275 DVSS.n3523 DVSS.t48 10.6405
R29276 DVSS.n3523 DVSS.t42 10.6405
R29277 DVSS.n3539 DVSS.t46 10.6405
R29278 DVSS.n3539 DVSS.t50 10.6405
R29279 DVSS.n5072 DVSS.t102 10.6405
R29280 DVSS.n5072 DVSS.t106 10.6405
R29281 DVSS.n6611 DVSS.t98 10.6405
R29282 DVSS.n6611 DVSS.t100 10.6405
R29283 DVSS.n5005 DVSS.t205 10.6405
R29284 DVSS.n5005 DVSS.t207 10.6405
R29285 DVSS.n5022 DVSS.t209 10.6405
R29286 DVSS.n5022 DVSS.t201 10.6405
R29287 DVSS.n1920 DVSS.t176 10.6405
R29288 DVSS.n1920 DVSS.t178 10.6405
R29289 DVSS.n1936 DVSS.t182 10.6405
R29290 DVSS.n1936 DVSS.t184 10.6405
R29291 DVSS.n3410 DVSS.t16 10.6405
R29292 DVSS.n3410 DVSS.t10 10.6405
R29293 DVSS.n3427 DVSS.t8 10.6405
R29294 DVSS.n3427 DVSS.t14 10.6405
R29295 DVSS.n6473 DVSS.t219 10.6405
R29296 DVSS.n6473 DVSS.t221 10.6405
R29297 DVSS.n6490 DVSS.t211 10.6405
R29298 DVSS.n6490 DVSS.t215 10.6405
R29299 DVSS.n3902 DVSS.n3779 10.4252
R29300 DVSS.n4367 DVSS.n4244 10.4252
R29301 DVSS.n2306 DVSS.n2183 10.4252
R29302 DVSS.n2771 DVSS.n2648 10.4252
R29303 DVSS.n5370 DVSS.n5247 10.4252
R29304 DVSS.n5835 DVSS.n5712 10.4252
R29305 DVSS.n305 DVSS.n182 10.4252
R29306 DVSS.n770 DVSS.n647 10.4252
R29307 DVSS.n6070 DVSS.n6068 10.2212
R29308 DVSS.n6098 DVSS.n6097 10.2212
R29309 DVSS.n6320 DVSS.n6318 10.2212
R29310 DVSS.n6348 DVSS.n6347 10.2212
R29311 DVSS.n4602 DVSS.n4600 10.2212
R29312 DVSS.n4630 DVSS.n4629 10.2212
R29313 DVSS.n4852 DVSS.n4850 10.2212
R29314 DVSS.n4880 DVSS.n4879 10.2212
R29315 DVSS.n3006 DVSS.n3004 10.2212
R29316 DVSS.n3034 DVSS.n3033 10.2212
R29317 DVSS.n3256 DVSS.n3254 10.2212
R29318 DVSS.n3284 DVSS.n3283 10.2212
R29319 DVSS.n1389 DVSS.n1387 10.2212
R29320 DVSS.n1417 DVSS.n1416 10.2212
R29321 DVSS.n1639 DVSS.n1637 10.2212
R29322 DVSS.n1667 DVSS.n1666 10.2212
R29323 DVSS.n1509 DVSS.n1504 9.87981
R29324 DVSS.n1550 DVSS.n1545 9.87981
R29325 DVSS.n4722 DVSS.n4717 9.87981
R29326 DVSS.n4763 DVSS.n4758 9.87981
R29327 DVSS.n6190 DVSS.n6185 9.87981
R29328 DVSS.n6231 DVSS.n6226 9.87981
R29329 DVSS.n3126 DVSS.n3121 9.87981
R29330 DVSS.n3167 DVSS.n3162 9.87981
R29331 DVSS.n3560 DVSS.n3559 9.56928
R29332 DVSS.n1957 DVSS.n1956 9.56793
R29333 DVSS.n6805 DVSS.n6804 9.56793
R29334 DVSS.n4537 DVSS.n4536 9.31763
R29335 DVSS.n2941 DVSS.n2940 9.31763
R29336 DVSS.n6005 DVSS.n6004 9.31763
R29337 DVSS.n940 DVSS.n939 9.31763
R29338 DVSS.n1836 DVSS.n1835 9.3005
R29339 DVSS.n5048 DVSS.n5047 9.3005
R29340 DVSS.n3737 DVSS.n3736 9.3005
R29341 DVSS.n3744 DVSS.n3740 9.3005
R29342 DVSS.n3745 DVSS.n3743 9.3005
R29343 DVSS.n3750 DVSS.n3742 9.3005
R29344 DVSS.n3750 DVSS.n3749 9.3005
R29345 DVSS.n3741 DVSS.n3739 9.3005
R29346 DVSS.n3755 DVSS.n3754 9.3005
R29347 DVSS.n3716 DVSS.n3715 9.3005
R29348 DVSS.n3723 DVSS.n3719 9.3005
R29349 DVSS.n3724 DVSS.n3722 9.3005
R29350 DVSS.n3729 DVSS.n3721 9.3005
R29351 DVSS.n3729 DVSS.n3728 9.3005
R29352 DVSS.n3720 DVSS.n3718 9.3005
R29353 DVSS.n3734 DVSS.n3733 9.3005
R29354 DVSS.n3950 DVSS.n3949 9.3005
R29355 DVSS.n3953 DVSS.n3952 9.3005
R29356 DVSS.n3954 DVSS.n3685 9.3005
R29357 DVSS.n3959 DVSS.n3958 9.3005
R29358 DVSS.n3957 DVSS.n3686 9.3005
R29359 DVSS.n3956 DVSS.n3955 9.3005
R29360 DVSS.n3652 DVSS.n3651 9.3005
R29361 DVSS.n3970 DVSS.n3969 9.3005
R29362 DVSS.n3971 DVSS.n3649 9.3005
R29363 DVSS.n3979 DVSS.n3978 9.3005
R29364 DVSS.n3977 DVSS.n3650 9.3005
R29365 DVSS.n3974 DVSS.n3973 9.3005
R29366 DVSS.n3972 DVSS.n3638 9.3005
R29367 DVSS.n3990 DVSS.n3637 9.3005
R29368 DVSS.n3992 DVSS.n3991 9.3005
R29369 DVSS.n3993 DVSS.n3636 9.3005
R29370 DVSS.n3996 DVSS.n3635 9.3005
R29371 DVSS.n3998 DVSS.n3997 9.3005
R29372 DVSS.n3999 DVSS.n3633 9.3005
R29373 DVSS.n4027 DVSS.n4026 9.3005
R29374 DVSS.n4025 DVSS.n3634 9.3005
R29375 DVSS.n4024 DVSS.n4023 9.3005
R29376 DVSS.n4000 DVSS.n3618 9.3005
R29377 DVSS.n4061 DVSS.n3619 9.3005
R29378 DVSS.n4062 DVSS.n3617 9.3005
R29379 DVSS.n4064 DVSS.n4063 9.3005
R29380 DVSS.n4065 DVSS.n3616 9.3005
R29381 DVSS.n4068 DVSS.n4067 9.3005
R29382 DVSS.n4073 DVSS.n4072 9.3005
R29383 DVSS.n4202 DVSS.n4201 9.3005
R29384 DVSS.n4209 DVSS.n4205 9.3005
R29385 DVSS.n4210 DVSS.n4208 9.3005
R29386 DVSS.n4215 DVSS.n4207 9.3005
R29387 DVSS.n4215 DVSS.n4214 9.3005
R29388 DVSS.n4206 DVSS.n4204 9.3005
R29389 DVSS.n4220 DVSS.n4219 9.3005
R29390 DVSS.n4181 DVSS.n4180 9.3005
R29391 DVSS.n4188 DVSS.n4184 9.3005
R29392 DVSS.n4189 DVSS.n4187 9.3005
R29393 DVSS.n4194 DVSS.n4186 9.3005
R29394 DVSS.n4194 DVSS.n4193 9.3005
R29395 DVSS.n4185 DVSS.n4183 9.3005
R29396 DVSS.n4199 DVSS.n4198 9.3005
R29397 DVSS.n4415 DVSS.n4414 9.3005
R29398 DVSS.n4418 DVSS.n4417 9.3005
R29399 DVSS.n4419 DVSS.n4150 9.3005
R29400 DVSS.n4424 DVSS.n4423 9.3005
R29401 DVSS.n4422 DVSS.n4151 9.3005
R29402 DVSS.n4421 DVSS.n4420 9.3005
R29403 DVSS.n4117 DVSS.n4116 9.3005
R29404 DVSS.n4435 DVSS.n4434 9.3005
R29405 DVSS.n4436 DVSS.n4114 9.3005
R29406 DVSS.n4444 DVSS.n4443 9.3005
R29407 DVSS.n4442 DVSS.n4115 9.3005
R29408 DVSS.n4439 DVSS.n4438 9.3005
R29409 DVSS.n4437 DVSS.n4103 9.3005
R29410 DVSS.n4455 DVSS.n4102 9.3005
R29411 DVSS.n4457 DVSS.n4456 9.3005
R29412 DVSS.n4458 DVSS.n4101 9.3005
R29413 DVSS.n4461 DVSS.n4100 9.3005
R29414 DVSS.n4463 DVSS.n4462 9.3005
R29415 DVSS.n4464 DVSS.n4098 9.3005
R29416 DVSS.n4492 DVSS.n4491 9.3005
R29417 DVSS.n4490 DVSS.n4099 9.3005
R29418 DVSS.n4489 DVSS.n4488 9.3005
R29419 DVSS.n4465 DVSS.n4083 9.3005
R29420 DVSS.n4526 DVSS.n4084 9.3005
R29421 DVSS.n4527 DVSS.n4082 9.3005
R29422 DVSS.n4529 DVSS.n4528 9.3005
R29423 DVSS.n4530 DVSS.n4081 9.3005
R29424 DVSS.n4532 DVSS.n4531 9.3005
R29425 DVSS.n4577 DVSS.n4576 9.3005
R29426 DVSS.n4592 DVSS.n4591 9.3005
R29427 DVSS.n4610 DVSS.n4609 9.3005
R29428 DVSS.n4620 DVSS.n4619 9.3005
R29429 DVSS.n4638 DVSS.n4637 9.3005
R29430 DVSS.n4653 DVSS.n4652 9.3005
R29431 DVSS.n4668 DVSS.n4667 9.3005
R29432 DVSS.n4683 DVSS.n4682 9.3005
R29433 DVSS.n4698 DVSS.n4697 9.3005
R29434 DVSS.n4713 DVSS.n4712 9.3005
R29435 DVSS.n4728 DVSS.n4727 9.3005
R29436 DVSS.n4752 DVSS.n4751 9.3005
R29437 DVSS.n4767 DVSS.n4766 9.3005
R29438 DVSS.n4782 DVSS.n4781 9.3005
R29439 DVSS.n4797 DVSS.n4796 9.3005
R29440 DVSS.n4812 DVSS.n4811 9.3005
R29441 DVSS.n4827 DVSS.n4826 9.3005
R29442 DVSS.n4842 DVSS.n4841 9.3005
R29443 DVSS.n4860 DVSS.n4859 9.3005
R29444 DVSS.n4870 DVSS.n4869 9.3005
R29445 DVSS.n4888 DVSS.n4887 9.3005
R29446 DVSS.n4903 DVSS.n4902 9.3005
R29447 DVSS.n4901 DVSS.n4900 9.3005
R29448 DVSS.n4868 DVSS.n4867 9.3005
R29449 DVSS.n4862 DVSS.n4861 9.3005
R29450 DVSS.n4829 DVSS.n4828 9.3005
R29451 DVSS.n4799 DVSS.n4798 9.3005
R29452 DVSS.n4769 DVSS.n4768 9.3005
R29453 DVSS.n4711 DVSS.n4710 9.3005
R29454 DVSS.n4681 DVSS.n4680 9.3005
R29455 DVSS.n4651 DVSS.n4650 9.3005
R29456 DVSS.n4618 DVSS.n4617 9.3005
R29457 DVSS.n4612 DVSS.n4611 9.3005
R29458 DVSS.n4579 DVSS.n4578 9.3005
R29459 DVSS.n4594 DVSS.n4593 9.3005
R29460 DVSS.n4636 DVSS.n4635 9.3005
R29461 DVSS.n4666 DVSS.n4665 9.3005
R29462 DVSS.n4696 DVSS.n4695 9.3005
R29463 DVSS.n4726 DVSS.n4725 9.3005
R29464 DVSS.n4754 DVSS.n4753 9.3005
R29465 DVSS.n4784 DVSS.n4783 9.3005
R29466 DVSS.n4814 DVSS.n4813 9.3005
R29467 DVSS.n4844 DVSS.n4843 9.3005
R29468 DVSS.n4886 DVSS.n4885 9.3005
R29469 DVSS.n6045 DVSS.n6044 9.3005
R29470 DVSS.n6060 DVSS.n6059 9.3005
R29471 DVSS.n6078 DVSS.n6077 9.3005
R29472 DVSS.n6088 DVSS.n6087 9.3005
R29473 DVSS.n6106 DVSS.n6105 9.3005
R29474 DVSS.n6121 DVSS.n6120 9.3005
R29475 DVSS.n6136 DVSS.n6135 9.3005
R29476 DVSS.n6151 DVSS.n6150 9.3005
R29477 DVSS.n6166 DVSS.n6165 9.3005
R29478 DVSS.n6181 DVSS.n6180 9.3005
R29479 DVSS.n6196 DVSS.n6195 9.3005
R29480 DVSS.n6220 DVSS.n6219 9.3005
R29481 DVSS.n6235 DVSS.n6234 9.3005
R29482 DVSS.n6250 DVSS.n6249 9.3005
R29483 DVSS.n6265 DVSS.n6264 9.3005
R29484 DVSS.n6280 DVSS.n6279 9.3005
R29485 DVSS.n6295 DVSS.n6294 9.3005
R29486 DVSS.n6310 DVSS.n6309 9.3005
R29487 DVSS.n6328 DVSS.n6327 9.3005
R29488 DVSS.n6338 DVSS.n6337 9.3005
R29489 DVSS.n6356 DVSS.n6355 9.3005
R29490 DVSS.n6371 DVSS.n6370 9.3005
R29491 DVSS.n6369 DVSS.n6368 9.3005
R29492 DVSS.n6336 DVSS.n6335 9.3005
R29493 DVSS.n6330 DVSS.n6329 9.3005
R29494 DVSS.n6297 DVSS.n6296 9.3005
R29495 DVSS.n6267 DVSS.n6266 9.3005
R29496 DVSS.n6237 DVSS.n6236 9.3005
R29497 DVSS.n6179 DVSS.n6178 9.3005
R29498 DVSS.n6149 DVSS.n6148 9.3005
R29499 DVSS.n6119 DVSS.n6118 9.3005
R29500 DVSS.n6086 DVSS.n6085 9.3005
R29501 DVSS.n6080 DVSS.n6079 9.3005
R29502 DVSS.n6047 DVSS.n6046 9.3005
R29503 DVSS.n6062 DVSS.n6061 9.3005
R29504 DVSS.n6104 DVSS.n6103 9.3005
R29505 DVSS.n6134 DVSS.n6133 9.3005
R29506 DVSS.n6164 DVSS.n6163 9.3005
R29507 DVSS.n6194 DVSS.n6193 9.3005
R29508 DVSS.n6222 DVSS.n6221 9.3005
R29509 DVSS.n6252 DVSS.n6251 9.3005
R29510 DVSS.n6282 DVSS.n6281 9.3005
R29511 DVSS.n6312 DVSS.n6311 9.3005
R29512 DVSS.n6354 DVSS.n6353 9.3005
R29513 DVSS.n6382 DVSS.n6381 9.3005
R29514 DVSS.n6381 DVSS.n6380 9.3005
R29515 DVSS.n6380 DVSS.n6379 9.3005
R29516 DVSS.n6352 DVSS.n6351 9.3005
R29517 DVSS.n6351 DVSS.n6350 9.3005
R29518 DVSS.n6350 DVSS.n6349 9.3005
R29519 DVSS.n6192 DVSS.n6191 9.3005
R29520 DVSS.n6191 DVSS.n6190 9.3005
R29521 DVSS.n6190 DVSS.n6189 9.3005
R29522 DVSS.n6162 DVSS.n6161 9.3005
R29523 DVSS.n6161 DVSS.n6160 9.3005
R29524 DVSS.n6160 DVSS.n6159 9.3005
R29525 DVSS.n6132 DVSS.n6131 9.3005
R29526 DVSS.n6131 DVSS.n6130 9.3005
R29527 DVSS.n6130 DVSS.n6129 9.3005
R29528 DVSS.n6102 DVSS.n6101 9.3005
R29529 DVSS.n6101 DVSS.n6100 9.3005
R29530 DVSS.n6100 DVSS.n6099 9.3005
R29531 DVSS.n6043 DVSS.n6042 9.3005
R29532 DVSS.n6042 DVSS.n6041 9.3005
R29533 DVSS.n6041 DVSS.n6040 9.3005
R29534 DVSS.n6058 DVSS.n6057 9.3005
R29535 DVSS.n6057 DVSS.n6056 9.3005
R29536 DVSS.n6056 DVSS.n6055 9.3005
R29537 DVSS.n6076 DVSS.n6075 9.3005
R29538 DVSS.n6075 DVSS.n6074 9.3005
R29539 DVSS.n6074 DVSS.n6073 9.3005
R29540 DVSS.n6117 DVSS.n6116 9.3005
R29541 DVSS.n6116 DVSS.n6115 9.3005
R29542 DVSS.n6115 DVSS.n6114 9.3005
R29543 DVSS.n6147 DVSS.n6146 9.3005
R29544 DVSS.n6146 DVSS.n6145 9.3005
R29545 DVSS.n6145 DVSS.n6144 9.3005
R29546 DVSS.n6177 DVSS.n6176 9.3005
R29547 DVSS.n6176 DVSS.n6175 9.3005
R29548 DVSS.n6175 DVSS.n6174 9.3005
R29549 DVSS.n6207 DVSS.n6206 9.3005
R29550 DVSS.n6206 DVSS.n6205 9.3005
R29551 DVSS.n6205 DVSS.n6204 9.3005
R29552 DVSS.n6218 DVSS.n6217 9.3005
R29553 DVSS.n6217 DVSS.n6216 9.3005
R29554 DVSS.n6216 DVSS.n6215 9.3005
R29555 DVSS.n6233 DVSS.n6232 9.3005
R29556 DVSS.n6232 DVSS.n6231 9.3005
R29557 DVSS.n6231 DVSS.n6230 9.3005
R29558 DVSS.n6248 DVSS.n6247 9.3005
R29559 DVSS.n6247 DVSS.n6246 9.3005
R29560 DVSS.n6246 DVSS.n6245 9.3005
R29561 DVSS.n6263 DVSS.n6262 9.3005
R29562 DVSS.n6262 DVSS.n6261 9.3005
R29563 DVSS.n6261 DVSS.n6260 9.3005
R29564 DVSS.n6278 DVSS.n6277 9.3005
R29565 DVSS.n6277 DVSS.n6276 9.3005
R29566 DVSS.n6276 DVSS.n6275 9.3005
R29567 DVSS.n6293 DVSS.n6292 9.3005
R29568 DVSS.n6292 DVSS.n6291 9.3005
R29569 DVSS.n6291 DVSS.n6290 9.3005
R29570 DVSS.n6308 DVSS.n6307 9.3005
R29571 DVSS.n6307 DVSS.n6306 9.3005
R29572 DVSS.n6306 DVSS.n6305 9.3005
R29573 DVSS.n6326 DVSS.n6325 9.3005
R29574 DVSS.n6325 DVSS.n6324 9.3005
R29575 DVSS.n6324 DVSS.n6323 9.3005
R29576 DVSS.n6367 DVSS.n6366 9.3005
R29577 DVSS.n6366 DVSS.n6365 9.3005
R29578 DVSS.n6365 DVSS.n6364 9.3005
R29579 DVSS.n4914 DVSS.n4913 9.3005
R29580 DVSS.n4913 DVSS.n4912 9.3005
R29581 DVSS.n4912 DVSS.n4911 9.3005
R29582 DVSS.n4884 DVSS.n4883 9.3005
R29583 DVSS.n4883 DVSS.n4882 9.3005
R29584 DVSS.n4882 DVSS.n4881 9.3005
R29585 DVSS.n4724 DVSS.n4723 9.3005
R29586 DVSS.n4723 DVSS.n4722 9.3005
R29587 DVSS.n4722 DVSS.n4721 9.3005
R29588 DVSS.n4694 DVSS.n4693 9.3005
R29589 DVSS.n4693 DVSS.n4692 9.3005
R29590 DVSS.n4692 DVSS.n4691 9.3005
R29591 DVSS.n4664 DVSS.n4663 9.3005
R29592 DVSS.n4663 DVSS.n4662 9.3005
R29593 DVSS.n4662 DVSS.n4661 9.3005
R29594 DVSS.n4634 DVSS.n4633 9.3005
R29595 DVSS.n4633 DVSS.n4632 9.3005
R29596 DVSS.n4632 DVSS.n4631 9.3005
R29597 DVSS.n4575 DVSS.n4574 9.3005
R29598 DVSS.n4574 DVSS.n4573 9.3005
R29599 DVSS.n4573 DVSS.n4572 9.3005
R29600 DVSS.n4590 DVSS.n4589 9.3005
R29601 DVSS.n4589 DVSS.n4588 9.3005
R29602 DVSS.n4588 DVSS.n4587 9.3005
R29603 DVSS.n4608 DVSS.n4607 9.3005
R29604 DVSS.n4607 DVSS.n4606 9.3005
R29605 DVSS.n4606 DVSS.n4605 9.3005
R29606 DVSS.n4649 DVSS.n4648 9.3005
R29607 DVSS.n4648 DVSS.n4647 9.3005
R29608 DVSS.n4647 DVSS.n4646 9.3005
R29609 DVSS.n4679 DVSS.n4678 9.3005
R29610 DVSS.n4678 DVSS.n4677 9.3005
R29611 DVSS.n4677 DVSS.n4676 9.3005
R29612 DVSS.n4709 DVSS.n4708 9.3005
R29613 DVSS.n4708 DVSS.n4707 9.3005
R29614 DVSS.n4707 DVSS.n4706 9.3005
R29615 DVSS.n4739 DVSS.n4738 9.3005
R29616 DVSS.n4738 DVSS.n4737 9.3005
R29617 DVSS.n4737 DVSS.n4736 9.3005
R29618 DVSS.n4750 DVSS.n4749 9.3005
R29619 DVSS.n4749 DVSS.n4748 9.3005
R29620 DVSS.n4748 DVSS.n4747 9.3005
R29621 DVSS.n4765 DVSS.n4764 9.3005
R29622 DVSS.n4764 DVSS.n4763 9.3005
R29623 DVSS.n4763 DVSS.n4762 9.3005
R29624 DVSS.n4780 DVSS.n4779 9.3005
R29625 DVSS.n4779 DVSS.n4778 9.3005
R29626 DVSS.n4778 DVSS.n4777 9.3005
R29627 DVSS.n4795 DVSS.n4794 9.3005
R29628 DVSS.n4794 DVSS.n4793 9.3005
R29629 DVSS.n4793 DVSS.n4792 9.3005
R29630 DVSS.n4810 DVSS.n4809 9.3005
R29631 DVSS.n4809 DVSS.n4808 9.3005
R29632 DVSS.n4808 DVSS.n4807 9.3005
R29633 DVSS.n4825 DVSS.n4824 9.3005
R29634 DVSS.n4824 DVSS.n4823 9.3005
R29635 DVSS.n4823 DVSS.n4822 9.3005
R29636 DVSS.n4840 DVSS.n4839 9.3005
R29637 DVSS.n4839 DVSS.n4838 9.3005
R29638 DVSS.n4838 DVSS.n4837 9.3005
R29639 DVSS.n4858 DVSS.n4857 9.3005
R29640 DVSS.n4857 DVSS.n4856 9.3005
R29641 DVSS.n4856 DVSS.n4855 9.3005
R29642 DVSS.n4899 DVSS.n4898 9.3005
R29643 DVSS.n4898 DVSS.n4897 9.3005
R29644 DVSS.n4897 DVSS.n4896 9.3005
R29645 DVSS.n3453 DVSS.n3452 9.3005
R29646 DVSS.n2004 DVSS.n2003 9.3005
R29647 DVSS.n2141 DVSS.n2140 9.3005
R29648 DVSS.n2148 DVSS.n2144 9.3005
R29649 DVSS.n2149 DVSS.n2147 9.3005
R29650 DVSS.n2154 DVSS.n2146 9.3005
R29651 DVSS.n2154 DVSS.n2153 9.3005
R29652 DVSS.n2145 DVSS.n2143 9.3005
R29653 DVSS.n2159 DVSS.n2158 9.3005
R29654 DVSS.n2120 DVSS.n2119 9.3005
R29655 DVSS.n2127 DVSS.n2123 9.3005
R29656 DVSS.n2128 DVSS.n2126 9.3005
R29657 DVSS.n2133 DVSS.n2125 9.3005
R29658 DVSS.n2133 DVSS.n2132 9.3005
R29659 DVSS.n2124 DVSS.n2122 9.3005
R29660 DVSS.n2138 DVSS.n2137 9.3005
R29661 DVSS.n2354 DVSS.n2353 9.3005
R29662 DVSS.n2357 DVSS.n2356 9.3005
R29663 DVSS.n2358 DVSS.n2089 9.3005
R29664 DVSS.n2363 DVSS.n2362 9.3005
R29665 DVSS.n2361 DVSS.n2090 9.3005
R29666 DVSS.n2360 DVSS.n2359 9.3005
R29667 DVSS.n2056 DVSS.n2055 9.3005
R29668 DVSS.n2374 DVSS.n2373 9.3005
R29669 DVSS.n2375 DVSS.n2053 9.3005
R29670 DVSS.n2383 DVSS.n2382 9.3005
R29671 DVSS.n2381 DVSS.n2054 9.3005
R29672 DVSS.n2378 DVSS.n2377 9.3005
R29673 DVSS.n2376 DVSS.n2042 9.3005
R29674 DVSS.n2394 DVSS.n2041 9.3005
R29675 DVSS.n2396 DVSS.n2395 9.3005
R29676 DVSS.n2397 DVSS.n2040 9.3005
R29677 DVSS.n2400 DVSS.n2039 9.3005
R29678 DVSS.n2402 DVSS.n2401 9.3005
R29679 DVSS.n2403 DVSS.n2037 9.3005
R29680 DVSS.n2431 DVSS.n2430 9.3005
R29681 DVSS.n2429 DVSS.n2038 9.3005
R29682 DVSS.n2428 DVSS.n2427 9.3005
R29683 DVSS.n2404 DVSS.n2022 9.3005
R29684 DVSS.n2465 DVSS.n2023 9.3005
R29685 DVSS.n2466 DVSS.n2021 9.3005
R29686 DVSS.n2468 DVSS.n2467 9.3005
R29687 DVSS.n2469 DVSS.n2020 9.3005
R29688 DVSS.n2472 DVSS.n2471 9.3005
R29689 DVSS.n2477 DVSS.n2476 9.3005
R29690 DVSS.n2606 DVSS.n2605 9.3005
R29691 DVSS.n2613 DVSS.n2609 9.3005
R29692 DVSS.n2614 DVSS.n2612 9.3005
R29693 DVSS.n2619 DVSS.n2611 9.3005
R29694 DVSS.n2619 DVSS.n2618 9.3005
R29695 DVSS.n2610 DVSS.n2608 9.3005
R29696 DVSS.n2624 DVSS.n2623 9.3005
R29697 DVSS.n2585 DVSS.n2584 9.3005
R29698 DVSS.n2592 DVSS.n2588 9.3005
R29699 DVSS.n2593 DVSS.n2591 9.3005
R29700 DVSS.n2598 DVSS.n2590 9.3005
R29701 DVSS.n2598 DVSS.n2597 9.3005
R29702 DVSS.n2589 DVSS.n2587 9.3005
R29703 DVSS.n2603 DVSS.n2602 9.3005
R29704 DVSS.n2819 DVSS.n2818 9.3005
R29705 DVSS.n2822 DVSS.n2821 9.3005
R29706 DVSS.n2823 DVSS.n2554 9.3005
R29707 DVSS.n2828 DVSS.n2827 9.3005
R29708 DVSS.n2826 DVSS.n2555 9.3005
R29709 DVSS.n2825 DVSS.n2824 9.3005
R29710 DVSS.n2521 DVSS.n2520 9.3005
R29711 DVSS.n2839 DVSS.n2838 9.3005
R29712 DVSS.n2840 DVSS.n2518 9.3005
R29713 DVSS.n2848 DVSS.n2847 9.3005
R29714 DVSS.n2846 DVSS.n2519 9.3005
R29715 DVSS.n2843 DVSS.n2842 9.3005
R29716 DVSS.n2841 DVSS.n2507 9.3005
R29717 DVSS.n2859 DVSS.n2506 9.3005
R29718 DVSS.n2861 DVSS.n2860 9.3005
R29719 DVSS.n2862 DVSS.n2505 9.3005
R29720 DVSS.n2865 DVSS.n2504 9.3005
R29721 DVSS.n2867 DVSS.n2866 9.3005
R29722 DVSS.n2868 DVSS.n2502 9.3005
R29723 DVSS.n2896 DVSS.n2895 9.3005
R29724 DVSS.n2894 DVSS.n2503 9.3005
R29725 DVSS.n2893 DVSS.n2892 9.3005
R29726 DVSS.n2869 DVSS.n2487 9.3005
R29727 DVSS.n2930 DVSS.n2488 9.3005
R29728 DVSS.n2931 DVSS.n2486 9.3005
R29729 DVSS.n2933 DVSS.n2932 9.3005
R29730 DVSS.n2934 DVSS.n2485 9.3005
R29731 DVSS.n2936 DVSS.n2935 9.3005
R29732 DVSS.n2981 DVSS.n2980 9.3005
R29733 DVSS.n2996 DVSS.n2995 9.3005
R29734 DVSS.n3014 DVSS.n3013 9.3005
R29735 DVSS.n3024 DVSS.n3023 9.3005
R29736 DVSS.n3042 DVSS.n3041 9.3005
R29737 DVSS.n3057 DVSS.n3056 9.3005
R29738 DVSS.n3072 DVSS.n3071 9.3005
R29739 DVSS.n3087 DVSS.n3086 9.3005
R29740 DVSS.n3102 DVSS.n3101 9.3005
R29741 DVSS.n3117 DVSS.n3116 9.3005
R29742 DVSS.n3132 DVSS.n3131 9.3005
R29743 DVSS.n3156 DVSS.n3155 9.3005
R29744 DVSS.n3171 DVSS.n3170 9.3005
R29745 DVSS.n3186 DVSS.n3185 9.3005
R29746 DVSS.n3201 DVSS.n3200 9.3005
R29747 DVSS.n3216 DVSS.n3215 9.3005
R29748 DVSS.n3231 DVSS.n3230 9.3005
R29749 DVSS.n3246 DVSS.n3245 9.3005
R29750 DVSS.n3264 DVSS.n3263 9.3005
R29751 DVSS.n3274 DVSS.n3273 9.3005
R29752 DVSS.n3292 DVSS.n3291 9.3005
R29753 DVSS.n3307 DVSS.n3306 9.3005
R29754 DVSS.n3305 DVSS.n3304 9.3005
R29755 DVSS.n3272 DVSS.n3271 9.3005
R29756 DVSS.n3266 DVSS.n3265 9.3005
R29757 DVSS.n3233 DVSS.n3232 9.3005
R29758 DVSS.n3203 DVSS.n3202 9.3005
R29759 DVSS.n3173 DVSS.n3172 9.3005
R29760 DVSS.n3115 DVSS.n3114 9.3005
R29761 DVSS.n3085 DVSS.n3084 9.3005
R29762 DVSS.n3055 DVSS.n3054 9.3005
R29763 DVSS.n3022 DVSS.n3021 9.3005
R29764 DVSS.n3016 DVSS.n3015 9.3005
R29765 DVSS.n2983 DVSS.n2982 9.3005
R29766 DVSS.n2998 DVSS.n2997 9.3005
R29767 DVSS.n3040 DVSS.n3039 9.3005
R29768 DVSS.n3070 DVSS.n3069 9.3005
R29769 DVSS.n3100 DVSS.n3099 9.3005
R29770 DVSS.n3130 DVSS.n3129 9.3005
R29771 DVSS.n3158 DVSS.n3157 9.3005
R29772 DVSS.n3188 DVSS.n3187 9.3005
R29773 DVSS.n3218 DVSS.n3217 9.3005
R29774 DVSS.n3248 DVSS.n3247 9.3005
R29775 DVSS.n3290 DVSS.n3289 9.3005
R29776 DVSS.n3318 DVSS.n3317 9.3005
R29777 DVSS.n3317 DVSS.n3316 9.3005
R29778 DVSS.n3316 DVSS.n3315 9.3005
R29779 DVSS.n3288 DVSS.n3287 9.3005
R29780 DVSS.n3287 DVSS.n3286 9.3005
R29781 DVSS.n3286 DVSS.n3285 9.3005
R29782 DVSS.n3128 DVSS.n3127 9.3005
R29783 DVSS.n3127 DVSS.n3126 9.3005
R29784 DVSS.n3126 DVSS.n3125 9.3005
R29785 DVSS.n3098 DVSS.n3097 9.3005
R29786 DVSS.n3097 DVSS.n3096 9.3005
R29787 DVSS.n3096 DVSS.n3095 9.3005
R29788 DVSS.n3068 DVSS.n3067 9.3005
R29789 DVSS.n3067 DVSS.n3066 9.3005
R29790 DVSS.n3066 DVSS.n3065 9.3005
R29791 DVSS.n3038 DVSS.n3037 9.3005
R29792 DVSS.n3037 DVSS.n3036 9.3005
R29793 DVSS.n3036 DVSS.n3035 9.3005
R29794 DVSS.n2979 DVSS.n2978 9.3005
R29795 DVSS.n2978 DVSS.n2977 9.3005
R29796 DVSS.n2977 DVSS.n2976 9.3005
R29797 DVSS.n2994 DVSS.n2993 9.3005
R29798 DVSS.n2993 DVSS.n2992 9.3005
R29799 DVSS.n2992 DVSS.n2991 9.3005
R29800 DVSS.n3012 DVSS.n3011 9.3005
R29801 DVSS.n3011 DVSS.n3010 9.3005
R29802 DVSS.n3010 DVSS.n3009 9.3005
R29803 DVSS.n3053 DVSS.n3052 9.3005
R29804 DVSS.n3052 DVSS.n3051 9.3005
R29805 DVSS.n3051 DVSS.n3050 9.3005
R29806 DVSS.n3083 DVSS.n3082 9.3005
R29807 DVSS.n3082 DVSS.n3081 9.3005
R29808 DVSS.n3081 DVSS.n3080 9.3005
R29809 DVSS.n3113 DVSS.n3112 9.3005
R29810 DVSS.n3112 DVSS.n3111 9.3005
R29811 DVSS.n3111 DVSS.n3110 9.3005
R29812 DVSS.n3143 DVSS.n3142 9.3005
R29813 DVSS.n3142 DVSS.n3141 9.3005
R29814 DVSS.n3141 DVSS.n3140 9.3005
R29815 DVSS.n3154 DVSS.n3153 9.3005
R29816 DVSS.n3153 DVSS.n3152 9.3005
R29817 DVSS.n3152 DVSS.n3151 9.3005
R29818 DVSS.n3169 DVSS.n3168 9.3005
R29819 DVSS.n3168 DVSS.n3167 9.3005
R29820 DVSS.n3167 DVSS.n3166 9.3005
R29821 DVSS.n3184 DVSS.n3183 9.3005
R29822 DVSS.n3183 DVSS.n3182 9.3005
R29823 DVSS.n3182 DVSS.n3181 9.3005
R29824 DVSS.n3199 DVSS.n3198 9.3005
R29825 DVSS.n3198 DVSS.n3197 9.3005
R29826 DVSS.n3197 DVSS.n3196 9.3005
R29827 DVSS.n3214 DVSS.n3213 9.3005
R29828 DVSS.n3213 DVSS.n3212 9.3005
R29829 DVSS.n3212 DVSS.n3211 9.3005
R29830 DVSS.n3229 DVSS.n3228 9.3005
R29831 DVSS.n3228 DVSS.n3227 9.3005
R29832 DVSS.n3227 DVSS.n3226 9.3005
R29833 DVSS.n3244 DVSS.n3243 9.3005
R29834 DVSS.n3243 DVSS.n3242 9.3005
R29835 DVSS.n3242 DVSS.n3241 9.3005
R29836 DVSS.n3262 DVSS.n3261 9.3005
R29837 DVSS.n3261 DVSS.n3260 9.3005
R29838 DVSS.n3260 DVSS.n3259 9.3005
R29839 DVSS.n3303 DVSS.n3302 9.3005
R29840 DVSS.n3302 DVSS.n3301 9.3005
R29841 DVSS.n3301 DVSS.n3300 9.3005
R29842 DVSS.n3457 DVSS.n3456 9.3005
R29843 DVSS.n2008 DVSS.n2007 9.3005
R29844 DVSS.n5052 DVSS.n5051 9.3005
R29845 DVSS.n6518 DVSS.n6517 9.3005
R29846 DVSS.n6515 DVSS.n6514 9.3005
R29847 DVSS.n5205 DVSS.n5204 9.3005
R29848 DVSS.n5212 DVSS.n5208 9.3005
R29849 DVSS.n5213 DVSS.n5211 9.3005
R29850 DVSS.n5218 DVSS.n5210 9.3005
R29851 DVSS.n5218 DVSS.n5217 9.3005
R29852 DVSS.n5209 DVSS.n5207 9.3005
R29853 DVSS.n5223 DVSS.n5222 9.3005
R29854 DVSS.n5184 DVSS.n5183 9.3005
R29855 DVSS.n5191 DVSS.n5187 9.3005
R29856 DVSS.n5192 DVSS.n5190 9.3005
R29857 DVSS.n5197 DVSS.n5189 9.3005
R29858 DVSS.n5197 DVSS.n5196 9.3005
R29859 DVSS.n5188 DVSS.n5186 9.3005
R29860 DVSS.n5202 DVSS.n5201 9.3005
R29861 DVSS.n5418 DVSS.n5417 9.3005
R29862 DVSS.n5421 DVSS.n5420 9.3005
R29863 DVSS.n5422 DVSS.n5153 9.3005
R29864 DVSS.n5427 DVSS.n5426 9.3005
R29865 DVSS.n5425 DVSS.n5154 9.3005
R29866 DVSS.n5424 DVSS.n5423 9.3005
R29867 DVSS.n5120 DVSS.n5119 9.3005
R29868 DVSS.n5438 DVSS.n5437 9.3005
R29869 DVSS.n5439 DVSS.n5117 9.3005
R29870 DVSS.n5447 DVSS.n5446 9.3005
R29871 DVSS.n5445 DVSS.n5118 9.3005
R29872 DVSS.n5442 DVSS.n5441 9.3005
R29873 DVSS.n5440 DVSS.n5106 9.3005
R29874 DVSS.n5458 DVSS.n5105 9.3005
R29875 DVSS.n5460 DVSS.n5459 9.3005
R29876 DVSS.n5461 DVSS.n5104 9.3005
R29877 DVSS.n5464 DVSS.n5103 9.3005
R29878 DVSS.n5466 DVSS.n5465 9.3005
R29879 DVSS.n5467 DVSS.n5101 9.3005
R29880 DVSS.n5495 DVSS.n5494 9.3005
R29881 DVSS.n5493 DVSS.n5102 9.3005
R29882 DVSS.n5492 DVSS.n5491 9.3005
R29883 DVSS.n5468 DVSS.n5086 9.3005
R29884 DVSS.n5529 DVSS.n5087 9.3005
R29885 DVSS.n5530 DVSS.n5085 9.3005
R29886 DVSS.n5532 DVSS.n5531 9.3005
R29887 DVSS.n5533 DVSS.n5084 9.3005
R29888 DVSS.n5536 DVSS.n5535 9.3005
R29889 DVSS.n5541 DVSS.n5540 9.3005
R29890 DVSS.n5670 DVSS.n5669 9.3005
R29891 DVSS.n5677 DVSS.n5673 9.3005
R29892 DVSS.n5678 DVSS.n5676 9.3005
R29893 DVSS.n5683 DVSS.n5675 9.3005
R29894 DVSS.n5683 DVSS.n5682 9.3005
R29895 DVSS.n5674 DVSS.n5672 9.3005
R29896 DVSS.n5688 DVSS.n5687 9.3005
R29897 DVSS.n5649 DVSS.n5648 9.3005
R29898 DVSS.n5656 DVSS.n5652 9.3005
R29899 DVSS.n5657 DVSS.n5655 9.3005
R29900 DVSS.n5662 DVSS.n5654 9.3005
R29901 DVSS.n5662 DVSS.n5661 9.3005
R29902 DVSS.n5653 DVSS.n5651 9.3005
R29903 DVSS.n5667 DVSS.n5666 9.3005
R29904 DVSS.n5883 DVSS.n5882 9.3005
R29905 DVSS.n5886 DVSS.n5885 9.3005
R29906 DVSS.n5887 DVSS.n5618 9.3005
R29907 DVSS.n5892 DVSS.n5891 9.3005
R29908 DVSS.n5890 DVSS.n5619 9.3005
R29909 DVSS.n5889 DVSS.n5888 9.3005
R29910 DVSS.n5585 DVSS.n5584 9.3005
R29911 DVSS.n5903 DVSS.n5902 9.3005
R29912 DVSS.n5904 DVSS.n5582 9.3005
R29913 DVSS.n5912 DVSS.n5911 9.3005
R29914 DVSS.n5910 DVSS.n5583 9.3005
R29915 DVSS.n5907 DVSS.n5906 9.3005
R29916 DVSS.n5905 DVSS.n5571 9.3005
R29917 DVSS.n5923 DVSS.n5570 9.3005
R29918 DVSS.n5925 DVSS.n5924 9.3005
R29919 DVSS.n5926 DVSS.n5569 9.3005
R29920 DVSS.n5929 DVSS.n5568 9.3005
R29921 DVSS.n5931 DVSS.n5930 9.3005
R29922 DVSS.n5932 DVSS.n5566 9.3005
R29923 DVSS.n5960 DVSS.n5959 9.3005
R29924 DVSS.n5958 DVSS.n5567 9.3005
R29925 DVSS.n5957 DVSS.n5956 9.3005
R29926 DVSS.n5933 DVSS.n5551 9.3005
R29927 DVSS.n5994 DVSS.n5552 9.3005
R29928 DVSS.n5995 DVSS.n5550 9.3005
R29929 DVSS.n5997 DVSS.n5996 9.3005
R29930 DVSS.n5998 DVSS.n5549 9.3005
R29931 DVSS.n6000 DVSS.n5999 9.3005
R29932 DVSS.n6546 DVSS.n6545 9.3005
R29933 DVSS.n6544 DVSS.n6543 9.3005
R29934 DVSS.n6714 DVSS.n6713 9.3005
R29935 DVSS.n140 DVSS.n139 9.3005
R29936 DVSS.n147 DVSS.n143 9.3005
R29937 DVSS.n148 DVSS.n146 9.3005
R29938 DVSS.n153 DVSS.n145 9.3005
R29939 DVSS.n153 DVSS.n152 9.3005
R29940 DVSS.n144 DVSS.n142 9.3005
R29941 DVSS.n158 DVSS.n157 9.3005
R29942 DVSS.n119 DVSS.n118 9.3005
R29943 DVSS.n126 DVSS.n122 9.3005
R29944 DVSS.n127 DVSS.n125 9.3005
R29945 DVSS.n132 DVSS.n124 9.3005
R29946 DVSS.n132 DVSS.n131 9.3005
R29947 DVSS.n123 DVSS.n121 9.3005
R29948 DVSS.n137 DVSS.n136 9.3005
R29949 DVSS.n353 DVSS.n352 9.3005
R29950 DVSS.n356 DVSS.n355 9.3005
R29951 DVSS.n357 DVSS.n88 9.3005
R29952 DVSS.n362 DVSS.n361 9.3005
R29953 DVSS.n360 DVSS.n89 9.3005
R29954 DVSS.n359 DVSS.n358 9.3005
R29955 DVSS.n55 DVSS.n54 9.3005
R29956 DVSS.n373 DVSS.n372 9.3005
R29957 DVSS.n374 DVSS.n52 9.3005
R29958 DVSS.n382 DVSS.n381 9.3005
R29959 DVSS.n380 DVSS.n53 9.3005
R29960 DVSS.n377 DVSS.n376 9.3005
R29961 DVSS.n375 DVSS.n41 9.3005
R29962 DVSS.n393 DVSS.n40 9.3005
R29963 DVSS.n395 DVSS.n394 9.3005
R29964 DVSS.n396 DVSS.n39 9.3005
R29965 DVSS.n399 DVSS.n38 9.3005
R29966 DVSS.n401 DVSS.n400 9.3005
R29967 DVSS.n402 DVSS.n36 9.3005
R29968 DVSS.n430 DVSS.n429 9.3005
R29969 DVSS.n428 DVSS.n37 9.3005
R29970 DVSS.n427 DVSS.n426 9.3005
R29971 DVSS.n403 DVSS.n21 9.3005
R29972 DVSS.n464 DVSS.n22 9.3005
R29973 DVSS.n465 DVSS.n20 9.3005
R29974 DVSS.n467 DVSS.n466 9.3005
R29975 DVSS.n468 DVSS.n19 9.3005
R29976 DVSS.n471 DVSS.n470 9.3005
R29977 DVSS.n476 DVSS.n475 9.3005
R29978 DVSS.n605 DVSS.n604 9.3005
R29979 DVSS.n612 DVSS.n608 9.3005
R29980 DVSS.n613 DVSS.n611 9.3005
R29981 DVSS.n618 DVSS.n610 9.3005
R29982 DVSS.n618 DVSS.n617 9.3005
R29983 DVSS.n609 DVSS.n607 9.3005
R29984 DVSS.n623 DVSS.n622 9.3005
R29985 DVSS.n584 DVSS.n583 9.3005
R29986 DVSS.n591 DVSS.n587 9.3005
R29987 DVSS.n592 DVSS.n590 9.3005
R29988 DVSS.n597 DVSS.n589 9.3005
R29989 DVSS.n597 DVSS.n596 9.3005
R29990 DVSS.n588 DVSS.n586 9.3005
R29991 DVSS.n602 DVSS.n601 9.3005
R29992 DVSS.n818 DVSS.n817 9.3005
R29993 DVSS.n821 DVSS.n820 9.3005
R29994 DVSS.n822 DVSS.n553 9.3005
R29995 DVSS.n827 DVSS.n826 9.3005
R29996 DVSS.n825 DVSS.n554 9.3005
R29997 DVSS.n824 DVSS.n823 9.3005
R29998 DVSS.n520 DVSS.n519 9.3005
R29999 DVSS.n838 DVSS.n837 9.3005
R30000 DVSS.n839 DVSS.n517 9.3005
R30001 DVSS.n847 DVSS.n846 9.3005
R30002 DVSS.n845 DVSS.n518 9.3005
R30003 DVSS.n842 DVSS.n841 9.3005
R30004 DVSS.n840 DVSS.n506 9.3005
R30005 DVSS.n858 DVSS.n505 9.3005
R30006 DVSS.n860 DVSS.n859 9.3005
R30007 DVSS.n861 DVSS.n504 9.3005
R30008 DVSS.n864 DVSS.n503 9.3005
R30009 DVSS.n866 DVSS.n865 9.3005
R30010 DVSS.n867 DVSS.n501 9.3005
R30011 DVSS.n895 DVSS.n894 9.3005
R30012 DVSS.n893 DVSS.n502 9.3005
R30013 DVSS.n892 DVSS.n891 9.3005
R30014 DVSS.n868 DVSS.n486 9.3005
R30015 DVSS.n929 DVSS.n487 9.3005
R30016 DVSS.n930 DVSS.n485 9.3005
R30017 DVSS.n932 DVSS.n931 9.3005
R30018 DVSS.n933 DVSS.n484 9.3005
R30019 DVSS.n935 DVSS.n934 9.3005
R30020 DVSS.n1364 DVSS.n1363 9.3005
R30021 DVSS.n1379 DVSS.n1378 9.3005
R30022 DVSS.n1397 DVSS.n1396 9.3005
R30023 DVSS.n1407 DVSS.n1406 9.3005
R30024 DVSS.n1425 DVSS.n1424 9.3005
R30025 DVSS.n1440 DVSS.n1439 9.3005
R30026 DVSS.n1455 DVSS.n1454 9.3005
R30027 DVSS.n1470 DVSS.n1469 9.3005
R30028 DVSS.n1485 DVSS.n1484 9.3005
R30029 DVSS.n1500 DVSS.n1499 9.3005
R30030 DVSS.n1515 DVSS.n1514 9.3005
R30031 DVSS.n1539 DVSS.n1538 9.3005
R30032 DVSS.n1554 DVSS.n1553 9.3005
R30033 DVSS.n1569 DVSS.n1568 9.3005
R30034 DVSS.n1584 DVSS.n1583 9.3005
R30035 DVSS.n1599 DVSS.n1598 9.3005
R30036 DVSS.n1614 DVSS.n1613 9.3005
R30037 DVSS.n1629 DVSS.n1628 9.3005
R30038 DVSS.n1647 DVSS.n1646 9.3005
R30039 DVSS.n1657 DVSS.n1656 9.3005
R30040 DVSS.n1675 DVSS.n1674 9.3005
R30041 DVSS.n1690 DVSS.n1689 9.3005
R30042 DVSS.n1688 DVSS.n1687 9.3005
R30043 DVSS.n1655 DVSS.n1654 9.3005
R30044 DVSS.n1649 DVSS.n1648 9.3005
R30045 DVSS.n1616 DVSS.n1615 9.3005
R30046 DVSS.n1586 DVSS.n1585 9.3005
R30047 DVSS.n1556 DVSS.n1555 9.3005
R30048 DVSS.n1498 DVSS.n1497 9.3005
R30049 DVSS.n1468 DVSS.n1467 9.3005
R30050 DVSS.n1438 DVSS.n1437 9.3005
R30051 DVSS.n1405 DVSS.n1404 9.3005
R30052 DVSS.n1399 DVSS.n1398 9.3005
R30053 DVSS.n1366 DVSS.n1365 9.3005
R30054 DVSS.n1381 DVSS.n1380 9.3005
R30055 DVSS.n1423 DVSS.n1422 9.3005
R30056 DVSS.n1453 DVSS.n1452 9.3005
R30057 DVSS.n1483 DVSS.n1482 9.3005
R30058 DVSS.n1513 DVSS.n1512 9.3005
R30059 DVSS.n1541 DVSS.n1540 9.3005
R30060 DVSS.n1571 DVSS.n1570 9.3005
R30061 DVSS.n1601 DVSS.n1600 9.3005
R30062 DVSS.n1631 DVSS.n1630 9.3005
R30063 DVSS.n1673 DVSS.n1672 9.3005
R30064 DVSS.n1701 DVSS.n1700 9.3005
R30065 DVSS.n1700 DVSS.n1699 9.3005
R30066 DVSS.n1699 DVSS.n1698 9.3005
R30067 DVSS.n1671 DVSS.n1670 9.3005
R30068 DVSS.n1670 DVSS.n1669 9.3005
R30069 DVSS.n1669 DVSS.n1668 9.3005
R30070 DVSS.n1511 DVSS.n1510 9.3005
R30071 DVSS.n1510 DVSS.n1509 9.3005
R30072 DVSS.n1509 DVSS.n1508 9.3005
R30073 DVSS.n1481 DVSS.n1480 9.3005
R30074 DVSS.n1480 DVSS.n1479 9.3005
R30075 DVSS.n1479 DVSS.n1478 9.3005
R30076 DVSS.n1451 DVSS.n1450 9.3005
R30077 DVSS.n1450 DVSS.n1449 9.3005
R30078 DVSS.n1449 DVSS.n1448 9.3005
R30079 DVSS.n1421 DVSS.n1420 9.3005
R30080 DVSS.n1420 DVSS.n1419 9.3005
R30081 DVSS.n1419 DVSS.n1418 9.3005
R30082 DVSS.n1362 DVSS.n1361 9.3005
R30083 DVSS.n1361 DVSS.n1360 9.3005
R30084 DVSS.n1360 DVSS.n1359 9.3005
R30085 DVSS.n1377 DVSS.n1376 9.3005
R30086 DVSS.n1376 DVSS.n1375 9.3005
R30087 DVSS.n1375 DVSS.n1374 9.3005
R30088 DVSS.n1395 DVSS.n1394 9.3005
R30089 DVSS.n1394 DVSS.n1393 9.3005
R30090 DVSS.n1393 DVSS.n1392 9.3005
R30091 DVSS.n1436 DVSS.n1435 9.3005
R30092 DVSS.n1435 DVSS.n1434 9.3005
R30093 DVSS.n1434 DVSS.n1433 9.3005
R30094 DVSS.n1466 DVSS.n1465 9.3005
R30095 DVSS.n1465 DVSS.n1464 9.3005
R30096 DVSS.n1464 DVSS.n1463 9.3005
R30097 DVSS.n1496 DVSS.n1495 9.3005
R30098 DVSS.n1495 DVSS.n1494 9.3005
R30099 DVSS.n1494 DVSS.n1493 9.3005
R30100 DVSS.n1526 DVSS.n1525 9.3005
R30101 DVSS.n1525 DVSS.n1524 9.3005
R30102 DVSS.n1524 DVSS.n1523 9.3005
R30103 DVSS.n1537 DVSS.n1536 9.3005
R30104 DVSS.n1536 DVSS.n1535 9.3005
R30105 DVSS.n1535 DVSS.n1534 9.3005
R30106 DVSS.n1552 DVSS.n1551 9.3005
R30107 DVSS.n1551 DVSS.n1550 9.3005
R30108 DVSS.n1550 DVSS.n1549 9.3005
R30109 DVSS.n1567 DVSS.n1566 9.3005
R30110 DVSS.n1566 DVSS.n1565 9.3005
R30111 DVSS.n1565 DVSS.n1564 9.3005
R30112 DVSS.n1582 DVSS.n1581 9.3005
R30113 DVSS.n1581 DVSS.n1580 9.3005
R30114 DVSS.n1580 DVSS.n1579 9.3005
R30115 DVSS.n1597 DVSS.n1596 9.3005
R30116 DVSS.n1596 DVSS.n1595 9.3005
R30117 DVSS.n1595 DVSS.n1594 9.3005
R30118 DVSS.n1612 DVSS.n1611 9.3005
R30119 DVSS.n1611 DVSS.n1610 9.3005
R30120 DVSS.n1610 DVSS.n1609 9.3005
R30121 DVSS.n1627 DVSS.n1626 9.3005
R30122 DVSS.n1626 DVSS.n1625 9.3005
R30123 DVSS.n1625 DVSS.n1624 9.3005
R30124 DVSS.n1645 DVSS.n1644 9.3005
R30125 DVSS.n1644 DVSS.n1643 9.3005
R30126 DVSS.n1643 DVSS.n1642 9.3005
R30127 DVSS.n1686 DVSS.n1685 9.3005
R30128 DVSS.n1685 DVSS.n1684 9.3005
R30129 DVSS.n1684 DVSS.n1683 9.3005
R30130 DVSS.n6757 DVSS.n6756 9.3005
R30131 DVSS.n1840 DVSS.n1839 9.3005
R30132 DVSS.n3963 DVSS.n3681 9.26007
R30133 DVSS.n3964 DVSS.n3963 9.26007
R30134 DVSS.n3965 DVSS.n3964 9.26007
R30135 DVSS.n3984 DVSS.n3983 9.26007
R30136 DVSS.n3986 DVSS.n3984 9.26007
R30137 DVSS.n3986 DVSS.n3985 9.26007
R30138 DVSS.n3985 DVSS.n3626 9.26007
R30139 DVSS.n4031 DVSS.n3626 9.26007
R30140 DVSS.n4057 DVSS.n4033 9.26007
R30141 DVSS.n4057 DVSS.n4056 9.26007
R30142 DVSS.n4056 DVSS.n4055 9.26007
R30143 DVSS.n4428 DVSS.n4146 9.26007
R30144 DVSS.n4429 DVSS.n4428 9.26007
R30145 DVSS.n4430 DVSS.n4429 9.26007
R30146 DVSS.n4449 DVSS.n4448 9.26007
R30147 DVSS.n4451 DVSS.n4449 9.26007
R30148 DVSS.n4451 DVSS.n4450 9.26007
R30149 DVSS.n4450 DVSS.n4091 9.26007
R30150 DVSS.n4496 DVSS.n4091 9.26007
R30151 DVSS.n4522 DVSS.n4498 9.26007
R30152 DVSS.n4522 DVSS.n4521 9.26007
R30153 DVSS.n4521 DVSS.n4520 9.26007
R30154 DVSS.n2367 DVSS.n2085 9.26007
R30155 DVSS.n2368 DVSS.n2367 9.26007
R30156 DVSS.n2369 DVSS.n2368 9.26007
R30157 DVSS.n2388 DVSS.n2387 9.26007
R30158 DVSS.n2390 DVSS.n2388 9.26007
R30159 DVSS.n2390 DVSS.n2389 9.26007
R30160 DVSS.n2389 DVSS.n2030 9.26007
R30161 DVSS.n2435 DVSS.n2030 9.26007
R30162 DVSS.n2461 DVSS.n2437 9.26007
R30163 DVSS.n2461 DVSS.n2460 9.26007
R30164 DVSS.n2460 DVSS.n2459 9.26007
R30165 DVSS.n2832 DVSS.n2550 9.26007
R30166 DVSS.n2833 DVSS.n2832 9.26007
R30167 DVSS.n2834 DVSS.n2833 9.26007
R30168 DVSS.n2853 DVSS.n2852 9.26007
R30169 DVSS.n2855 DVSS.n2853 9.26007
R30170 DVSS.n2855 DVSS.n2854 9.26007
R30171 DVSS.n2854 DVSS.n2495 9.26007
R30172 DVSS.n2900 DVSS.n2495 9.26007
R30173 DVSS.n2926 DVSS.n2902 9.26007
R30174 DVSS.n2926 DVSS.n2925 9.26007
R30175 DVSS.n2925 DVSS.n2924 9.26007
R30176 DVSS.n5431 DVSS.n5149 9.26007
R30177 DVSS.n5432 DVSS.n5431 9.26007
R30178 DVSS.n5433 DVSS.n5432 9.26007
R30179 DVSS.n5452 DVSS.n5451 9.26007
R30180 DVSS.n5454 DVSS.n5452 9.26007
R30181 DVSS.n5454 DVSS.n5453 9.26007
R30182 DVSS.n5453 DVSS.n5094 9.26007
R30183 DVSS.n5499 DVSS.n5094 9.26007
R30184 DVSS.n5525 DVSS.n5501 9.26007
R30185 DVSS.n5525 DVSS.n5524 9.26007
R30186 DVSS.n5524 DVSS.n5523 9.26007
R30187 DVSS.n5896 DVSS.n5614 9.26007
R30188 DVSS.n5897 DVSS.n5896 9.26007
R30189 DVSS.n5898 DVSS.n5897 9.26007
R30190 DVSS.n5917 DVSS.n5916 9.26007
R30191 DVSS.n5919 DVSS.n5917 9.26007
R30192 DVSS.n5919 DVSS.n5918 9.26007
R30193 DVSS.n5918 DVSS.n5559 9.26007
R30194 DVSS.n5964 DVSS.n5559 9.26007
R30195 DVSS.n5990 DVSS.n5966 9.26007
R30196 DVSS.n5990 DVSS.n5989 9.26007
R30197 DVSS.n5989 DVSS.n5988 9.26007
R30198 DVSS.n366 DVSS.n84 9.26007
R30199 DVSS.n367 DVSS.n366 9.26007
R30200 DVSS.n368 DVSS.n367 9.26007
R30201 DVSS.n387 DVSS.n386 9.26007
R30202 DVSS.n389 DVSS.n387 9.26007
R30203 DVSS.n389 DVSS.n388 9.26007
R30204 DVSS.n388 DVSS.n29 9.26007
R30205 DVSS.n434 DVSS.n29 9.26007
R30206 DVSS.n460 DVSS.n436 9.26007
R30207 DVSS.n460 DVSS.n459 9.26007
R30208 DVSS.n459 DVSS.n458 9.26007
R30209 DVSS.n831 DVSS.n549 9.26007
R30210 DVSS.n832 DVSS.n831 9.26007
R30211 DVSS.n833 DVSS.n832 9.26007
R30212 DVSS.n852 DVSS.n851 9.26007
R30213 DVSS.n854 DVSS.n852 9.26007
R30214 DVSS.n854 DVSS.n853 9.26007
R30215 DVSS.n853 DVSS.n494 9.26007
R30216 DVSS.n899 DVSS.n494 9.26007
R30217 DVSS.n925 DVSS.n901 9.26007
R30218 DVSS.n925 DVSS.n924 9.26007
R30219 DVSS.n924 DVSS.n923 9.26007
R30220 DVSS.n1232 DVSS.n1231 9.15497
R30221 DVSS.n1231 DVSS.n1230 9.15497
R30222 DVSS.n1742 DVSS.n1741 9.15497
R30223 DVSS.n1745 DVSS.n1744 9.15497
R30224 DVSS.n1744 DVSS.n1743 9.15497
R30225 DVSS.n1750 DVSS.n1749 9.15497
R30226 DVSS.n1749 DVSS.n1748 9.15497
R30227 DVSS.n1757 DVSS.n1756 9.15497
R30228 DVSS.n1756 DVSS.n1755 9.15497
R30229 DVSS.n1761 DVSS.n1760 9.15497
R30230 DVSS.n1760 DVSS.n1759 9.15497
R30231 DVSS.n1765 DVSS.n1764 9.15497
R30232 DVSS.n1764 DVSS.n1763 9.15497
R30233 DVSS.n1769 DVSS.n1768 9.15497
R30234 DVSS.n1768 DVSS.n1767 9.15497
R30235 DVSS.n1773 DVSS.n1772 9.15497
R30236 DVSS.n1772 DVSS.n1771 9.15497
R30237 DVSS.n1777 DVSS.n1776 9.15497
R30238 DVSS.n1776 DVSS.n1775 9.15497
R30239 DVSS.n5068 DVSS.n5067 9.15497
R30240 DVSS.n5067 DVSS.n5066 9.15497
R30241 DVSS.n6691 DVSS.n6690 9.15497
R30242 DVSS.n6692 DVSS.n6691 9.15497
R30243 DVSS.n6684 DVSS.n6683 9.15497
R30244 DVSS.n6683 DVSS.n6682 9.15497
R30245 DVSS.n6680 DVSS.n6679 9.15497
R30246 DVSS.n6679 DVSS.n6678 9.15497
R30247 DVSS.n6675 DVSS.n6674 9.15497
R30248 DVSS.n6674 DVSS.n6673 9.15497
R30249 DVSS.n6667 DVSS.n6666 9.15497
R30250 DVSS.n6666 DVSS.n6665 9.15497
R30251 DVSS.n6662 DVSS.n6661 9.15497
R30252 DVSS.n6661 DVSS.n6660 9.15497
R30253 DVSS.n6658 DVSS.n6657 9.15497
R30254 DVSS.n6657 DVSS.n6656 9.15497
R30255 DVSS.n6720 DVSS.n6719 9.15497
R30256 DVSS.n6719 DVSS.n6718 9.15497
R30257 DVSS.n4954 DVSS.n4953 9.15497
R30258 DVSS.n4957 DVSS.n4956 9.15497
R30259 DVSS.n4956 DVSS.n4955 9.15497
R30260 DVSS.n4962 DVSS.n4961 9.15497
R30261 DVSS.n4961 DVSS.n4960 9.15497
R30262 DVSS.n4969 DVSS.n4968 9.15497
R30263 DVSS.n4968 DVSS.n4967 9.15497
R30264 DVSS.n4973 DVSS.n4972 9.15497
R30265 DVSS.n4972 DVSS.n4971 9.15497
R30266 DVSS.n4977 DVSS.n4976 9.15497
R30267 DVSS.n4976 DVSS.n4975 9.15497
R30268 DVSS.n4981 DVSS.n4980 9.15497
R30269 DVSS.n4980 DVSS.n4979 9.15497
R30270 DVSS.n4985 DVSS.n4984 9.15497
R30271 DVSS.n4984 DVSS.n4983 9.15497
R30272 DVSS.n4989 DVSS.n4988 9.15497
R30273 DVSS.n4988 DVSS.n4987 9.15497
R30274 DVSS.n1856 DVSS.n1855 9.15497
R30275 DVSS.n1855 DVSS.n1854 9.15497
R30276 DVSS.n6726 DVSS.n6725 9.15497
R30277 DVSS.n6727 DVSS.n6726 9.15497
R30278 DVSS.n3362 DVSS.n3361 9.15497
R30279 DVSS.n3360 DVSS.n3359 9.15497
R30280 DVSS.n3359 DVSS.n3358 9.15497
R30281 DVSS.n3367 DVSS.n3366 9.15497
R30282 DVSS.n3366 DVSS.n3365 9.15497
R30283 DVSS.n3374 DVSS.n3373 9.15497
R30284 DVSS.n3373 DVSS.n3372 9.15497
R30285 DVSS.n3378 DVSS.n3377 9.15497
R30286 DVSS.n3377 DVSS.n3376 9.15497
R30287 DVSS.n3382 DVSS.n3381 9.15497
R30288 DVSS.n3381 DVSS.n3380 9.15497
R30289 DVSS.n3386 DVSS.n3385 9.15497
R30290 DVSS.n3385 DVSS.n3384 9.15497
R30291 DVSS.n3390 DVSS.n3389 9.15497
R30292 DVSS.n3389 DVSS.n3388 9.15497
R30293 DVSS.n3394 DVSS.n3393 9.15497
R30294 DVSS.n3393 DVSS.n3392 9.15497
R30295 DVSS.n6737 DVSS.n6736 9.15497
R30296 DVSS.n3466 DVSS.n3465 9.15497
R30297 DVSS.n3465 DVSS.n3464 9.15497
R30298 DVSS.n3398 DVSS.n3397 9.15497
R30299 DVSS.n3397 DVSS.n3396 9.15497
R30300 DVSS.n3403 DVSS.n3402 9.15497
R30301 DVSS.n3402 DVSS.n3401 9.15497
R30302 DVSS.n3408 DVSS.n3407 9.15497
R30303 DVSS.n3407 DVSS.n3406 9.15497
R30304 DVSS.n3415 DVSS.n3414 9.15497
R30305 DVSS.n3414 DVSS.n3413 9.15497
R30306 DVSS.n3419 DVSS.n3418 9.15497
R30307 DVSS.n3418 DVSS.n3417 9.15497
R30308 DVSS.n3424 DVSS.n3423 9.15497
R30309 DVSS.n3432 DVSS.n3431 9.15497
R30310 DVSS.n3436 DVSS.n3435 9.15497
R30311 DVSS.n3440 DVSS.n3439 9.15497
R30312 DVSS.n3439 DVSS.n3438 9.15497
R30313 DVSS.n3446 DVSS.n3445 9.15497
R30314 DVSS.n3445 DVSS.n3444 9.15497
R30315 DVSS.n3450 DVSS.n3449 9.15497
R30316 DVSS.n3449 DVSS.n3448 9.15497
R30317 DVSS.n3456 DVSS.n3455 9.15497
R30318 DVSS.n3455 DVSS.n3454 9.15497
R30319 DVSS.n6731 DVSS.n6730 9.15497
R30320 DVSS.n6730 DVSS.n6729 9.15497
R30321 DVSS.n1895 DVSS.n1894 9.15497
R30322 DVSS.n1894 DVSS.n1893 9.15497
R30323 DVSS.n1902 DVSS.n1901 9.15497
R30324 DVSS.n1903 DVSS.n1902 9.15497
R30325 DVSS.n1906 DVSS.n1905 9.15497
R30326 DVSS.n1905 DVSS.n1904 9.15497
R30327 DVSS.n1910 DVSS.n1909 9.15497
R30328 DVSS.n1909 DVSS.n1908 9.15497
R30329 DVSS.n1914 DVSS.n1913 9.15497
R30330 DVSS.n1913 DVSS.n1912 9.15497
R30331 DVSS.n1918 DVSS.n1917 9.15497
R30332 DVSS.n1917 DVSS.n1916 9.15497
R30333 DVSS.n1925 DVSS.n1924 9.15497
R30334 DVSS.n1930 DVSS.n1929 9.15497
R30335 DVSS.n1929 DVSS.n1928 9.15497
R30336 DVSS.n1934 DVSS.n1933 9.15497
R30337 DVSS.n1933 DVSS.n1932 9.15497
R30338 DVSS.n1942 DVSS.n1941 9.15497
R30339 DVSS.n1947 DVSS.n1946 9.15497
R30340 DVSS.n1946 DVSS.n1945 9.15497
R30341 DVSS.n1951 DVSS.n1950 9.15497
R30342 DVSS.n1950 DVSS.n1949 9.15497
R30343 DVSS.n1958 DVSS.n1957 9.15497
R30344 DVSS.n1963 DVSS.n1962 9.15497
R30345 DVSS.n1962 DVSS.n1961 9.15497
R30346 DVSS.n1967 DVSS.n1966 9.15497
R30347 DVSS.n1966 DVSS.n1965 9.15497
R30348 DVSS.n1971 DVSS.n1970 9.15497
R30349 DVSS.n1970 DVSS.n1969 9.15497
R30350 DVSS.n1976 DVSS.n1975 9.15497
R30351 DVSS.n1975 DVSS.n1974 9.15497
R30352 DVSS.n1985 DVSS.n1984 9.15497
R30353 DVSS.n1984 DVSS.n1983 9.15497
R30354 DVSS.n1989 DVSS.n1988 9.15497
R30355 DVSS.n1988 DVSS.n1987 9.15497
R30356 DVSS.n1994 DVSS.n1993 9.15497
R30357 DVSS.n1993 DVSS.n1992 9.15497
R30358 DVSS.n1997 DVSS.n1996 9.15497
R30359 DVSS.n1996 DVSS.n1995 9.15497
R30360 DVSS.n2001 DVSS.n2000 9.15497
R30361 DVSS.n2000 DVSS.n1999 9.15497
R30362 DVSS.n2007 DVSS.n2006 9.15497
R30363 DVSS.n2006 DVSS.n2005 9.15497
R30364 DVSS.n3475 DVSS.n3474 9.15497
R30365 DVSS.n3476 DVSS.n3475 9.15497
R30366 DVSS.n3480 DVSS.n3479 9.15497
R30367 DVSS.n3479 DVSS.n3478 9.15497
R30368 DVSS.n5061 DVSS.n5060 9.15497
R30369 DVSS.n5060 DVSS.n5059 9.15497
R30370 DVSS.n4993 DVSS.n4992 9.15497
R30371 DVSS.n4992 DVSS.n4991 9.15497
R30372 DVSS.n4998 DVSS.n4997 9.15497
R30373 DVSS.n4997 DVSS.n4996 9.15497
R30374 DVSS.n5003 DVSS.n5002 9.15497
R30375 DVSS.n5002 DVSS.n5001 9.15497
R30376 DVSS.n5010 DVSS.n5009 9.15497
R30377 DVSS.n5009 DVSS.n5008 9.15497
R30378 DVSS.n5014 DVSS.n5013 9.15497
R30379 DVSS.n5013 DVSS.n5012 9.15497
R30380 DVSS.n5019 DVSS.n5018 9.15497
R30381 DVSS.n5027 DVSS.n5026 9.15497
R30382 DVSS.n5031 DVSS.n5030 9.15497
R30383 DVSS.n5035 DVSS.n5034 9.15497
R30384 DVSS.n5034 DVSS.n5033 9.15497
R30385 DVSS.n5041 DVSS.n5040 9.15497
R30386 DVSS.n5040 DVSS.n5039 9.15497
R30387 DVSS.n5045 DVSS.n5044 9.15497
R30388 DVSS.n5044 DVSS.n5043 9.15497
R30389 DVSS.n5051 DVSS.n5050 9.15497
R30390 DVSS.n5050 DVSS.n5049 9.15497
R30391 DVSS.n6643 DVSS.n6642 9.15497
R30392 DVSS.n6644 DVSS.n6643 9.15497
R30393 DVSS.n6527 DVSS.n6526 9.15497
R30394 DVSS.n6526 DVSS.n6525 9.15497
R30395 DVSS.n6422 DVSS.n6421 9.15497
R30396 DVSS.n6425 DVSS.n6424 9.15497
R30397 DVSS.n6424 DVSS.n6423 9.15497
R30398 DVSS.n6430 DVSS.n6429 9.15497
R30399 DVSS.n6429 DVSS.n6428 9.15497
R30400 DVSS.n6437 DVSS.n6436 9.15497
R30401 DVSS.n6436 DVSS.n6435 9.15497
R30402 DVSS.n6441 DVSS.n6440 9.15497
R30403 DVSS.n6440 DVSS.n6439 9.15497
R30404 DVSS.n6445 DVSS.n6444 9.15497
R30405 DVSS.n6444 DVSS.n6443 9.15497
R30406 DVSS.n6449 DVSS.n6448 9.15497
R30407 DVSS.n6448 DVSS.n6447 9.15497
R30408 DVSS.n6453 DVSS.n6452 9.15497
R30409 DVSS.n6452 DVSS.n6451 9.15497
R30410 DVSS.n6457 DVSS.n6456 9.15497
R30411 DVSS.n6456 DVSS.n6455 9.15497
R30412 DVSS.n6461 DVSS.n6460 9.15497
R30413 DVSS.n6460 DVSS.n6459 9.15497
R30414 DVSS.n6466 DVSS.n6465 9.15497
R30415 DVSS.n6465 DVSS.n6464 9.15497
R30416 DVSS.n6471 DVSS.n6470 9.15497
R30417 DVSS.n6470 DVSS.n6469 9.15497
R30418 DVSS.n6478 DVSS.n6477 9.15497
R30419 DVSS.n6477 DVSS.n6476 9.15497
R30420 DVSS.n6482 DVSS.n6481 9.15497
R30421 DVSS.n6481 DVSS.n6480 9.15497
R30422 DVSS.n6487 DVSS.n6486 9.15497
R30423 DVSS.n6486 DVSS.n6485 9.15497
R30424 DVSS.n6495 DVSS.n6494 9.15497
R30425 DVSS.n6494 DVSS.n6493 9.15497
R30426 DVSS.n6499 DVSS.n6498 9.15497
R30427 DVSS.n6498 DVSS.n6497 9.15497
R30428 DVSS.n6504 DVSS.n6503 9.15497
R30429 DVSS.n6503 DVSS.n6502 9.15497
R30430 DVSS.n6509 DVSS.n6508 9.15497
R30431 DVSS.n6512 DVSS.n6511 9.15497
R30432 DVSS.n6517 DVSS.n6516 9.15497
R30433 DVSS.n6639 DVSS.n6638 9.15497
R30434 DVSS.n6638 DVSS.n6637 9.15497
R30435 DVSS.n6635 DVSS.n6634 9.15497
R30436 DVSS.n6634 DVSS.n6633 9.15497
R30437 DVSS.n6631 DVSS.n6630 9.15497
R30438 DVSS.n6630 DVSS.n6629 9.15497
R30439 DVSS.n6626 DVSS.n6625 9.15497
R30440 DVSS.n6621 DVSS.n6620 9.15497
R30441 DVSS.n6620 DVSS.n6619 9.15497
R30442 DVSS.n6617 DVSS.n6616 9.15497
R30443 DVSS.n6616 DVSS.n6615 9.15497
R30444 DVSS.n6609 DVSS.n6608 9.15497
R30445 DVSS.n6604 DVSS.n6603 9.15497
R30446 DVSS.n6603 DVSS.n6602 9.15497
R30447 DVSS.n6600 DVSS.n6599 9.15497
R30448 DVSS.n6599 DVSS.n6598 9.15497
R30449 DVSS.n6593 DVSS.n6592 9.15497
R30450 DVSS.n6592 DVSS.n6591 9.15497
R30451 DVSS.n6588 DVSS.n6587 9.15497
R30452 DVSS.n6587 DVSS.n6586 9.15497
R30453 DVSS.n6584 DVSS.n6583 9.15497
R30454 DVSS.n6583 DVSS.n6582 9.15497
R30455 DVSS.n6580 DVSS.n6579 9.15497
R30456 DVSS.n6579 DVSS.n6578 9.15497
R30457 DVSS.n6575 DVSS.n6574 9.15497
R30458 DVSS.n6574 DVSS.n6573 9.15497
R30459 DVSS.n6566 DVSS.n6565 9.15497
R30460 DVSS.n6565 DVSS.n6564 9.15497
R30461 DVSS.n6562 DVSS.n6561 9.15497
R30462 DVSS.n6561 DVSS.n6560 9.15497
R30463 DVSS.n6558 DVSS.n5075 9.15497
R30464 DVSS.n5075 DVSS.n5074 9.15497
R30465 DVSS.n6557 DVSS.n6556 9.15497
R30466 DVSS.n6556 DVSS.n6555 9.15497
R30467 DVSS.n6552 DVSS.n6551 9.15497
R30468 DVSS.n6551 DVSS.n6550 9.15497
R30469 DVSS.n6543 DVSS.n6542 9.15497
R30470 DVSS.n6542 DVSS.n6541 9.15497
R30471 DVSS.n6535 DVSS.n6534 9.15497
R30472 DVSS.n6534 DVSS.n6533 9.15497
R30473 DVSS.n6702 DVSS.n6701 9.15497
R30474 DVSS.n6696 DVSS.n6695 9.15497
R30475 DVSS.n6695 DVSS.n6694 9.15497
R30476 DVSS.n6653 DVSS.n6652 9.15497
R30477 DVSS.n6652 DVSS.n6651 9.15497
R30478 DVSS.n6647 DVSS.n6646 9.15497
R30479 DVSS.n6646 DVSS.n6645 9.15497
R30480 DVSS.n6715 DVSS.n6714 9.15497
R30481 DVSS.n6716 DVSS.n6715 9.15497
R30482 DVSS.n3513 DVSS.n3512 9.15497
R30483 DVSS.n3512 DVSS.n3511 9.15497
R30484 DVSS.n3517 DVSS.n3516 9.15497
R30485 DVSS.n3516 DVSS.n3515 9.15497
R30486 DVSS.n3521 DVSS.n3520 9.15497
R30487 DVSS.n3520 DVSS.n3519 9.15497
R30488 DVSS.n3528 DVSS.n3527 9.15497
R30489 DVSS.n3533 DVSS.n3532 9.15497
R30490 DVSS.n3532 DVSS.n3531 9.15497
R30491 DVSS.n3537 DVSS.n3536 9.15497
R30492 DVSS.n3536 DVSS.n3535 9.15497
R30493 DVSS.n3545 DVSS.n3544 9.15497
R30494 DVSS.n3550 DVSS.n3549 9.15497
R30495 DVSS.n3549 DVSS.n3548 9.15497
R30496 DVSS.n3554 DVSS.n3553 9.15497
R30497 DVSS.n3553 DVSS.n3552 9.15497
R30498 DVSS.n3561 DVSS.n3560 9.15497
R30499 DVSS.n3566 DVSS.n3565 9.15497
R30500 DVSS.n3565 DVSS.n3564 9.15497
R30501 DVSS.n3570 DVSS.n3569 9.15497
R30502 DVSS.n3569 DVSS.n3568 9.15497
R30503 DVSS.n3574 DVSS.n3573 9.15497
R30504 DVSS.n3573 DVSS.n3572 9.15497
R30505 DVSS.n3579 DVSS.n3578 9.15497
R30506 DVSS.n3578 DVSS.n3577 9.15497
R30507 DVSS.n3588 DVSS.n3587 9.15497
R30508 DVSS.n3587 DVSS.n3586 9.15497
R30509 DVSS.n3592 DVSS.n3591 9.15497
R30510 DVSS.n3591 DVSS.n3590 9.15497
R30511 DVSS.n3599 DVSS.n3595 9.15497
R30512 DVSS.n3595 DVSS.n3594 9.15497
R30513 DVSS.n3598 DVSS.n3597 9.15497
R30514 DVSS.n3597 DVSS.n3596 9.15497
R30515 DVSS.n3604 DVSS.n3603 9.15497
R30516 DVSS.n3603 DVSS.n3602 9.15497
R30517 DVSS.n3508 DVSS.n3507 9.15497
R30518 DVSS.n3507 DVSS.n3506 9.15497
R30519 DVSS.n3488 DVSS.n3487 9.15497
R30520 DVSS.n3487 DVSS.n3486 9.15497
R30521 DVSS.n3492 DVSS.n3491 9.15497
R30522 DVSS.n3491 DVSS.n3490 9.15497
R30523 DVSS.n3497 DVSS.n3496 9.15497
R30524 DVSS.n3496 DVSS.n3495 9.15497
R30525 DVSS.n3504 DVSS.n3503 9.15497
R30526 DVSS.n3505 DVSS.n3504 9.15497
R30527 DVSS.n1888 DVSS.n1887 9.15497
R30528 DVSS.n1887 DVSS.n1886 9.15497
R30529 DVSS.n1884 DVSS.n1883 9.15497
R30530 DVSS.n1883 DVSS.n1882 9.15497
R30531 DVSS.n1879 DVSS.n1878 9.15497
R30532 DVSS.n1878 DVSS.n1877 9.15497
R30533 DVSS.n1871 DVSS.n1870 9.15497
R30534 DVSS.n1870 DVSS.n1869 9.15497
R30535 DVSS.n1866 DVSS.n1865 9.15497
R30536 DVSS.n1865 DVSS.n1864 9.15497
R30537 DVSS.n1862 DVSS.n1861 9.15497
R30538 DVSS.n1861 DVSS.n1860 9.15497
R30539 DVSS.n6751 DVSS.n6750 9.15497
R30540 DVSS.n6752 DVSS.n6751 9.15497
R30541 DVSS.n6 DVSS.n5 9.15497
R30542 DVSS.n5 DVSS.n4 9.15497
R30543 DVSS.n6875 DVSS.n6874 9.15497
R30544 DVSS.n6874 DVSS.n6873 9.15497
R30545 DVSS.n6871 DVSS.n6870 9.15497
R30546 DVSS.n6870 DVSS.n6869 9.15497
R30547 DVSS.n6866 DVSS.n6865 9.15497
R30548 DVSS.n6865 DVSS.n6864 9.15497
R30549 DVSS.n6861 DVSS.n6860 9.15497
R30550 DVSS.n6860 DVSS.n6859 9.15497
R30551 DVSS.n6857 DVSS.n6856 9.15497
R30552 DVSS.n6858 DVSS.n6857 9.15497
R30553 DVSS.n6852 DVSS.n6851 9.15497
R30554 DVSS.n6851 DVSS.n6850 9.15497
R30555 DVSS.n6848 DVSS.n6847 9.15497
R30556 DVSS.n6847 DVSS.n6846 9.15497
R30557 DVSS.n6844 DVSS.n6843 9.15497
R30558 DVSS.n6843 DVSS.n6842 9.15497
R30559 DVSS.n6837 DVSS.n6836 9.15497
R30560 DVSS.n6832 DVSS.n6831 9.15497
R30561 DVSS.n6831 DVSS.n6830 9.15497
R30562 DVSS.n6828 DVSS.n6827 9.15497
R30563 DVSS.n6827 DVSS.n6826 9.15497
R30564 DVSS.n6820 DVSS.n6819 9.15497
R30565 DVSS.n6815 DVSS.n6814 9.15497
R30566 DVSS.n6814 DVSS.n6813 9.15497
R30567 DVSS.n6811 DVSS.n6810 9.15497
R30568 DVSS.n6810 DVSS.n6809 9.15497
R30569 DVSS.n6806 DVSS.n6805 9.15497
R30570 DVSS.n6800 DVSS.n6799 9.15497
R30571 DVSS.n6799 DVSS.n6798 9.15497
R30572 DVSS.n6796 DVSS.n6795 9.15497
R30573 DVSS.n6795 DVSS.n6794 9.15497
R30574 DVSS.n6792 DVSS.n6791 9.15497
R30575 DVSS.n6791 DVSS.n6790 9.15497
R30576 DVSS.n6787 DVSS.n6786 9.15497
R30577 DVSS.n6786 DVSS.n6785 9.15497
R30578 DVSS.n6778 DVSS.n6777 9.15497
R30579 DVSS.n6777 DVSS.n6776 9.15497
R30580 DVSS.n6774 DVSS.n6773 9.15497
R30581 DVSS.n6773 DVSS.n6772 9.15497
R30582 DVSS.n6770 DVSS.n6769 9.15497
R30583 DVSS.n6769 DVSS.n6768 9.15497
R30584 DVSS.n6767 DVSS.n6766 9.15497
R30585 DVSS.n6766 DVSS.n6765 9.15497
R30586 DVSS.n6762 DVSS.n6761 9.15497
R30587 DVSS.n6761 DVSS.n6760 9.15497
R30588 DVSS.n6756 DVSS.n6755 9.15497
R30589 DVSS.n6755 DVSS.n6754 9.15497
R30590 DVSS.n1849 DVSS.n1848 9.15497
R30591 DVSS.n1848 DVSS.n1847 9.15497
R30592 DVSS.n1781 DVSS.n1780 9.15497
R30593 DVSS.n1780 DVSS.n1779 9.15497
R30594 DVSS.n1786 DVSS.n1785 9.15497
R30595 DVSS.n1785 DVSS.n1784 9.15497
R30596 DVSS.n1791 DVSS.n1790 9.15497
R30597 DVSS.n1790 DVSS.n1789 9.15497
R30598 DVSS.n1798 DVSS.n1797 9.15497
R30599 DVSS.n1797 DVSS.n1796 9.15497
R30600 DVSS.n1802 DVSS.n1801 9.15497
R30601 DVSS.n1801 DVSS.n1800 9.15497
R30602 DVSS.n1807 DVSS.n1806 9.15497
R30603 DVSS.n1815 DVSS.n1814 9.15497
R30604 DVSS.n1819 DVSS.n1818 9.15497
R30605 DVSS.n1823 DVSS.n1822 9.15497
R30606 DVSS.n1822 DVSS.n1821 9.15497
R30607 DVSS.n1829 DVSS.n1828 9.15497
R30608 DVSS.n1828 DVSS.n1827 9.15497
R30609 DVSS.n1833 DVSS.n1832 9.15497
R30610 DVSS.n1832 DVSS.n1831 9.15497
R30611 DVSS.n1839 DVSS.n1838 9.15497
R30612 DVSS.n1838 DVSS.n1837 9.15497
R30613 DVSS.n1328 DVSS.n1327 9.15497
R30614 DVSS.n1049 DVSS.n1048 9.15497
R30615 DVSS.n1045 DVSS.n1044 9.15497
R30616 DVSS.n1033 DVSS.n1032 9.15497
R30617 DVSS.n1029 DVSS.n1028 9.15497
R30618 DVSS.n1025 DVSS.n1024 9.15497
R30619 DVSS.n1017 DVSS.n1016 9.15497
R30620 DVSS.n1036 DVSS.n1035 9.15497
R30621 DVSS.n1042 DVSS.n1041 9.15497
R30622 DVSS.n1014 DVSS.n1013 9.15497
R30623 DVSS.n968 DVSS.n967 9.15497
R30624 DVSS.n975 DVSS.n974 9.15497
R30625 DVSS.n978 DVSS.n977 9.15497
R30626 DVSS.n982 DVSS.n981 9.15497
R30627 DVSS.n985 DVSS.n984 9.15497
R30628 DVSS.n989 DVSS.n988 9.15497
R30629 DVSS.n992 DVSS.n991 9.15497
R30630 DVSS.n996 DVSS.n995 9.15497
R30631 DVSS.n999 DVSS.n998 9.15497
R30632 DVSS.n1003 DVSS.n1002 9.15497
R30633 DVSS.n1010 DVSS.n1009 9.15497
R30634 DVSS.n1059 DVSS.n1058 9.15497
R30635 DVSS.n1057 DVSS.n1056 9.15497
R30636 DVSS.n1094 DVSS.n1093 9.15497
R30637 DVSS.n1092 DVSS.n1091 9.15497
R30638 DVSS.n1100 DVSS.n1099 9.15497
R30639 DVSS.n1097 DVSS.n1096 9.15497
R30640 DVSS.n1106 DVSS.n1105 9.15497
R30641 DVSS.n1103 DVSS.n1102 9.15497
R30642 DVSS.n1089 DVSS.n1088 9.15497
R30643 DVSS.n1052 DVSS.n1051 9.15497
R30644 DVSS.n1069 DVSS.n1068 9.15497
R30645 DVSS.n1072 DVSS.n1071 9.15497
R30646 DVSS.n1076 DVSS.n1075 9.15497
R30647 DVSS.n1082 DVSS.n1081 9.15497
R30648 DVSS.n1086 DVSS.n1085 9.15497
R30649 DVSS.n1221 DVSS.n1220 9.15497
R30650 DVSS.n1220 DVSS.n1219 9.15497
R30651 DVSS.n1225 DVSS.n1224 9.15497
R30652 DVSS.n1216 DVSS.n1215 9.15497
R30653 DVSS.n1212 DVSS.n1211 9.15497
R30654 DVSS.n1209 DVSS.n1208 9.15497
R30655 DVSS.n1205 DVSS.n1204 9.15497
R30656 DVSS.n1202 DVSS.n1201 9.15497
R30657 DVSS.n1196 DVSS.n1195 9.15497
R30658 DVSS.n1192 DVSS.n1191 9.15497
R30659 DVSS.n1188 DVSS.n1187 9.15497
R30660 DVSS.n1185 DVSS.n1184 9.15497
R30661 DVSS.n1178 DVSS.n1177 9.15497
R30662 DVSS.n1175 DVSS.n1174 9.15497
R30663 DVSS.n1170 DVSS.n1169 9.15497
R30664 DVSS.n1164 DVSS.n1163 9.15497
R30665 DVSS.n1218 DVSS.n1217 9.15497
R30666 DVSS.n1236 DVSS.n1235 9.15497
R30667 DVSS.n1235 DVSS.n1234 9.15497
R30668 DVSS.n1240 DVSS.n1239 9.15497
R30669 DVSS.n1239 DVSS.n1238 9.15497
R30670 DVSS.n1245 DVSS.n1244 9.15497
R30671 DVSS.n1244 DVSS.n1243 9.15497
R30672 DVSS.n1249 DVSS.n1248 9.15497
R30673 DVSS.n1248 DVSS.n1247 9.15497
R30674 DVSS.n1253 DVSS.n1252 9.15497
R30675 DVSS.n1252 DVSS.n1251 9.15497
R30676 DVSS.n1257 DVSS.n1256 9.15497
R30677 DVSS.n1256 DVSS.n1255 9.15497
R30678 DVSS.n1266 DVSS.n1265 9.15497
R30679 DVSS.n1265 DVSS.n1264 9.15497
R30680 DVSS.n1271 DVSS.n1270 9.15497
R30681 DVSS.n1270 DVSS.n1269 9.15497
R30682 DVSS.n1275 DVSS.n1274 9.15497
R30683 DVSS.n1278 DVSS.n1277 9.15497
R30684 DVSS.n1282 DVSS.n1281 9.15497
R30685 DVSS.n1287 DVSS.n1286 9.15497
R30686 DVSS.n1291 DVSS.n1290 9.15497
R30687 DVSS.n1295 DVSS.n1294 9.15497
R30688 DVSS.n1303 DVSS.n1302 9.15497
R30689 DVSS.n1306 DVSS.n1305 9.15497
R30690 DVSS.n1311 DVSS.n1310 9.15497
R30691 DVSS.n1317 DVSS.n1316 9.15497
R30692 DVSS.n1324 DVSS.n1323 9.15497
R30693 DVSS.n1327 DVSS.n1326 9.15497
R30694 DVSS.n1341 DVSS.n1340 9.15497
R30695 DVSS.n1342 DVSS.n1341 9.15497
R30696 DVSS.n1334 DVSS.n1333 9.15497
R30697 DVSS.n1154 DVSS.n1153 9.15497
R30698 DVSS.n1151 DVSS.n1150 9.15497
R30699 DVSS.n1146 DVSS.n1145 9.15497
R30700 DVSS.n1138 DVSS.n1137 9.15497
R30701 DVSS.n1134 DVSS.n1133 9.15497
R30702 DVSS.n3519 DVSS.t47 9.02059
R30703 DVSS.n6629 DVSS.t101 9.02059
R30704 DVSS.n4069 DVSS.n3615 9.01392
R30705 DVSS.n3623 DVSS.n3614 9.01392
R30706 DVSS.n4060 DVSS.n4059 9.01392
R30707 DVSS.n3621 DVSS.n3620 9.01392
R30708 DVSS.n4029 DVSS.n4028 9.01392
R30709 DVSS.n3631 DVSS.n3629 9.01392
R30710 DVSS.n3641 DVSS.n3640 9.01392
R30711 DVSS.n3989 DVSS.n3988 9.01392
R30712 DVSS.n3647 DVSS.n3639 9.01392
R30713 DVSS.n3981 DVSS.n3980 9.01392
R30714 DVSS.n3968 DVSS.n3967 9.01392
R30715 DVSS.n3679 DVSS.n3678 9.01392
R30716 DVSS.n3961 DVSS.n3960 9.01392
R30717 DVSS.n3684 DVSS.n3683 9.01392
R30718 DVSS.n4533 DVSS.n4080 9.01392
R30719 DVSS.n4088 DVSS.n4079 9.01392
R30720 DVSS.n4525 DVSS.n4524 9.01392
R30721 DVSS.n4086 DVSS.n4085 9.01392
R30722 DVSS.n4494 DVSS.n4493 9.01392
R30723 DVSS.n4096 DVSS.n4094 9.01392
R30724 DVSS.n4106 DVSS.n4105 9.01392
R30725 DVSS.n4454 DVSS.n4453 9.01392
R30726 DVSS.n4112 DVSS.n4104 9.01392
R30727 DVSS.n4446 DVSS.n4445 9.01392
R30728 DVSS.n4433 DVSS.n4432 9.01392
R30729 DVSS.n4144 DVSS.n4143 9.01392
R30730 DVSS.n4426 DVSS.n4425 9.01392
R30731 DVSS.n4149 DVSS.n4148 9.01392
R30732 DVSS.n2473 DVSS.n2019 9.01392
R30733 DVSS.n2027 DVSS.n2018 9.01392
R30734 DVSS.n2464 DVSS.n2463 9.01392
R30735 DVSS.n2025 DVSS.n2024 9.01392
R30736 DVSS.n2433 DVSS.n2432 9.01392
R30737 DVSS.n2035 DVSS.n2033 9.01392
R30738 DVSS.n2045 DVSS.n2044 9.01392
R30739 DVSS.n2393 DVSS.n2392 9.01392
R30740 DVSS.n2051 DVSS.n2043 9.01392
R30741 DVSS.n2385 DVSS.n2384 9.01392
R30742 DVSS.n2372 DVSS.n2371 9.01392
R30743 DVSS.n2083 DVSS.n2082 9.01392
R30744 DVSS.n2365 DVSS.n2364 9.01392
R30745 DVSS.n2088 DVSS.n2087 9.01392
R30746 DVSS.n2937 DVSS.n2484 9.01392
R30747 DVSS.n2492 DVSS.n2483 9.01392
R30748 DVSS.n2929 DVSS.n2928 9.01392
R30749 DVSS.n2490 DVSS.n2489 9.01392
R30750 DVSS.n2898 DVSS.n2897 9.01392
R30751 DVSS.n2500 DVSS.n2498 9.01392
R30752 DVSS.n2510 DVSS.n2509 9.01392
R30753 DVSS.n2858 DVSS.n2857 9.01392
R30754 DVSS.n2516 DVSS.n2508 9.01392
R30755 DVSS.n2850 DVSS.n2849 9.01392
R30756 DVSS.n2837 DVSS.n2836 9.01392
R30757 DVSS.n2548 DVSS.n2547 9.01392
R30758 DVSS.n2830 DVSS.n2829 9.01392
R30759 DVSS.n2553 DVSS.n2552 9.01392
R30760 DVSS.n5537 DVSS.n5083 9.01392
R30761 DVSS.n5091 DVSS.n5082 9.01392
R30762 DVSS.n5528 DVSS.n5527 9.01392
R30763 DVSS.n5089 DVSS.n5088 9.01392
R30764 DVSS.n5497 DVSS.n5496 9.01392
R30765 DVSS.n5099 DVSS.n5097 9.01392
R30766 DVSS.n5109 DVSS.n5108 9.01392
R30767 DVSS.n5457 DVSS.n5456 9.01392
R30768 DVSS.n5115 DVSS.n5107 9.01392
R30769 DVSS.n5449 DVSS.n5448 9.01392
R30770 DVSS.n5436 DVSS.n5435 9.01392
R30771 DVSS.n5147 DVSS.n5146 9.01392
R30772 DVSS.n5429 DVSS.n5428 9.01392
R30773 DVSS.n5152 DVSS.n5151 9.01392
R30774 DVSS.n6001 DVSS.n5548 9.01392
R30775 DVSS.n5556 DVSS.n5547 9.01392
R30776 DVSS.n5993 DVSS.n5992 9.01392
R30777 DVSS.n5554 DVSS.n5553 9.01392
R30778 DVSS.n5962 DVSS.n5961 9.01392
R30779 DVSS.n5564 DVSS.n5562 9.01392
R30780 DVSS.n5574 DVSS.n5573 9.01392
R30781 DVSS.n5922 DVSS.n5921 9.01392
R30782 DVSS.n5580 DVSS.n5572 9.01392
R30783 DVSS.n5914 DVSS.n5913 9.01392
R30784 DVSS.n5901 DVSS.n5900 9.01392
R30785 DVSS.n5612 DVSS.n5611 9.01392
R30786 DVSS.n5894 DVSS.n5893 9.01392
R30787 DVSS.n5617 DVSS.n5616 9.01392
R30788 DVSS.n472 DVSS.n18 9.01392
R30789 DVSS.n26 DVSS.n17 9.01392
R30790 DVSS.n463 DVSS.n462 9.01392
R30791 DVSS.n24 DVSS.n23 9.01392
R30792 DVSS.n432 DVSS.n431 9.01392
R30793 DVSS.n34 DVSS.n32 9.01392
R30794 DVSS.n44 DVSS.n43 9.01392
R30795 DVSS.n392 DVSS.n391 9.01392
R30796 DVSS.n50 DVSS.n42 9.01392
R30797 DVSS.n384 DVSS.n383 9.01392
R30798 DVSS.n371 DVSS.n370 9.01392
R30799 DVSS.n82 DVSS.n81 9.01392
R30800 DVSS.n364 DVSS.n363 9.01392
R30801 DVSS.n87 DVSS.n86 9.01392
R30802 DVSS.n936 DVSS.n483 9.01392
R30803 DVSS.n491 DVSS.n482 9.01392
R30804 DVSS.n928 DVSS.n927 9.01392
R30805 DVSS.n489 DVSS.n488 9.01392
R30806 DVSS.n897 DVSS.n896 9.01392
R30807 DVSS.n499 DVSS.n497 9.01392
R30808 DVSS.n509 DVSS.n508 9.01392
R30809 DVSS.n857 DVSS.n856 9.01392
R30810 DVSS.n515 DVSS.n507 9.01392
R30811 DVSS.n849 DVSS.n848 9.01392
R30812 DVSS.n836 DVSS.n835 9.01392
R30813 DVSS.n547 DVSS.n546 9.01392
R30814 DVSS.n829 DVSS.n828 9.01392
R30815 DVSS.n552 DVSS.n551 9.01392
R30816 DVSS.n3952 DVSS.n3684 9.01392
R30817 DVSS.n3960 DVSS.n3959 9.01392
R30818 DVSS.n3955 DVSS.n3678 9.01392
R30819 DVSS.n3969 DVSS.n3968 9.01392
R30820 DVSS.n3980 DVSS.n3979 9.01392
R30821 DVSS.n3974 DVSS.n3639 9.01392
R30822 DVSS.n3990 DVSS.n3989 9.01392
R30823 DVSS.n3640 DVSS.n3636 9.01392
R30824 DVSS.n3997 DVSS.n3631 9.01392
R30825 DVSS.n4028 DVSS.n4027 9.01392
R30826 DVSS.n4023 DVSS.n3620 9.01392
R30827 DVSS.n4061 DVSS.n4060 9.01392
R30828 DVSS.n4063 DVSS.n3614 9.01392
R30829 DVSS.n4069 DVSS.n4068 9.01392
R30830 DVSS.n4417 DVSS.n4149 9.01392
R30831 DVSS.n4425 DVSS.n4424 9.01392
R30832 DVSS.n4420 DVSS.n4143 9.01392
R30833 DVSS.n4434 DVSS.n4433 9.01392
R30834 DVSS.n4445 DVSS.n4444 9.01392
R30835 DVSS.n4439 DVSS.n4104 9.01392
R30836 DVSS.n4455 DVSS.n4454 9.01392
R30837 DVSS.n4105 DVSS.n4101 9.01392
R30838 DVSS.n4462 DVSS.n4096 9.01392
R30839 DVSS.n4493 DVSS.n4492 9.01392
R30840 DVSS.n4488 DVSS.n4085 9.01392
R30841 DVSS.n4526 DVSS.n4525 9.01392
R30842 DVSS.n4528 DVSS.n4079 9.01392
R30843 DVSS.n4533 DVSS.n4532 9.01392
R30844 DVSS.n2356 DVSS.n2088 9.01392
R30845 DVSS.n2364 DVSS.n2363 9.01392
R30846 DVSS.n2359 DVSS.n2082 9.01392
R30847 DVSS.n2373 DVSS.n2372 9.01392
R30848 DVSS.n2384 DVSS.n2383 9.01392
R30849 DVSS.n2378 DVSS.n2043 9.01392
R30850 DVSS.n2394 DVSS.n2393 9.01392
R30851 DVSS.n2044 DVSS.n2040 9.01392
R30852 DVSS.n2401 DVSS.n2035 9.01392
R30853 DVSS.n2432 DVSS.n2431 9.01392
R30854 DVSS.n2427 DVSS.n2024 9.01392
R30855 DVSS.n2465 DVSS.n2464 9.01392
R30856 DVSS.n2467 DVSS.n2018 9.01392
R30857 DVSS.n2473 DVSS.n2472 9.01392
R30858 DVSS.n2821 DVSS.n2553 9.01392
R30859 DVSS.n2829 DVSS.n2828 9.01392
R30860 DVSS.n2824 DVSS.n2547 9.01392
R30861 DVSS.n2838 DVSS.n2837 9.01392
R30862 DVSS.n2849 DVSS.n2848 9.01392
R30863 DVSS.n2843 DVSS.n2508 9.01392
R30864 DVSS.n2859 DVSS.n2858 9.01392
R30865 DVSS.n2509 DVSS.n2505 9.01392
R30866 DVSS.n2866 DVSS.n2500 9.01392
R30867 DVSS.n2897 DVSS.n2896 9.01392
R30868 DVSS.n2892 DVSS.n2489 9.01392
R30869 DVSS.n2930 DVSS.n2929 9.01392
R30870 DVSS.n2932 DVSS.n2483 9.01392
R30871 DVSS.n2937 DVSS.n2936 9.01392
R30872 DVSS.n5420 DVSS.n5152 9.01392
R30873 DVSS.n5428 DVSS.n5427 9.01392
R30874 DVSS.n5423 DVSS.n5146 9.01392
R30875 DVSS.n5437 DVSS.n5436 9.01392
R30876 DVSS.n5448 DVSS.n5447 9.01392
R30877 DVSS.n5442 DVSS.n5107 9.01392
R30878 DVSS.n5458 DVSS.n5457 9.01392
R30879 DVSS.n5108 DVSS.n5104 9.01392
R30880 DVSS.n5465 DVSS.n5099 9.01392
R30881 DVSS.n5496 DVSS.n5495 9.01392
R30882 DVSS.n5491 DVSS.n5088 9.01392
R30883 DVSS.n5529 DVSS.n5528 9.01392
R30884 DVSS.n5531 DVSS.n5082 9.01392
R30885 DVSS.n5537 DVSS.n5536 9.01392
R30886 DVSS.n5885 DVSS.n5617 9.01392
R30887 DVSS.n5893 DVSS.n5892 9.01392
R30888 DVSS.n5888 DVSS.n5611 9.01392
R30889 DVSS.n5902 DVSS.n5901 9.01392
R30890 DVSS.n5913 DVSS.n5912 9.01392
R30891 DVSS.n5907 DVSS.n5572 9.01392
R30892 DVSS.n5923 DVSS.n5922 9.01392
R30893 DVSS.n5573 DVSS.n5569 9.01392
R30894 DVSS.n5930 DVSS.n5564 9.01392
R30895 DVSS.n5961 DVSS.n5960 9.01392
R30896 DVSS.n5956 DVSS.n5553 9.01392
R30897 DVSS.n5994 DVSS.n5993 9.01392
R30898 DVSS.n5996 DVSS.n5547 9.01392
R30899 DVSS.n6001 DVSS.n6000 9.01392
R30900 DVSS.n355 DVSS.n87 9.01392
R30901 DVSS.n363 DVSS.n362 9.01392
R30902 DVSS.n358 DVSS.n81 9.01392
R30903 DVSS.n372 DVSS.n371 9.01392
R30904 DVSS.n383 DVSS.n382 9.01392
R30905 DVSS.n377 DVSS.n42 9.01392
R30906 DVSS.n393 DVSS.n392 9.01392
R30907 DVSS.n43 DVSS.n39 9.01392
R30908 DVSS.n400 DVSS.n34 9.01392
R30909 DVSS.n431 DVSS.n430 9.01392
R30910 DVSS.n426 DVSS.n23 9.01392
R30911 DVSS.n464 DVSS.n463 9.01392
R30912 DVSS.n466 DVSS.n17 9.01392
R30913 DVSS.n472 DVSS.n471 9.01392
R30914 DVSS.n820 DVSS.n552 9.01392
R30915 DVSS.n828 DVSS.n827 9.01392
R30916 DVSS.n823 DVSS.n546 9.01392
R30917 DVSS.n837 DVSS.n836 9.01392
R30918 DVSS.n848 DVSS.n847 9.01392
R30919 DVSS.n842 DVSS.n507 9.01392
R30920 DVSS.n858 DVSS.n857 9.01392
R30921 DVSS.n508 DVSS.n504 9.01392
R30922 DVSS.n865 DVSS.n499 9.01392
R30923 DVSS.n896 DVSS.n895 9.01392
R30924 DVSS.n891 DVSS.n488 9.01392
R30925 DVSS.n929 DVSS.n928 9.01392
R30926 DVSS.n931 DVSS.n482 9.01392
R30927 DVSS.n936 DVSS.n935 9.01392
R30928 DVSS.n1916 DVSS.t175 9.00582
R30929 DVSS.n6842 DVSS.t35 9.00582
R30930 DVSS.n1060 DVSS.n1057 8.99329
R30931 DVSS.n1107 DVSS.n1106 8.99094
R30932 DVSS.n1101 DVSS.n1100 8.99094
R30933 DVSS.n1095 DVSS.n1094 8.99094
R30934 DVSS.n1095 DVSS.n1092 8.99094
R30935 DVSS.n1101 DVSS.n1097 8.99094
R30936 DVSS.n1107 DVSS.n1103 8.99094
R30937 DVSS.n3910 DVSS.n3902 8.9737
R30938 DVSS.n4375 DVSS.n4367 8.9737
R30939 DVSS.n2314 DVSS.n2306 8.9737
R30940 DVSS.n2779 DVSS.n2771 8.9737
R30941 DVSS.n5378 DVSS.n5370 8.9737
R30942 DVSS.n5843 DVSS.n5835 8.9737
R30943 DVSS.n313 DVSS.n305 8.9737
R30944 DVSS.n778 DVSS.n770 8.9737
R30945 DVSS.n3950 DVSS.n3713 8.8706
R30946 DVSS.n4415 DVSS.n4178 8.8706
R30947 DVSS.n2354 DVSS.n2117 8.8706
R30948 DVSS.n2819 DVSS.n2582 8.8706
R30949 DVSS.n5418 DVSS.n5181 8.8706
R30950 DVSS.n5883 DVSS.n5646 8.8706
R30951 DVSS.n353 DVSS.n116 8.8706
R30952 DVSS.n818 DVSS.n581 8.8706
R30953 DVSS.n1123 DVSS.n1049 8.85585
R30954 DVSS.n1226 DVSS.n1225 8.85585
R30955 DVSS.n1090 DVSS.n1086 8.85488
R30956 DVSS.n1083 DVSS.n1076 8.85488
R30957 DVSS.n1073 DVSS.n1069 8.85488
R30958 DVSS.n1046 DVSS.n1042 8.85488
R30959 DVSS.n1037 DVSS.n1033 8.85488
R30960 DVSS.n1030 DVSS.n1025 8.85488
R30961 DVSS.n1018 DVSS.n1014 8.85488
R30962 DVSS.n1011 DVSS.n1003 8.85488
R30963 DVSS.n1000 DVSS.n996 8.85488
R30964 DVSS.n993 DVSS.n989 8.85488
R30965 DVSS.n986 DVSS.n982 8.85488
R30966 DVSS.n979 DVSS.n975 8.85488
R30967 DVSS.n1290 DVSS.n1289 8.85488
R30968 DVSS.n1302 DVSS.n1301 8.85488
R30969 DVSS.n1310 DVSS.n1309 8.85488
R30970 DVSS.n1323 DVSS.n1322 8.85488
R30971 DVSS.n1155 DVSS.n1151 8.85488
R30972 DVSS.n1147 DVSS.n1138 8.85488
R30973 DVSS.n6736 DVSS.n6735 8.85488
R30974 DVSS.n1046 DVSS.n1045 8.85488
R30975 DVSS.n1030 DVSS.n1029 8.85488
R30976 DVSS.n1018 DVSS.n1017 8.85488
R30977 DVSS.n1037 DVSS.n1036 8.85488
R30978 DVSS.n1125 DVSS.n968 8.85488
R30979 DVSS.n979 DVSS.n978 8.85488
R30980 DVSS.n986 DVSS.n985 8.85488
R30981 DVSS.n993 DVSS.n992 8.85488
R30982 DVSS.n1000 DVSS.n999 8.85488
R30983 DVSS.n1011 DVSS.n1010 8.85488
R30984 DVSS.n1090 DVSS.n1089 8.85488
R30985 DVSS.n1118 DVSS.n1052 8.85488
R30986 DVSS.n1073 DVSS.n1072 8.85488
R30987 DVSS.n1083 DVSS.n1082 8.85488
R30988 DVSS.n1213 DVSS.n1209 8.85488
R30989 DVSS.n1206 DVSS.n1202 8.85488
R30990 DVSS.n1197 DVSS.n1192 8.85488
R30991 DVSS.n1189 DVSS.n1185 8.85488
R30992 DVSS.n1179 DVSS.n1175 8.85488
R30993 DVSS.n1213 DVSS.n1212 8.85488
R30994 DVSS.n1206 DVSS.n1205 8.85488
R30995 DVSS.n1197 DVSS.n1196 8.85488
R30996 DVSS.n1189 DVSS.n1188 8.85488
R30997 DVSS.n1179 DVSS.n1178 8.85488
R30998 DVSS.n1155 DVSS.n1154 8.85488
R30999 DVSS.n1147 DVSS.n1146 8.85488
R31000 DVSS.n1135 DVSS.n1134 8.85488
R31001 DVSS.n6701 DVSS.n6700 8.85487
R31002 DVSS.n1226 DVSS.n1216 8.85487
R31003 DVSS.n1335 DVSS.n1334 8.85487
R31004 DVSS.n1060 DVSS.n1059 8.85257
R31005 DVSS.n3887 DVSS.n3886 8.15208
R31006 DVSS.n4352 DVSS.n4351 8.15208
R31007 DVSS.n2291 DVSS.n2290 8.15208
R31008 DVSS.n2756 DVSS.n2755 8.15208
R31009 DVSS.n5355 DVSS.n5354 8.15208
R31010 DVSS.n5820 DVSS.n5819 8.15208
R31011 DVSS.n290 DVSS.n289 8.15208
R31012 DVSS.n755 DVSS.n754 8.15208
R31013 DVSS.n3699 DVSS.n3698 7.5692
R31014 DVSS.n3708 DVSS.n3699 7.5692
R31015 DVSS.n3708 DVSS.n3707 7.5692
R31016 DVSS.n3707 DVSS.n3705 7.5692
R31017 DVSS.n3705 DVSS.n3703 7.5692
R31018 DVSS.n3703 DVSS.n3701 7.5692
R31019 DVSS.n3701 DVSS.n3688 7.5692
R31020 DVSS.n3713 DVSS.n3688 7.5692
R31021 DVSS.n4039 DVSS.n4034 7.5692
R31022 DVSS.n4048 DVSS.n4039 7.5692
R31023 DVSS.n4048 DVSS.n4047 7.5692
R31024 DVSS.n4047 DVSS.n4046 7.5692
R31025 DVSS.n4046 DVSS.n4043 7.5692
R31026 DVSS.n4043 DVSS.n4042 7.5692
R31027 DVSS.n4042 DVSS.n3612 7.5692
R31028 DVSS.n4071 DVSS.n3612 7.5692
R31029 DVSS.n4164 DVSS.n4163 7.5692
R31030 DVSS.n4173 DVSS.n4164 7.5692
R31031 DVSS.n4173 DVSS.n4172 7.5692
R31032 DVSS.n4172 DVSS.n4170 7.5692
R31033 DVSS.n4170 DVSS.n4168 7.5692
R31034 DVSS.n4168 DVSS.n4166 7.5692
R31035 DVSS.n4166 DVSS.n4153 7.5692
R31036 DVSS.n4178 DVSS.n4153 7.5692
R31037 DVSS.n4504 DVSS.n4499 7.5692
R31038 DVSS.n4513 DVSS.n4504 7.5692
R31039 DVSS.n4513 DVSS.n4512 7.5692
R31040 DVSS.n4512 DVSS.n4511 7.5692
R31041 DVSS.n4511 DVSS.n4508 7.5692
R31042 DVSS.n4508 DVSS.n4507 7.5692
R31043 DVSS.n4507 DVSS.n4077 7.5692
R31044 DVSS.n4535 DVSS.n4077 7.5692
R31045 DVSS.n2103 DVSS.n2102 7.5692
R31046 DVSS.n2112 DVSS.n2103 7.5692
R31047 DVSS.n2112 DVSS.n2111 7.5692
R31048 DVSS.n2111 DVSS.n2109 7.5692
R31049 DVSS.n2109 DVSS.n2107 7.5692
R31050 DVSS.n2107 DVSS.n2105 7.5692
R31051 DVSS.n2105 DVSS.n2092 7.5692
R31052 DVSS.n2117 DVSS.n2092 7.5692
R31053 DVSS.n2443 DVSS.n2438 7.5692
R31054 DVSS.n2452 DVSS.n2443 7.5692
R31055 DVSS.n2452 DVSS.n2451 7.5692
R31056 DVSS.n2451 DVSS.n2450 7.5692
R31057 DVSS.n2450 DVSS.n2447 7.5692
R31058 DVSS.n2447 DVSS.n2446 7.5692
R31059 DVSS.n2446 DVSS.n2016 7.5692
R31060 DVSS.n2475 DVSS.n2016 7.5692
R31061 DVSS.n2568 DVSS.n2567 7.5692
R31062 DVSS.n2577 DVSS.n2568 7.5692
R31063 DVSS.n2577 DVSS.n2576 7.5692
R31064 DVSS.n2576 DVSS.n2574 7.5692
R31065 DVSS.n2574 DVSS.n2572 7.5692
R31066 DVSS.n2572 DVSS.n2570 7.5692
R31067 DVSS.n2570 DVSS.n2557 7.5692
R31068 DVSS.n2582 DVSS.n2557 7.5692
R31069 DVSS.n2908 DVSS.n2903 7.5692
R31070 DVSS.n2917 DVSS.n2908 7.5692
R31071 DVSS.n2917 DVSS.n2916 7.5692
R31072 DVSS.n2916 DVSS.n2915 7.5692
R31073 DVSS.n2915 DVSS.n2912 7.5692
R31074 DVSS.n2912 DVSS.n2911 7.5692
R31075 DVSS.n2911 DVSS.n2481 7.5692
R31076 DVSS.n2939 DVSS.n2481 7.5692
R31077 DVSS.n5167 DVSS.n5166 7.5692
R31078 DVSS.n5176 DVSS.n5167 7.5692
R31079 DVSS.n5176 DVSS.n5175 7.5692
R31080 DVSS.n5175 DVSS.n5173 7.5692
R31081 DVSS.n5173 DVSS.n5171 7.5692
R31082 DVSS.n5171 DVSS.n5169 7.5692
R31083 DVSS.n5169 DVSS.n5156 7.5692
R31084 DVSS.n5181 DVSS.n5156 7.5692
R31085 DVSS.n5507 DVSS.n5502 7.5692
R31086 DVSS.n5516 DVSS.n5507 7.5692
R31087 DVSS.n5516 DVSS.n5515 7.5692
R31088 DVSS.n5515 DVSS.n5514 7.5692
R31089 DVSS.n5514 DVSS.n5511 7.5692
R31090 DVSS.n5511 DVSS.n5510 7.5692
R31091 DVSS.n5510 DVSS.n5080 7.5692
R31092 DVSS.n5539 DVSS.n5080 7.5692
R31093 DVSS.n5632 DVSS.n5631 7.5692
R31094 DVSS.n5641 DVSS.n5632 7.5692
R31095 DVSS.n5641 DVSS.n5640 7.5692
R31096 DVSS.n5640 DVSS.n5638 7.5692
R31097 DVSS.n5638 DVSS.n5636 7.5692
R31098 DVSS.n5636 DVSS.n5634 7.5692
R31099 DVSS.n5634 DVSS.n5621 7.5692
R31100 DVSS.n5646 DVSS.n5621 7.5692
R31101 DVSS.n5972 DVSS.n5967 7.5692
R31102 DVSS.n5981 DVSS.n5972 7.5692
R31103 DVSS.n5981 DVSS.n5980 7.5692
R31104 DVSS.n5980 DVSS.n5979 7.5692
R31105 DVSS.n5979 DVSS.n5976 7.5692
R31106 DVSS.n5976 DVSS.n5975 7.5692
R31107 DVSS.n5975 DVSS.n5545 7.5692
R31108 DVSS.n6003 DVSS.n5545 7.5692
R31109 DVSS.n102 DVSS.n101 7.5692
R31110 DVSS.n111 DVSS.n102 7.5692
R31111 DVSS.n111 DVSS.n110 7.5692
R31112 DVSS.n110 DVSS.n108 7.5692
R31113 DVSS.n108 DVSS.n106 7.5692
R31114 DVSS.n106 DVSS.n104 7.5692
R31115 DVSS.n104 DVSS.n91 7.5692
R31116 DVSS.n116 DVSS.n91 7.5692
R31117 DVSS.n442 DVSS.n437 7.5692
R31118 DVSS.n451 DVSS.n442 7.5692
R31119 DVSS.n451 DVSS.n450 7.5692
R31120 DVSS.n450 DVSS.n449 7.5692
R31121 DVSS.n449 DVSS.n446 7.5692
R31122 DVSS.n446 DVSS.n445 7.5692
R31123 DVSS.n445 DVSS.n15 7.5692
R31124 DVSS.n474 DVSS.n15 7.5692
R31125 DVSS.n567 DVSS.n566 7.5692
R31126 DVSS.n576 DVSS.n567 7.5692
R31127 DVSS.n576 DVSS.n575 7.5692
R31128 DVSS.n575 DVSS.n573 7.5692
R31129 DVSS.n573 DVSS.n571 7.5692
R31130 DVSS.n571 DVSS.n569 7.5692
R31131 DVSS.n569 DVSS.n556 7.5692
R31132 DVSS.n581 DVSS.n556 7.5692
R31133 DVSS.n907 DVSS.n902 7.5692
R31134 DVSS.n916 DVSS.n907 7.5692
R31135 DVSS.n916 DVSS.n915 7.5692
R31136 DVSS.n915 DVSS.n914 7.5692
R31137 DVSS.n914 DVSS.n911 7.5692
R31138 DVSS.n911 DVSS.n910 7.5692
R31139 DVSS.n910 DVSS.n480 7.5692
R31140 DVSS.n938 DVSS.n480 7.5692
R31141 DVSS.n4072 DVSS.n4071 7.1358
R31142 DVSS.n4536 DVSS.n4535 7.1358
R31143 DVSS.n2476 DVSS.n2475 7.1358
R31144 DVSS.n2940 DVSS.n2939 7.1358
R31145 DVSS.n5540 DVSS.n5539 7.1358
R31146 DVSS.n6004 DVSS.n6003 7.1358
R31147 DVSS.n475 DVSS.n474 7.1358
R31148 DVSS.n939 DVSS.n938 7.1358
R31149 DVSS.n4072 DVSS.n3611 6.65838
R31150 DVSS.n4536 DVSS.n4076 6.65838
R31151 DVSS.n2476 DVSS.n2015 6.65838
R31152 DVSS.n2940 DVSS.n2480 6.65838
R31153 DVSS.n5540 DVSS.n5079 6.65838
R31154 DVSS.n6004 DVSS.n5544 6.65838
R31155 DVSS.n475 DVSS.n14 6.65838
R31156 DVSS.n939 DVSS.n479 6.65838
R31157 DVSS.n1385 DVSS.n1384 6.58671
R31158 DVSS.n1412 DVSS.n1411 6.58671
R31159 DVSS.n1635 DVSS.n1634 6.58671
R31160 DVSS.n1662 DVSS.n1661 6.58671
R31161 DVSS.n4598 DVSS.n4597 6.58671
R31162 DVSS.n4625 DVSS.n4624 6.58671
R31163 DVSS.n4848 DVSS.n4847 6.58671
R31164 DVSS.n4875 DVSS.n4874 6.58671
R31165 DVSS.n6066 DVSS.n6065 6.58671
R31166 DVSS.n6093 DVSS.n6092 6.58671
R31167 DVSS.n6316 DVSS.n6315 6.58671
R31168 DVSS.n6343 DVSS.n6342 6.58671
R31169 DVSS.n3002 DVSS.n3001 6.58671
R31170 DVSS.n3029 DVSS.n3028 6.58671
R31171 DVSS.n3252 DVSS.n3251 6.58671
R31172 DVSS.n3279 DVSS.n3278 6.58671
R31173 DVSS.n3914 DVSS.n3913 6.46787
R31174 DVSS.n4379 DVSS.n4378 6.46787
R31175 DVSS.n2318 DVSS.n2317 6.46787
R31176 DVSS.n2783 DVSS.n2782 6.46787
R31177 DVSS.n5382 DVSS.n5381 6.46787
R31178 DVSS.n5847 DVSS.n5846 6.46787
R31179 DVSS.n317 DVSS.n316 6.46787
R31180 DVSS.n782 DVSS.n781 6.46787
R31181 DVSS.n1517 DVSS.n1516 6.02403
R31182 DVSS.n1528 DVSS.n1527 6.02403
R31183 DVSS.n4730 DVSS.n4729 6.02403
R31184 DVSS.n4741 DVSS.n4740 6.02403
R31185 DVSS.n6198 DVSS.n6197 6.02403
R31186 DVSS.n6209 DVSS.n6208 6.02403
R31187 DVSS.n3134 DVSS.n3133 6.02403
R31188 DVSS.n3145 DVSS.n3144 6.02403
R31189 DVSS.n3866 DVSS.n3865 5.72682
R31190 DVSS.n3865 DVSS.n3864 5.72682
R31191 DVSS.n3864 DVSS.n3861 5.72682
R31192 DVSS.n3861 DVSS.n3860 5.72682
R31193 DVSS.n3860 DVSS.n3857 5.72682
R31194 DVSS.n3857 DVSS.n3856 5.72682
R31195 DVSS.n3856 DVSS.n3849 5.72682
R31196 DVSS.n3872 DVSS.n3849 5.72682
R31197 DVSS.n4331 DVSS.n4330 5.72682
R31198 DVSS.n4330 DVSS.n4329 5.72682
R31199 DVSS.n4329 DVSS.n4326 5.72682
R31200 DVSS.n4326 DVSS.n4325 5.72682
R31201 DVSS.n4325 DVSS.n4322 5.72682
R31202 DVSS.n4322 DVSS.n4321 5.72682
R31203 DVSS.n4321 DVSS.n4314 5.72682
R31204 DVSS.n4337 DVSS.n4314 5.72682
R31205 DVSS.n2270 DVSS.n2269 5.72682
R31206 DVSS.n2269 DVSS.n2268 5.72682
R31207 DVSS.n2268 DVSS.n2265 5.72682
R31208 DVSS.n2265 DVSS.n2264 5.72682
R31209 DVSS.n2264 DVSS.n2261 5.72682
R31210 DVSS.n2261 DVSS.n2260 5.72682
R31211 DVSS.n2260 DVSS.n2253 5.72682
R31212 DVSS.n2276 DVSS.n2253 5.72682
R31213 DVSS.n2735 DVSS.n2734 5.72682
R31214 DVSS.n2734 DVSS.n2733 5.72682
R31215 DVSS.n2733 DVSS.n2730 5.72682
R31216 DVSS.n2730 DVSS.n2729 5.72682
R31217 DVSS.n2729 DVSS.n2726 5.72682
R31218 DVSS.n2726 DVSS.n2725 5.72682
R31219 DVSS.n2725 DVSS.n2718 5.72682
R31220 DVSS.n2741 DVSS.n2718 5.72682
R31221 DVSS.n5334 DVSS.n5333 5.72682
R31222 DVSS.n5333 DVSS.n5332 5.72682
R31223 DVSS.n5332 DVSS.n5329 5.72682
R31224 DVSS.n5329 DVSS.n5328 5.72682
R31225 DVSS.n5328 DVSS.n5325 5.72682
R31226 DVSS.n5325 DVSS.n5324 5.72682
R31227 DVSS.n5324 DVSS.n5317 5.72682
R31228 DVSS.n5340 DVSS.n5317 5.72682
R31229 DVSS.n5799 DVSS.n5798 5.72682
R31230 DVSS.n5798 DVSS.n5797 5.72682
R31231 DVSS.n5797 DVSS.n5794 5.72682
R31232 DVSS.n5794 DVSS.n5793 5.72682
R31233 DVSS.n5793 DVSS.n5790 5.72682
R31234 DVSS.n5790 DVSS.n5789 5.72682
R31235 DVSS.n5789 DVSS.n5782 5.72682
R31236 DVSS.n5805 DVSS.n5782 5.72682
R31237 DVSS.n269 DVSS.n268 5.72682
R31238 DVSS.n268 DVSS.n267 5.72682
R31239 DVSS.n267 DVSS.n264 5.72682
R31240 DVSS.n264 DVSS.n263 5.72682
R31241 DVSS.n263 DVSS.n260 5.72682
R31242 DVSS.n260 DVSS.n259 5.72682
R31243 DVSS.n259 DVSS.n252 5.72682
R31244 DVSS.n275 DVSS.n252 5.72682
R31245 DVSS.n734 DVSS.n733 5.72682
R31246 DVSS.n733 DVSS.n732 5.72682
R31247 DVSS.n732 DVSS.n729 5.72682
R31248 DVSS.n729 DVSS.n728 5.72682
R31249 DVSS.n728 DVSS.n725 5.72682
R31250 DVSS.n725 DVSS.n724 5.72682
R31251 DVSS.n724 DVSS.n717 5.72682
R31252 DVSS.n740 DVSS.n717 5.72682
R31253 DVSS.n1394 DVSS.n1383 5.64756
R31254 DVSS.n1420 DVSS.n1409 5.64756
R31255 DVSS.n1644 DVSS.n1633 5.64756
R31256 DVSS.n1670 DVSS.n1659 5.64756
R31257 DVSS.n6714 DVSS.n3485 5.64756
R31258 DVSS.n4607 DVSS.n4596 5.64756
R31259 DVSS.n4633 DVSS.n4622 5.64756
R31260 DVSS.n4857 DVSS.n4846 5.64756
R31261 DVSS.n4883 DVSS.n4872 5.64756
R31262 DVSS.n3751 DVSS.n3750 5.64756
R31263 DVSS.n3750 DVSS.n3740 5.64756
R31264 DVSS.n3730 DVSS.n3729 5.64756
R31265 DVSS.n3729 DVSS.n3719 5.64756
R31266 DVSS.n4216 DVSS.n4215 5.64756
R31267 DVSS.n4215 DVSS.n4205 5.64756
R31268 DVSS.n4195 DVSS.n4194 5.64756
R31269 DVSS.n4194 DVSS.n4184 5.64756
R31270 DVSS.n6075 DVSS.n6064 5.64756
R31271 DVSS.n6101 DVSS.n6090 5.64756
R31272 DVSS.n6325 DVSS.n6314 5.64756
R31273 DVSS.n6351 DVSS.n6340 5.64756
R31274 DVSS.n3011 DVSS.n3000 5.64756
R31275 DVSS.n3037 DVSS.n3026 5.64756
R31276 DVSS.n3261 DVSS.n3250 5.64756
R31277 DVSS.n3287 DVSS.n3276 5.64756
R31278 DVSS.n6756 DVSS.n6749 5.64756
R31279 DVSS.n2155 DVSS.n2154 5.64756
R31280 DVSS.n2154 DVSS.n2144 5.64756
R31281 DVSS.n2134 DVSS.n2133 5.64756
R31282 DVSS.n2133 DVSS.n2123 5.64756
R31283 DVSS.n2620 DVSS.n2619 5.64756
R31284 DVSS.n2619 DVSS.n2609 5.64756
R31285 DVSS.n2599 DVSS.n2598 5.64756
R31286 DVSS.n2598 DVSS.n2588 5.64756
R31287 DVSS.n5219 DVSS.n5218 5.64756
R31288 DVSS.n5218 DVSS.n5208 5.64756
R31289 DVSS.n5198 DVSS.n5197 5.64756
R31290 DVSS.n5197 DVSS.n5187 5.64756
R31291 DVSS.n5684 DVSS.n5683 5.64756
R31292 DVSS.n5683 DVSS.n5673 5.64756
R31293 DVSS.n5663 DVSS.n5662 5.64756
R31294 DVSS.n5662 DVSS.n5652 5.64756
R31295 DVSS.n154 DVSS.n153 5.64756
R31296 DVSS.n153 DVSS.n143 5.64756
R31297 DVSS.n133 DVSS.n132 5.64756
R31298 DVSS.n132 DVSS.n122 5.64756
R31299 DVSS.n619 DVSS.n618 5.64756
R31300 DVSS.n618 DVSS.n608 5.64756
R31301 DVSS.n598 DVSS.n597 5.64756
R31302 DVSS.n597 DVSS.n587 5.64756
R31303 DVSS.n3979 DVSS.n3649 5.57999
R31304 DVSS.n4027 DVSS.n3634 5.57999
R31305 DVSS.n4444 DVSS.n4114 5.57999
R31306 DVSS.n4492 DVSS.n4099 5.57999
R31307 DVSS.n2383 DVSS.n2053 5.57999
R31308 DVSS.n2431 DVSS.n2038 5.57999
R31309 DVSS.n2848 DVSS.n2518 5.57999
R31310 DVSS.n2896 DVSS.n2503 5.57999
R31311 DVSS.n5447 DVSS.n5117 5.57999
R31312 DVSS.n5495 DVSS.n5102 5.57999
R31313 DVSS.n5912 DVSS.n5582 5.57999
R31314 DVSS.n5960 DVSS.n5567 5.57999
R31315 DVSS.n382 DVSS.n52 5.57999
R31316 DVSS.n430 DVSS.n37 5.57999
R31317 DVSS.n847 DVSS.n517 5.57999
R31318 DVSS.n895 DVSS.n502 5.57999
R31319 DVSS.n3969 DVSS.n3677 5.34556
R31320 DVSS.n4434 DVSS.n4142 5.34556
R31321 DVSS.n2373 DVSS.n2081 5.34556
R31322 DVSS.n2838 DVSS.n2546 5.34556
R31323 DVSS.n5437 DVSS.n5145 5.34556
R31324 DVSS.n5902 DVSS.n5610 5.34556
R31325 DVSS.n372 DVSS.n80 5.34556
R31326 DVSS.n837 DVSS.n545 5.34556
R31327 DVSS.n4023 DVSS.n4022 5.29867
R31328 DVSS.n4488 DVSS.n4487 5.29867
R31329 DVSS.n2427 DVSS.n2426 5.29867
R31330 DVSS.n2892 DVSS.n2891 5.29867
R31331 DVSS.n5491 DVSS.n5490 5.29867
R31332 DVSS.n5956 DVSS.n5955 5.29867
R31333 DVSS.n426 DVSS.n425 5.29867
R31334 DVSS.n891 DVSS.n890 5.29867
R31335 DVSS.n1502 DVSS.n1501 5.27109
R31336 DVSS.n1543 DVSS.n1542 5.27109
R31337 DVSS.n4715 DVSS.n4714 5.27109
R31338 DVSS.n4756 DVSS.n4755 5.27109
R31339 DVSS.n6183 DVSS.n6182 5.27109
R31340 DVSS.n6224 DVSS.n6223 5.27109
R31341 DVSS.n3119 DVSS.n3118 5.27109
R31342 DVSS.n3160 DVSS.n3159 5.27109
R31343 DVSS.n6204 DVSS.n6203 5.11084
R31344 DVSS.n6215 DVSS.n6214 5.11084
R31345 DVSS.n4736 DVSS.n4735 5.11084
R31346 DVSS.n4747 DVSS.n4746 5.11084
R31347 DVSS.n3140 DVSS.n3139 5.11084
R31348 DVSS.n3151 DVSS.n3150 5.11084
R31349 DVSS.n1523 DVSS.n1522 5.11084
R31350 DVSS.n1534 DVSS.n1533 5.11084
R31351 DVSS.n1376 DVSS.n1368 4.89462
R31352 DVSS.n1435 DVSS.n1427 4.89462
R31353 DVSS.n1626 DVSS.n1618 4.89462
R31354 DVSS.n1685 DVSS.n1677 4.89462
R31355 DVSS.n4589 DVSS.n4581 4.89462
R31356 DVSS.n4648 DVSS.n4640 4.89462
R31357 DVSS.n4839 DVSS.n4831 4.89462
R31358 DVSS.n4898 DVSS.n4890 4.89462
R31359 DVSS.n3754 DVSS.n3737 4.89462
R31360 DVSS.n3733 DVSS.n3716 4.89462
R31361 DVSS.n4219 DVSS.n4202 4.89462
R31362 DVSS.n4198 DVSS.n4181 4.89462
R31363 DVSS.n6057 DVSS.n6049 4.89462
R31364 DVSS.n6116 DVSS.n6108 4.89462
R31365 DVSS.n6307 DVSS.n6299 4.89462
R31366 DVSS.n6366 DVSS.n6358 4.89462
R31367 DVSS.n2993 DVSS.n2985 4.89462
R31368 DVSS.n3052 DVSS.n3044 4.89462
R31369 DVSS.n3243 DVSS.n3235 4.89462
R31370 DVSS.n3302 DVSS.n3294 4.89462
R31371 DVSS.n2158 DVSS.n2141 4.89462
R31372 DVSS.n2137 DVSS.n2120 4.89462
R31373 DVSS.n2623 DVSS.n2606 4.89462
R31374 DVSS.n2602 DVSS.n2585 4.89462
R31375 DVSS.n5222 DVSS.n5205 4.89462
R31376 DVSS.n5201 DVSS.n5184 4.89462
R31377 DVSS.n5687 DVSS.n5670 4.89462
R31378 DVSS.n5666 DVSS.n5649 4.89462
R31379 DVSS.n157 DVSS.n140 4.89462
R31380 DVSS.n136 DVSS.n119 4.89462
R31381 DVSS.n622 DVSS.n605 4.89462
R31382 DVSS.n601 DVSS.n584 4.89462
R31383 DVSS.n3922 DVSS.n3776 4.74328
R31384 DVSS.n3817 DVSS.n3792 4.74328
R31385 DVSS.n4387 DVSS.n4241 4.74328
R31386 DVSS.n4282 DVSS.n4257 4.74328
R31387 DVSS.n2326 DVSS.n2180 4.74328
R31388 DVSS.n2221 DVSS.n2196 4.74328
R31389 DVSS.n2791 DVSS.n2645 4.74328
R31390 DVSS.n2686 DVSS.n2661 4.74328
R31391 DVSS.n5390 DVSS.n5244 4.74328
R31392 DVSS.n5285 DVSS.n5260 4.74328
R31393 DVSS.n5855 DVSS.n5709 4.74328
R31394 DVSS.n5750 DVSS.n5725 4.74328
R31395 DVSS.n325 DVSS.n179 4.74328
R31396 DVSS.n220 DVSS.n195 4.74328
R31397 DVSS.n790 DVSS.n644 4.74328
R31398 DVSS.n685 DVSS.n660 4.74328
R31399 DVSS.n1168 DVSS.n1167 4.72584
R31400 DVSS.n1117 DVSS.n1116 4.72584
R31401 DVSS.n4575 DVSS.n4564 4.71739
R31402 DVSS.n6043 DVSS.n6032 4.71739
R31403 DVSS.n2979 DVSS.n2968 4.71739
R31404 DVSS.n1362 DVSS.n1351 4.71739
R31405 DVSS.n3481 DVSS.n3480 4.65375
R31406 DVSS.n7 DVSS.n6 4.65375
R31407 DVSS.n1120 DVSS.n1119 4.6505
R31408 DVSS.n1065 DVSS.n1064 4.6505
R31409 DVSS.n1127 DVSS.n1126 4.6505
R31410 DVSS.n972 DVSS.n971 4.6505
R31411 DVSS.n1007 DVSS.n1006 4.6505
R31412 DVSS.n1022 DVSS.n1021 4.6505
R31413 DVSS.n1812 DVSS.n1811 4.6505
R31414 DVSS.n1795 DVSS.n1794 4.6505
R31415 DVSS.n1754 DVSS.n1753 4.6505
R31416 DVSS.n1751 DVSS.n1750 4.6505
R31417 DVSS.n1758 DVSS.n1757 4.6505
R31418 DVSS.n1762 DVSS.n1761 4.6505
R31419 DVSS.n1766 DVSS.n1765 4.6505
R31420 DVSS.n1770 DVSS.n1769 4.6505
R31421 DVSS.n1774 DVSS.n1773 4.6505
R31422 DVSS.n1778 DVSS.n1777 4.6505
R31423 DVSS.n6690 DVSS.n6689 4.6505
R31424 DVSS.n6687 DVSS.n6686 4.6505
R31425 DVSS.n6672 DVSS.n6671 4.6505
R31426 DVSS.n6685 DVSS.n6684 4.6505
R31427 DVSS.n6681 DVSS.n6680 4.6505
R31428 DVSS.n6676 DVSS.n6675 4.6505
R31429 DVSS.n6668 DVSS.n6667 4.6505
R31430 DVSS.n6663 DVSS.n6662 4.6505
R31431 DVSS.n6659 DVSS.n6658 4.6505
R31432 DVSS.n6721 DVSS.n6720 4.6505
R31433 DVSS.n5024 DVSS.n5023 4.6505
R31434 DVSS.n5007 DVSS.n5006 4.6505
R31435 DVSS.n4966 DVSS.n4965 4.6505
R31436 DVSS.n4963 DVSS.n4962 4.6505
R31437 DVSS.n4970 DVSS.n4969 4.6505
R31438 DVSS.n4974 DVSS.n4973 4.6505
R31439 DVSS.n4978 DVSS.n4977 4.6505
R31440 DVSS.n4982 DVSS.n4981 4.6505
R31441 DVSS.n4986 DVSS.n4985 4.6505
R31442 DVSS.n4990 DVSS.n4989 4.6505
R31443 DVSS.n3922 DVSS.n3921 4.6505
R31444 DVSS.n3942 DVSS.n3941 4.6505
R31445 DVSS.n3924 DVSS.n3923 4.6505
R31446 DVSS.n3927 DVSS.n3774 4.6505
R31447 DVSS.n3931 DVSS.n3930 4.6505
R31448 DVSS.n3933 DVSS.n3932 4.6505
R31449 DVSS.n3773 DVSS.n3770 4.6505
R31450 DVSS.n3758 DVSS.n3756 4.6505
R31451 DVSS.n3799 DVSS.n3735 4.6505
R31452 DVSS.n3830 DVSS.n3829 4.6505
R31453 DVSS.n3832 DVSS.n3831 4.6505
R31454 DVSS.n3816 DVSS.n3811 4.6505
R31455 DVSS.n3805 DVSS.n3801 4.6505
R31456 DVSS.n3840 DVSS.n3839 4.6505
R31457 DVSS.n3842 DVSS.n3841 4.6505
R31458 DVSS.n3818 DVSS.n3817 4.6505
R31459 DVSS.n4387 DVSS.n4386 4.6505
R31460 DVSS.n4407 DVSS.n4406 4.6505
R31461 DVSS.n4389 DVSS.n4388 4.6505
R31462 DVSS.n4392 DVSS.n4239 4.6505
R31463 DVSS.n4396 DVSS.n4395 4.6505
R31464 DVSS.n4398 DVSS.n4397 4.6505
R31465 DVSS.n4238 DVSS.n4235 4.6505
R31466 DVSS.n4223 DVSS.n4221 4.6505
R31467 DVSS.n4264 DVSS.n4200 4.6505
R31468 DVSS.n4295 DVSS.n4294 4.6505
R31469 DVSS.n4297 DVSS.n4296 4.6505
R31470 DVSS.n4281 DVSS.n4276 4.6505
R31471 DVSS.n4270 DVSS.n4266 4.6505
R31472 DVSS.n4305 DVSS.n4304 4.6505
R31473 DVSS.n4307 DVSS.n4306 4.6505
R31474 DVSS.n4283 DVSS.n4282 4.6505
R31475 DVSS.n4616 DVSS.n4615 4.6505
R31476 DVSS.n4866 DVSS.n4865 4.6505
R31477 DVSS.n4945 DVSS.n4944 4.6505
R31478 DVSS.n6084 DVSS.n6083 4.6505
R31479 DVSS.n6334 DVSS.n6333 4.6505
R31480 DVSS.n6413 DVSS.n6412 4.6505
R31481 DVSS.n3429 DVSS.n3428 4.6505
R31482 DVSS.n3412 DVSS.n3411 4.6505
R31483 DVSS.n3371 DVSS.n3370 4.6505
R31484 DVSS.n3368 DVSS.n3367 4.6505
R31485 DVSS.n3375 DVSS.n3374 4.6505
R31486 DVSS.n3379 DVSS.n3378 4.6505
R31487 DVSS.n3383 DVSS.n3382 4.6505
R31488 DVSS.n3387 DVSS.n3386 4.6505
R31489 DVSS.n3391 DVSS.n3390 4.6505
R31490 DVSS.n3395 DVSS.n3394 4.6505
R31491 DVSS.n6741 DVSS.n1857 4.6505
R31492 DVSS.n6738 DVSS.n6737 4.6505
R31493 DVSS.n1898 DVSS.n1858 4.6505
R31494 DVSS.n1899 DVSS.n1898 4.6505
R31495 DVSS.n1922 DVSS.n1921 4.6505
R31496 DVSS.n1939 DVSS.n1938 4.6505
R31497 DVSS.n1954 DVSS.n1953 4.6505
R31498 DVSS.n1981 DVSS.n1980 4.6505
R31499 DVSS.n1907 DVSS.n1906 4.6505
R31500 DVSS.n2326 DVSS.n2325 4.6505
R31501 DVSS.n2346 DVSS.n2345 4.6505
R31502 DVSS.n2328 DVSS.n2327 4.6505
R31503 DVSS.n2331 DVSS.n2178 4.6505
R31504 DVSS.n2335 DVSS.n2334 4.6505
R31505 DVSS.n2337 DVSS.n2336 4.6505
R31506 DVSS.n2177 DVSS.n2174 4.6505
R31507 DVSS.n2162 DVSS.n2160 4.6505
R31508 DVSS.n2203 DVSS.n2139 4.6505
R31509 DVSS.n2234 DVSS.n2233 4.6505
R31510 DVSS.n2236 DVSS.n2235 4.6505
R31511 DVSS.n2220 DVSS.n2215 4.6505
R31512 DVSS.n2209 DVSS.n2205 4.6505
R31513 DVSS.n2244 DVSS.n2243 4.6505
R31514 DVSS.n2246 DVSS.n2245 4.6505
R31515 DVSS.n2222 DVSS.n2221 4.6505
R31516 DVSS.n2791 DVSS.n2790 4.6505
R31517 DVSS.n2811 DVSS.n2810 4.6505
R31518 DVSS.n2793 DVSS.n2792 4.6505
R31519 DVSS.n2796 DVSS.n2643 4.6505
R31520 DVSS.n2800 DVSS.n2799 4.6505
R31521 DVSS.n2802 DVSS.n2801 4.6505
R31522 DVSS.n2642 DVSS.n2639 4.6505
R31523 DVSS.n2627 DVSS.n2625 4.6505
R31524 DVSS.n2668 DVSS.n2604 4.6505
R31525 DVSS.n2699 DVSS.n2698 4.6505
R31526 DVSS.n2701 DVSS.n2700 4.6505
R31527 DVSS.n2685 DVSS.n2680 4.6505
R31528 DVSS.n2674 DVSS.n2670 4.6505
R31529 DVSS.n2709 DVSS.n2708 4.6505
R31530 DVSS.n2711 DVSS.n2710 4.6505
R31531 DVSS.n2687 DVSS.n2686 4.6505
R31532 DVSS.n3020 DVSS.n3019 4.6505
R31533 DVSS.n3270 DVSS.n3269 4.6505
R31534 DVSS.n3350 DVSS.n3349 4.6505
R31535 DVSS.n3399 DVSS.n3398 4.6505
R31536 DVSS.n3404 DVSS.n3403 4.6505
R31537 DVSS.n3409 DVSS.n3408 4.6505
R31538 DVSS.n3416 DVSS.n3415 4.6505
R31539 DVSS.n3420 DVSS.n3419 4.6505
R31540 DVSS.n3425 DVSS.n3424 4.6505
R31541 DVSS.n3433 DVSS.n3432 4.6505
R31542 DVSS.n3437 DVSS.n3436 4.6505
R31543 DVSS.n3441 DVSS.n3440 4.6505
R31544 DVSS.n3447 DVSS.n3446 4.6505
R31545 DVSS.n3451 DVSS.n3450 4.6505
R31546 DVSS.n6732 DVSS.n6731 4.6505
R31547 DVSS.n1896 DVSS.n1895 4.6505
R31548 DVSS.n1901 DVSS.n1900 4.6505
R31549 DVSS.n1911 DVSS.n1910 4.6505
R31550 DVSS.n1915 DVSS.n1914 4.6505
R31551 DVSS.n1919 DVSS.n1918 4.6505
R31552 DVSS.n1926 DVSS.n1925 4.6505
R31553 DVSS.n1931 DVSS.n1930 4.6505
R31554 DVSS.n1935 DVSS.n1934 4.6505
R31555 DVSS.n1943 DVSS.n1942 4.6505
R31556 DVSS.n1948 DVSS.n1947 4.6505
R31557 DVSS.n1952 DVSS.n1951 4.6505
R31558 DVSS.n1959 DVSS.n1958 4.6505
R31559 DVSS.n1964 DVSS.n1963 4.6505
R31560 DVSS.n1968 DVSS.n1967 4.6505
R31561 DVSS.n1972 DVSS.n1971 4.6505
R31562 DVSS.n1977 DVSS.n1976 4.6505
R31563 DVSS.n1986 DVSS.n1985 4.6505
R31564 DVSS.n1990 DVSS.n1989 4.6505
R31565 DVSS.n1994 DVSS.n1991 4.6505
R31566 DVSS.n1998 DVSS.n1997 4.6505
R31567 DVSS.n2002 DVSS.n2001 4.6505
R31568 DVSS.n4994 DVSS.n4993 4.6505
R31569 DVSS.n4999 DVSS.n4998 4.6505
R31570 DVSS.n5004 DVSS.n5003 4.6505
R31571 DVSS.n5011 DVSS.n5010 4.6505
R31572 DVSS.n5015 DVSS.n5014 4.6505
R31573 DVSS.n5020 DVSS.n5019 4.6505
R31574 DVSS.n5028 DVSS.n5027 4.6505
R31575 DVSS.n5032 DVSS.n5031 4.6505
R31576 DVSS.n5036 DVSS.n5035 4.6505
R31577 DVSS.n5042 DVSS.n5041 4.6505
R31578 DVSS.n5046 DVSS.n5045 4.6505
R31579 DVSS.n6492 DVSS.n6491 4.6505
R31580 DVSS.n6475 DVSS.n6474 4.6505
R31581 DVSS.n6434 DVSS.n6433 4.6505
R31582 DVSS.n6431 DVSS.n6430 4.6505
R31583 DVSS.n6438 DVSS.n6437 4.6505
R31584 DVSS.n6442 DVSS.n6441 4.6505
R31585 DVSS.n6446 DVSS.n6445 4.6505
R31586 DVSS.n6450 DVSS.n6449 4.6505
R31587 DVSS.n6454 DVSS.n6453 4.6505
R31588 DVSS.n6458 DVSS.n6457 4.6505
R31589 DVSS.n6462 DVSS.n6461 4.6505
R31590 DVSS.n6467 DVSS.n6466 4.6505
R31591 DVSS.n6472 DVSS.n6471 4.6505
R31592 DVSS.n6479 DVSS.n6478 4.6505
R31593 DVSS.n6483 DVSS.n6482 4.6505
R31594 DVSS.n6488 DVSS.n6487 4.6505
R31595 DVSS.n6496 DVSS.n6495 4.6505
R31596 DVSS.n6500 DVSS.n6499 4.6505
R31597 DVSS.n6505 DVSS.n6504 4.6505
R31598 DVSS.n6510 DVSS.n6509 4.6505
R31599 DVSS.n6513 DVSS.n6512 4.6505
R31600 DVSS.n5390 DVSS.n5389 4.6505
R31601 DVSS.n5410 DVSS.n5409 4.6505
R31602 DVSS.n5392 DVSS.n5391 4.6505
R31603 DVSS.n5395 DVSS.n5242 4.6505
R31604 DVSS.n5399 DVSS.n5398 4.6505
R31605 DVSS.n5401 DVSS.n5400 4.6505
R31606 DVSS.n5241 DVSS.n5238 4.6505
R31607 DVSS.n5226 DVSS.n5224 4.6505
R31608 DVSS.n5267 DVSS.n5203 4.6505
R31609 DVSS.n5298 DVSS.n5297 4.6505
R31610 DVSS.n5300 DVSS.n5299 4.6505
R31611 DVSS.n5284 DVSS.n5279 4.6505
R31612 DVSS.n5273 DVSS.n5269 4.6505
R31613 DVSS.n5308 DVSS.n5307 4.6505
R31614 DVSS.n5310 DVSS.n5309 4.6505
R31615 DVSS.n5286 DVSS.n5285 4.6505
R31616 DVSS.n5855 DVSS.n5854 4.6505
R31617 DVSS.n5875 DVSS.n5874 4.6505
R31618 DVSS.n5857 DVSS.n5856 4.6505
R31619 DVSS.n5860 DVSS.n5707 4.6505
R31620 DVSS.n5864 DVSS.n5863 4.6505
R31621 DVSS.n5866 DVSS.n5865 4.6505
R31622 DVSS.n5706 DVSS.n5703 4.6505
R31623 DVSS.n5691 DVSS.n5689 4.6505
R31624 DVSS.n5732 DVSS.n5668 4.6505
R31625 DVSS.n5763 DVSS.n5762 4.6505
R31626 DVSS.n5765 DVSS.n5764 4.6505
R31627 DVSS.n5749 DVSS.n5744 4.6505
R31628 DVSS.n5738 DVSS.n5734 4.6505
R31629 DVSS.n5773 DVSS.n5772 4.6505
R31630 DVSS.n5775 DVSS.n5774 4.6505
R31631 DVSS.n5751 DVSS.n5750 4.6505
R31632 DVSS.n6628 DVSS.n5073 4.6505
R31633 DVSS.n6614 DVSS.n6613 4.6505
R31634 DVSS.n6596 DVSS.n6595 4.6505
R31635 DVSS.n6572 DVSS.n6571 4.6505
R31636 DVSS.n6642 DVSS.n6641 4.6505
R31637 DVSS.n6640 DVSS.n6639 4.6505
R31638 DVSS.n6636 DVSS.n6635 4.6505
R31639 DVSS.n6632 DVSS.n6631 4.6505
R31640 DVSS.n6627 DVSS.n6626 4.6505
R31641 DVSS.n6622 DVSS.n6621 4.6505
R31642 DVSS.n6618 DVSS.n6617 4.6505
R31643 DVSS.n6610 DVSS.n6609 4.6505
R31644 DVSS.n6605 DVSS.n6604 4.6505
R31645 DVSS.n6601 DVSS.n6600 4.6505
R31646 DVSS.n6594 DVSS.n6593 4.6505
R31647 DVSS.n6589 DVSS.n6588 4.6505
R31648 DVSS.n6585 DVSS.n6584 4.6505
R31649 DVSS.n6581 DVSS.n6580 4.6505
R31650 DVSS.n6576 DVSS.n6575 4.6505
R31651 DVSS.n6567 DVSS.n6566 4.6505
R31652 DVSS.n6563 DVSS.n6562 4.6505
R31653 DVSS.n6559 DVSS.n6558 4.6505
R31654 DVSS.n6557 DVSS.n6554 4.6505
R31655 DVSS.n6553 DVSS.n6552 4.6505
R31656 DVSS.n6706 DVSS.n5069 4.6505
R31657 DVSS.n6703 DVSS.n6702 4.6505
R31658 DVSS.n6697 DVSS.n6696 4.6505
R31659 DVSS.n6654 DVSS.n6653 4.6505
R31660 DVSS.n6648 DVSS.n6647 4.6505
R31661 DVSS.n6655 DVSS.n5070 4.6505
R31662 DVSS.n5071 DVSS.n5070 4.6505
R31663 DVSS.n3584 DVSS.n3583 4.6505
R31664 DVSS.n3557 DVSS.n3556 4.6505
R31665 DVSS.n3542 DVSS.n3541 4.6505
R31666 DVSS.n3525 DVSS.n3524 4.6505
R31667 DVSS.n3514 DVSS.n3513 4.6505
R31668 DVSS.n3518 DVSS.n3517 4.6505
R31669 DVSS.n3522 DVSS.n3521 4.6505
R31670 DVSS.n3529 DVSS.n3528 4.6505
R31671 DVSS.n3534 DVSS.n3533 4.6505
R31672 DVSS.n3538 DVSS.n3537 4.6505
R31673 DVSS.n3546 DVSS.n3545 4.6505
R31674 DVSS.n3551 DVSS.n3550 4.6505
R31675 DVSS.n3555 DVSS.n3554 4.6505
R31676 DVSS.n3562 DVSS.n3561 4.6505
R31677 DVSS.n3567 DVSS.n3566 4.6505
R31678 DVSS.n3571 DVSS.n3570 4.6505
R31679 DVSS.n3575 DVSS.n3574 4.6505
R31680 DVSS.n3580 DVSS.n3579 4.6505
R31681 DVSS.n3589 DVSS.n3588 4.6505
R31682 DVSS.n3593 DVSS.n3592 4.6505
R31683 DVSS.n3600 DVSS.n3599 4.6505
R31684 DVSS.n3605 DVSS.n3604 4.6505
R31685 DVSS.n3509 DVSS.n3508 4.6505
R31686 DVSS.n3489 DVSS.n3488 4.6505
R31687 DVSS.n3493 DVSS.n3492 4.6505
R31688 DVSS.n3498 DVSS.n3497 4.6505
R31689 DVSS.n3503 DVSS.n3502 4.6505
R31690 DVSS.n3500 DVSS.n3499 4.6505
R31691 DVSS.n3501 DVSS.n3500 4.6505
R31692 DVSS.n6725 DVSS.n6724 4.6505
R31693 DVSS.n1889 DVSS.n1888 4.6505
R31694 DVSS.n1885 DVSS.n1884 4.6505
R31695 DVSS.n1880 DVSS.n1879 4.6505
R31696 DVSS.n1872 DVSS.n1871 4.6505
R31697 DVSS.n1867 DVSS.n1866 4.6505
R31698 DVSS.n1863 DVSS.n1862 4.6505
R31699 DVSS.n6750 DVSS.n2 4.6505
R31700 DVSS.n1876 DVSS.n1875 4.6505
R31701 DVSS.n1891 DVSS.n1890 4.6505
R31702 DVSS.n6868 DVSS.n8 4.6505
R31703 DVSS.n9 DVSS.n8 4.6505
R31704 DVSS.n6784 DVSS.n6783 4.6505
R31705 DVSS.n6808 DVSS.n10 4.6505
R31706 DVSS.n6825 DVSS.n6824 4.6505
R31707 DVSS.n6841 DVSS.n6840 4.6505
R31708 DVSS.n325 DVSS.n324 4.6505
R31709 DVSS.n345 DVSS.n344 4.6505
R31710 DVSS.n327 DVSS.n326 4.6505
R31711 DVSS.n330 DVSS.n177 4.6505
R31712 DVSS.n334 DVSS.n333 4.6505
R31713 DVSS.n336 DVSS.n335 4.6505
R31714 DVSS.n176 DVSS.n173 4.6505
R31715 DVSS.n161 DVSS.n159 4.6505
R31716 DVSS.n202 DVSS.n138 4.6505
R31717 DVSS.n233 DVSS.n232 4.6505
R31718 DVSS.n235 DVSS.n234 4.6505
R31719 DVSS.n219 DVSS.n214 4.6505
R31720 DVSS.n208 DVSS.n204 4.6505
R31721 DVSS.n243 DVSS.n242 4.6505
R31722 DVSS.n245 DVSS.n244 4.6505
R31723 DVSS.n221 DVSS.n220 4.6505
R31724 DVSS.n790 DVSS.n789 4.6505
R31725 DVSS.n810 DVSS.n809 4.6505
R31726 DVSS.n792 DVSS.n791 4.6505
R31727 DVSS.n795 DVSS.n642 4.6505
R31728 DVSS.n799 DVSS.n798 4.6505
R31729 DVSS.n801 DVSS.n800 4.6505
R31730 DVSS.n641 DVSS.n638 4.6505
R31731 DVSS.n626 DVSS.n624 4.6505
R31732 DVSS.n667 DVSS.n603 4.6505
R31733 DVSS.n698 DVSS.n697 4.6505
R31734 DVSS.n700 DVSS.n699 4.6505
R31735 DVSS.n684 DVSS.n679 4.6505
R31736 DVSS.n673 DVSS.n669 4.6505
R31737 DVSS.n708 DVSS.n707 4.6505
R31738 DVSS.n710 DVSS.n709 4.6505
R31739 DVSS.n686 DVSS.n685 4.6505
R31740 DVSS.n1403 DVSS.n1402 4.6505
R31741 DVSS.n1653 DVSS.n1652 4.6505
R31742 DVSS.n1732 DVSS.n1731 4.6505
R31743 DVSS.n6876 DVSS.n6875 4.6505
R31744 DVSS.n6872 DVSS.n6871 4.6505
R31745 DVSS.n6867 DVSS.n6866 4.6505
R31746 DVSS.n6862 DVSS.n6861 4.6505
R31747 DVSS.n6856 DVSS.n6855 4.6505
R31748 DVSS.n6853 DVSS.n6852 4.6505
R31749 DVSS.n6849 DVSS.n6848 4.6505
R31750 DVSS.n6845 DVSS.n6844 4.6505
R31751 DVSS.n6838 DVSS.n6837 4.6505
R31752 DVSS.n6833 DVSS.n6832 4.6505
R31753 DVSS.n6829 DVSS.n6828 4.6505
R31754 DVSS.n6821 DVSS.n6820 4.6505
R31755 DVSS.n6816 DVSS.n6815 4.6505
R31756 DVSS.n6812 DVSS.n6811 4.6505
R31757 DVSS.n6807 DVSS.n6806 4.6505
R31758 DVSS.n6801 DVSS.n6800 4.6505
R31759 DVSS.n6797 DVSS.n6796 4.6505
R31760 DVSS.n6793 DVSS.n6792 4.6505
R31761 DVSS.n6788 DVSS.n6787 4.6505
R31762 DVSS.n6779 DVSS.n6778 4.6505
R31763 DVSS.n6775 DVSS.n6774 4.6505
R31764 DVSS.n6771 DVSS.n6770 4.6505
R31765 DVSS.n6763 DVSS.n6762 4.6505
R31766 DVSS.n1782 DVSS.n1781 4.6505
R31767 DVSS.n1787 DVSS.n1786 4.6505
R31768 DVSS.n1792 DVSS.n1791 4.6505
R31769 DVSS.n1799 DVSS.n1798 4.6505
R31770 DVSS.n1803 DVSS.n1802 4.6505
R31771 DVSS.n1808 DVSS.n1807 4.6505
R31772 DVSS.n1816 DVSS.n1815 4.6505
R31773 DVSS.n1820 DVSS.n1819 4.6505
R31774 DVSS.n1824 DVSS.n1823 4.6505
R31775 DVSS.n1830 DVSS.n1829 4.6505
R31776 DVSS.n1834 DVSS.n1833 4.6505
R31777 DVSS.n1048 DVSS.n1047 4.6505
R31778 DVSS.n1122 DVSS.n1121 4.6505
R31779 DVSS.n1044 DVSS.n1043 4.6505
R31780 DVSS.n1032 DVSS.n1031 4.6505
R31781 DVSS.n1028 DVSS.n1027 4.6505
R31782 DVSS.n1024 DVSS.n1023 4.6505
R31783 DVSS.n1016 DVSS.n1015 4.6505
R31784 DVSS.n1035 DVSS.n1034 4.6505
R31785 DVSS.n1041 DVSS.n1040 4.6505
R31786 DVSS.n1013 DVSS.n1012 4.6505
R31787 DVSS.n967 DVSS.n966 4.6505
R31788 DVSS.n974 DVSS.n973 4.6505
R31789 DVSS.n977 DVSS.n976 4.6505
R31790 DVSS.n981 DVSS.n980 4.6505
R31791 DVSS.n984 DVSS.n983 4.6505
R31792 DVSS.n988 DVSS.n987 4.6505
R31793 DVSS.n991 DVSS.n990 4.6505
R31794 DVSS.n995 DVSS.n994 4.6505
R31795 DVSS.n998 DVSS.n997 4.6505
R31796 DVSS.n1002 DVSS.n1001 4.6505
R31797 DVSS.n1009 DVSS.n1008 4.6505
R31798 DVSS.n1088 DVSS.n1087 4.6505
R31799 DVSS.n1051 DVSS.n1050 4.6505
R31800 DVSS.n1068 DVSS.n1067 4.6505
R31801 DVSS.n1071 DVSS.n1070 4.6505
R31802 DVSS.n1075 DVSS.n1074 4.6505
R31803 DVSS.n1081 DVSS.n1080 4.6505
R31804 DVSS.n1085 DVSS.n1084 4.6505
R31805 DVSS.n1199 DVSS.n1198 4.6505
R31806 DVSS.n1172 DVSS.n1159 4.6505
R31807 DVSS.n1224 DVSS.n1223 4.6505
R31808 DVSS.n1215 DVSS.n1214 4.6505
R31809 DVSS.n1211 DVSS.n1210 4.6505
R31810 DVSS.n1208 DVSS.n1207 4.6505
R31811 DVSS.n1204 DVSS.n1203 4.6505
R31812 DVSS.n1201 DVSS.n1200 4.6505
R31813 DVSS.n1195 DVSS.n1194 4.6505
R31814 DVSS.n1191 DVSS.n1190 4.6505
R31815 DVSS.n1187 DVSS.n1186 4.6505
R31816 DVSS.n1184 DVSS.n1183 4.6505
R31817 DVSS.n1177 DVSS.n1176 4.6505
R31818 DVSS.n1174 DVSS.n1173 4.6505
R31819 DVSS.n1171 DVSS.n1170 4.6505
R31820 DVSS.n1165 DVSS.n1164 4.6505
R31821 DVSS.n1162 DVSS.n1161 4.6505
R31822 DVSS.n1263 DVSS.n1262 4.6505
R31823 DVSS.n1285 DVSS.n1284 4.6505
R31824 DVSS.n1300 DVSS.n1299 4.6505
R31825 DVSS.n1315 DVSS.n1314 4.6505
R31826 DVSS.n1329 DVSS.n1328 4.6505
R31827 DVSS.n1233 DVSS.n1232 4.6505
R31828 DVSS.n1237 DVSS.n1236 4.6505
R31829 DVSS.n1241 DVSS.n1240 4.6505
R31830 DVSS.n1246 DVSS.n1245 4.6505
R31831 DVSS.n1250 DVSS.n1249 4.6505
R31832 DVSS.n1254 DVSS.n1253 4.6505
R31833 DVSS.n1258 DVSS.n1257 4.6505
R31834 DVSS.n1267 DVSS.n1266 4.6505
R31835 DVSS.n1272 DVSS.n1271 4.6505
R31836 DVSS.n1276 DVSS.n1275 4.6505
R31837 DVSS.n1279 DVSS.n1278 4.6505
R31838 DVSS.n1283 DVSS.n1282 4.6505
R31839 DVSS.n1288 DVSS.n1287 4.6505
R31840 DVSS.n1292 DVSS.n1291 4.6505
R31841 DVSS.n1296 DVSS.n1295 4.6505
R31842 DVSS.n1304 DVSS.n1303 4.6505
R31843 DVSS.n1307 DVSS.n1306 4.6505
R31844 DVSS.n1312 DVSS.n1311 4.6505
R31845 DVSS.n1318 DVSS.n1317 4.6505
R31846 DVSS.n1325 DVSS.n1324 4.6505
R31847 DVSS.n1340 DVSS.n1339 4.6505
R31848 DVSS.n1338 DVSS.n1330 4.6505
R31849 DVSS.n1337 DVSS.n1336 4.6505
R31850 DVSS.n1142 DVSS.n1141 4.6505
R31851 DVSS.n1333 DVSS.n1332 4.6505
R31852 DVSS.n1153 DVSS.n1152 4.6505
R31853 DVSS.n1150 DVSS.n1149 4.6505
R31854 DVSS.n1145 DVSS.n1144 4.6505
R31855 DVSS.n1137 DVSS.n1136 4.6505
R31856 DVSS.n1133 DVSS.n1132 4.6505
R31857 DVSS.n1131 DVSS.n1130 4.6505
R31858 DVSS.n1487 DVSS.n1486 4.51815
R31859 DVSS.n1558 DVSS.n1557 4.51815
R31860 DVSS.n4700 DVSS.n4699 4.51815
R31861 DVSS.n4771 DVSS.n4770 4.51815
R31862 DVSS.n6168 DVSS.n6167 4.51815
R31863 DVSS.n6239 DVSS.n6238 4.51815
R31864 DVSS.n3104 DVSS.n3103 4.51815
R31865 DVSS.n3175 DVSS.n3174 4.51815
R31866 DVSS.n3946 DVSS.n3714 4.5005
R31867 DVSS.n4411 DVSS.n4179 4.5005
R31868 DVSS.n5054 DVSS.n5053 4.5005
R31869 DVSS.n2350 DVSS.n2118 4.5005
R31870 DVSS.n2815 DVSS.n2583 4.5005
R31871 DVSS.n2010 DVSS.n2009 4.5005
R31872 DVSS.n3459 DVSS.n3458 4.5005
R31873 DVSS.n5414 DVSS.n5182 4.5005
R31874 DVSS.n5879 DVSS.n5647 4.5005
R31875 DVSS.n6520 DVSS.n6519 4.5005
R31876 DVSS.n6540 DVSS.n6539 4.5005
R31877 DVSS.n349 DVSS.n117 4.5005
R31878 DVSS.n814 DVSS.n582 4.5005
R31879 DVSS.n1842 DVSS.n1841 4.5005
R31880 DVSS.n3952 DVSS.n3951 4.40783
R31881 DVSS.n4417 DVSS.n4416 4.40783
R31882 DVSS.n2356 DVSS.n2355 4.40783
R31883 DVSS.n2821 DVSS.n2820 4.40783
R31884 DVSS.n5420 DVSS.n5419 4.40783
R31885 DVSS.n5885 DVSS.n5884 4.40783
R31886 DVSS.n355 DVSS.n354 4.40783
R31887 DVSS.n820 DVSS.n819 4.40783
R31888 DVSS.n1274 DVSS.n1273 4.35669
R31889 DVSS.n1169 DVSS.n1168 4.35669
R31890 DVSS.n3843 DVSS.n3799 4.31208
R31891 DVSS.n4308 DVSS.n4264 4.31208
R31892 DVSS.n2247 DVSS.n2203 4.31208
R31893 DVSS.n2712 DVSS.n2668 4.31208
R31894 DVSS.n5311 DVSS.n5267 4.31208
R31895 DVSS.n5776 DVSS.n5732 4.31208
R31896 DVSS.n246 DVSS.n202 4.31208
R31897 DVSS.n711 DVSS.n667 4.31208
R31898 DVSS.n1361 DVSS.n1353 4.14168
R31899 DVSS.n1450 DVSS.n1442 4.14168
R31900 DVSS.n1611 DVSS.n1603 4.14168
R31901 DVSS.n1700 DVSS.n1692 4.14168
R31902 DVSS.n4574 DVSS.n4566 4.14168
R31903 DVSS.n4663 DVSS.n4655 4.14168
R31904 DVSS.n4824 DVSS.n4816 4.14168
R31905 DVSS.n4913 DVSS.n4905 4.14168
R31906 DVSS.n6042 DVSS.n6034 4.14168
R31907 DVSS.n6131 DVSS.n6123 4.14168
R31908 DVSS.n6292 DVSS.n6284 4.14168
R31909 DVSS.n6381 DVSS.n6373 4.14168
R31910 DVSS.n2978 DVSS.n2970 4.14168
R31911 DVSS.n3067 DVSS.n3059 4.14168
R31912 DVSS.n3228 DVSS.n3220 4.14168
R31913 DVSS.n3317 DVSS.n3309 4.14168
R31914 DVSS.n3842 DVSS.n3800 4.04261
R31915 DVSS.n4307 DVSS.n4265 4.04261
R31916 DVSS.n2246 DVSS.n2204 4.04261
R31917 DVSS.n2711 DVSS.n2669 4.04261
R31918 DVSS.n5310 DVSS.n5268 4.04261
R31919 DVSS.n5775 DVSS.n5733 4.04261
R31920 DVSS.n245 DVSS.n203 4.04261
R31921 DVSS.n710 DVSS.n668 4.04261
R31922 DVSS.n3753 DVSS.n3738 3.93153
R31923 DVSS.n3732 DVSS.n3717 3.93153
R31924 DVSS.n4218 DVSS.n4203 3.93153
R31925 DVSS.n4197 DVSS.n4182 3.93153
R31926 DVSS.n2157 DVSS.n2142 3.93153
R31927 DVSS.n2136 DVSS.n2121 3.93153
R31928 DVSS.n2622 DVSS.n2607 3.93153
R31929 DVSS.n2601 DVSS.n2586 3.93153
R31930 DVSS.n5221 DVSS.n5206 3.93153
R31931 DVSS.n5200 DVSS.n5185 3.93153
R31932 DVSS.n5686 DVSS.n5671 3.93153
R31933 DVSS.n5665 DVSS.n5650 3.93153
R31934 DVSS.n156 DVSS.n141 3.93153
R31935 DVSS.n135 DVSS.n120 3.93153
R31936 DVSS.n621 DVSS.n606 3.93153
R31937 DVSS.n600 DVSS.n585 3.93153
R31938 DVSS.n3799 DVSS.n3786 3.8405
R31939 DVSS.n4264 DVSS.n4251 3.8405
R31940 DVSS.n2203 DVSS.n2190 3.8405
R31941 DVSS.n2668 DVSS.n2655 3.8405
R31942 DVSS.n5267 DVSS.n5254 3.8405
R31943 DVSS.n5732 DVSS.n5719 3.8405
R31944 DVSS.n202 DVSS.n189 3.8405
R31945 DVSS.n667 DVSS.n654 3.8405
R31946 DVSS.n3839 DVSS.n3838 3.77313
R31947 DVSS.n4304 DVSS.n4303 3.77313
R31948 DVSS.n2243 DVSS.n2242 3.77313
R31949 DVSS.n2708 DVSS.n2707 3.77313
R31950 DVSS.n5307 DVSS.n5306 3.77313
R31951 DVSS.n5772 DVSS.n5771 3.77313
R31952 DVSS.n242 DVSS.n241 3.77313
R31953 DVSS.n707 DVSS.n706 3.77313
R31954 DVSS.n1472 DVSS.n1471 3.76521
R31955 DVSS.n1573 DVSS.n1572 3.76521
R31956 DVSS.n4685 DVSS.n4684 3.76521
R31957 DVSS.n4786 DVSS.n4785 3.76521
R31958 DVSS.n6153 DVSS.n6152 3.76521
R31959 DVSS.n6254 DVSS.n6253 3.76521
R31960 DVSS.n3089 DVSS.n3088 3.76521
R31961 DVSS.n3190 DVSS.n3189 3.76521
R31962 DVSS.n1222 DVSS.n1221 3.69563
R31963 DVSS.n1746 DVSS.n1745 3.69446
R31964 DVSS.n4958 DVSS.n4957 3.69446
R31965 DVSS.n3363 DVSS.n3360 3.69446
R31966 DVSS.n6426 DVSS.n6425 3.69446
R31967 DVSS.n1299 DVSS.n1298 3.68864
R31968 DVSS.n1021 DVSS.n1019 3.68864
R31969 DVSS.n1811 DVSS.n1809 3.68864
R31970 DVSS.n6824 DVSS.n6823 3.68864
R31971 DVSS.n3541 DVSS.n3540 3.68864
R31972 DVSS.n6613 DVSS.n6612 3.68864
R31973 DVSS.n5023 DVSS.n5021 3.68864
R31974 DVSS.n1938 DVSS.n1937 3.68864
R31975 DVSS.n3428 DVSS.n3426 3.68864
R31976 DVSS.n6491 DVSS.n6489 3.68864
R31977 DVSS.n3809 DVSS.n3805 3.50366
R31978 DVSS.n4274 DVSS.n4270 3.50366
R31979 DVSS.n2213 DVSS.n2209 3.50366
R31980 DVSS.n2678 DVSS.n2674 3.50366
R31981 DVSS.n5277 DVSS.n5273 3.50366
R31982 DVSS.n5742 DVSS.n5738 3.50366
R31983 DVSS.n212 DVSS.n208 3.50366
R31984 DVSS.n677 DVSS.n673 3.50366
R31985 DVSS.n1465 DVSS.n1457 3.38874
R31986 DVSS.n1596 DVSS.n1588 3.38874
R31987 DVSS.n4678 DVSS.n4670 3.38874
R31988 DVSS.n4809 DVSS.n4801 3.38874
R31989 DVSS.n6146 DVSS.n6138 3.38874
R31990 DVSS.n6277 DVSS.n6269 3.38874
R31991 DVSS.n3082 DVSS.n3074 3.38874
R31992 DVSS.n3213 DVSS.n3205 3.38874
R31993 DVSS.n1524 DVSS.n1519 3.2936
R31994 DVSS.n1535 DVSS.n1530 3.2936
R31995 DVSS.n4737 DVSS.n4732 3.2936
R31996 DVSS.n4748 DVSS.n4743 3.2936
R31997 DVSS.n6205 DVSS.n6200 3.2936
R31998 DVSS.n6216 DVSS.n6211 3.2936
R31999 DVSS.n3141 DVSS.n3136 3.2936
R32000 DVSS.n3152 DVSS.n3147 3.2936
R32001 DVSS.n3833 DVSS.n3811 3.23418
R32002 DVSS.n4298 DVSS.n4276 3.23418
R32003 DVSS.n2237 DVSS.n2215 3.23418
R32004 DVSS.n2702 DVSS.n2680 3.23418
R32005 DVSS.n5301 DVSS.n5279 3.23418
R32006 DVSS.n5766 DVSS.n5744 3.23418
R32007 DVSS.n236 DVSS.n214 3.23418
R32008 DVSS.n701 DVSS.n679 3.23418
R32009 DVSS.n3947 DVSS.n3945 3.20387
R32010 DVSS.n4412 DVSS.n4410 3.20387
R32011 DVSS.n2351 DVSS.n2349 3.20387
R32012 DVSS.n2816 DVSS.n2814 3.20387
R32013 DVSS.n5415 DVSS.n5413 3.20387
R32014 DVSS.n5880 DVSS.n5878 3.20387
R32015 DVSS.n350 DVSS.n348 3.20387
R32016 DVSS.n815 DVSS.n813 3.20387
R32017 DVSS.n4950 DVSS.n4949 3.0928
R32018 DVSS.n3355 DVSS.n3354 3.0928
R32019 DVSS.n6418 DVSS.n6417 3.0928
R32020 DVSS.n1737 DVSS.n1736 3.0928
R32021 DVSS.n6884 DVSS.n6883 3.07616
R32022 DVSS.n3467 DVSS.n3466 3.03311
R32023 DVSS.n3474 DVSS.n3473 3.03311
R32024 DVSS.n5062 DVSS.n5061 3.03311
R32025 DVSS.n6528 DVSS.n6527 3.03311
R32026 DVSS.n6536 DVSS.n6535 3.03311
R32027 DVSS.n6709 DVSS.n5068 3.03311
R32028 DVSS.n6744 DVSS.n1856 3.03311
R32029 DVSS.n1850 DVSS.n1849 3.03311
R32030 DVSS.n1457 DVSS.n1456 3.01226
R32031 DVSS.n1588 DVSS.n1587 3.01226
R32032 DVSS.n4670 DVSS.n4669 3.01226
R32033 DVSS.n4801 DVSS.n4800 3.01226
R32034 DVSS.n6138 DVSS.n6137 3.01226
R32035 DVSS.n6269 DVSS.n6268 3.01226
R32036 DVSS.n3074 DVSS.n3073 3.01226
R32037 DVSS.n3205 DVSS.n3204 3.01226
R32038 DVSS.n3832 DVSS.n3815 2.96471
R32039 DVSS.n4297 DVSS.n4280 2.96471
R32040 DVSS.n2236 DVSS.n2219 2.96471
R32041 DVSS.n2701 DVSS.n2684 2.96471
R32042 DVSS.n5300 DVSS.n5283 2.96471
R32043 DVSS.n5765 DVSS.n5748 2.96471
R32044 DVSS.n235 DVSS.n218 2.96471
R32045 DVSS.n700 DVSS.n683 2.96471
R32046 DVSS.n1262 DVSS.n1261 2.84494
R32047 DVSS.n6783 DVSS.n6782 2.84494
R32048 DVSS.n3583 DVSS.n3582 2.84494
R32049 DVSS.n6571 DVSS.n6570 2.84494
R32050 DVSS.n1980 DVSS.n1979 2.84494
R32051 DVSS.n3829 DVSS.n3828 2.69524
R32052 DVSS.n4294 DVSS.n4293 2.69524
R32053 DVSS.n2233 DVSS.n2232 2.69524
R32054 DVSS.n2698 DVSS.n2697 2.69524
R32055 DVSS.n5297 DVSS.n5296 2.69524
R32056 DVSS.n5762 DVSS.n5761 2.69524
R32057 DVSS.n232 DVSS.n231 2.69524
R32058 DVSS.n697 DVSS.n696 2.69524
R32059 DVSS.n1480 DVSS.n1472 2.63579
R32060 DVSS.n1581 DVSS.n1573 2.63579
R32061 DVSS.n4693 DVSS.n4685 2.63579
R32062 DVSS.n4794 DVSS.n4786 2.63579
R32063 DVSS.n6161 DVSS.n6153 2.63579
R32064 DVSS.n6262 DVSS.n6254 2.63579
R32065 DVSS.n3097 DVSS.n3089 2.63579
R32066 DVSS.n3198 DVSS.n3190 2.63579
R32067 DVSS.n3921 DVSS.n3920 2.5605
R32068 DVSS.n4386 DVSS.n4385 2.5605
R32069 DVSS.n2325 DVSS.n2324 2.5605
R32070 DVSS.n2790 DVSS.n2789 2.5605
R32071 DVSS.n5389 DVSS.n5388 2.5605
R32072 DVSS.n5854 DVSS.n5853 2.5605
R32073 DVSS.n324 DVSS.n323 2.5605
R32074 DVSS.n789 DVSS.n788 2.5605
R32075 DVSS.n3824 DVSS.n3818 2.42576
R32076 DVSS.n3824 DVSS.n3792 2.42576
R32077 DVSS.n4289 DVSS.n4283 2.42576
R32078 DVSS.n4289 DVSS.n4257 2.42576
R32079 DVSS.n2228 DVSS.n2222 2.42576
R32080 DVSS.n2228 DVSS.n2196 2.42576
R32081 DVSS.n2693 DVSS.n2687 2.42576
R32082 DVSS.n2693 DVSS.n2661 2.42576
R32083 DVSS.n5292 DVSS.n5286 2.42576
R32084 DVSS.n5292 DVSS.n5260 2.42576
R32085 DVSS.n5757 DVSS.n5751 2.42576
R32086 DVSS.n5757 DVSS.n5725 2.42576
R32087 DVSS.n227 DVSS.n221 2.42576
R32088 DVSS.n227 DVSS.n195 2.42576
R32089 DVSS.n692 DVSS.n686 2.42576
R32090 DVSS.n692 DVSS.n660 2.42576
R32091 DVSS.n1039 DVSS.n1038 2.31779
R32092 DVSS.n1826 DVSS.n1825 2.31469
R32093 DVSS.n5038 DVSS.n5037 2.31469
R32094 DVSS.n3443 DVSS.n3442 2.31469
R32095 DVSS.n6507 DVSS.n6506 2.31469
R32096 DVSS.n3782 DVSS.n3776 2.29103
R32097 DVSS.n4247 DVSS.n4241 2.29103
R32098 DVSS.n2186 DVSS.n2180 2.29103
R32099 DVSS.n2651 DVSS.n2645 2.29103
R32100 DVSS.n5250 DVSS.n5244 2.29103
R32101 DVSS.n5715 DVSS.n5709 2.29103
R32102 DVSS.n185 DVSS.n179 2.29103
R32103 DVSS.n650 DVSS.n644 2.29103
R32104 DVSS.n1353 DVSS.n1352 2.25932
R32105 DVSS.n1442 DVSS.n1441 2.25932
R32106 DVSS.n1603 DVSS.n1602 2.25932
R32107 DVSS.n1692 DVSS.n1691 2.25932
R32108 DVSS.n4566 DVSS.n4565 2.25932
R32109 DVSS.n4655 DVSS.n4654 2.25932
R32110 DVSS.n4816 DVSS.n4815 2.25932
R32111 DVSS.n4905 DVSS.n4904 2.25932
R32112 DVSS.n6034 DVSS.n6033 2.25932
R32113 DVSS.n6123 DVSS.n6122 2.25932
R32114 DVSS.n6284 DVSS.n6283 2.25932
R32115 DVSS.n6373 DVSS.n6372 2.25932
R32116 DVSS.n2970 DVSS.n2969 2.25932
R32117 DVSS.n3059 DVSS.n3058 2.25932
R32118 DVSS.n3220 DVSS.n3219 2.25932
R32119 DVSS.n3309 DVSS.n3308 2.25932
R32120 DVSS.n1054 DVSS.n969 2.16799
R32121 DVSS.n3828 DVSS.n3818 2.15629
R32122 DVSS.n3886 DVSS.n3792 2.15629
R32123 DVSS.n4293 DVSS.n4283 2.15629
R32124 DVSS.n4351 DVSS.n4257 2.15629
R32125 DVSS.n2232 DVSS.n2222 2.15629
R32126 DVSS.n2290 DVSS.n2196 2.15629
R32127 DVSS.n2697 DVSS.n2687 2.15629
R32128 DVSS.n2755 DVSS.n2661 2.15629
R32129 DVSS.n5296 DVSS.n5286 2.15629
R32130 DVSS.n5354 DVSS.n5260 2.15629
R32131 DVSS.n5761 DVSS.n5751 2.15629
R32132 DVSS.n5819 DVSS.n5725 2.15629
R32133 DVSS.n231 DVSS.n221 2.15629
R32134 DVSS.n289 DVSS.n195 2.15629
R32135 DVSS.n696 DVSS.n686 2.15629
R32136 DVSS.n754 DVSS.n660 2.15629
R32137 DVSS.n3829 DVSS.n3815 1.88682
R32138 DVSS.n4294 DVSS.n4280 1.88682
R32139 DVSS.n2233 DVSS.n2219 1.88682
R32140 DVSS.n2698 DVSS.n2684 1.88682
R32141 DVSS.n5297 DVSS.n5283 1.88682
R32142 DVSS.n5762 DVSS.n5748 1.88682
R32143 DVSS.n232 DVSS.n218 1.88682
R32144 DVSS.n697 DVSS.n683 1.88682
R32145 DVSS.n1495 DVSS.n1487 1.88285
R32146 DVSS.n1566 DVSS.n1558 1.88285
R32147 DVSS.n4708 DVSS.n4700 1.88285
R32148 DVSS.n4779 DVSS.n4771 1.88285
R32149 DVSS.n6176 DVSS.n6168 1.88285
R32150 DVSS.n6247 DVSS.n6239 1.88285
R32151 DVSS.n3112 DVSS.n3104 1.88285
R32152 DVSS.n3183 DVSS.n3175 1.88285
R32153 DVSS DVSS.n6722 1.77928
R32154 DVSS.n3920 DVSS.n3918 1.68471
R32155 DVSS.n3914 DVSS.n3782 1.68471
R32156 DVSS.n4385 DVSS.n4383 1.68471
R32157 DVSS.n4379 DVSS.n4247 1.68471
R32158 DVSS.n2324 DVSS.n2322 1.68471
R32159 DVSS.n2318 DVSS.n2186 1.68471
R32160 DVSS.n2789 DVSS.n2787 1.68471
R32161 DVSS.n2783 DVSS.n2651 1.68471
R32162 DVSS.n5388 DVSS.n5386 1.68471
R32163 DVSS.n5382 DVSS.n5250 1.68471
R32164 DVSS.n5853 DVSS.n5851 1.68471
R32165 DVSS.n5847 DVSS.n5715 1.68471
R32166 DVSS.n323 DVSS.n321 1.68471
R32167 DVSS.n317 DVSS.n185 1.68471
R32168 DVSS.n788 DVSS.n786 1.68471
R32169 DVSS.n782 DVSS.n650 1.68471
R32170 DVSS.n3941 DVSS.n3940 1.64728
R32171 DVSS.n4406 DVSS.n4405 1.64728
R32172 DVSS.n2345 DVSS.n2344 1.64728
R32173 DVSS.n2810 DVSS.n2809 1.64728
R32174 DVSS.n5409 DVSS.n5408 1.64728
R32175 DVSS.n5874 DVSS.n5873 1.64728
R32176 DVSS.n344 DVSS.n343 1.64728
R32177 DVSS.n809 DVSS.n808 1.64728
R32178 DVSS.n3833 DVSS.n3832 1.61734
R32179 DVSS.n4298 DVSS.n4297 1.61734
R32180 DVSS.n2237 DVSS.n2236 1.61734
R32181 DVSS.n2702 DVSS.n2701 1.61734
R32182 DVSS.n5301 DVSS.n5300 1.61734
R32183 DVSS.n5766 DVSS.n5765 1.61734
R32184 DVSS.n236 DVSS.n235 1.61734
R32185 DVSS.n701 DVSS.n700 1.61734
R32186 DVSS.n3952 DVSS.n3685 1.59464
R32187 DVSS.n3959 DVSS.n3685 1.59464
R32188 DVSS.n3959 DVSS.n3686 1.59464
R32189 DVSS.n3955 DVSS.n3686 1.59464
R32190 DVSS.n3955 DVSS.n3652 1.59464
R32191 DVSS.n3969 DVSS.n3652 1.59464
R32192 DVSS.n3979 DVSS.n3650 1.59464
R32193 DVSS.n3974 DVSS.n3638 1.59464
R32194 DVSS.n3990 DVSS.n3638 1.59464
R32195 DVSS.n3991 DVSS.n3990 1.59464
R32196 DVSS.n3991 DVSS.n3636 1.59464
R32197 DVSS.n3997 DVSS.n3996 1.59464
R32198 DVSS.n3997 DVSS.n3633 1.59464
R32199 DVSS.n4027 DVSS.n3633 1.59464
R32200 DVSS.n4023 DVSS.n3618 1.59464
R32201 DVSS.n4061 DVSS.n3618 1.59464
R32202 DVSS.n4062 DVSS.n4061 1.59464
R32203 DVSS.n4063 DVSS.n4062 1.59464
R32204 DVSS.n4063 DVSS.n3616 1.59464
R32205 DVSS.n4068 DVSS.n3616 1.59464
R32206 DVSS.n4417 DVSS.n4150 1.59464
R32207 DVSS.n4424 DVSS.n4150 1.59464
R32208 DVSS.n4424 DVSS.n4151 1.59464
R32209 DVSS.n4420 DVSS.n4151 1.59464
R32210 DVSS.n4420 DVSS.n4117 1.59464
R32211 DVSS.n4434 DVSS.n4117 1.59464
R32212 DVSS.n4444 DVSS.n4115 1.59464
R32213 DVSS.n4439 DVSS.n4103 1.59464
R32214 DVSS.n4455 DVSS.n4103 1.59464
R32215 DVSS.n4456 DVSS.n4455 1.59464
R32216 DVSS.n4456 DVSS.n4101 1.59464
R32217 DVSS.n4462 DVSS.n4461 1.59464
R32218 DVSS.n4462 DVSS.n4098 1.59464
R32219 DVSS.n4492 DVSS.n4098 1.59464
R32220 DVSS.n4488 DVSS.n4083 1.59464
R32221 DVSS.n4526 DVSS.n4083 1.59464
R32222 DVSS.n4527 DVSS.n4526 1.59464
R32223 DVSS.n4528 DVSS.n4527 1.59464
R32224 DVSS.n4528 DVSS.n4081 1.59464
R32225 DVSS.n4532 DVSS.n4081 1.59464
R32226 DVSS.n2356 DVSS.n2089 1.59464
R32227 DVSS.n2363 DVSS.n2089 1.59464
R32228 DVSS.n2363 DVSS.n2090 1.59464
R32229 DVSS.n2359 DVSS.n2090 1.59464
R32230 DVSS.n2359 DVSS.n2056 1.59464
R32231 DVSS.n2373 DVSS.n2056 1.59464
R32232 DVSS.n2383 DVSS.n2054 1.59464
R32233 DVSS.n2378 DVSS.n2042 1.59464
R32234 DVSS.n2394 DVSS.n2042 1.59464
R32235 DVSS.n2395 DVSS.n2394 1.59464
R32236 DVSS.n2395 DVSS.n2040 1.59464
R32237 DVSS.n2401 DVSS.n2400 1.59464
R32238 DVSS.n2401 DVSS.n2037 1.59464
R32239 DVSS.n2431 DVSS.n2037 1.59464
R32240 DVSS.n2427 DVSS.n2022 1.59464
R32241 DVSS.n2465 DVSS.n2022 1.59464
R32242 DVSS.n2466 DVSS.n2465 1.59464
R32243 DVSS.n2467 DVSS.n2466 1.59464
R32244 DVSS.n2467 DVSS.n2020 1.59464
R32245 DVSS.n2472 DVSS.n2020 1.59464
R32246 DVSS.n2821 DVSS.n2554 1.59464
R32247 DVSS.n2828 DVSS.n2554 1.59464
R32248 DVSS.n2828 DVSS.n2555 1.59464
R32249 DVSS.n2824 DVSS.n2555 1.59464
R32250 DVSS.n2824 DVSS.n2521 1.59464
R32251 DVSS.n2838 DVSS.n2521 1.59464
R32252 DVSS.n2848 DVSS.n2519 1.59464
R32253 DVSS.n2843 DVSS.n2507 1.59464
R32254 DVSS.n2859 DVSS.n2507 1.59464
R32255 DVSS.n2860 DVSS.n2859 1.59464
R32256 DVSS.n2860 DVSS.n2505 1.59464
R32257 DVSS.n2866 DVSS.n2865 1.59464
R32258 DVSS.n2866 DVSS.n2502 1.59464
R32259 DVSS.n2896 DVSS.n2502 1.59464
R32260 DVSS.n2892 DVSS.n2487 1.59464
R32261 DVSS.n2930 DVSS.n2487 1.59464
R32262 DVSS.n2931 DVSS.n2930 1.59464
R32263 DVSS.n2932 DVSS.n2931 1.59464
R32264 DVSS.n2932 DVSS.n2485 1.59464
R32265 DVSS.n2936 DVSS.n2485 1.59464
R32266 DVSS.n5420 DVSS.n5153 1.59464
R32267 DVSS.n5427 DVSS.n5153 1.59464
R32268 DVSS.n5427 DVSS.n5154 1.59464
R32269 DVSS.n5423 DVSS.n5154 1.59464
R32270 DVSS.n5423 DVSS.n5120 1.59464
R32271 DVSS.n5437 DVSS.n5120 1.59464
R32272 DVSS.n5447 DVSS.n5118 1.59464
R32273 DVSS.n5442 DVSS.n5106 1.59464
R32274 DVSS.n5458 DVSS.n5106 1.59464
R32275 DVSS.n5459 DVSS.n5458 1.59464
R32276 DVSS.n5459 DVSS.n5104 1.59464
R32277 DVSS.n5465 DVSS.n5464 1.59464
R32278 DVSS.n5465 DVSS.n5101 1.59464
R32279 DVSS.n5495 DVSS.n5101 1.59464
R32280 DVSS.n5491 DVSS.n5086 1.59464
R32281 DVSS.n5529 DVSS.n5086 1.59464
R32282 DVSS.n5530 DVSS.n5529 1.59464
R32283 DVSS.n5531 DVSS.n5530 1.59464
R32284 DVSS.n5531 DVSS.n5084 1.59464
R32285 DVSS.n5536 DVSS.n5084 1.59464
R32286 DVSS.n5885 DVSS.n5618 1.59464
R32287 DVSS.n5892 DVSS.n5618 1.59464
R32288 DVSS.n5892 DVSS.n5619 1.59464
R32289 DVSS.n5888 DVSS.n5619 1.59464
R32290 DVSS.n5888 DVSS.n5585 1.59464
R32291 DVSS.n5902 DVSS.n5585 1.59464
R32292 DVSS.n5912 DVSS.n5583 1.59464
R32293 DVSS.n5907 DVSS.n5571 1.59464
R32294 DVSS.n5923 DVSS.n5571 1.59464
R32295 DVSS.n5924 DVSS.n5923 1.59464
R32296 DVSS.n5924 DVSS.n5569 1.59464
R32297 DVSS.n5930 DVSS.n5929 1.59464
R32298 DVSS.n5930 DVSS.n5566 1.59464
R32299 DVSS.n5960 DVSS.n5566 1.59464
R32300 DVSS.n5956 DVSS.n5551 1.59464
R32301 DVSS.n5994 DVSS.n5551 1.59464
R32302 DVSS.n5995 DVSS.n5994 1.59464
R32303 DVSS.n5996 DVSS.n5995 1.59464
R32304 DVSS.n5996 DVSS.n5549 1.59464
R32305 DVSS.n6000 DVSS.n5549 1.59464
R32306 DVSS.n355 DVSS.n88 1.59464
R32307 DVSS.n362 DVSS.n88 1.59464
R32308 DVSS.n362 DVSS.n89 1.59464
R32309 DVSS.n358 DVSS.n89 1.59464
R32310 DVSS.n358 DVSS.n55 1.59464
R32311 DVSS.n372 DVSS.n55 1.59464
R32312 DVSS.n382 DVSS.n53 1.59464
R32313 DVSS.n377 DVSS.n41 1.59464
R32314 DVSS.n393 DVSS.n41 1.59464
R32315 DVSS.n394 DVSS.n393 1.59464
R32316 DVSS.n394 DVSS.n39 1.59464
R32317 DVSS.n400 DVSS.n399 1.59464
R32318 DVSS.n400 DVSS.n36 1.59464
R32319 DVSS.n430 DVSS.n36 1.59464
R32320 DVSS.n426 DVSS.n21 1.59464
R32321 DVSS.n464 DVSS.n21 1.59464
R32322 DVSS.n465 DVSS.n464 1.59464
R32323 DVSS.n466 DVSS.n465 1.59464
R32324 DVSS.n466 DVSS.n19 1.59464
R32325 DVSS.n471 DVSS.n19 1.59464
R32326 DVSS.n820 DVSS.n553 1.59464
R32327 DVSS.n827 DVSS.n553 1.59464
R32328 DVSS.n827 DVSS.n554 1.59464
R32329 DVSS.n823 DVSS.n554 1.59464
R32330 DVSS.n823 DVSS.n520 1.59464
R32331 DVSS.n837 DVSS.n520 1.59464
R32332 DVSS.n847 DVSS.n518 1.59464
R32333 DVSS.n842 DVSS.n506 1.59464
R32334 DVSS.n858 DVSS.n506 1.59464
R32335 DVSS.n859 DVSS.n858 1.59464
R32336 DVSS.n859 DVSS.n504 1.59464
R32337 DVSS.n865 DVSS.n864 1.59464
R32338 DVSS.n865 DVSS.n501 1.59464
R32339 DVSS.n895 DVSS.n501 1.59464
R32340 DVSS.n891 DVSS.n486 1.59464
R32341 DVSS.n929 DVSS.n486 1.59464
R32342 DVSS.n930 DVSS.n929 1.59464
R32343 DVSS.n931 DVSS.n930 1.59464
R32344 DVSS.n931 DVSS.n484 1.59464
R32345 DVSS.n935 DVSS.n484 1.59464
R32346 DVSS.n3769 DVSS.n3758 1.54748
R32347 DVSS.n4234 DVSS.n4223 1.54748
R32348 DVSS.n2173 DVSS.n2162 1.54748
R32349 DVSS.n2638 DVSS.n2627 1.54748
R32350 DVSS.n5237 DVSS.n5226 1.54748
R32351 DVSS.n5702 DVSS.n5691 1.54748
R32352 DVSS.n172 DVSS.n161 1.54748
R32353 DVSS.n637 DVSS.n626 1.54748
R32354 DVSS.n1368 DVSS.n1367 1.50638
R32355 DVSS.n1427 DVSS.n1426 1.50638
R32356 DVSS.n1618 DVSS.n1617 1.50638
R32357 DVSS.n1677 DVSS.n1676 1.50638
R32358 DVSS.n4581 DVSS.n4580 1.50638
R32359 DVSS.n4640 DVSS.n4639 1.50638
R32360 DVSS.n4831 DVSS.n4830 1.50638
R32361 DVSS.n4890 DVSS.n4889 1.50638
R32362 DVSS.n3739 DVSS.n3737 1.50638
R32363 DVSS.n3718 DVSS.n3716 1.50638
R32364 DVSS.n4204 DVSS.n4202 1.50638
R32365 DVSS.n4183 DVSS.n4181 1.50638
R32366 DVSS.n6049 DVSS.n6048 1.50638
R32367 DVSS.n6108 DVSS.n6107 1.50638
R32368 DVSS.n6299 DVSS.n6298 1.50638
R32369 DVSS.n6358 DVSS.n6357 1.50638
R32370 DVSS.n2985 DVSS.n2984 1.50638
R32371 DVSS.n3044 DVSS.n3043 1.50638
R32372 DVSS.n3235 DVSS.n3234 1.50638
R32373 DVSS.n3294 DVSS.n3293 1.50638
R32374 DVSS.n2143 DVSS.n2141 1.50638
R32375 DVSS.n2122 DVSS.n2120 1.50638
R32376 DVSS.n2608 DVSS.n2606 1.50638
R32377 DVSS.n2587 DVSS.n2585 1.50638
R32378 DVSS.n5207 DVSS.n5205 1.50638
R32379 DVSS.n5186 DVSS.n5184 1.50638
R32380 DVSS.n5672 DVSS.n5670 1.50638
R32381 DVSS.n5651 DVSS.n5649 1.50638
R32382 DVSS.n142 DVSS.n140 1.50638
R32383 DVSS.n121 DVSS.n119 1.50638
R32384 DVSS.n607 DVSS.n605 1.50638
R32385 DVSS.n586 DVSS.n584 1.50638
R32386 DVSS.n6878 DVSS.n2 1.47174
R32387 DVSS.n6722 DVSS.n6721 1.46851
R32388 DVSS.n3996 DVSS.n3995 1.45398
R32389 DVSS.n4461 DVSS.n4460 1.45398
R32390 DVSS.n2400 DVSS.n2399 1.45398
R32391 DVSS.n2865 DVSS.n2864 1.45398
R32392 DVSS.n5464 DVSS.n5463 1.45398
R32393 DVSS.n5929 DVSS.n5928 1.45398
R32394 DVSS.n399 DVSS.n398 1.45398
R32395 DVSS.n864 DVSS.n863 1.45398
R32396 DVSS.n3746 DVSS.n3745 1.45108
R32397 DVSS.n3725 DVSS.n3724 1.45108
R32398 DVSS.n4211 DVSS.n4210 1.45108
R32399 DVSS.n4190 DVSS.n4189 1.45108
R32400 DVSS.n2150 DVSS.n2149 1.45108
R32401 DVSS.n2129 DVSS.n2128 1.45108
R32402 DVSS.n2615 DVSS.n2614 1.45108
R32403 DVSS.n2594 DVSS.n2593 1.45108
R32404 DVSS.n5214 DVSS.n5213 1.45108
R32405 DVSS.n5193 DVSS.n5192 1.45108
R32406 DVSS.n5679 DVSS.n5678 1.45108
R32407 DVSS.n5658 DVSS.n5657 1.45108
R32408 DVSS.n149 DVSS.n148 1.45108
R32409 DVSS.n128 DVSS.n127 1.45108
R32410 DVSS.n614 DVSS.n613 1.45108
R32411 DVSS.n593 DVSS.n592 1.45108
R32412 DVSS.n3934 DVSS.n3770 1.44767
R32413 DVSS.n4399 DVSS.n4235 1.44767
R32414 DVSS.n2338 DVSS.n2174 1.44767
R32415 DVSS.n2803 DVSS.n2639 1.44767
R32416 DVSS.n5402 DVSS.n5238 1.44767
R32417 DVSS.n5867 DVSS.n5703 1.44767
R32418 DVSS.n337 DVSS.n173 1.44767
R32419 DVSS.n802 DVSS.n638 1.44767
R32420 DVSS.n3933 DVSS.n3772 1.34787
R32421 DVSS.n3811 DVSS.n3809 1.34787
R32422 DVSS.n4398 DVSS.n4237 1.34787
R32423 DVSS.n4276 DVSS.n4274 1.34787
R32424 DVSS.n2337 DVSS.n2176 1.34787
R32425 DVSS.n2215 DVSS.n2213 1.34787
R32426 DVSS.n2802 DVSS.n2641 1.34787
R32427 DVSS.n2680 DVSS.n2678 1.34787
R32428 DVSS.n5401 DVSS.n5240 1.34787
R32429 DVSS.n5279 DVSS.n5277 1.34787
R32430 DVSS.n5866 DVSS.n5705 1.34787
R32431 DVSS.n5744 DVSS.n5742 1.34787
R32432 DVSS.n336 DVSS.n175 1.34787
R32433 DVSS.n214 DVSS.n212 1.34787
R32434 DVSS.n801 DVSS.n640 1.34787
R32435 DVSS.n679 DVSS.n677 1.34787
R32436 DVSS.n3975 DVSS.n3974 1.26643
R32437 DVSS.n4440 DVSS.n4439 1.26643
R32438 DVSS.n2379 DVSS.n2378 1.26643
R32439 DVSS.n2844 DVSS.n2843 1.26643
R32440 DVSS.n5443 DVSS.n5442 1.26643
R32441 DVSS.n5908 DVSS.n5907 1.26643
R32442 DVSS.n378 DVSS.n377 1.26643
R32443 DVSS.n843 DVSS.n842 1.26643
R32444 DVSS.n3510 DVSS 1.2505
R32445 DVSS.n6854 DVSS 1.2505
R32446 DVSS.n3930 DVSS.n3929 1.24806
R32447 DVSS.n4395 DVSS.n4394 1.24806
R32448 DVSS.n2334 DVSS.n2333 1.24806
R32449 DVSS.n2799 DVSS.n2798 1.24806
R32450 DVSS.n5398 DVSS.n5397 1.24806
R32451 DVSS.n5863 DVSS.n5862 1.24806
R32452 DVSS.n333 DVSS.n332 1.24806
R32453 DVSS.n798 DVSS.n797 1.24806
R32454 DVSS.n3927 DVSS.n3926 1.14826
R32455 DVSS.n4392 DVSS.n4391 1.14826
R32456 DVSS.n2331 DVSS.n2330 1.14826
R32457 DVSS.n2796 DVSS.n2795 1.14826
R32458 DVSS.n5395 DVSS.n5394 1.14826
R32459 DVSS.n5860 DVSS.n5859 1.14826
R32460 DVSS.n330 DVSS.n329 1.14826
R32461 DVSS.n795 DVSS.n794 1.14826
R32462 DVSS.n1129 DVSS 1.13082
R32463 DVSS.n1510 DVSS.n1502 1.12991
R32464 DVSS.n1551 DVSS.n1543 1.12991
R32465 DVSS.n4723 DVSS.n4715 1.12991
R32466 DVSS.n4764 DVSS.n4756 1.12991
R32467 DVSS.n6191 DVSS.n6183 1.12991
R32468 DVSS.n6232 DVSS.n6224 1.12991
R32469 DVSS.n3127 DVSS.n3119 1.12991
R32470 DVSS.n3168 DVSS.n3160 1.12991
R32471 DVSS.n5065 DVSS.n5064 1.10762
R32472 DVSS.n3470 DVSS.n3469 1.10762
R32473 DVSS.n6531 DVSS.n6530 1.10762
R32474 DVSS.n1853 DVSS.n1852 1.10762
R32475 DVSS.n3921 DVSS.n3779 1.07839
R32476 DVSS.n3838 DVSS.n3805 1.07839
R32477 DVSS.n4386 DVSS.n4244 1.07839
R32478 DVSS.n4303 DVSS.n4270 1.07839
R32479 DVSS.n2325 DVSS.n2183 1.07839
R32480 DVSS.n2242 DVSS.n2209 1.07839
R32481 DVSS.n2790 DVSS.n2648 1.07839
R32482 DVSS.n2707 DVSS.n2674 1.07839
R32483 DVSS.n5389 DVSS.n5247 1.07839
R32484 DVSS.n5306 DVSS.n5273 1.07839
R32485 DVSS.n5854 DVSS.n5712 1.07839
R32486 DVSS.n5771 DVSS.n5738 1.07839
R32487 DVSS.n324 DVSS.n182 1.07839
R32488 DVSS.n241 DVSS.n208 1.07839
R32489 DVSS.n789 DVSS.n647 1.07839
R32490 DVSS.n706 DVSS.n673 1.07839
R32491 DVSS.n3924 DVSS.n3775 0.973599
R32492 DVSS.n4389 DVSS.n4240 0.973599
R32493 DVSS.n2328 DVSS.n2179 0.973599
R32494 DVSS.n2793 DVSS.n2644 0.973599
R32495 DVSS.n5392 DVSS.n5243 0.973599
R32496 DVSS.n5857 DVSS.n5708 0.973599
R32497 DVSS.n327 DVSS.n178 0.973599
R32498 DVSS.n792 DVSS.n643 0.973599
R32499 DVSS.n3839 DVSS.n3800 0.808921
R32500 DVSS.n4304 DVSS.n4265 0.808921
R32501 DVSS.n2243 DVSS.n2204 0.808921
R32502 DVSS.n2708 DVSS.n2669 0.808921
R32503 DVSS.n5307 DVSS.n5268 0.808921
R32504 DVSS.n5772 DVSS.n5733 0.808921
R32505 DVSS.n242 DVSS.n203 0.808921
R32506 DVSS.n707 DVSS.n668 0.808921
R32507 DVSS.n1383 DVSS.n1382 0.753441
R32508 DVSS.n1409 DVSS.n1408 0.753441
R32509 DVSS.n1633 DVSS.n1632 0.753441
R32510 DVSS.n1659 DVSS.n1658 0.753441
R32511 DVSS.n6714 DVSS.n3484 0.753441
R32512 DVSS.n4596 DVSS.n4595 0.753441
R32513 DVSS.n4622 DVSS.n4621 0.753441
R32514 DVSS.n4846 DVSS.n4845 0.753441
R32515 DVSS.n4872 DVSS.n4871 0.753441
R32516 DVSS.n3752 DVSS.n3751 0.753441
R32517 DVSS.n3743 DVSS.n3740 0.753441
R32518 DVSS.n3731 DVSS.n3730 0.753441
R32519 DVSS.n3722 DVSS.n3719 0.753441
R32520 DVSS.n4217 DVSS.n4216 0.753441
R32521 DVSS.n4208 DVSS.n4205 0.753441
R32522 DVSS.n4196 DVSS.n4195 0.753441
R32523 DVSS.n4187 DVSS.n4184 0.753441
R32524 DVSS.n6064 DVSS.n6063 0.753441
R32525 DVSS.n6090 DVSS.n6089 0.753441
R32526 DVSS.n6314 DVSS.n6313 0.753441
R32527 DVSS.n6340 DVSS.n6339 0.753441
R32528 DVSS.n3000 DVSS.n2999 0.753441
R32529 DVSS.n3026 DVSS.n3025 0.753441
R32530 DVSS.n3250 DVSS.n3249 0.753441
R32531 DVSS.n3276 DVSS.n3275 0.753441
R32532 DVSS.n6756 DVSS.n6748 0.753441
R32533 DVSS.n2156 DVSS.n2155 0.753441
R32534 DVSS.n2147 DVSS.n2144 0.753441
R32535 DVSS.n2135 DVSS.n2134 0.753441
R32536 DVSS.n2126 DVSS.n2123 0.753441
R32537 DVSS.n2621 DVSS.n2620 0.753441
R32538 DVSS.n2612 DVSS.n2609 0.753441
R32539 DVSS.n2600 DVSS.n2599 0.753441
R32540 DVSS.n2591 DVSS.n2588 0.753441
R32541 DVSS.n5220 DVSS.n5219 0.753441
R32542 DVSS.n5211 DVSS.n5208 0.753441
R32543 DVSS.n5199 DVSS.n5198 0.753441
R32544 DVSS.n5190 DVSS.n5187 0.753441
R32545 DVSS.n5685 DVSS.n5684 0.753441
R32546 DVSS.n5676 DVSS.n5673 0.753441
R32547 DVSS.n5664 DVSS.n5663 0.753441
R32548 DVSS.n5655 DVSS.n5652 0.753441
R32549 DVSS.n155 DVSS.n154 0.753441
R32550 DVSS.n146 DVSS.n143 0.753441
R32551 DVSS.n134 DVSS.n133 0.753441
R32552 DVSS.n125 DVSS.n122 0.753441
R32553 DVSS.n620 DVSS.n619 0.753441
R32554 DVSS.n611 DVSS.n608 0.753441
R32555 DVSS.n599 DVSS.n598 0.753441
R32556 DVSS.n590 DVSS.n587 0.753441
R32557 DVSS.n1141 DVSS.n1140 0.747945
R32558 DVSS.n1875 DVSS.n1874 0.747945
R32559 DVSS.n6671 DVSS.n6670 0.747945
R32560 DVSS.n4948 DVSS 0.681041
R32561 DVSS.n3353 DVSS 0.681041
R32562 DVSS.n6416 DVSS 0.681041
R32563 DVSS.n1735 DVSS 0.681041
R32564 DVSS.n3926 DVSS.n3924 0.649233
R32565 DVSS.n4391 DVSS.n4389 0.649233
R32566 DVSS.n2330 DVSS.n2328 0.649233
R32567 DVSS.n2795 DVSS.n2793 0.649233
R32568 DVSS.n5394 DVSS.n5392 0.649233
R32569 DVSS.n5859 DVSS.n5857 0.649233
R32570 DVSS.n329 DVSS.n327 0.649233
R32571 DVSS.n794 DVSS.n792 0.649233
R32572 DVSS.n3918 DVSS.n3776 0.606816
R32573 DVSS.n4383 DVSS.n4241 0.606816
R32574 DVSS.n2322 DVSS.n2180 0.606816
R32575 DVSS.n2787 DVSS.n2645 0.606816
R32576 DVSS.n5386 DVSS.n5244 0.606816
R32577 DVSS.n5851 DVSS.n5709 0.606816
R32578 DVSS.n321 DVSS.n179 0.606816
R32579 DVSS.n786 DVSS.n644 0.606816
R32580 DVSS DVSS.n1129 0.574303
R32581 DVSS.n3951 DVSS.n3950 0.563137
R32582 DVSS.n4416 DVSS.n4415 0.563137
R32583 DVSS.n2355 DVSS.n2354 0.563137
R32584 DVSS.n2820 DVSS.n2819 0.563137
R32585 DVSS.n5419 DVSS.n5418 0.563137
R32586 DVSS.n5884 DVSS.n5883 0.563137
R32587 DVSS.n354 DVSS.n353 0.563137
R32588 DVSS.n819 DVSS.n818 0.563137
R32589 DVSS.n3929 DVSS.n3927 0.549428
R32590 DVSS.n4394 DVSS.n4392 0.549428
R32591 DVSS.n2333 DVSS.n2331 0.549428
R32592 DVSS.n2798 DVSS.n2796 0.549428
R32593 DVSS.n5397 DVSS.n5395 0.549428
R32594 DVSS.n5862 DVSS.n5860 0.549428
R32595 DVSS.n332 DVSS.n330 0.549428
R32596 DVSS.n797 DVSS.n795 0.549428
R32597 DVSS.n3843 DVSS.n3842 0.539447
R32598 DVSS.n4308 DVSS.n4307 0.539447
R32599 DVSS.n2247 DVSS.n2246 0.539447
R32600 DVSS.n2712 DVSS.n2711 0.539447
R32601 DVSS.n5311 DVSS.n5310 0.539447
R32602 DVSS.n5776 DVSS.n5775 0.539447
R32603 DVSS.n246 DVSS.n245 0.539447
R32604 DVSS.n711 DVSS.n710 0.539447
R32605 DVSS.n6878 DVSS.n6877 0.537004
R32606 DVSS.n6722 DVSS.n3482 0.534792
R32607 DVSS.n1223 DVSS.n1222 0.526461
R32608 DVSS.n1115 DVSS.n1114 0.526088
R32609 DVSS.n1734 DVSS.n1732 0.509446
R32610 DVSS.n4947 DVSS.n4945 0.507079
R32611 DVSS.n6415 DVSS.n6413 0.507079
R32612 DVSS.n3352 DVSS.n3350 0.507079
R32613 DVSS.n1747 DVSS.n1746 0.502212
R32614 DVSS.n4959 DVSS.n4958 0.502212
R32615 DVSS.n3364 DVSS.n3363 0.502212
R32616 DVSS.n6427 DVSS.n6426 0.502212
R32617 DVSS.n3930 DVSS.n3772 0.449623
R32618 DVSS.n4395 DVSS.n4237 0.449623
R32619 DVSS.n2334 DVSS.n2176 0.449623
R32620 DVSS.n2799 DVSS.n2641 0.449623
R32621 DVSS.n5398 DVSS.n5240 0.449623
R32622 DVSS.n5863 DVSS.n5705 0.449623
R32623 DVSS.n333 DVSS.n175 0.449623
R32624 DVSS.n798 DVSS.n640 0.449623
R32625 DVSS.n1525 DVSS.n1517 0.376971
R32626 DVSS.n1536 DVSS.n1528 0.376971
R32627 DVSS.n4738 DVSS.n4730 0.376971
R32628 DVSS.n4749 DVSS.n4741 0.376971
R32629 DVSS.n6206 DVSS.n6198 0.376971
R32630 DVSS.n6217 DVSS.n6209 0.376971
R32631 DVSS.n3142 DVSS.n3134 0.376971
R32632 DVSS.n3153 DVSS.n3145 0.376971
R32633 DVSS.n3934 DVSS.n3933 0.349818
R32634 DVSS.n3779 DVSS.n3778 0.349818
R32635 DVSS.n4399 DVSS.n4398 0.349818
R32636 DVSS.n4244 DVSS.n4243 0.349818
R32637 DVSS.n2338 DVSS.n2337 0.349818
R32638 DVSS.n2183 DVSS.n2182 0.349818
R32639 DVSS.n2803 DVSS.n2802 0.349818
R32640 DVSS.n2648 DVSS.n2647 0.349818
R32641 DVSS.n5402 DVSS.n5401 0.349818
R32642 DVSS.n5247 DVSS.n5246 0.349818
R32643 DVSS.n5867 DVSS.n5866 0.349818
R32644 DVSS.n5712 DVSS.n5711 0.349818
R32645 DVSS.n337 DVSS.n336 0.349818
R32646 DVSS.n182 DVSS.n181 0.349818
R32647 DVSS.n802 DVSS.n801 0.349818
R32648 DVSS.n647 DVSS.n646 0.349818
R32649 DVSS.n3943 DVSS.n3755 0.337926
R32650 DVSS.n3945 DVSS.n3734 0.337926
R32651 DVSS.n4408 DVSS.n4220 0.337926
R32652 DVSS.n4410 DVSS.n4199 0.337926
R32653 DVSS.n2347 DVSS.n2159 0.337926
R32654 DVSS.n2349 DVSS.n2138 0.337926
R32655 DVSS.n2812 DVSS.n2624 0.337926
R32656 DVSS.n2814 DVSS.n2603 0.337926
R32657 DVSS.n5411 DVSS.n5223 0.337926
R32658 DVSS.n5413 DVSS.n5202 0.337926
R32659 DVSS.n5876 DVSS.n5688 0.337926
R32660 DVSS.n5878 DVSS.n5667 0.337926
R32661 DVSS.n346 DVSS.n158 0.337926
R32662 DVSS.n348 DVSS.n137 0.337926
R32663 DVSS.n811 DVSS.n623 0.337926
R32664 DVSS.n813 DVSS.n602 0.337926
R32665 DVSS.n6879 DVSS.n6878 0.33789
R32666 DVSS.n3975 DVSS.n3650 0.328705
R32667 DVSS.n4440 DVSS.n4115 0.328705
R32668 DVSS.n2379 DVSS.n2054 0.328705
R32669 DVSS.n2844 DVSS.n2519 0.328705
R32670 DVSS.n5443 DVSS.n5118 0.328705
R32671 DVSS.n5908 DVSS.n5583 0.328705
R32672 DVSS.n378 DVSS.n53 0.328705
R32673 DVSS.n843 DVSS.n518 0.328705
R32674 DVSS.n4951 DVSS.n4950 0.298465
R32675 DVSS.n3356 DVSS.n3355 0.298465
R32676 DVSS.n6419 DVSS.n6418 0.298465
R32677 DVSS.n1738 DVSS.n1737 0.298465
R32678 DVSS.n4950 DVSS 0.285841
R32679 DVSS.n3355 DVSS 0.285841
R32680 DVSS.n6418 DVSS 0.285841
R32681 DVSS.n1737 DVSS 0.285841
R32682 DVSS.n4022 DVSS.n3634 0.281819
R32683 DVSS.n4487 DVSS.n4099 0.281819
R32684 DVSS.n2426 DVSS.n2038 0.281819
R32685 DVSS.n2891 DVSS.n2503 0.281819
R32686 DVSS.n5490 DVSS.n5102 0.281819
R32687 DVSS.n5955 DVSS.n5567 0.281819
R32688 DVSS.n425 DVSS.n37 0.281819
R32689 DVSS.n890 DVSS.n502 0.281819
R32690 DVSS.n3770 DVSS.n3769 0.250013
R32691 DVSS.n4235 DVSS.n4234 0.250013
R32692 DVSS.n2174 DVSS.n2173 0.250013
R32693 DVSS.n2639 DVSS.n2638 0.250013
R32694 DVSS.n5238 DVSS.n5237 0.250013
R32695 DVSS.n5703 DVSS.n5702 0.250013
R32696 DVSS.n173 DVSS.n172 0.250013
R32697 DVSS.n638 DVSS.n637 0.250013
R32698 DVSS.n3677 DVSS.n3649 0.234932
R32699 DVSS.n4142 DVSS.n4114 0.234932
R32700 DVSS.n2081 DVSS.n2053 0.234932
R32701 DVSS.n2546 DVSS.n2518 0.234932
R32702 DVSS.n5145 DVSS.n5117 0.234932
R32703 DVSS.n5610 DVSS.n5582 0.234932
R32704 DVSS.n80 DVSS.n52 0.234932
R32705 DVSS.n545 DVSS.n517 0.234932
R32706 DVSS.n1233 DVSS 0.212305
R32707 DVSS.n1121 DVSS 0.212135
R32708 DVSS DVSS.n1338 0.199538
R32709 DVSS.n3943 DVSS.n3942 0.198603
R32710 DVSS.n4408 DVSS.n4407 0.198603
R32711 DVSS.n2347 DVSS.n2346 0.198603
R32712 DVSS.n2812 DVSS.n2811 0.198603
R32713 DVSS.n5411 DVSS.n5410 0.198603
R32714 DVSS.n5876 DVSS.n5875 0.198603
R32715 DVSS.n346 DVSS.n345 0.198603
R32716 DVSS.n811 DVSS.n810 0.198603
R32717 DVSS.n3945 DVSS.n3944 0.196998
R32718 DVSS.n4410 DVSS.n4409 0.196998
R32719 DVSS.n2349 DVSS.n2348 0.196998
R32720 DVSS.n2814 DVSS.n2813 0.196998
R32721 DVSS.n5413 DVSS.n5412 0.196998
R32722 DVSS.n5878 DVSS.n5877 0.196998
R32723 DVSS.n348 DVSS.n347 0.196998
R32724 DVSS.n813 DVSS.n812 0.196998
R32725 DVSS DVSS.n6885 0.170371
R32726 DVSS.n1117 DVSS.n1095 0.156029
R32727 DVSS.n1117 DVSS.n1101 0.156029
R32728 DVSS.n1117 DVSS.n1107 0.156029
R32729 DVSS.n1117 DVSS.n1060 0.153643
R32730 DVSS.n1321 DVSS.n1320 0.153643
R32731 DVSS.n6700 DVSS.n6699 0.151309
R32732 DVSS.n1335 DVSS.n1156 0.151309
R32733 DVSS.n1124 DVSS.n1123 0.151309
R32734 DVSS.n1227 DVSS.n1226 0.151309
R32735 DVSS.n6735 DVSS.n6734 0.151294
R32736 DVSS.n6525 DVSS.n6523 0.151294
R32737 DVSS.n1124 DVSS.n1037 0.151294
R32738 DVSS.n1124 DVSS.n1030 0.151294
R32739 DVSS.n1124 DVSS.n1046 0.151294
R32740 DVSS.n1124 DVSS.n1018 0.151294
R32741 DVSS.n1125 DVSS.n1124 0.151294
R32742 DVSS.n1124 DVSS.n979 0.151294
R32743 DVSS.n1124 DVSS.n986 0.151294
R32744 DVSS.n1124 DVSS.n993 0.151294
R32745 DVSS.n1124 DVSS.n1000 0.151294
R32746 DVSS.n1124 DVSS.n1011 0.151294
R32747 DVSS.n1118 DVSS.n1117 0.151294
R32748 DVSS.n1117 DVSS.n1073 0.151294
R32749 DVSS.n1117 DVSS.n1083 0.151294
R32750 DVSS.n1117 DVSS.n1090 0.151294
R32751 DVSS.n1227 DVSS.n1213 0.151294
R32752 DVSS.n1227 DVSS.n1206 0.151294
R32753 DVSS.n1227 DVSS.n1197 0.151294
R32754 DVSS.n1227 DVSS.n1189 0.151294
R32755 DVSS.n1227 DVSS.n1179 0.151294
R32756 DVSS.n1322 DVSS.n1321 0.151294
R32757 DVSS.n1156 DVSS.n1155 0.151294
R32758 DVSS.n1156 DVSS.n1147 0.151294
R32759 DVSS.n1156 DVSS.n1135 0.151294
R32760 DVSS.n0 DVSS 0.15024
R32761 DVSS.n3940 DVSS.n3758 0.150208
R32762 DVSS.n4405 DVSS.n4223 0.150208
R32763 DVSS.n2344 DVSS.n2162 0.150208
R32764 DVSS.n2809 DVSS.n2627 0.150208
R32765 DVSS.n5408 DVSS.n5226 0.150208
R32766 DVSS.n5873 DVSS.n5691 0.150208
R32767 DVSS.n343 DVSS.n161 0.150208
R32768 DVSS.n808 DVSS.n626 0.150208
R32769 DVSS.n4074 DVSS.n3609 0.142979
R32770 DVSS.n2478 DVSS.n2013 0.142979
R32771 DVSS.n5542 DVSS.n5077 0.142979
R32772 DVSS.n477 DVSS.n12 0.142979
R32773 DVSS.n3995 DVSS.n3636 0.141159
R32774 DVSS.n4460 DVSS.n4101 0.141159
R32775 DVSS.n2399 DVSS.n2040 0.141159
R32776 DVSS.n2864 DVSS.n2505 0.141159
R32777 DVSS.n5463 DVSS.n5104 0.141159
R32778 DVSS.n5928 DVSS.n5569 0.141159
R32779 DVSS.n398 DVSS.n39 0.141159
R32780 DVSS.n863 DVSS.n504 0.141159
R32781 DVSS.n3606 DVSS 0.13698
R32782 DVSS.n6759 DVSS 0.13698
R32783 DVSS DVSS.n6707 0.13045
R32784 DVSS DVSS.n6742 0.13045
R32785 DVSS.n4949 DVSS.n4948 0.128407
R32786 DVSS.n3354 DVSS.n3353 0.128407
R32787 DVSS.n6417 DVSS.n6416 0.128407
R32788 DVSS.n1736 DVSS.n1735 0.128407
R32789 DVSS.n1734 DVSS.n1733 0.1255
R32790 DVSS.n4947 DVSS.n4946 0.11623
R32791 DVSS.n6415 DVSS.n6414 0.11623
R32792 DVSS.n3352 DVSS.n3351 0.11623
R32793 DVSS.n6885 DVSS.n6884 0.115146
R32794 DVSS.n1128 DVSS.n0 0.110861
R32795 DVSS.n4068 DVSS.n3611 0.0942729
R32796 DVSS.n4532 DVSS.n4076 0.0942729
R32797 DVSS.n2472 DVSS.n2015 0.0942729
R32798 DVSS.n2936 DVSS.n2480 0.0942729
R32799 DVSS.n5536 DVSS.n5079 0.0942729
R32800 DVSS.n6000 DVSS.n5544 0.0942729
R32801 DVSS.n471 DVSS.n14 0.0942729
R32802 DVSS.n935 DVSS.n479 0.0942729
R32803 DVSS.n3942 DVSS.n3756 0.0932835
R32804 DVSS.n3773 DVSS.n3756 0.0932835
R32805 DVSS.n3932 DVSS.n3773 0.0932835
R32806 DVSS.n3932 DVSS.n3931 0.0932835
R32807 DVSS.n3931 DVSS.n3774 0.0932835
R32808 DVSS.n3923 DVSS.n3774 0.0932835
R32809 DVSS.n3923 DVSS.n3922 0.0932835
R32810 DVSS.n3841 DVSS.n3735 0.0932835
R32811 DVSS.n3841 DVSS.n3840 0.0932835
R32812 DVSS.n3840 DVSS.n3801 0.0932835
R32813 DVSS.n3816 DVSS.n3801 0.0932835
R32814 DVSS.n3831 DVSS.n3816 0.0932835
R32815 DVSS.n3831 DVSS.n3830 0.0932835
R32816 DVSS.n3830 DVSS.n3817 0.0932835
R32817 DVSS.n4407 DVSS.n4221 0.0932835
R32818 DVSS.n4238 DVSS.n4221 0.0932835
R32819 DVSS.n4397 DVSS.n4238 0.0932835
R32820 DVSS.n4397 DVSS.n4396 0.0932835
R32821 DVSS.n4396 DVSS.n4239 0.0932835
R32822 DVSS.n4388 DVSS.n4239 0.0932835
R32823 DVSS.n4388 DVSS.n4387 0.0932835
R32824 DVSS.n4306 DVSS.n4200 0.0932835
R32825 DVSS.n4306 DVSS.n4305 0.0932835
R32826 DVSS.n4305 DVSS.n4266 0.0932835
R32827 DVSS.n4281 DVSS.n4266 0.0932835
R32828 DVSS.n4296 DVSS.n4281 0.0932835
R32829 DVSS.n4296 DVSS.n4295 0.0932835
R32830 DVSS.n4295 DVSS.n4282 0.0932835
R32831 DVSS.n2346 DVSS.n2160 0.0932835
R32832 DVSS.n2177 DVSS.n2160 0.0932835
R32833 DVSS.n2336 DVSS.n2177 0.0932835
R32834 DVSS.n2336 DVSS.n2335 0.0932835
R32835 DVSS.n2335 DVSS.n2178 0.0932835
R32836 DVSS.n2327 DVSS.n2178 0.0932835
R32837 DVSS.n2327 DVSS.n2326 0.0932835
R32838 DVSS.n2245 DVSS.n2139 0.0932835
R32839 DVSS.n2245 DVSS.n2244 0.0932835
R32840 DVSS.n2244 DVSS.n2205 0.0932835
R32841 DVSS.n2220 DVSS.n2205 0.0932835
R32842 DVSS.n2235 DVSS.n2220 0.0932835
R32843 DVSS.n2235 DVSS.n2234 0.0932835
R32844 DVSS.n2234 DVSS.n2221 0.0932835
R32845 DVSS.n2811 DVSS.n2625 0.0932835
R32846 DVSS.n2642 DVSS.n2625 0.0932835
R32847 DVSS.n2801 DVSS.n2642 0.0932835
R32848 DVSS.n2801 DVSS.n2800 0.0932835
R32849 DVSS.n2800 DVSS.n2643 0.0932835
R32850 DVSS.n2792 DVSS.n2643 0.0932835
R32851 DVSS.n2792 DVSS.n2791 0.0932835
R32852 DVSS.n2710 DVSS.n2604 0.0932835
R32853 DVSS.n2710 DVSS.n2709 0.0932835
R32854 DVSS.n2709 DVSS.n2670 0.0932835
R32855 DVSS.n2685 DVSS.n2670 0.0932835
R32856 DVSS.n2700 DVSS.n2685 0.0932835
R32857 DVSS.n2700 DVSS.n2699 0.0932835
R32858 DVSS.n2699 DVSS.n2686 0.0932835
R32859 DVSS.n5410 DVSS.n5224 0.0932835
R32860 DVSS.n5241 DVSS.n5224 0.0932835
R32861 DVSS.n5400 DVSS.n5241 0.0932835
R32862 DVSS.n5400 DVSS.n5399 0.0932835
R32863 DVSS.n5399 DVSS.n5242 0.0932835
R32864 DVSS.n5391 DVSS.n5242 0.0932835
R32865 DVSS.n5391 DVSS.n5390 0.0932835
R32866 DVSS.n5309 DVSS.n5203 0.0932835
R32867 DVSS.n5309 DVSS.n5308 0.0932835
R32868 DVSS.n5308 DVSS.n5269 0.0932835
R32869 DVSS.n5284 DVSS.n5269 0.0932835
R32870 DVSS.n5299 DVSS.n5284 0.0932835
R32871 DVSS.n5299 DVSS.n5298 0.0932835
R32872 DVSS.n5298 DVSS.n5285 0.0932835
R32873 DVSS.n5875 DVSS.n5689 0.0932835
R32874 DVSS.n5706 DVSS.n5689 0.0932835
R32875 DVSS.n5865 DVSS.n5706 0.0932835
R32876 DVSS.n5865 DVSS.n5864 0.0932835
R32877 DVSS.n5864 DVSS.n5707 0.0932835
R32878 DVSS.n5856 DVSS.n5707 0.0932835
R32879 DVSS.n5856 DVSS.n5855 0.0932835
R32880 DVSS.n5774 DVSS.n5668 0.0932835
R32881 DVSS.n5774 DVSS.n5773 0.0932835
R32882 DVSS.n5773 DVSS.n5734 0.0932835
R32883 DVSS.n5749 DVSS.n5734 0.0932835
R32884 DVSS.n5764 DVSS.n5749 0.0932835
R32885 DVSS.n5764 DVSS.n5763 0.0932835
R32886 DVSS.n5763 DVSS.n5750 0.0932835
R32887 DVSS.n345 DVSS.n159 0.0932835
R32888 DVSS.n176 DVSS.n159 0.0932835
R32889 DVSS.n335 DVSS.n176 0.0932835
R32890 DVSS.n335 DVSS.n334 0.0932835
R32891 DVSS.n334 DVSS.n177 0.0932835
R32892 DVSS.n326 DVSS.n177 0.0932835
R32893 DVSS.n326 DVSS.n325 0.0932835
R32894 DVSS.n244 DVSS.n138 0.0932835
R32895 DVSS.n244 DVSS.n243 0.0932835
R32896 DVSS.n243 DVSS.n204 0.0932835
R32897 DVSS.n219 DVSS.n204 0.0932835
R32898 DVSS.n234 DVSS.n219 0.0932835
R32899 DVSS.n234 DVSS.n233 0.0932835
R32900 DVSS.n233 DVSS.n220 0.0932835
R32901 DVSS.n810 DVSS.n624 0.0932835
R32902 DVSS.n641 DVSS.n624 0.0932835
R32903 DVSS.n800 DVSS.n641 0.0932835
R32904 DVSS.n800 DVSS.n799 0.0932835
R32905 DVSS.n799 DVSS.n642 0.0932835
R32906 DVSS.n791 DVSS.n642 0.0932835
R32907 DVSS.n791 DVSS.n790 0.0932835
R32908 DVSS.n709 DVSS.n603 0.0932835
R32909 DVSS.n709 DVSS.n708 0.0932835
R32910 DVSS.n708 DVSS.n669 0.0932835
R32911 DVSS.n684 DVSS.n669 0.0932835
R32912 DVSS.n699 DVSS.n684 0.0932835
R32913 DVSS.n699 DVSS.n698 0.0932835
R32914 DVSS.n698 DVSS.n685 0.0932835
R32915 DVSS.n4074 DVSS.n4073 0.0919929
R32916 DVSS.n2478 DVSS.n2477 0.0919929
R32917 DVSS.n5542 DVSS.n5541 0.0919929
R32918 DVSS.n477 DVSS.n476 0.0919929
R32919 DVSS.n6884 DVSS 0.0919821
R32920 DVSS.n3944 DVSS.n3943 0.0870759
R32921 DVSS.n4409 DVSS.n4408 0.0870759
R32922 DVSS.n2348 DVSS.n2347 0.0870759
R32923 DVSS.n2813 DVSS.n2812 0.0870759
R32924 DVSS.n5412 DVSS.n5411 0.0870759
R32925 DVSS.n5877 DVSS.n5876 0.0870759
R32926 DVSS.n347 DVSS.n346 0.0870759
R32927 DVSS.n812 DVSS.n811 0.0870759
R32928 DVSS.n1907 DVSS 0.0862219
R32929 DVSS.n6641 DVSS 0.0862219
R32930 DVSS.n3509 DVSS 0.0854216
R32931 DVSS.n6855 DVSS 0.0854216
R32932 DVSS.n3742 DVSS.n3741 0.0793691
R32933 DVSS.n3721 DVSS.n3720 0.0793691
R32934 DVSS.n4207 DVSS.n4206 0.0793691
R32935 DVSS.n4186 DVSS.n4185 0.0793691
R32936 DVSS.n2146 DVSS.n2145 0.0793691
R32937 DVSS.n2125 DVSS.n2124 0.0793691
R32938 DVSS.n2611 DVSS.n2610 0.0793691
R32939 DVSS.n2590 DVSS.n2589 0.0793691
R32940 DVSS.n5210 DVSS.n5209 0.0793691
R32941 DVSS.n5189 DVSS.n5188 0.0793691
R32942 DVSS.n5675 DVSS.n5674 0.0793691
R32943 DVSS.n5654 DVSS.n5653 0.0793691
R32944 DVSS.n145 DVSS.n144 0.0793691
R32945 DVSS.n124 DVSS.n123 0.0793691
R32946 DVSS.n610 DVSS.n609 0.0793691
R32947 DVSS.n589 DVSS.n588 0.0793691
R32948 DVSS.n4616 DVSS.n4612 0.0772544
R32949 DVSS.n4618 DVSS.n4616 0.0772544
R32950 DVSS.n4750 DVSS.n4739 0.0772544
R32951 DVSS.n4866 DVSS.n4862 0.0772544
R32952 DVSS.n4868 DVSS.n4866 0.0772544
R32953 DVSS.n6084 DVSS.n6080 0.0772544
R32954 DVSS.n6086 DVSS.n6084 0.0772544
R32955 DVSS.n6218 DVSS.n6207 0.0772544
R32956 DVSS.n6334 DVSS.n6330 0.0772544
R32957 DVSS.n6336 DVSS.n6334 0.0772544
R32958 DVSS.n3020 DVSS.n3016 0.0772544
R32959 DVSS.n3022 DVSS.n3020 0.0772544
R32960 DVSS.n3154 DVSS.n3143 0.0772544
R32961 DVSS.n3270 DVSS.n3266 0.0772544
R32962 DVSS.n3272 DVSS.n3270 0.0772544
R32963 DVSS.n1403 DVSS.n1399 0.0772544
R32964 DVSS.n1405 DVSS.n1403 0.0772544
R32965 DVSS.n1537 DVSS.n1526 0.0772544
R32966 DVSS.n1653 DVSS.n1649 0.0772544
R32967 DVSS.n1655 DVSS.n1653 0.0772544
R32968 DVSS.n3778 DVSS.n3775 0.0753538
R32969 DVSS.n4243 DVSS.n4240 0.0753538
R32970 DVSS.n2182 DVSS.n2179 0.0753538
R32971 DVSS.n2647 DVSS.n2644 0.0753538
R32972 DVSS.n5246 DVSS.n5243 0.0753538
R32973 DVSS.n5711 DVSS.n5708 0.0753538
R32974 DVSS.n181 DVSS.n178 0.0753538
R32975 DVSS.n646 DVSS.n643 0.0753538
R32976 DVSS.n4945 DVSS.n4914 0.067386
R32977 DVSS.n6413 DVSS.n6382 0.067386
R32978 DVSS.n3350 DVSS.n3318 0.067386
R32979 DVSS.n1732 DVSS.n1701 0.067386
R32980 DVSS.n3971 DVSS.n3970 0.0637979
R32981 DVSS.n3978 DVSS.n3971 0.0637979
R32982 DVSS.n4026 DVSS.n4025 0.0637979
R32983 DVSS.n4025 DVSS.n4024 0.0637979
R32984 DVSS.n4436 DVSS.n4435 0.0637979
R32985 DVSS.n4443 DVSS.n4436 0.0637979
R32986 DVSS.n4491 DVSS.n4490 0.0637979
R32987 DVSS.n4490 DVSS.n4489 0.0637979
R32988 DVSS.n2375 DVSS.n2374 0.0637979
R32989 DVSS.n2382 DVSS.n2375 0.0637979
R32990 DVSS.n2430 DVSS.n2429 0.0637979
R32991 DVSS.n2429 DVSS.n2428 0.0637979
R32992 DVSS.n2840 DVSS.n2839 0.0637979
R32993 DVSS.n2847 DVSS.n2840 0.0637979
R32994 DVSS.n2895 DVSS.n2894 0.0637979
R32995 DVSS.n2894 DVSS.n2893 0.0637979
R32996 DVSS.n5439 DVSS.n5438 0.0637979
R32997 DVSS.n5446 DVSS.n5439 0.0637979
R32998 DVSS.n5494 DVSS.n5493 0.0637979
R32999 DVSS.n5493 DVSS.n5492 0.0637979
R33000 DVSS.n5904 DVSS.n5903 0.0637979
R33001 DVSS.n5911 DVSS.n5904 0.0637979
R33002 DVSS.n5959 DVSS.n5958 0.0637979
R33003 DVSS.n5958 DVSS.n5957 0.0637979
R33004 DVSS.n374 DVSS.n373 0.0637979
R33005 DVSS.n381 DVSS.n374 0.0637979
R33006 DVSS.n429 DVSS.n428 0.0637979
R33007 DVSS.n428 DVSS.n427 0.0637979
R33008 DVSS.n839 DVSS.n838 0.0637979
R33009 DVSS.n846 DVSS.n839 0.0637979
R33010 DVSS.n894 DVSS.n893 0.0637979
R33011 DVSS.n893 DVSS.n892 0.0637979
R33012 DVSS.n1911 DVSS.n1907 0.0617245
R33013 DVSS.n1915 DVSS.n1911 0.0617245
R33014 DVSS.n1919 DVSS.n1915 0.0617245
R33015 DVSS.n1935 DVSS.n1931 0.0617245
R33016 DVSS.n1952 DVSS.n1948 0.0617245
R33017 DVSS.n1968 DVSS.n1964 0.0617245
R33018 DVSS.n1972 DVSS.n1968 0.0617245
R33019 DVSS.n1990 DVSS.n1986 0.0617245
R33020 DVSS.n1991 DVSS.n1990 0.0617245
R33021 DVSS.n2002 DVSS.n1998 0.0617245
R33022 DVSS.n6641 DVSS.n6640 0.0617245
R33023 DVSS.n6640 DVSS.n6636 0.0617245
R33024 DVSS.n6636 DVSS.n6632 0.0617245
R33025 DVSS.n6622 DVSS.n6618 0.0617245
R33026 DVSS.n6605 DVSS.n6601 0.0617245
R33027 DVSS.n6589 DVSS.n6585 0.0617245
R33028 DVSS.n6585 DVSS.n6581 0.0617245
R33029 DVSS.n6567 DVSS.n6563 0.0617245
R33030 DVSS.n6563 DVSS.n6559 0.0617245
R33031 DVSS.n6554 DVSS.n6553 0.0617245
R33032 DVSS.n3518 DVSS.n3514 0.0617245
R33033 DVSS.n3522 DVSS.n3518 0.0617245
R33034 DVSS.n3538 DVSS.n3534 0.0617245
R33035 DVSS.n3555 DVSS.n3551 0.0617245
R33036 DVSS.n3571 DVSS.n3567 0.0617245
R33037 DVSS.n3575 DVSS.n3571 0.0617245
R33038 DVSS.n3593 DVSS.n3589 0.0617245
R33039 DVSS.n3600 DVSS.n3593 0.0617245
R33040 DVSS.n3605 DVSS.n3601 0.0617245
R33041 DVSS.n6853 DVSS.n6849 0.0617245
R33042 DVSS.n6849 DVSS.n6845 0.0617245
R33043 DVSS.n6833 DVSS.n6829 0.0617245
R33044 DVSS.n6816 DVSS.n6812 0.0617245
R33045 DVSS.n6801 DVSS.n6797 0.0617245
R33046 DVSS.n6797 DVSS.n6793 0.0617245
R33047 DVSS.n6779 DVSS.n6775 0.0617245
R33048 DVSS.n6775 DVSS.n6771 0.0617245
R33049 DVSS.n6764 DVSS.n6763 0.0617245
R33050 DVSS.n1762 DVSS.n1758 0.0611061
R33051 DVSS.n1766 DVSS.n1762 0.0611061
R33052 DVSS.n1770 DVSS.n1766 0.0611061
R33053 DVSS.n1774 DVSS.n1770 0.0611061
R33054 DVSS.n1778 DVSS.n1774 0.0611061
R33055 DVSS.n1782 DVSS.n1778 0.0611061
R33056 DVSS.n1787 DVSS.n1782 0.0611061
R33057 DVSS.n1803 DVSS.n1799 0.0611061
R33058 DVSS.n1820 DVSS.n1816 0.0611061
R33059 DVSS.n1824 DVSS.n1820 0.0611061
R33060 DVSS.n1834 DVSS.n1830 0.0611061
R33061 DVSS.n4974 DVSS.n4970 0.0611061
R33062 DVSS.n4978 DVSS.n4974 0.0611061
R33063 DVSS.n4982 DVSS.n4978 0.0611061
R33064 DVSS.n4986 DVSS.n4982 0.0611061
R33065 DVSS.n4990 DVSS.n4986 0.0611061
R33066 DVSS.n4994 DVSS.n4990 0.0611061
R33067 DVSS.n4999 DVSS.n4994 0.0611061
R33068 DVSS.n5015 DVSS.n5011 0.0611061
R33069 DVSS.n5032 DVSS.n5028 0.0611061
R33070 DVSS.n5036 DVSS.n5032 0.0611061
R33071 DVSS.n5046 DVSS.n5042 0.0611061
R33072 DVSS.n3379 DVSS.n3375 0.0611061
R33073 DVSS.n3383 DVSS.n3379 0.0611061
R33074 DVSS.n3387 DVSS.n3383 0.0611061
R33075 DVSS.n3391 DVSS.n3387 0.0611061
R33076 DVSS.n3395 DVSS.n3391 0.0611061
R33077 DVSS.n3399 DVSS.n3395 0.0611061
R33078 DVSS.n3404 DVSS.n3399 0.0611061
R33079 DVSS.n3420 DVSS.n3416 0.0611061
R33080 DVSS.n3437 DVSS.n3433 0.0611061
R33081 DVSS.n3441 DVSS.n3437 0.0611061
R33082 DVSS.n3451 DVSS.n3447 0.0611061
R33083 DVSS.n6442 DVSS.n6438 0.0611061
R33084 DVSS.n6446 DVSS.n6442 0.0611061
R33085 DVSS.n6450 DVSS.n6446 0.0611061
R33086 DVSS.n6454 DVSS.n6450 0.0611061
R33087 DVSS.n6458 DVSS.n6454 0.0611061
R33088 DVSS.n6462 DVSS.n6458 0.0611061
R33089 DVSS.n6467 DVSS.n6462 0.0611061
R33090 DVSS.n6483 DVSS.n6479 0.0611061
R33091 DVSS.n6500 DVSS.n6496 0.0611061
R33092 DVSS.n6505 DVSS.n6500 0.0611061
R33093 DVSS.n6513 DVSS.n6510 0.0611061
R33094 DVSS.n1954 DVSS.n1952 0.0610867
R33095 DVSS.n6601 DVSS.n6596 0.0610867
R33096 DVSS.n3557 DVSS.n3555 0.0610867
R33097 DVSS.n6812 DVSS.n6808 0.0610867
R33098 DVSS.n2004 DVSS.n2002 0.060449
R33099 DVSS.n6553 DVSS.n6546 0.060449
R33100 DVSS.n1836 DVSS.n1834 0.0592121
R33101 DVSS.n5048 DVSS.n5046 0.0592121
R33102 DVSS.n3453 DVSS.n3451 0.0592121
R33103 DVSS.n6515 DVSS.n6513 0.0592121
R33104 DVSS.n4590 DVSS.n4579 0.058614
R33105 DVSS.n4608 DVSS.n4594 0.058614
R33106 DVSS.n4636 DVSS.n4634 0.058614
R33107 DVSS.n4651 DVSS.n4649 0.058614
R33108 DVSS.n4666 DVSS.n4664 0.058614
R33109 DVSS.n4681 DVSS.n4679 0.058614
R33110 DVSS.n4696 DVSS.n4694 0.058614
R33111 DVSS.n4711 DVSS.n4709 0.058614
R33112 DVSS.n4726 DVSS.n4724 0.058614
R33113 DVSS.n4765 DVSS.n4754 0.058614
R33114 DVSS.n4780 DVSS.n4769 0.058614
R33115 DVSS.n4795 DVSS.n4784 0.058614
R33116 DVSS.n4810 DVSS.n4799 0.058614
R33117 DVSS.n4825 DVSS.n4814 0.058614
R33118 DVSS.n4840 DVSS.n4829 0.058614
R33119 DVSS.n4858 DVSS.n4844 0.058614
R33120 DVSS.n4886 DVSS.n4884 0.058614
R33121 DVSS.n4901 DVSS.n4899 0.058614
R33122 DVSS.n6058 DVSS.n6047 0.058614
R33123 DVSS.n6076 DVSS.n6062 0.058614
R33124 DVSS.n6104 DVSS.n6102 0.058614
R33125 DVSS.n6119 DVSS.n6117 0.058614
R33126 DVSS.n6134 DVSS.n6132 0.058614
R33127 DVSS.n6149 DVSS.n6147 0.058614
R33128 DVSS.n6164 DVSS.n6162 0.058614
R33129 DVSS.n6179 DVSS.n6177 0.058614
R33130 DVSS.n6194 DVSS.n6192 0.058614
R33131 DVSS.n6233 DVSS.n6222 0.058614
R33132 DVSS.n6248 DVSS.n6237 0.058614
R33133 DVSS.n6263 DVSS.n6252 0.058614
R33134 DVSS.n6278 DVSS.n6267 0.058614
R33135 DVSS.n6293 DVSS.n6282 0.058614
R33136 DVSS.n6308 DVSS.n6297 0.058614
R33137 DVSS.n6326 DVSS.n6312 0.058614
R33138 DVSS.n6354 DVSS.n6352 0.058614
R33139 DVSS.n6369 DVSS.n6367 0.058614
R33140 DVSS.n2994 DVSS.n2983 0.058614
R33141 DVSS.n3012 DVSS.n2998 0.058614
R33142 DVSS.n3040 DVSS.n3038 0.058614
R33143 DVSS.n3055 DVSS.n3053 0.058614
R33144 DVSS.n3070 DVSS.n3068 0.058614
R33145 DVSS.n3085 DVSS.n3083 0.058614
R33146 DVSS.n3100 DVSS.n3098 0.058614
R33147 DVSS.n3115 DVSS.n3113 0.058614
R33148 DVSS.n3130 DVSS.n3128 0.058614
R33149 DVSS.n3169 DVSS.n3158 0.058614
R33150 DVSS.n3184 DVSS.n3173 0.058614
R33151 DVSS.n3199 DVSS.n3188 0.058614
R33152 DVSS.n3214 DVSS.n3203 0.058614
R33153 DVSS.n3229 DVSS.n3218 0.058614
R33154 DVSS.n3244 DVSS.n3233 0.058614
R33155 DVSS.n3262 DVSS.n3248 0.058614
R33156 DVSS.n3290 DVSS.n3288 0.058614
R33157 DVSS.n3305 DVSS.n3303 0.058614
R33158 DVSS.n1377 DVSS.n1366 0.058614
R33159 DVSS.n1395 DVSS.n1381 0.058614
R33160 DVSS.n1423 DVSS.n1421 0.058614
R33161 DVSS.n1438 DVSS.n1436 0.058614
R33162 DVSS.n1453 DVSS.n1451 0.058614
R33163 DVSS.n1468 DVSS.n1466 0.058614
R33164 DVSS.n1483 DVSS.n1481 0.058614
R33165 DVSS.n1498 DVSS.n1496 0.058614
R33166 DVSS.n1513 DVSS.n1511 0.058614
R33167 DVSS.n1552 DVSS.n1541 0.058614
R33168 DVSS.n1567 DVSS.n1556 0.058614
R33169 DVSS.n1582 DVSS.n1571 0.058614
R33170 DVSS.n1597 DVSS.n1586 0.058614
R33171 DVSS.n1612 DVSS.n1601 0.058614
R33172 DVSS.n1627 DVSS.n1616 0.058614
R33173 DVSS.n1645 DVSS.n1631 0.058614
R33174 DVSS.n1673 DVSS.n1671 0.058614
R33175 DVSS.n1688 DVSS.n1686 0.058614
R33176 DVSS.n1804 DVSS.n1803 0.0585808
R33177 DVSS.n5016 DVSS.n5015 0.0585808
R33178 DVSS.n3421 DVSS.n3420 0.0585808
R33179 DVSS.n6484 DVSS.n6483 0.0585808
R33180 DVSS.n1758 DVSS.n1754 0.0566869
R33181 DVSS.n4970 DVSS.n4966 0.0566869
R33182 DVSS.n3375 DVSS.n3371 0.0566869
R33183 DVSS.n6438 DVSS.n6434 0.0566869
R33184 DVSS.n3948 DVSS.n3714 0.0547553
R33185 DVSS.n4413 DVSS.n4179 0.0547553
R33186 DVSS.n2352 DVSS.n2118 0.0547553
R33187 DVSS.n2817 DVSS.n2583 0.0547553
R33188 DVSS.n5416 DVSS.n5182 0.0547553
R33189 DVSS.n5881 DVSS.n5647 0.0547553
R33190 DVSS.n351 DVSS.n117 0.0547553
R33191 DVSS.n816 DVSS.n582 0.0547553
R33192 DVSS.n6663 DVSS.n6659 0.0535973
R33193 DVSS.n6685 DVSS.n6681 0.0535973
R33194 DVSS.n1867 DVSS.n1863 0.0535973
R33195 DVSS.n1889 DVSS.n1885 0.0535973
R33196 DVSS.n4073 DVSS.n3610 0.0520957
R33197 DVSS.n2477 DVSS.n2014 0.0520957
R33198 DVSS.n5541 DVSS.n5078 0.0520957
R33199 DVSS.n476 DVSS.n13 0.0520957
R33200 DVSS.n3953 DVSS.n3687 0.0505
R33201 DVSS.n4418 DVSS.n4152 0.0505
R33202 DVSS.n2357 DVSS.n2091 0.0505
R33203 DVSS.n2822 DVSS.n2556 0.0505
R33204 DVSS.n5421 DVSS.n5155 0.0505
R33205 DVSS.n5886 DVSS.n5620 0.0505
R33206 DVSS.n356 DVSS.n90 0.0505
R33207 DVSS.n821 DVSS.n555 0.0505
R33208 DVSS DVSS.n4537 0.0487678
R33209 DVSS DVSS.n2941 0.0487678
R33210 DVSS DVSS.n6005 0.0487678
R33211 DVSS DVSS.n940 0.0487678
R33212 DVSS.n1991 DVSS 0.0476939
R33213 DVSS.n6559 DVSS 0.0476939
R33214 DVSS DVSS.n3600 0.0476939
R33215 DVSS.n6771 DVSS 0.0476939
R33216 DVSS.n1931 DVSS.n1927 0.0470561
R33217 DVSS.n6623 DVSS.n6622 0.0470561
R33218 DVSS.n3534 DVSS.n3530 0.0470561
R33219 DVSS.n6834 DVSS.n6833 0.0470561
R33220 DVSS.n1982 DVSS.n1981 0.0464184
R33221 DVSS.n6572 DVSS.n6568 0.0464184
R33222 DVSS.n3514 DVSS.n3510 0.0464184
R33223 DVSS.n3585 DVSS.n3584 0.0464184
R33224 DVSS.n6854 DVSS.n6853 0.0464184
R33225 DVSS.n6784 DVSS.n6780 0.0464184
R33226 DVSS.n1165 DVSS.n1162 0.0459545
R33227 DVSS.n1237 DVSS.n1233 0.045783
R33228 DVSS.n1241 DVSS.n1237 0.045783
R33229 DVSS.n1246 DVSS.n1241 0.045783
R33230 DVSS.n1250 DVSS.n1246 0.045783
R33231 DVSS.n1254 DVSS.n1250 0.045783
R33232 DVSS.n1258 DVSS.n1254 0.045783
R33233 DVSS.n1276 DVSS.n1272 0.045783
R33234 DVSS.n1279 DVSS.n1276 0.045783
R33235 DVSS.n1292 DVSS.n1288 0.045783
R33236 DVSS.n1307 DVSS.n1304 0.045783
R33237 DVSS.n1325 DVSS.n1318 0.045783
R33238 DVSS.n1329 DVSS.n1325 0.045783
R33239 DVSS.n1339 DVSS.n1329 0.045783
R33240 DVSS.n1939 DVSS.n1935 0.0457806
R33241 DVSS.n1960 DVSS.n1959 0.0457806
R33242 DVSS.n6618 DVSS.n6614 0.0457806
R33243 DVSS.n6594 DVSS.n6590 0.0457806
R33244 DVSS.n3542 DVSS.n3538 0.0457806
R33245 DVSS.n3563 DVSS.n3562 0.0457806
R33246 DVSS.n6829 DVSS.n6825 0.0457806
R33247 DVSS.n6807 DVSS.n6802 0.0457806
R33248 DVSS.n1114 DVSS.n1113 0.0456128
R33249 DVSS.n1113 DVSS.n1112 0.0456128
R33250 DVSS.n1112 DVSS.n1111 0.0456128
R33251 DVSS.n1111 DVSS.n1110 0.0456128
R33252 DVSS.n1110 DVSS.n1109 0.0456128
R33253 DVSS.n1109 DVSS.n1108 0.0456128
R33254 DVSS.n1288 DVSS.n1285 0.0453113
R33255 DVSS.n1788 DVSS.n1787 0.0434293
R33256 DVSS.n1812 DVSS.n1808 0.0434293
R33257 DVSS.n5000 DVSS.n4999 0.0434293
R33258 DVSS.n5024 DVSS.n5020 0.0434293
R33259 DVSS.n3405 DVSS.n3404 0.0434293
R33260 DVSS.n3429 DVSS.n3425 0.0434293
R33261 DVSS.n6468 DVSS.n6467 0.0434293
R33262 DVSS.n6492 DVSS.n6488 0.0434293
R33263 DVSS.n6681 DVSS.n6677 0.0430885
R33264 DVSS.n1885 DVSS.n1881 0.0430885
R33265 DVSS.n1977 DVSS.n1973 0.0425918
R33266 DVSS.n6577 DVSS.n6576 0.0425918
R33267 DVSS.n3580 DVSS.n3576 0.0425918
R33268 DVSS.n6789 DVSS.n6788 0.0425918
R33269 DVSS.n3607 DVSS.n3606 0.0425792
R33270 DVSS.n6759 DVSS.n6758 0.0425792
R33271 DVSS.n6659 DVSS.n3483 0.0419823
R33272 DVSS.n1863 DVSS.n1859 0.0419823
R33273 DVSS.n1751 DVSS.n1747 0.0415354
R33274 DVSS.n4963 DVSS.n4959 0.0415354
R33275 DVSS.n3368 DVSS.n3364 0.0415354
R33276 DVSS.n6431 DVSS.n6427 0.0415354
R33277 DVSS.n4537 DVSS.n4075 0.0401852
R33278 DVSS.n2941 DVSS.n2479 0.0401852
R33279 DVSS.n6005 DVSS.n5543 0.0401852
R33280 DVSS.n940 DVSS.n478 0.0401852
R33281 DVSS.n6664 DVSS.n6663 0.0375575
R33282 DVSS.n1868 DVSS.n1867 0.0375575
R33283 DVSS.n6689 DVSS.n6687 0.0364513
R33284 DVSS.n6724 DVSS.n1891 0.0364513
R33285 DVSS.n1826 DVSS.n1824 0.036243
R33286 DVSS.n5038 DVSS.n5036 0.036243
R33287 DVSS.n3443 DVSS.n3441 0.036243
R33288 DVSS.n6507 DVSS.n6505 0.036243
R33289 DVSS.n1308 DVSS.n1307 0.034934
R33290 DVSS.n1263 DVSS.n1259 0.0344623
R33291 DVSS.n1283 DVSS.n1280 0.0339906
R33292 DVSS.n1304 DVSS.n1300 0.0339906
R33293 DVSS.n1799 DVSS.n1795 0.0333283
R33294 DVSS.n5011 DVSS.n5007 0.0333283
R33295 DVSS.n3416 DVSS.n3412 0.0333283
R33296 DVSS.n6479 DVSS.n6475 0.0333283
R33297 DVSS.n1926 DVSS.n1922 0.03175
R33298 DVSS.n1948 DVSS.n1944 0.03175
R33299 DVSS.n6628 DVSS.n6627 0.03175
R33300 DVSS.n6606 DVSS.n6605 0.03175
R33301 DVSS.n3529 DVSS.n3525 0.03175
R33302 DVSS.n3551 DVSS.n3547 0.03175
R33303 DVSS.n6841 DVSS.n6838 0.03175
R33304 DVSS.n6817 DVSS.n6816 0.03175
R33305 DVSS.n1268 DVSS.n1267 0.0316321
R33306 DVSS.n1922 DVSS.n1919 0.0304745
R33307 DVSS.n1944 DVSS.n1943 0.0304745
R33308 DVSS.n6632 DVSS.n6628 0.0304745
R33309 DVSS.n6610 DVSS.n6606 0.0304745
R33310 DVSS.n3525 DVSS.n3522 0.0304745
R33311 DVSS.n3547 DVSS.n3546 0.0304745
R33312 DVSS.n6845 DVSS.n6841 0.0304745
R33313 DVSS.n6821 DVSS.n6817 0.0304745
R33314 DVSS.n1173 DVSS.n1172 0.0298561
R33315 DVSS.n6676 DVSS.n6672 0.0298142
R33316 DVSS.n1880 DVSS.n1876 0.0298142
R33317 DVSS.n3714 DVSS 0.0286915
R33318 DVSS.n4179 DVSS 0.0286915
R33319 DVSS.n2118 DVSS 0.0286915
R33320 DVSS.n2583 DVSS 0.0286915
R33321 DVSS.n5182 DVSS 0.0286915
R33322 DVSS.n5647 DVSS 0.0286915
R33323 DVSS.n117 DVSS 0.0286915
R33324 DVSS.n582 DVSS 0.0286915
R33325 DVSS.n1795 DVSS.n1792 0.0282778
R33326 DVSS.n5007 DVSS.n5004 0.0282778
R33327 DVSS.n3412 DVSS.n3409 0.0282778
R33328 DVSS.n6475 DVSS.n6472 0.0282778
R33329 DVSS.n1166 DVSS.n1165 0.0279621
R33330 DVSS.n5065 DVSS.n3608 0.0271646
R33331 DVSS.n3470 DVSS.n2012 0.0271646
R33332 DVSS.n6531 DVSS.n5076 0.0271646
R33333 DVSS.n1853 DVSS.n11 0.0271646
R33334 DVSS.n1830 DVSS.n1826 0.026142
R33335 DVSS.n5042 DVSS.n5038 0.026142
R33336 DVSS.n3447 DVSS.n3443 0.026142
R33337 DVSS.n6510 DVSS.n6507 0.026142
R33338 DVSS.n1851 DVSS.n1843 0.0249644
R33339 DVSS.n5063 DVSS.n5055 0.0249644
R33340 DVSS.n3468 DVSS.n3460 0.0249644
R33341 DVSS.n6529 DVSS.n6521 0.0249644
R33342 DVSS.n6738 DVSS.n6732 0.0245
R33343 DVSS.n6703 DVSS.n6697 0.0245
R33344 DVSS.n3493 DVSS.n3489 0.0245
R33345 DVSS.n6876 DVSS.n6872 0.0245
R33346 DVSS.n4066 DVSS.n3610 0.0244362
R33347 DVSS.n2470 DVSS.n2014 0.0244362
R33348 DVSS.n5534 DVSS.n5078 0.0244362
R33349 DVSS.n469 DVSS.n13 0.0244362
R33350 DVSS.n6672 DVSS.n6668 0.0242832
R33351 DVSS.n1876 DVSS.n1872 0.0242832
R33352 DVSS.n1844 DVSS 0.0237145
R33353 DVSS.n5056 DVSS 0.0237145
R33354 DVSS.n3461 DVSS 0.0237145
R33355 DVSS.n6522 DVSS 0.0237145
R33356 DVSS.n6532 DVSS 0.0236262
R33357 DVSS.n3472 DVSS 0.0236262
R33358 DVSS.n1293 DVSS.n1292 0.0236132
R33359 DVSS.n1315 DVSS.n1312 0.0236132
R33360 DVSS.n1162 DVSS 0.0232273
R33361 DVSS.n6688 DVSS 0.023177
R33362 DVSS.n6723 DVSS 0.023177
R33363 DVSS.n1339 DVSS 0.0231415
R33364 DVSS DVSS.n1120 0.0230564
R33365 DVSS DVSS.n1127 0.0229719
R33366 DVSS.n6708 DVSS 0.0229545
R33367 DVSS.n6743 DVSS 0.0229545
R33368 DVSS.n3744 DVSS.n3742 0.0228214
R33369 DVSS.n3723 DVSS.n3721 0.0228214
R33370 DVSS.n4209 DVSS.n4207 0.0228214
R33371 DVSS.n4188 DVSS.n4186 0.0228214
R33372 DVSS.n2148 DVSS.n2146 0.0228214
R33373 DVSS.n2127 DVSS.n2125 0.0228214
R33374 DVSS.n2613 DVSS.n2611 0.0228214
R33375 DVSS.n2592 DVSS.n2590 0.0228214
R33376 DVSS.n5212 DVSS.n5210 0.0228214
R33377 DVSS.n5191 DVSS.n5189 0.0228214
R33378 DVSS.n5677 DVSS.n5675 0.0228214
R33379 DVSS.n5656 DVSS.n5654 0.0228214
R33380 DVSS.n147 DVSS.n145 0.0228214
R33381 DVSS.n126 DVSS.n124 0.0228214
R33382 DVSS.n612 DVSS.n610 0.0228214
R33383 DVSS.n591 DVSS.n589 0.0228214
R33384 DVSS.n1296 DVSS.n1293 0.0226698
R33385 DVSS.n1318 DVSS.n1315 0.0226698
R33386 DVSS.n1183 DVSS.n1182 0.0222446
R33387 DVSS.n1008 DVSS.n1004 0.0210993
R33388 DVSS.n6540 DVSS.n6538 0.0204913
R33389 DVSS.n2011 DVSS.n2010 0.0201544
R33390 DVSS.n1040 DVSS.n1039 0.0200389
R33391 DVSS.n6712 DVSS.n6711 0.0199344
R33392 DVSS.n5064 DVSS.n4952 0.0198972
R33393 DVSS.n3469 DVSS.n3357 0.0198972
R33394 DVSS.n6530 DVSS.n6420 0.0198972
R33395 DVSS.n1852 DVSS.n1739 0.0198972
R33396 DVSS.n3755 DVSS.n3736 0.0198452
R33397 DVSS.n3734 DVSS.n3715 0.0198452
R33398 DVSS.n4220 DVSS.n4201 0.0198452
R33399 DVSS.n4199 DVSS.n4180 0.0198452
R33400 DVSS.n2159 DVSS.n2140 0.0198452
R33401 DVSS.n2138 DVSS.n2119 0.0198452
R33402 DVSS.n2624 DVSS.n2605 0.0198452
R33403 DVSS.n2603 DVSS.n2584 0.0198452
R33404 DVSS.n5223 DVSS.n5204 0.0198452
R33405 DVSS.n5202 DVSS.n5183 0.0198452
R33406 DVSS.n5688 DVSS.n5669 0.0198452
R33407 DVSS.n5667 DVSS.n5648 0.0198452
R33408 DVSS.n158 DVSS.n139 0.0198452
R33409 DVSS.n137 DVSS.n118 0.0198452
R33410 DVSS.n623 DVSS.n604 0.0198452
R33411 DVSS.n602 DVSS.n583 0.0198452
R33412 DVSS.n1973 DVSS.n1972 0.0196327
R33413 DVSS.n6581 DVSS.n6577 0.0196327
R33414 DVSS.n3576 DVSS.n3575 0.0196327
R33415 DVSS.n6793 DVSS.n6789 0.0196327
R33416 DVSS.n6747 DVSS.n6746 0.0195975
R33417 DVSS.n3482 DVSS.n3481 0.01875
R33418 DVSS.n6877 DVSS.n7 0.01875
R33419 DVSS.n1130 DVSS 0.0187371
R33420 DVSS.n3954 DVSS.n3953 0.0185851
R33421 DVSS.n3958 DVSS.n3954 0.0185851
R33422 DVSS.n3958 DVSS.n3957 0.0185851
R33423 DVSS.n3957 DVSS.n3956 0.0185851
R33424 DVSS.n3956 DVSS.n3651 0.0185851
R33425 DVSS.n3970 DVSS.n3651 0.0185851
R33426 DVSS.n3978 DVSS.n3977 0.0185851
R33427 DVSS.n3973 DVSS.n3972 0.0185851
R33428 DVSS.n3972 DVSS.n3637 0.0185851
R33429 DVSS.n3992 DVSS.n3637 0.0185851
R33430 DVSS.n3993 DVSS.n3992 0.0185851
R33431 DVSS.n3998 DVSS.n3635 0.0185851
R33432 DVSS.n3999 DVSS.n3998 0.0185851
R33433 DVSS.n4026 DVSS.n3999 0.0185851
R33434 DVSS.n4024 DVSS.n4000 0.0185851
R33435 DVSS.n4000 DVSS.n3619 0.0185851
R33436 DVSS.n3619 DVSS.n3617 0.0185851
R33437 DVSS.n4064 DVSS.n3617 0.0185851
R33438 DVSS.n4065 DVSS.n4064 0.0185851
R33439 DVSS.n4067 DVSS.n4065 0.0185851
R33440 DVSS.n4419 DVSS.n4418 0.0185851
R33441 DVSS.n4423 DVSS.n4419 0.0185851
R33442 DVSS.n4423 DVSS.n4422 0.0185851
R33443 DVSS.n4422 DVSS.n4421 0.0185851
R33444 DVSS.n4421 DVSS.n4116 0.0185851
R33445 DVSS.n4435 DVSS.n4116 0.0185851
R33446 DVSS.n4443 DVSS.n4442 0.0185851
R33447 DVSS.n4438 DVSS.n4437 0.0185851
R33448 DVSS.n4437 DVSS.n4102 0.0185851
R33449 DVSS.n4457 DVSS.n4102 0.0185851
R33450 DVSS.n4458 DVSS.n4457 0.0185851
R33451 DVSS.n4463 DVSS.n4100 0.0185851
R33452 DVSS.n4464 DVSS.n4463 0.0185851
R33453 DVSS.n4491 DVSS.n4464 0.0185851
R33454 DVSS.n4489 DVSS.n4465 0.0185851
R33455 DVSS.n4465 DVSS.n4084 0.0185851
R33456 DVSS.n4084 DVSS.n4082 0.0185851
R33457 DVSS.n4529 DVSS.n4082 0.0185851
R33458 DVSS.n4530 DVSS.n4529 0.0185851
R33459 DVSS.n4531 DVSS.n4530 0.0185851
R33460 DVSS.n2358 DVSS.n2357 0.0185851
R33461 DVSS.n2362 DVSS.n2358 0.0185851
R33462 DVSS.n2362 DVSS.n2361 0.0185851
R33463 DVSS.n2361 DVSS.n2360 0.0185851
R33464 DVSS.n2360 DVSS.n2055 0.0185851
R33465 DVSS.n2374 DVSS.n2055 0.0185851
R33466 DVSS.n2382 DVSS.n2381 0.0185851
R33467 DVSS.n2377 DVSS.n2376 0.0185851
R33468 DVSS.n2376 DVSS.n2041 0.0185851
R33469 DVSS.n2396 DVSS.n2041 0.0185851
R33470 DVSS.n2397 DVSS.n2396 0.0185851
R33471 DVSS.n2402 DVSS.n2039 0.0185851
R33472 DVSS.n2403 DVSS.n2402 0.0185851
R33473 DVSS.n2430 DVSS.n2403 0.0185851
R33474 DVSS.n2428 DVSS.n2404 0.0185851
R33475 DVSS.n2404 DVSS.n2023 0.0185851
R33476 DVSS.n2023 DVSS.n2021 0.0185851
R33477 DVSS.n2468 DVSS.n2021 0.0185851
R33478 DVSS.n2469 DVSS.n2468 0.0185851
R33479 DVSS.n2471 DVSS.n2469 0.0185851
R33480 DVSS.n2823 DVSS.n2822 0.0185851
R33481 DVSS.n2827 DVSS.n2823 0.0185851
R33482 DVSS.n2827 DVSS.n2826 0.0185851
R33483 DVSS.n2826 DVSS.n2825 0.0185851
R33484 DVSS.n2825 DVSS.n2520 0.0185851
R33485 DVSS.n2839 DVSS.n2520 0.0185851
R33486 DVSS.n2847 DVSS.n2846 0.0185851
R33487 DVSS.n2842 DVSS.n2841 0.0185851
R33488 DVSS.n2841 DVSS.n2506 0.0185851
R33489 DVSS.n2861 DVSS.n2506 0.0185851
R33490 DVSS.n2862 DVSS.n2861 0.0185851
R33491 DVSS.n2867 DVSS.n2504 0.0185851
R33492 DVSS.n2868 DVSS.n2867 0.0185851
R33493 DVSS.n2895 DVSS.n2868 0.0185851
R33494 DVSS.n2893 DVSS.n2869 0.0185851
R33495 DVSS.n2869 DVSS.n2488 0.0185851
R33496 DVSS.n2488 DVSS.n2486 0.0185851
R33497 DVSS.n2933 DVSS.n2486 0.0185851
R33498 DVSS.n2934 DVSS.n2933 0.0185851
R33499 DVSS.n2935 DVSS.n2934 0.0185851
R33500 DVSS.n5422 DVSS.n5421 0.0185851
R33501 DVSS.n5426 DVSS.n5422 0.0185851
R33502 DVSS.n5426 DVSS.n5425 0.0185851
R33503 DVSS.n5425 DVSS.n5424 0.0185851
R33504 DVSS.n5424 DVSS.n5119 0.0185851
R33505 DVSS.n5438 DVSS.n5119 0.0185851
R33506 DVSS.n5446 DVSS.n5445 0.0185851
R33507 DVSS.n5441 DVSS.n5440 0.0185851
R33508 DVSS.n5440 DVSS.n5105 0.0185851
R33509 DVSS.n5460 DVSS.n5105 0.0185851
R33510 DVSS.n5461 DVSS.n5460 0.0185851
R33511 DVSS.n5466 DVSS.n5103 0.0185851
R33512 DVSS.n5467 DVSS.n5466 0.0185851
R33513 DVSS.n5494 DVSS.n5467 0.0185851
R33514 DVSS.n5492 DVSS.n5468 0.0185851
R33515 DVSS.n5468 DVSS.n5087 0.0185851
R33516 DVSS.n5087 DVSS.n5085 0.0185851
R33517 DVSS.n5532 DVSS.n5085 0.0185851
R33518 DVSS.n5533 DVSS.n5532 0.0185851
R33519 DVSS.n5535 DVSS.n5533 0.0185851
R33520 DVSS.n5887 DVSS.n5886 0.0185851
R33521 DVSS.n5891 DVSS.n5887 0.0185851
R33522 DVSS.n5891 DVSS.n5890 0.0185851
R33523 DVSS.n5890 DVSS.n5889 0.0185851
R33524 DVSS.n5889 DVSS.n5584 0.0185851
R33525 DVSS.n5903 DVSS.n5584 0.0185851
R33526 DVSS.n5911 DVSS.n5910 0.0185851
R33527 DVSS.n5906 DVSS.n5905 0.0185851
R33528 DVSS.n5905 DVSS.n5570 0.0185851
R33529 DVSS.n5925 DVSS.n5570 0.0185851
R33530 DVSS.n5926 DVSS.n5925 0.0185851
R33531 DVSS.n5931 DVSS.n5568 0.0185851
R33532 DVSS.n5932 DVSS.n5931 0.0185851
R33533 DVSS.n5959 DVSS.n5932 0.0185851
R33534 DVSS.n5957 DVSS.n5933 0.0185851
R33535 DVSS.n5933 DVSS.n5552 0.0185851
R33536 DVSS.n5552 DVSS.n5550 0.0185851
R33537 DVSS.n5997 DVSS.n5550 0.0185851
R33538 DVSS.n5998 DVSS.n5997 0.0185851
R33539 DVSS.n5999 DVSS.n5998 0.0185851
R33540 DVSS.n357 DVSS.n356 0.0185851
R33541 DVSS.n361 DVSS.n357 0.0185851
R33542 DVSS.n361 DVSS.n360 0.0185851
R33543 DVSS.n360 DVSS.n359 0.0185851
R33544 DVSS.n359 DVSS.n54 0.0185851
R33545 DVSS.n373 DVSS.n54 0.0185851
R33546 DVSS.n381 DVSS.n380 0.0185851
R33547 DVSS.n376 DVSS.n375 0.0185851
R33548 DVSS.n375 DVSS.n40 0.0185851
R33549 DVSS.n395 DVSS.n40 0.0185851
R33550 DVSS.n396 DVSS.n395 0.0185851
R33551 DVSS.n401 DVSS.n38 0.0185851
R33552 DVSS.n402 DVSS.n401 0.0185851
R33553 DVSS.n429 DVSS.n402 0.0185851
R33554 DVSS.n427 DVSS.n403 0.0185851
R33555 DVSS.n403 DVSS.n22 0.0185851
R33556 DVSS.n22 DVSS.n20 0.0185851
R33557 DVSS.n467 DVSS.n20 0.0185851
R33558 DVSS.n468 DVSS.n467 0.0185851
R33559 DVSS.n470 DVSS.n468 0.0185851
R33560 DVSS.n822 DVSS.n821 0.0185851
R33561 DVSS.n826 DVSS.n822 0.0185851
R33562 DVSS.n826 DVSS.n825 0.0185851
R33563 DVSS.n825 DVSS.n824 0.0185851
R33564 DVSS.n824 DVSS.n519 0.0185851
R33565 DVSS.n838 DVSS.n519 0.0185851
R33566 DVSS.n846 DVSS.n845 0.0185851
R33567 DVSS.n841 DVSS.n840 0.0185851
R33568 DVSS.n840 DVSS.n505 0.0185851
R33569 DVSS.n860 DVSS.n505 0.0185851
R33570 DVSS.n861 DVSS.n860 0.0185851
R33571 DVSS.n866 DVSS.n503 0.0185851
R33572 DVSS.n867 DVSS.n866 0.0185851
R33573 DVSS.n894 DVSS.n867 0.0185851
R33574 DVSS.n892 DVSS.n868 0.0185851
R33575 DVSS.n868 DVSS.n487 0.0185851
R33576 DVSS.n487 DVSS.n485 0.0185851
R33577 DVSS.n932 DVSS.n485 0.0185851
R33578 DVSS.n933 DVSS.n932 0.0185851
R33579 DVSS.n934 DVSS.n933 0.0185851
R33580 DVSS.n1171 DVSS.n1166 0.0184924
R33581 DVSS.n3471 DVSS.n2011 0.0184133
R33582 DVSS.n1067 DVSS.n1066 0.0183571
R33583 DVSS.n1080 DVSS.n1079 0.0183259
R33584 DVSS.n1792 DVSS.n1788 0.0181768
R33585 DVSS.n1816 DVSS.n1812 0.0181768
R33586 DVSS.n5004 DVSS.n5000 0.0181768
R33587 DVSS.n5028 DVSS.n5024 0.0181768
R33588 DVSS.n3409 DVSS.n3405 0.0181768
R33589 DVSS.n3433 DVSS.n3429 0.0181768
R33590 DVSS.n6472 DVSS.n6468 0.0181768
R33591 DVSS.n6496 DVSS.n6492 0.0181768
R33592 DVSS.n6538 DVSS.n6537 0.0180768
R33593 DVSS.n4728 DVSS.n4726 0.0180439
R33594 DVSS.n4754 DVSS.n4752 0.0180439
R33595 DVSS.n6196 DVSS.n6194 0.0180439
R33596 DVSS.n6222 DVSS.n6220 0.0180439
R33597 DVSS.n3132 DVSS.n3130 0.0180439
R33598 DVSS.n3158 DVSS.n3156 0.0180439
R33599 DVSS.n1515 DVSS.n1513 0.0180439
R33600 DVSS.n1541 DVSS.n1539 0.0180439
R33601 DVSS.n4952 DVSS.n4951 0.0179419
R33602 DVSS.n3357 DVSS.n3356 0.0179419
R33603 DVSS.n6420 DVSS.n6419 0.0179419
R33604 DVSS.n1739 DVSS.n1738 0.0179419
R33605 DVSS.n6746 DVSS.n6745 0.0179177
R33606 DVSS.n6885 DVSS.n0 0.0176509
R33607 DVSS.n6687 DVSS.n6685 0.017646
R33608 DVSS.n1891 DVSS.n1889 0.017646
R33609 DVSS.n6711 DVSS.n6710 0.0175813
R33610 DVSS.n1851 DVSS.n1850 0.0175455
R33611 DVSS.n5063 DVSS.n5062 0.0175455
R33612 DVSS.n3468 DVSS.n3467 0.0175455
R33613 DVSS.n6529 DVSS.n6528 0.0175455
R33614 DVSS.n3606 DVSS.n3605 0.0170816
R33615 DVSS.n6763 DVSS.n6759 0.0170816
R33616 DVSS.n3994 DVSS.n3635 0.0169894
R33617 DVSS.n4459 DVSS.n4100 0.0169894
R33618 DVSS.n2398 DVSS.n2039 0.0169894
R33619 DVSS.n2863 DVSS.n2504 0.0169894
R33620 DVSS.n5462 DVSS.n5103 0.0169894
R33621 DVSS.n5927 DVSS.n5568 0.0169894
R33622 DVSS.n397 DVSS.n38 0.0169894
R33623 DVSS.n862 DVSS.n503 0.0169894
R33624 DVSS.n4610 DVSS.n4608 0.0169474
R33625 DVSS.n4634 DVSS.n4620 0.0169474
R33626 DVSS.n4860 DVSS.n4858 0.0169474
R33627 DVSS.n4884 DVSS.n4870 0.0169474
R33628 DVSS.n6078 DVSS.n6076 0.0169474
R33629 DVSS.n6102 DVSS.n6088 0.0169474
R33630 DVSS.n6328 DVSS.n6326 0.0169474
R33631 DVSS.n6352 DVSS.n6338 0.0169474
R33632 DVSS.n3014 DVSS.n3012 0.0169474
R33633 DVSS.n3038 DVSS.n3024 0.0169474
R33634 DVSS.n3264 DVSS.n3262 0.0169474
R33635 DVSS.n3288 DVSS.n3274 0.0169474
R33636 DVSS.n1397 DVSS.n1395 0.0169474
R33637 DVSS.n1421 DVSS.n1407 0.0169474
R33638 DVSS.n1647 DVSS.n1645 0.0169474
R33639 DVSS.n1671 DVSS.n1657 0.0169474
R33640 DVSS.n1144 DVSS.n1142 0.0168374
R33641 DVSS.n1172 DVSS.n1171 0.0165985
R33642 DVSS.n6668 DVSS.n6664 0.0165398
R33643 DVSS.n1872 DVSS.n1868 0.0165398
R33644 DVSS.n1067 DVSS.n1065 0.0164774
R33645 DVSS.n1943 DVSS.n1939 0.0164439
R33646 DVSS.n1964 DVSS.n1960 0.0164439
R33647 DVSS.n3473 DVSS.n3471 0.0164439
R33648 DVSS.n6614 DVSS.n6610 0.0164439
R33649 DVSS.n6590 DVSS.n6589 0.0164439
R33650 DVSS.n6537 DVSS.n6536 0.0164439
R33651 DVSS.n3546 DVSS.n3542 0.0164439
R33652 DVSS.n3567 DVSS.n3563 0.0164439
R33653 DVSS.n6825 DVSS.n6821 0.0164439
R33654 DVSS.n6802 DVSS.n6801 0.0164439
R33655 DVSS.n1194 DVSS.n1193 0.016125
R33656 DVSS.n6710 DVSS.n6709 0.0159703
R33657 DVSS.n6745 DVSS.n6744 0.0159703
R33658 DVSS.n4713 DVSS.n4711 0.0158509
R33659 DVSS.n4769 DVSS.n4767 0.0158509
R33660 DVSS.n6181 DVSS.n6179 0.0158509
R33661 DVSS.n6237 DVSS.n6235 0.0158509
R33662 DVSS.n3117 DVSS.n3115 0.0158509
R33663 DVSS.n3173 DVSS.n3171 0.0158509
R33664 DVSS.n1500 DVSS.n1498 0.0158509
R33665 DVSS.n1556 DVSS.n1554 0.0158509
R33666 DVSS.n4066 DVSS 0.0153308
R33667 DVSS.n2470 DVSS 0.0153308
R33668 DVSS.n5534 DVSS 0.0153308
R33669 DVSS.n469 DVSS 0.0153308
R33670 DVSS.n3510 DVSS.n3509 0.0152059
R33671 DVSS.n6855 DVSS.n6854 0.0152059
R33672 DVSS.n1927 DVSS.n1926 0.0151684
R33673 DVSS.n6627 DVSS.n6623 0.0151684
R33674 DVSS.n3530 DVSS.n3529 0.0151684
R33675 DVSS.n6838 DVSS.n6834 0.0151684
R33676 DVSS.n966 DVSS.n965 0.0150131
R33677 DVSS.n3976 DVSS.n3973 0.0148617
R33678 DVSS.n4441 DVSS.n4438 0.0148617
R33679 DVSS.n2380 DVSS.n2377 0.0148617
R33680 DVSS.n2845 DVSS.n2842 0.0148617
R33681 DVSS.n5444 DVSS.n5441 0.0148617
R33682 DVSS.n5909 DVSS.n5906 0.0148617
R33683 DVSS.n379 DVSS.n376 0.0148617
R33684 DVSS.n844 DVSS.n841 0.0148617
R33685 DVSS.n4592 DVSS.n4590 0.0147544
R33686 DVSS.n4649 DVSS.n4638 0.0147544
R33687 DVSS.n4842 DVSS.n4840 0.0147544
R33688 DVSS.n4899 DVSS.n4888 0.0147544
R33689 DVSS.n6060 DVSS.n6058 0.0147544
R33690 DVSS.n6117 DVSS.n6106 0.0147544
R33691 DVSS.n6310 DVSS.n6308 0.0147544
R33692 DVSS.n6367 DVSS.n6356 0.0147544
R33693 DVSS.n2996 DVSS.n2994 0.0147544
R33694 DVSS.n3053 DVSS.n3042 0.0147544
R33695 DVSS.n3246 DVSS.n3244 0.0147544
R33696 DVSS.n3303 DVSS.n3292 0.0147544
R33697 DVSS.n1379 DVSS.n1377 0.0147544
R33698 DVSS.n1436 DVSS.n1425 0.0147544
R33699 DVSS.n1629 DVSS.n1627 0.0147544
R33700 DVSS.n1686 DVSS.n1675 0.0147544
R33701 DVSS.n6732 DVSS.n1858 0.01475
R33702 DVSS.n6697 DVSS.n6655 0.01475
R33703 DVSS.n3499 DVSS.n3493 0.01475
R33704 DVSS.n6872 DVSS.n6868 0.01475
R33705 DVSS.n1272 DVSS.n1268 0.0146509
R33706 DVSS.n1998 DVSS 0.0145306
R33707 DVSS.n6554 DVSS 0.0145306
R33708 DVSS.n3601 DVSS 0.0145306
R33709 DVSS DVSS.n6764 0.0145306
R33710 DVSS.n6739 DVSS.n6738 0.0145
R33711 DVSS.n6704 DVSS.n6703 0.0145
R33712 DVSS.n6742 DVSS.n6741 0.014
R33713 DVSS.n6707 DVSS.n6706 0.014
R33714 DVSS.n4698 DVSS.n4696 0.0136579
R33715 DVSS.n4784 DVSS.n4782 0.0136579
R33716 DVSS.n6166 DVSS.n6164 0.0136579
R33717 DVSS.n6252 DVSS.n6250 0.0136579
R33718 DVSS.n3102 DVSS.n3100 0.0136579
R33719 DVSS.n3188 DVSS.n3186 0.0136579
R33720 DVSS.n1485 DVSS.n1483 0.0136579
R33721 DVSS.n1571 DVSS.n1569 0.0136579
R33722 DVSS.n1027 DVSS.n1026 0.0136086
R33723 DVSS.n1008 DVSS.n1007 0.0136086
R33724 DVSS.n6881 DVSS.n1 0.0133739
R33725 DVSS.n4577 DVSS.n4575 0.0125614
R33726 DVSS.n4664 DVSS.n4653 0.0125614
R33727 DVSS.n4827 DVSS.n4825 0.0125614
R33728 DVSS.n4914 DVSS.n4903 0.0125614
R33729 DVSS.n6045 DVSS.n6043 0.0125614
R33730 DVSS.n6132 DVSS.n6121 0.0125614
R33731 DVSS.n6295 DVSS.n6293 0.0125614
R33732 DVSS.n6382 DVSS.n6371 0.0125614
R33733 DVSS.n2981 DVSS.n2979 0.0125614
R33734 DVSS.n3068 DVSS.n3057 0.0125614
R33735 DVSS.n3231 DVSS.n3229 0.0125614
R33736 DVSS.n3318 DVSS.n3307 0.0125614
R33737 DVSS.n1364 DVSS.n1362 0.0125614
R33738 DVSS.n1451 DVSS.n1440 0.0125614
R33739 DVSS.n1614 DVSS.n1612 0.0125614
R33740 DVSS.n1701 DVSS.n1690 0.0125614
R33741 DVSS.n1280 DVSS.n1279 0.0122925
R33742 DVSS.n1300 DVSS.n1296 0.0122925
R33743 DVSS.n1332 DVSS.n1331 0.0122781
R33744 DVSS.n6721 DVSS.n3483 0.012115
R33745 DVSS.n1859 DVSS.n2 0.012115
R33746 DVSS.n1986 DVSS.n1982 0.0119796
R33747 DVSS.n6568 DVSS.n6567 0.0119796
R33748 DVSS.n3589 DVSS.n3585 0.0119796
R33749 DVSS.n6780 DVSS.n6779 0.0119796
R33750 DVSS.n1843 DVSS.n1842 0.0117068
R33751 DVSS.n5055 DVSS.n5054 0.0117068
R33752 DVSS.n3460 DVSS.n3459 0.0117068
R33753 DVSS.n6521 DVSS.n6520 0.0117068
R33754 DVSS.n1144 DVSS.n1143 0.0115182
R33755 DVSS.n4683 DVSS.n4681 0.0114649
R33756 DVSS.n4799 DVSS.n4797 0.0114649
R33757 DVSS.n6151 DVSS.n6149 0.0114649
R33758 DVSS.n6267 DVSS.n6265 0.0114649
R33759 DVSS.n3087 DVSS.n3085 0.0114649
R33760 DVSS.n3203 DVSS.n3201 0.0114649
R33761 DVSS.n1470 DVSS.n1468 0.0114649
R33762 DVSS.n1586 DVSS.n1584 0.0114649
R33763 DVSS.n1312 DVSS.n1308 0.0113491
R33764 DVSS.n6677 DVSS.n6676 0.0110088
R33765 DVSS.n1881 DVSS.n1880 0.0110088
R33766 DVSS.n4679 DVSS.n4668 0.0103684
R33767 DVSS.n4812 DVSS.n4810 0.0103684
R33768 DVSS.n6147 DVSS.n6136 0.0103684
R33769 DVSS.n6280 DVSS.n6278 0.0103684
R33770 DVSS.n3083 DVSS.n3072 0.0103684
R33771 DVSS.n3216 DVSS.n3214 0.0103684
R33772 DVSS.n1466 DVSS.n1455 0.0103684
R33773 DVSS.n1599 DVSS.n1597 0.0103684
R33774 DVSS.n1896 DVSS.n1858 0.01025
R33775 DVSS.n1899 DVSS 0.01025
R33776 DVSS.n6655 DVSS.n6654 0.01025
R33777 DVSS DVSS.n5071 0.01025
R33778 DVSS.n3499 DVSS.n3498 0.01025
R33779 DVSS.n3501 DVSS 0.01025
R33780 DVSS.n6868 DVSS.n6867 0.01025
R33781 DVSS DVSS.n9 0.01025
R33782 DVSS.n2010 DVSS.n2008 0.0100663
R33783 DVSS.n6544 DVSS.n6540 0.0100663
R33784 DVSS.n6713 DVSS.n6712 0.00978218
R33785 DVSS.n6757 DVSS.n6747 0.00978218
R33786 DVSS DVSS.n3609 0.00950424
R33787 DVSS DVSS.n2013 0.00950424
R33788 DVSS DVSS.n5077 0.00950424
R33789 DVSS DVSS.n12 0.00950424
R33790 DVSS.n1842 DVSS.n1840 0.00933838
R33791 DVSS.n5054 DVSS.n5052 0.00933838
R33792 DVSS.n3459 DVSS.n3457 0.00933838
R33793 DVSS.n6520 DVSS.n6518 0.00933838
R33794 DVSS.n4668 DVSS.n4666 0.00927193
R33795 DVSS.n4814 DVSS.n4812 0.00927193
R33796 DVSS.n6136 DVSS.n6134 0.00927193
R33797 DVSS.n6282 DVSS.n6280 0.00927193
R33798 DVSS.n3072 DVSS.n3070 0.00927193
R33799 DVSS.n3218 DVSS.n3216 0.00927193
R33800 DVSS.n1455 DVSS.n1453 0.00927193
R33801 DVSS.n1601 DVSS.n1599 0.00927193
R33802 DVSS.n1259 DVSS.n1258 0.00899057
R33803 DVSS.n6536 DVSS.n6532 0.00895784
R33804 DVSS.n3473 DVSS.n3472 0.00895784
R33805 DVSS.n1897 DVSS.n1896 0.00875
R33806 DVSS.n6654 DVSS.n6649 0.00875
R33807 DVSS.n3498 DVSS.n3494 0.00875
R33808 DVSS.n6867 DVSS.n6863 0.00875
R33809 DVSS.n6709 DVSS.n6708 0.00872187
R33810 DVSS.n6744 DVSS.n6743 0.00872187
R33811 DVSS.n1850 DVSS.n1844 0.00856303
R33812 DVSS.n5062 DVSS.n5056 0.00856303
R33813 DVSS.n3467 DVSS.n3461 0.00856303
R33814 DVSS.n6528 DVSS.n6522 0.00856303
R33815 DVSS.n1130 DVSS.n964 0.00847872
R33816 DVSS.n4694 DVSS.n4683 0.00817544
R33817 DVSS.n4797 DVSS.n4795 0.00817544
R33818 DVSS.n6162 DVSS.n6151 0.00817544
R33819 DVSS.n6265 DVSS.n6263 0.00817544
R33820 DVSS.n3098 DVSS.n3087 0.00817544
R33821 DVSS.n3201 DVSS.n3199 0.00817544
R33822 DVSS.n1481 DVSS.n1470 0.00817544
R33823 DVSS.n1584 DVSS.n1582 0.00817544
R33824 DVSS.n1149 DVSS.n1148 0.00771884
R33825 DVSS.n6740 DVSS.n6739 0.00725
R33826 DVSS.n6705 DVSS.n6704 0.00725
R33827 DVSS.n4579 DVSS.n4577 0.00707895
R33828 DVSS.n4653 DVSS.n4651 0.00707895
R33829 DVSS.n4829 DVSS.n4827 0.00707895
R33830 DVSS.n4903 DVSS.n4901 0.00707895
R33831 DVSS.n6047 DVSS.n6045 0.00707895
R33832 DVSS.n6121 DVSS.n6119 0.00707895
R33833 DVSS.n6297 DVSS.n6295 0.00707895
R33834 DVSS.n6371 DVSS.n6369 0.00707895
R33835 DVSS.n2983 DVSS.n2981 0.00707895
R33836 DVSS.n3057 DVSS.n3055 0.00707895
R33837 DVSS.n3233 DVSS.n3231 0.00707895
R33838 DVSS.n3307 DVSS.n3305 0.00707895
R33839 DVSS.n1366 DVSS.n1364 0.00707895
R33840 DVSS.n1440 DVSS.n1438 0.00707895
R33841 DVSS.n1616 DVSS.n1614 0.00707895
R33842 DVSS.n1690 DVSS.n1688 0.00707895
R33843 DVSS.n3949 DVSS.n3687 0.00688298
R33844 DVSS.n4414 DVSS.n4152 0.00688298
R33845 DVSS.n2353 DVSS.n2091 0.00688298
R33846 DVSS.n2818 DVSS.n2556 0.00688298
R33847 DVSS.n5417 DVSS.n5155 0.00688298
R33848 DVSS.n5882 DVSS.n5620 0.00688298
R33849 DVSS.n352 DVSS.n90 0.00688298
R33850 DVSS.n817 DVSS.n555 0.00688298
R33851 DVSS.n3741 DVSS.n3736 0.00645238
R33852 DVSS.n3720 DVSS.n3715 0.00645238
R33853 DVSS.n4206 DVSS.n4201 0.00645238
R33854 DVSS.n4185 DVSS.n4180 0.00645238
R33855 DVSS.n2145 DVSS.n2140 0.00645238
R33856 DVSS.n2124 DVSS.n2119 0.00645238
R33857 DVSS.n2610 DVSS.n2605 0.00645238
R33858 DVSS.n2589 DVSS.n2584 0.00645238
R33859 DVSS.n5209 DVSS.n5204 0.00645238
R33860 DVSS.n5188 DVSS.n5183 0.00645238
R33861 DVSS.n5674 DVSS.n5669 0.00645238
R33862 DVSS.n5653 DVSS.n5648 0.00645238
R33863 DVSS.n144 DVSS.n139 0.00645238
R33864 DVSS.n123 DVSS.n118 0.00645238
R33865 DVSS.n609 DVSS.n604 0.00645238
R33866 DVSS.n588 DVSS.n583 0.00645238
R33867 DVSS.n4709 DVSS.n4698 0.00598246
R33868 DVSS.n4782 DVSS.n4780 0.00598246
R33869 DVSS.n6177 DVSS.n6166 0.00598246
R33870 DVSS.n6250 DVSS.n6248 0.00598246
R33871 DVSS.n3113 DVSS.n3102 0.00598246
R33872 DVSS.n3186 DVSS.n3184 0.00598246
R33873 DVSS.n1496 DVSS.n1485 0.00598246
R33874 DVSS.n1569 DVSS.n1567 0.00598246
R33875 DVSS.n3944 DVSS.n3735 0.00565464
R33876 DVSS.n4409 DVSS.n4200 0.00565464
R33877 DVSS.n2348 DVSS.n2139 0.00565464
R33878 DVSS.n2813 DVSS.n2604 0.00565464
R33879 DVSS.n5412 DVSS.n5203 0.00565464
R33880 DVSS.n5877 DVSS.n5668 0.00565464
R33881 DVSS.n347 DVSS.n138 0.00565464
R33882 DVSS.n812 DVSS.n603 0.00565464
R33883 DVSS.n1754 DVSS.n1751 0.00491919
R33884 DVSS.n4966 DVSS.n4963 0.00491919
R33885 DVSS.n3371 DVSS.n3368 0.00491919
R33886 DVSS.n6434 DVSS.n6431 0.00491919
R33887 DVSS.n4594 DVSS.n4592 0.00488596
R33888 DVSS.n4638 DVSS.n4636 0.00488596
R33889 DVSS.n4844 DVSS.n4842 0.00488596
R33890 DVSS.n4888 DVSS.n4886 0.00488596
R33891 DVSS.n6062 DVSS.n6060 0.00488596
R33892 DVSS.n6106 DVSS.n6104 0.00488596
R33893 DVSS.n6312 DVSS.n6310 0.00488596
R33894 DVSS.n6356 DVSS.n6354 0.00488596
R33895 DVSS.n2998 DVSS.n2996 0.00488596
R33896 DVSS.n3042 DVSS.n3040 0.00488596
R33897 DVSS.n3248 DVSS.n3246 0.00488596
R33898 DVSS.n3292 DVSS.n3290 0.00488596
R33899 DVSS.n1381 DVSS.n1379 0.00488596
R33900 DVSS.n1425 DVSS.n1423 0.00488596
R33901 DVSS.n1631 DVSS.n1629 0.00488596
R33902 DVSS.n1675 DVSS.n1673 0.00488596
R33903 DVSS.n1200 DVSS.n1199 0.00476136
R33904 DVSS.n3949 DVSS.n3948 0.00475532
R33905 DVSS.n4414 DVSS.n4413 0.00475532
R33906 DVSS.n2353 DVSS.n2352 0.00475532
R33907 DVSS.n2818 DVSS.n2817 0.00475532
R33908 DVSS.n5417 DVSS.n5416 0.00475532
R33909 DVSS.n5882 DVSS.n5881 0.00475532
R33910 DVSS.n352 DVSS.n351 0.00475532
R33911 DVSS.n817 DVSS.n816 0.00475532
R33912 DVSS.n6689 DVSS.n6688 0.00437168
R33913 DVSS.n6724 DVSS.n6723 0.00437168
R33914 DVSS.n1981 DVSS.n1977 0.00432653
R33915 DVSS.n6576 DVSS.n6572 0.00432653
R33916 DVSS.n3584 DVSS.n3580 0.00432653
R33917 DVSS.n6788 DVSS.n6784 0.00432653
R33918 DVSS.n3947 DVSS.n3946 0.00423171
R33919 DVSS.n4412 DVSS.n4411 0.00423171
R33920 DVSS.n2351 DVSS.n2350 0.00423171
R33921 DVSS.n2816 DVSS.n2815 0.00423171
R33922 DVSS.n5415 DVSS.n5414 0.00423171
R33923 DVSS.n5880 DVSS.n5879 0.00423171
R33924 DVSS.n350 DVSS.n349 0.00423171
R33925 DVSS.n815 DVSS.n814 0.00423171
R33926 DVSS.n3977 DVSS.n3976 0.0042234
R33927 DVSS.n4442 DVSS.n4441 0.0042234
R33928 DVSS.n2381 DVSS.n2380 0.0042234
R33929 DVSS.n2846 DVSS.n2845 0.0042234
R33930 DVSS.n5445 DVSS.n5444 0.0042234
R33931 DVSS.n5910 DVSS.n5909 0.0042234
R33932 DVSS.n380 DVSS.n379 0.0042234
R33933 DVSS.n845 DVSS.n844 0.0042234
R33934 DVSS.n4724 DVSS.n4713 0.00378947
R33935 DVSS.n4767 DVSS.n4765 0.00378947
R33936 DVSS.n6192 DVSS.n6181 0.00378947
R33937 DVSS.n6235 DVSS.n6233 0.00378947
R33938 DVSS.n3128 DVSS.n3117 0.00378947
R33939 DVSS.n3171 DVSS.n3169 0.00378947
R33940 DVSS.n1511 DVSS.n1500 0.00378947
R33941 DVSS.n1554 DVSS.n1552 0.00378947
R33942 DVSS.n973 DVSS.n972 0.00377715
R33943 DVSS.n6741 DVSS.n6740 0.00375
R33944 DVSS.n6706 DVSS.n6705 0.00375
R33945 DVSS.n3745 DVSS.n3744 0.00347619
R33946 DVSS.n3724 DVSS.n3723 0.00347619
R33947 DVSS.n4210 DVSS.n4209 0.00347619
R33948 DVSS.n4189 DVSS.n4188 0.00347619
R33949 DVSS.n2149 DVSS.n2148 0.00347619
R33950 DVSS.n2128 DVSS.n2127 0.00347619
R33951 DVSS.n2614 DVSS.n2613 0.00347619
R33952 DVSS.n2593 DVSS.n2592 0.00347619
R33953 DVSS.n5213 DVSS.n5212 0.00347619
R33954 DVSS.n5192 DVSS.n5191 0.00347619
R33955 DVSS.n5678 DVSS.n5677 0.00347619
R33956 DVSS.n5657 DVSS.n5656 0.00347619
R33957 DVSS.n148 DVSS.n147 0.00347619
R33958 DVSS.n127 DVSS.n126 0.00347619
R33959 DVSS.n613 DVSS.n612 0.00347619
R33960 DVSS.n592 DVSS.n591 0.00347619
R33961 DVSS.n1267 DVSS.n1263 0.00333019
R33962 DVSS.n1338 DVSS.n1337 0.00315957
R33963 DVSS.n1808 DVSS.n1804 0.00302525
R33964 DVSS.n5020 DVSS.n5016 0.00302525
R33965 DVSS.n3425 DVSS.n3421 0.00302525
R33966 DVSS.n6488 DVSS.n6484 0.00302525
R33967 DVSS.n3489 DVSS.n3482 0.003
R33968 DVSS.n6877 DVSS.n6876 0.003
R33969 DVSS.n1900 DVSS.n1899 0.00275
R33970 DVSS.n6648 DVSS.n5071 0.00275
R33971 DVSS.n3502 DVSS.n3501 0.00275
R33972 DVSS.n6862 DVSS.n9 0.00275
R33973 DVSS.n4612 DVSS.n4610 0.00269298
R33974 DVSS.n4620 DVSS.n4618 0.00269298
R33975 DVSS.n4862 DVSS.n4860 0.00269298
R33976 DVSS.n4870 DVSS.n4868 0.00269298
R33977 DVSS.n6080 DVSS.n6078 0.00269298
R33978 DVSS.n6088 DVSS.n6086 0.00269298
R33979 DVSS.n6330 DVSS.n6328 0.00269298
R33980 DVSS.n6338 DVSS.n6336 0.00269298
R33981 DVSS.n3016 DVSS.n3014 0.00269298
R33982 DVSS.n3024 DVSS.n3022 0.00269298
R33983 DVSS.n3266 DVSS.n3264 0.00269298
R33984 DVSS.n3274 DVSS.n3272 0.00269298
R33985 DVSS.n1399 DVSS.n1397 0.00269298
R33986 DVSS.n1407 DVSS.n1405 0.00269298
R33987 DVSS.n1649 DVSS.n1647 0.00269298
R33988 DVSS.n1657 DVSS.n1655 0.00269298
R33989 DVSS DVSS.n4074 0.00261864
R33990 DVSS DVSS.n2478 0.00261864
R33991 DVSS DVSS.n5542 0.00261864
R33992 DVSS DVSS.n477 0.00261864
R33993 DVSS.n1900 DVSS 0.0025
R33994 DVSS DVSS.n6648 0.0025
R33995 DVSS.n3502 DVSS 0.0025
R33996 DVSS DVSS.n6862 0.0025
R33997 DVSS.n1840 DVSS.n1836 0.00239394
R33998 DVSS.n5052 DVSS.n5048 0.00239394
R33999 DVSS.n3457 DVSS.n3453 0.00239394
R34000 DVSS.n6518 DVSS.n6515 0.00239394
R34001 DVSS.n1023 DVSS.n1022 0.00237266
R34002 DVSS.n3994 DVSS.n3993 0.00209574
R34003 DVSS.n4459 DVSS.n4458 0.00209574
R34004 DVSS.n2398 DVSS.n2397 0.00209574
R34005 DVSS.n2863 DVSS.n2862 0.00209574
R34006 DVSS.n5462 DVSS.n5461 0.00209574
R34007 DVSS.n5927 DVSS.n5926 0.00209574
R34008 DVSS.n397 DVSS.n396 0.00209574
R34009 DVSS.n862 DVSS.n861 0.00209574
R34010 DVSS.n1129 DVSS.n1128 0.00181464
R34011 DVSS.n2008 DVSS.n2004 0.00177551
R34012 DVSS.n6546 DVSS.n6544 0.00177551
R34013 DVSS.n6713 DVSS.n3607 0.00173762
R34014 DVSS.n6758 DVSS.n6757 0.00173762
R34015 DVSS.n4739 DVSS.n4728 0.00159649
R34016 DVSS.n4752 DVSS.n4750 0.00159649
R34017 DVSS.n6207 DVSS.n6196 0.00159649
R34018 DVSS.n6220 DVSS.n6218 0.00159649
R34019 DVSS.n3143 DVSS.n3132 0.00159649
R34020 DVSS.n3156 DVSS.n3154 0.00159649
R34021 DVSS.n1526 DVSS.n1515 0.00159649
R34022 DVSS.n1539 DVSS.n1537 0.00159649
R34023 DVSS.n4067 DVSS.n4066 0.00156383
R34024 DVSS.n4531 DVSS.n4075 0.00156383
R34025 DVSS.n2471 DVSS.n2470 0.00156383
R34026 DVSS.n2935 DVSS.n2479 0.00156383
R34027 DVSS.n5535 DVSS.n5534 0.00156383
R34028 DVSS.n5999 DVSS.n5543 0.00156383
R34029 DVSS.n470 DVSS.n469 0.00156383
R34030 DVSS.n934 DVSS.n478 0.00156383
R34031 DVSS.n6883 DVSS.n6881 0.00150094
R34032 DVSS.n3948 DVSS.n3947 0.00149989
R34033 DVSS.n4413 DVSS.n4412 0.00149989
R34034 DVSS.n2352 DVSS.n2351 0.00149989
R34035 DVSS.n2817 DVSS.n2816 0.00149989
R34036 DVSS.n5416 DVSS.n5415 0.00149989
R34037 DVSS.n5881 DVSS.n5880 0.00149989
R34038 DVSS.n351 DVSS.n350 0.00149989
R34039 DVSS.n816 DVSS.n815 0.00149989
R34040 DVSS.n6883 DVSS.n6882 0.00149986
R34041 DVSS.n1128 DVSS 0.00127576
R34042 DVSS DVSS.n1897 0.00125
R34043 DVSS.n6649 DVSS 0.00125
R34044 DVSS.n3494 DVSS 0.00125
R34045 DVSS.n6863 DVSS 0.00125
R34046 DVSS.n1959 DVSS.n1954 0.00113776
R34047 DVSS.n6596 DVSS.n6594 0.00113776
R34048 DVSS.n3562 DVSS.n3557 0.00113776
R34049 DVSS.n6808 DVSS.n6807 0.00113776
R34050 DVSS.n6880 DVSS.n6879 0.00100053
R34051 DVSS.n6881 DVSS.n6880 0.00100053
R34052 DVSS.n5064 DVSS.n5063 0.001
R34053 DVSS.n3469 DVSS.n3468 0.001
R34054 DVSS.n6530 DVSS.n6529 0.001
R34055 DVSS.n1852 DVSS.n1851 0.001
R34056 DVSS.n3471 DVSS.n3470 0.001
R34057 DVSS.n6537 DVSS.n6531 0.001
R34058 DVSS.n6710 DVSS.n5065 0.001
R34059 DVSS.n6745 DVSS.n1853 0.001
R34060 DVSS.n1285 DVSS.n1283 0.000971698
R34061 DVSS.n3946 DVSS.n3687 0.000500988
R34062 DVSS.n3951 DVSS.n3687 0.000500988
R34063 DVSS.n4411 DVSS.n4152 0.000500988
R34064 DVSS.n4416 DVSS.n4152 0.000500988
R34065 DVSS.n2350 DVSS.n2091 0.000500988
R34066 DVSS.n2355 DVSS.n2091 0.000500988
R34067 DVSS.n2815 DVSS.n2556 0.000500988
R34068 DVSS.n2820 DVSS.n2556 0.000500988
R34069 DVSS.n5414 DVSS.n5155 0.000500988
R34070 DVSS.n5419 DVSS.n5155 0.000500988
R34071 DVSS.n5879 DVSS.n5620 0.000500988
R34072 DVSS.n5884 DVSS.n5620 0.000500988
R34073 DVSS.n349 DVSS.n90 0.000500988
R34074 DVSS.n354 DVSS.n90 0.000500988
R34075 DVSS.n814 DVSS.n555 0.000500988
R34076 DVSS.n819 DVSS.n555 0.000500988
R34077 DVSS.n4948 DVSS.n4947 0.000500921
R34078 DVSS.n3353 DVSS.n3352 0.000500921
R34079 DVSS.n6416 DVSS.n6415 0.000500921
R34080 DVSS.n1735 DVSS.n1734 0.000500921
R34081 DVSS.n3976 DVSS.n3975 0.000500379
R34082 DVSS.n4441 DVSS.n4440 0.000500379
R34083 DVSS.n2380 DVSS.n2379 0.000500379
R34084 DVSS.n2845 DVSS.n2844 0.000500379
R34085 DVSS.n5444 DVSS.n5443 0.000500379
R34086 DVSS.n5909 DVSS.n5908 0.000500379
R34087 DVSS.n379 DVSS.n378 0.000500379
R34088 DVSS.n844 DVSS.n843 0.000500379
R34089 DVSS.n4066 DVSS.n3611 0.000500334
R34090 DVSS.n4076 DVSS.n4075 0.000500334
R34091 DVSS.n2470 DVSS.n2015 0.000500334
R34092 DVSS.n2480 DVSS.n2479 0.000500334
R34093 DVSS.n5534 DVSS.n5079 0.000500334
R34094 DVSS.n5544 DVSS.n5543 0.000500334
R34095 DVSS.n469 DVSS.n14 0.000500334
R34096 DVSS.n479 DVSS.n478 0.000500334
R34097 DVSS.n3995 DVSS.n3994 0.000500219
R34098 DVSS.n4460 DVSS.n4459 0.000500219
R34099 DVSS.n2399 DVSS.n2398 0.000500219
R34100 DVSS.n2864 DVSS.n2863 0.000500219
R34101 DVSS.n5463 DVSS.n5462 0.000500219
R34102 DVSS.n5928 DVSS.n5927 0.000500219
R34103 DVSS.n398 DVSS.n397 0.000500219
R34104 DVSS.n863 DVSS.n862 0.000500219
R34105 DVSS.n3610 DVSS.n3609 0.000500102
R34106 DVSS.n2014 DVSS.n2013 0.000500102
R34107 DVSS.n5078 DVSS.n5077 0.000500102
R34108 DVSS.n13 DVSS.n12 0.000500102
R34109 a_10204_n8486.n5 a_10204_n8486.t8 136.804
R34110 a_10204_n8486.n5 a_10204_n8486.t6 136.325
R34111 a_10204_n8486.n20 a_10204_n8486.t2 119.999
R34112 a_10204_n8486.n11 a_10204_n8486.t3 93.9023
R34113 a_10204_n8486.n0 a_10204_n8486.t4 93.3044
R34114 a_10204_n8486.n0 a_10204_n8486.t7 93.0848
R34115 a_10204_n8486.n19 a_10204_n8486.n18 92.5005
R34116 a_10204_n8486.n12 a_10204_n8486.t9 92.4623
R34117 a_10204_n8486.n0 a_10204_n8486.t5 69.2281
R34118 a_10204_n8486.n27 a_10204_n8486.n26 29.4833
R34119 a_10204_n8486.n15 a_10204_n8486.t0 27.6955
R34120 a_10204_n8486.t1 a_10204_n8486.n46 27.6955
R34121 a_10204_n8486.n20 a_10204_n8486.n19 15.4626
R34122 a_10204_n8486.n2 a_10204_n8486.n30 9.3005
R34123 a_10204_n8486.n2 a_10204_n8486.n22 9.3005
R34124 a_10204_n8486.n2 a_10204_n8486.n21 9.3005
R34125 a_10204_n8486.n2 a_10204_n8486.n28 9.3005
R34126 a_10204_n8486.n28 a_10204_n8486.n27 9.3005
R34127 a_10204_n8486.n2 a_10204_n8486.n29 9.3005
R34128 a_10204_n8486.n2 a_10204_n8486.n31 9.3005
R34129 a_10204_n8486.n46 a_10204_n8486.n45 9.02061
R34130 a_10204_n8486.n46 a_10204_n8486.n41 9.02061
R34131 a_10204_n8486.n16 a_10204_n8486.n15 9.01961
R34132 a_10204_n8486.n35 a_10204_n8486.n33 8.28285
R34133 a_10204_n8486.n3 a_10204_n8486.n8 8.28285
R34134 a_10204_n8486.n28 a_10204_n8486.n24 5.64756
R34135 a_10204_n8486.n1 a_10204_n8486.n35 5.32328
R34136 a_10204_n8486.n13 a_10204_n8486.n17 4.14168
R34137 a_10204_n8486.n40 a_10204_n8486.n7 4.14168
R34138 a_10204_n8486.n1 a_10204_n8486.n12 4.06959
R34139 a_10204_n8486.n26 a_10204_n8486.n25 3.93153
R34140 a_10204_n8486.n38 a_10204_n8486.n36 3.76521
R34141 a_10204_n8486.n44 a_10204_n8486.n43 3.76521
R34142 a_10204_n8486.n35 a_10204_n8486.n34 3.38874
R34143 a_10204_n8486.n4 a_10204_n8486.n3 3.11016
R34144 a_10204_n8486.n14 a_10204_n8486.n13 3.07321
R34145 a_10204_n8486.n39 a_10204_n8486.n38 3.04543
R34146 a_10204_n8486.n40 a_10204_n8486.n4 3.03311
R34147 a_10204_n8486.n4 a_10204_n8486.n9 3.03311
R34148 a_10204_n8486.n38 a_10204_n8486.n37 2.63579
R34149 a_10204_n8486.n45 a_10204_n8486.n44 2.63579
R34150 a_10204_n8486.n4 a_10204_n8486.n1 2.43716
R34151 a_10204_n8486.n1 a_10204_n8486.n14 2.36361
R34152 a_10204_n8486.n1 a_10204_n8486.n39 2.27338
R34153 a_10204_n8486.n13 a_10204_n8486.n16 2.25932
R34154 a_10204_n8486.n41 a_10204_n8486.n40 2.25932
R34155 a_10204_n8486.n12 a_10204_n8486.n11 1.80772
R34156 a_10204_n8486.n5 a_10204_n8486.n10 1.61433
R34157 a_10204_n8486.n2 a_10204_n8486.n20 1.45534
R34158 a_10204_n8486.n11 a_10204_n8486.n5 1.19419
R34159 a_10204_n8486.n32 a_10204_n8486.n2 1.14499
R34160 a_10204_n8486.n43 a_10204_n8486.n42 1.12991
R34161 a_10204_n8486.n7 a_10204_n8486.n6 1.12991
R34162 a_10204_n8486.n32 a_10204_n8486.n0 1.12005
R34163 a_10204_n8486.n14 a_10204_n8486.n32 0.839613
R34164 a_10204_n8486.n24 a_10204_n8486.n23 0.753441
R34165 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n30 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t9 254.28
R34166 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n7 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n5 197.427
R34167 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n4 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n2 158.445
R34168 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n7 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n6 106.596
R34169 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n18 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t8 60.2505
R34170 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n4 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n3 52.2253
R34171 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n3 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t5 21.2805
R34172 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n3 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t7 21.2805
R34173 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n2 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t4 21.2805
R34174 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n2 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t6 21.2805
R34175 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n5 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t0 17.8272
R34176 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n5 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t2 17.8272
R34177 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n6 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t1 17.8272
R34178 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n6 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.t3 17.8272
R34179 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n8 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n4 12.778
R34180 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n27 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n26 9.3005
R34181 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n16 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n15 9.3005
R34182 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n19 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n18 8.76429
R34183 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n8 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n7 8.36086
R34184 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n14 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n13 8.21641
R34185 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n25 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n24 8.21641
R34186 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n31 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y 5.917
R34187 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n17 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n10 5.64756
R34188 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n12 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n11 5.64756
R34189 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n23 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n22 5.64756
R34190 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n29 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n28 5.64756
R34191 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n0 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n21 4.00441
R34192 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n1 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n9 3.69833
R34193 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n0 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n29 3.03311
R34194 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n1 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n17 3.03311
R34195 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n31 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n30 2.75704
R34196 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n8 2.42212
R34197 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n31 2.35727
R34198 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n0 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n19 2.28739
R34199 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n15 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n14 1.09595
R34200 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n26 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n25 1.09595
R34201 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n17 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n16 0.753441
R34202 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n16 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n12 0.753441
R34203 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n27 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n23 0.753441
R34204 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n29 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n27 0.753441
R34205 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n21 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n20 0.738413
R34206 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n30 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n0 0.313579
R34207 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n0 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y.n1 0.141649
R34208 a_6804_n8486.n3 a_6804_n8486.t9 136.804
R34209 a_6804_n8486.n3 a_6804_n8486.t7 136.325
R34210 a_6804_n8486.n10 a_6804_n8486.t2 119.999
R34211 a_6804_n8486.n26 a_6804_n8486.t6 93.9023
R34212 a_6804_n8486.n22 a_6804_n8486.t4 93.3044
R34213 a_6804_n8486.n22 a_6804_n8486.t8 93.0848
R34214 a_6804_n8486.n9 a_6804_n8486.n8 92.5005
R34215 a_6804_n8486.n27 a_6804_n8486.t3 92.4623
R34216 a_6804_n8486.n23 a_6804_n8486.t5 69.2281
R34217 a_6804_n8486.n17 a_6804_n8486.n16 29.4833
R34218 a_6804_n8486.n38 a_6804_n8486.t0 27.6955
R34219 a_6804_n8486.t1 a_6804_n8486.n49 27.6955
R34220 a_6804_n8486.n10 a_6804_n8486.n9 15.4626
R34221 a_6804_n8486.n0 a_6804_n8486.n20 9.3005
R34222 a_6804_n8486.n0 a_6804_n8486.n12 9.3005
R34223 a_6804_n8486.n0 a_6804_n8486.n11 9.3005
R34224 a_6804_n8486.n0 a_6804_n8486.n18 9.3005
R34225 a_6804_n8486.n18 a_6804_n8486.n17 9.3005
R34226 a_6804_n8486.n0 a_6804_n8486.n19 9.3005
R34227 a_6804_n8486.n0 a_6804_n8486.n21 9.3005
R34228 a_6804_n8486.n39 a_6804_n8486.n38 9.02061
R34229 a_6804_n8486.n49 a_6804_n8486.n48 9.02061
R34230 a_6804_n8486.n49 a_6804_n8486.n7 9.02061
R34231 a_6804_n8486.n30 a_6804_n8486.n29 8.28285
R34232 a_6804_n8486.n42 a_6804_n8486.n43 8.28285
R34233 a_6804_n8486.n18 a_6804_n8486.n14 5.64756
R34234 a_6804_n8486.n1 a_6804_n8486.n36 5.31864
R34235 a_6804_n8486.n40 a_6804_n8486.n37 4.14168
R34236 a_6804_n8486.n47 a_6804_n8486.n46 4.14168
R34237 a_6804_n8486.n1 a_6804_n8486.n27 4.06959
R34238 a_6804_n8486.n16 a_6804_n8486.n15 3.93153
R34239 a_6804_n8486.n36 a_6804_n8486.n35 3.76521
R34240 a_6804_n8486.n30 a_6804_n8486.n28 3.76521
R34241 a_6804_n8486.n6 a_6804_n8486.n5 3.76521
R34242 a_6804_n8486.n32 a_6804_n8486.n31 3.38874
R34243 a_6804_n8486.n2 a_6804_n8486.n42 3.11333
R34244 a_6804_n8486.n33 a_6804_n8486.n32 3.07249
R34245 a_6804_n8486.n33 a_6804_n8486.n30 3.07078
R34246 a_6804_n8486.n41 a_6804_n8486.n40 3.04338
R34247 a_6804_n8486.n47 a_6804_n8486.n2 3.03311
R34248 a_6804_n8486.n2 a_6804_n8486.n44 3.03311
R34249 a_6804_n8486.n36 a_6804_n8486.n34 2.63579
R34250 a_6804_n8486.n7 a_6804_n8486.n6 2.63579
R34251 a_6804_n8486.n1 a_6804_n8486.n41 2.27447
R34252 a_6804_n8486.n40 a_6804_n8486.n39 2.25932
R34253 a_6804_n8486.n48 a_6804_n8486.n47 2.25932
R34254 a_6804_n8486.n27 a_6804_n8486.n26 1.80772
R34255 a_6804_n8486.n3 a_6804_n8486.n25 1.61433
R34256 a_6804_n8486.n5 a_6804_n8486.n4 1.50638
R34257 a_6804_n8486.n0 a_6804_n8486.n10 1.45534
R34258 a_6804_n8486.n26 a_6804_n8486.n3 1.19419
R34259 a_6804_n8486.n24 a_6804_n8486.n23 0.944378
R34260 a_6804_n8486.n14 a_6804_n8486.n13 0.753441
R34261 a_6804_n8486.n46 a_6804_n8486.n45 0.753441
R34262 a_6804_n8486.n23 a_6804_n8486.n22 0.176176
R34263 a_6804_n8486.n2 a_6804_n8486.n1 2.36361
R34264 a_6804_n8486.n1 a_6804_n8486.n33 2.36353
R34265 a_6804_n8486.n24 a_6804_n8486.n0 1.14499
R34266 a_6804_n8486.n2 a_6804_n8486.n24 0.92021
R34267 SELB.n1 SELB.t1 186.374
R34268 SELB.n1 SELB.t2 170.308
R34269 SELB.n2 SELB.n1 139.876
R34270 SELB.n8 SELB.t6 84.8325
R34271 SELB.n9 SELB.t9 84.8325
R34272 SELB.n14 SELB.t4 84.8325
R34273 SELB.n22 SELB.t3 84.8325
R34274 SELB SELB.n10 84.6593
R34275 SELB.n11 SELB.n7 76.0005
R34276 SELB.n13 SELB.n12 76.0005
R34277 SELB.n16 SELB.n15 76.0005
R34278 SELB.n17 SELB.n6 76.0005
R34279 SELB.n21 SELB.n20 76.0005
R34280 SELB.n8 SELB.t8 48.6825
R34281 SELB.n9 SELB.t0 48.6825
R34282 SELB.n14 SELB.t7 48.6825
R34283 SELB.n22 SELB.t5 48.6825
R34284 SELB.n0 SELB 42.9181
R34285 SELB.n10 SELB.n8 34.8915
R34286 SELB.n13 SELB.n7 24.4602
R34287 SELB.n15 SELB.n13 24.4602
R34288 SELB.n21 SELB.n6 24.4602
R34289 SELB.n17 SELB 21.4593
R34290 SELB.n10 SELB.n9 21.2229
R34291 SELB.n14 SELB.n6 20.5035
R34292 SELB SELB.n11 19.2005
R34293 SELB.n20 SELB.n19 18.824
R34294 SELB.n11 SELB 16.9417
R34295 SELB SELB.n17 14.6829
R34296 SELB.n0 SELB 12.8005
R34297 SELB.n23 SELB.n22 12.2304
R34298 SELB.n22 SELB.n21 11.1512
R34299 SELB.n20 SELB 10.9181
R34300 SELB.n26 SELB.n25 9.3005
R34301 SELB.n30 SELB.n28 9.3005
R34302 SELB.n12 SELB 6.4005
R34303 SELB.n19 SELB 6.4005
R34304 SELB.n38 SELB 5.6255
R34305 SELB.n25 SELB.n24 5.20629
R34306 SELB.n3 SELB 4.98883
R34307 SELB.n37 SELB.n36 4.5005
R34308 SELB SELB.n16 4.14168
R34309 SELB.n15 SELB.n14 3.95722
R34310 SELB.n31 SELB 3.65919
R34311 SELB.n19 SELB.n18 3.42907
R34312 SELB.n9 SELB.n7 3.23781
R34313 SELB.n26 SELB.n5 3.2005
R34314 SELB.n32 SELB.n31 3.03171
R34315 SELB SELB.n30 2.51479
R34316 SELB.n27 SELB.n26 1.96244
R34317 SELB.n28 SELB.n27 1.83038
R34318 SELB SELB.n2 1.61978
R34319 SELB.n34 SELB 1.15796
R34320 SELB.n34 SELB.n33 1.10531
R34321 SELB.n36 SELB.n35 1.10429
R34322 SELB.n24 SELB.n23 1.0796
R34323 SELB.n30 SELB.n29 0.93044
R34324 SELB.n2 SELB.n0 0.925801
R34325 SELB.n33 SELB 0.592448
R34326 SELB.n18 SELB 0.457643
R34327 SELB.n3 SELB 0.232113
R34328 SELB SELB.n5 0.229071
R34329 SELB.n33 SELB.n32 0.128495
R34330 SELB.n31 SELB.n28 0.0395621
R34331 SELB.n4 SELB.n3 0.0278528
R34332 SELB.n37 SELB 0.0274737
R34333 SELB.n38 SELB.n37 0.0248421
R34334 SELB.n4 SELB 0.00479904
R34335 SELB.n35 SELB.n34 0.00434615
R34336 SELB SELB.n38 0.00181579
R34337 SELB.n36 SELB.n4 0.00100097
R34338 VO.n8 VO.n7 148.663
R34339 VO.n16 VO.t1 122.728
R34340 VO.n5 VO.t0 22.4191
R34341 VO.n9 VO.n8 10.5541
R34342 VO.n7 VO 9.62836
R34343 VO.n10 VO.n9 9.3005
R34344 VO VO.n12 7.00682
R34345 VO VO.n11 6.32867
R34346 VO.n15 VO.n14 5.92892
R34347 VO.n15 VO.n3 4.72813
R34348 VO.n16 VO 4.69453
R34349 VO.n12 VO.n2 4.6505
R34350 VO.n19 VO.n18 4.6505
R34351 VO.n12 VO 2.96471
R34352 VO.n22 VO.n21 2.68157
R34353 VO VO.n15 2.42576
R34354 VO.n8 VO.n5 2.19143
R34355 VO.n13 VO 2.15629
R34356 VO.n11 VO.n2 2.04091
R34357 VO.n18 VO.n17 1.75208
R34358 VO.n6 VO.n4 1.61734
R34359 VO.n14 VO 1.61734
R34360 VO.n11 VO.n10 0.816947
R34361 VO.n17 VO.n16 0.795743
R34362 VO.n10 VO.n4 0.674184
R34363 VO.n18 VO.n13 0.539447
R34364 VO.n24 VO.n23 0.480413
R34365 VO.n24 VO 0.449398
R34366 VO.n7 VO 0.343399
R34367 VO VO.n6 0.269974
R34368 VO.n21 VO.n20 0.0807632
R34369 VO.n23 VO.n22 0.0740294
R34370 VO VO.n25 0.067276
R34371 VO.n25 VO.n24 0.0391741
R34372 VO.n0 VO 0.0282247
R34373 VO.n1 VO.n0 0.0216236
R34374 VO.n25 VO.n1 0.0203034
R34375 VO.n19 VO.n3 0.0176053
R34376 VO.n21 VO.n2 0.00971053
R34377 VO.n20 VO.n19 0.00576316
R34378 a_3606_n8490.n3 a_3606_n8490.t9 136.804
R34379 a_3606_n8490.n3 a_3606_n8490.t6 136.325
R34380 a_3606_n8490.n10 a_3606_n8490.t2 119.999
R34381 a_3606_n8490.n26 a_3606_n8490.t7 93.9023
R34382 a_3606_n8490.n22 a_3606_n8490.t3 93.3044
R34383 a_3606_n8490.n22 a_3606_n8490.t8 93.0848
R34384 a_3606_n8490.n9 a_3606_n8490.n8 92.5005
R34385 a_3606_n8490.n27 a_3606_n8490.t4 92.4623
R34386 a_3606_n8490.n23 a_3606_n8490.t5 69.2281
R34387 a_3606_n8490.n17 a_3606_n8490.n16 29.4833
R34388 a_3606_n8490.n38 a_3606_n8490.t0 27.6955
R34389 a_3606_n8490.t1 a_3606_n8490.n49 27.6955
R34390 a_3606_n8490.n10 a_3606_n8490.n9 15.4626
R34391 a_3606_n8490.n0 a_3606_n8490.n20 9.3005
R34392 a_3606_n8490.n0 a_3606_n8490.n12 9.3005
R34393 a_3606_n8490.n0 a_3606_n8490.n11 9.3005
R34394 a_3606_n8490.n0 a_3606_n8490.n18 9.3005
R34395 a_3606_n8490.n18 a_3606_n8490.n17 9.3005
R34396 a_3606_n8490.n0 a_3606_n8490.n19 9.3005
R34397 a_3606_n8490.n0 a_3606_n8490.n21 9.3005
R34398 a_3606_n8490.n39 a_3606_n8490.n38 9.02061
R34399 a_3606_n8490.n49 a_3606_n8490.n48 9.02061
R34400 a_3606_n8490.n49 a_3606_n8490.n7 9.02061
R34401 a_3606_n8490.n30 a_3606_n8490.n29 8.28285
R34402 a_3606_n8490.n42 a_3606_n8490.n43 8.28285
R34403 a_3606_n8490.n18 a_3606_n8490.n14 5.64756
R34404 a_3606_n8490.n1 a_3606_n8490.n36 5.31864
R34405 a_3606_n8490.n40 a_3606_n8490.n37 4.14168
R34406 a_3606_n8490.n47 a_3606_n8490.n46 4.14168
R34407 a_3606_n8490.n1 a_3606_n8490.n27 4.06959
R34408 a_3606_n8490.n16 a_3606_n8490.n15 3.93153
R34409 a_3606_n8490.n36 a_3606_n8490.n35 3.76521
R34410 a_3606_n8490.n30 a_3606_n8490.n28 3.76521
R34411 a_3606_n8490.n6 a_3606_n8490.n5 3.76521
R34412 a_3606_n8490.n32 a_3606_n8490.n31 3.38874
R34413 a_3606_n8490.n2 a_3606_n8490.n42 3.11333
R34414 a_3606_n8490.n33 a_3606_n8490.n32 3.07249
R34415 a_3606_n8490.n33 a_3606_n8490.n30 3.07078
R34416 a_3606_n8490.n41 a_3606_n8490.n40 3.04338
R34417 a_3606_n8490.n47 a_3606_n8490.n2 3.03311
R34418 a_3606_n8490.n2 a_3606_n8490.n44 3.03311
R34419 a_3606_n8490.n36 a_3606_n8490.n34 2.63579
R34420 a_3606_n8490.n7 a_3606_n8490.n6 2.63579
R34421 a_3606_n8490.n1 a_3606_n8490.n41 2.27447
R34422 a_3606_n8490.n40 a_3606_n8490.n39 2.25932
R34423 a_3606_n8490.n48 a_3606_n8490.n47 2.25932
R34424 a_3606_n8490.n27 a_3606_n8490.n26 1.80772
R34425 a_3606_n8490.n3 a_3606_n8490.n25 1.61433
R34426 a_3606_n8490.n5 a_3606_n8490.n4 1.50638
R34427 a_3606_n8490.n0 a_3606_n8490.n10 1.45534
R34428 a_3606_n8490.n26 a_3606_n8490.n3 1.19419
R34429 a_3606_n8490.n24 a_3606_n8490.n23 0.944378
R34430 a_3606_n8490.n14 a_3606_n8490.n13 0.753441
R34431 a_3606_n8490.n46 a_3606_n8490.n45 0.753441
R34432 a_3606_n8490.n23 a_3606_n8490.n22 0.176176
R34433 a_3606_n8490.n2 a_3606_n8490.n1 2.36361
R34434 a_3606_n8490.n1 a_3606_n8490.n33 2.36353
R34435 a_3606_n8490.n24 a_3606_n8490.n0 1.14499
R34436 a_3606_n8490.n2 a_3606_n8490.n24 0.92021
R34437 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 356.022
R34438 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n64 292.5
R34439 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n28 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n23 152
R34440 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n33 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n22 152
R34441 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n38 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n21 152
R34442 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n43 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n20 152
R34443 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n19 152
R34444 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n53 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n18 152
R34445 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n58 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n17 152
R34446 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n60 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n59 152
R34447 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n55 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n54 152
R34448 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n50 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n49 152
R34449 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n45 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n44 152
R34450 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n40 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n39 152
R34451 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n34 152
R34452 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n30 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n29 152
R34453 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n64 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t0 147.756
R34454 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t1 105.415
R34455 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t4 84.8325
R34456 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t5 84.8325
R34457 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n13 60.1541
R34458 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n15 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 50.1642
R34459 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t2 48.6825
R34460 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t3 48.6825
R34461 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n62 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n61 45.1373
R34462 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 36.3683
R34463 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n1 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n60 33.7894
R34464 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n56 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n55 29.03
R34465 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n51 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n50 29.03
R34466 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n45 29.03
R34467 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n41 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n40 29.03
R34468 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n35 29.03
R34469 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n31 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n30 29.03
R34470 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n26 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n25 28.4823
R34471 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n25 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n24 26.4823
R34472 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n15 15.6972
R34473 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n59 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n11 16.3795
R34474 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n54 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n6 16.2631
R34475 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n49 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n8 16.1289
R34476 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n10 15.9761
R34477 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n65 10.4732
R34478 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n11 2.10258
R34479 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n6 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 2.08561
R34480 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n57 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n56 9.3005
R34481 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 2.07495
R34482 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n52 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n51 9.3005
R34483 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n10 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 2.07042
R34484 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n47 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n46 9.3005
R34485 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n9 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 2.07192
R34486 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n42 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n41 9.3005
R34487 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n7 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 2.0795
R34488 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n37 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n36 9.3005
R34489 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n32 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n5 2.77054
R34490 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n32 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n31 9.3005
R34491 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n5 2.09329
R34492 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n27 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n26 9.3005
R34493 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n2 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n1 18.3534
R34494 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n26 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n23 8.76414
R34495 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n31 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n22 7.66868
R34496 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n60 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n17 7.12095
R34497 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n63 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n62 6.98232
R34498 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n62 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 6.73734
R34499 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n21 6.57323
R34500 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n55 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n18 6.0255
R34501 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n28 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n27 6.02403
R34502 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n41 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n20 5.47777
R34503 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n33 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n32 5.27109
R34504 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n61 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 5.22977
R34505 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n63 5.04292
R34506 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n50 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n19 4.93005
R34507 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n59 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n58 4.89462
R34508 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 4.74124
R34509 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n2 4.55946
R34510 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n38 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n37 4.51815
R34511 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n37 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n7 2.64533
R34512 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n27 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n24 4.45253
R34513 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n19 4.38232
R34514 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n54 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n53 4.14168
R34515 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 3.87929
R34516 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 3.87929
R34517 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n45 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n20 3.83459
R34518 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n43 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n42 3.76521
R34519 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n42 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n9 2.50198
R34520 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n16 3.43953
R34521 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n49 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n48 3.38874
R34522 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n51 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n18 3.28686
R34523 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n47 3.01226
R34524 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n47 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n10 2.33997
R34525 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n40 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n21 2.73914
R34526 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n43 2.63579
R34527 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n39 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n9 15.804
R34528 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n53 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n52 2.25932
R34529 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n52 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n8 2.15681
R34530 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n56 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n17 2.19141
R34531 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n39 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n38 1.88285
R34532 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n34 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n7 15.6099
R34533 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n22 1.64368
R34534 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 1.52175
R34535 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n25 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.t6 1.50675
R34536 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n58 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n57 1.50638
R34537 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n57 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n6 1.95132
R34538 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 1.37511
R34539 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n15 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 1.1768
R34540 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n34 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n33 1.12991
R34541 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n29 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n5 15.3925
R34542 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n11 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n1 4.58496
R34543 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 0.679754
R34544 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n30 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n23 0.548227
R34545 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n61 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH 0.546841
R34546 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n24 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 0.471686
R34547 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 0.468612
R34548 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n29 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n28 0.376971
R34549 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n2 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 0.310701
R34550 a_6804_n3484.n3 a_6804_n3484.t4 136.804
R34551 a_6804_n3484.n3 a_6804_n3484.t3 136.325
R34552 a_6804_n3484.n10 a_6804_n3484.t2 119.999
R34553 a_6804_n3484.n26 a_6804_n3484.t8 93.9023
R34554 a_6804_n3484.n22 a_6804_n3484.t5 93.3044
R34555 a_6804_n3484.n22 a_6804_n3484.t9 93.0848
R34556 a_6804_n3484.n9 a_6804_n3484.n8 92.5005
R34557 a_6804_n3484.n27 a_6804_n3484.t7 92.4623
R34558 a_6804_n3484.n23 a_6804_n3484.t6 69.2281
R34559 a_6804_n3484.n17 a_6804_n3484.n16 29.4833
R34560 a_6804_n3484.n38 a_6804_n3484.t0 27.6955
R34561 a_6804_n3484.t1 a_6804_n3484.n49 27.6955
R34562 a_6804_n3484.n10 a_6804_n3484.n9 15.4626
R34563 a_6804_n3484.n0 a_6804_n3484.n20 9.3005
R34564 a_6804_n3484.n0 a_6804_n3484.n12 9.3005
R34565 a_6804_n3484.n0 a_6804_n3484.n11 9.3005
R34566 a_6804_n3484.n0 a_6804_n3484.n18 9.3005
R34567 a_6804_n3484.n18 a_6804_n3484.n17 9.3005
R34568 a_6804_n3484.n0 a_6804_n3484.n19 9.3005
R34569 a_6804_n3484.n0 a_6804_n3484.n21 9.3005
R34570 a_6804_n3484.n39 a_6804_n3484.n38 9.02061
R34571 a_6804_n3484.n49 a_6804_n3484.n48 9.02061
R34572 a_6804_n3484.n49 a_6804_n3484.n7 9.02061
R34573 a_6804_n3484.n30 a_6804_n3484.n29 8.28285
R34574 a_6804_n3484.n42 a_6804_n3484.n43 8.28285
R34575 a_6804_n3484.n18 a_6804_n3484.n14 5.64756
R34576 a_6804_n3484.n1 a_6804_n3484.n36 5.31864
R34577 a_6804_n3484.n40 a_6804_n3484.n37 4.14168
R34578 a_6804_n3484.n47 a_6804_n3484.n46 4.14168
R34579 a_6804_n3484.n1 a_6804_n3484.n27 4.06959
R34580 a_6804_n3484.n16 a_6804_n3484.n15 3.93153
R34581 a_6804_n3484.n36 a_6804_n3484.n35 3.76521
R34582 a_6804_n3484.n30 a_6804_n3484.n28 3.76521
R34583 a_6804_n3484.n6 a_6804_n3484.n5 3.76521
R34584 a_6804_n3484.n32 a_6804_n3484.n31 3.38874
R34585 a_6804_n3484.n2 a_6804_n3484.n42 3.11333
R34586 a_6804_n3484.n33 a_6804_n3484.n32 3.07249
R34587 a_6804_n3484.n33 a_6804_n3484.n30 3.07078
R34588 a_6804_n3484.n41 a_6804_n3484.n40 3.04338
R34589 a_6804_n3484.n47 a_6804_n3484.n2 3.03311
R34590 a_6804_n3484.n2 a_6804_n3484.n44 3.03311
R34591 a_6804_n3484.n36 a_6804_n3484.n34 2.63579
R34592 a_6804_n3484.n7 a_6804_n3484.n6 2.63579
R34593 a_6804_n3484.n1 a_6804_n3484.n41 2.27447
R34594 a_6804_n3484.n40 a_6804_n3484.n39 2.25932
R34595 a_6804_n3484.n48 a_6804_n3484.n47 2.25932
R34596 a_6804_n3484.n27 a_6804_n3484.n26 1.80772
R34597 a_6804_n3484.n3 a_6804_n3484.n25 1.61433
R34598 a_6804_n3484.n5 a_6804_n3484.n4 1.50638
R34599 a_6804_n3484.n0 a_6804_n3484.n10 1.45534
R34600 a_6804_n3484.n26 a_6804_n3484.n3 1.19419
R34601 a_6804_n3484.n24 a_6804_n3484.n23 0.944378
R34602 a_6804_n3484.n14 a_6804_n3484.n13 0.753441
R34603 a_6804_n3484.n46 a_6804_n3484.n45 0.753441
R34604 a_6804_n3484.n23 a_6804_n3484.n22 0.176176
R34605 a_6804_n3484.n2 a_6804_n3484.n1 2.36361
R34606 a_6804_n3484.n1 a_6804_n3484.n33 2.36353
R34607 a_6804_n3484.n24 a_6804_n3484.n0 1.14499
R34608 a_6804_n3484.n2 a_6804_n3484.n24 0.92021
R34609 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n31 185
R34610 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n43 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n42 185
R34611 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n63 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n50 185
R34612 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n62 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n61 185
R34613 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n83 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n70 185
R34614 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n82 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n81 185
R34615 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n105 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n91 185
R34616 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n104 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n103 185
R34617 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n120 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t4 120.037
R34618 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n149 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t5 120.037
R34619 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n32 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t15 120.037
R34620 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n51 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t16 120.037
R34621 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n71 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t9 120.037
R34622 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n92 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t10 120.037
R34623 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n43 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n37 112.831
R34624 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n62 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n57 112.831
R34625 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n82 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n76 112.831
R34626 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n104 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n99 112.831
R34627 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n45 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n36 104.172
R34628 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n64 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n56 104.172
R34629 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n84 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n75 104.172
R34630 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n106 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n97 104.172
R34631 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n119 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n118 92.5005
R34632 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n148 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n147 92.5005
R34633 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n35 92.5005
R34634 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n56 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n55 92.5005
R34635 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n75 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n74 92.5005
R34636 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n97 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n96 92.5005
R34637 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t15 66.8281
R34638 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n56 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t16 66.8281
R34639 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n75 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t9 66.8281
R34640 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n97 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t10 66.8281
R34641 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n112 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t8 47.0064
R34642 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t1 36.328
R34643 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n7 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t12 35.7839
R34644 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n114 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t0 35.2053
R34645 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n126 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n125 29.4833
R34646 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n142 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n141 29.4833
R34647 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n45 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n44 29.4833
R34648 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n64 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n63 29.4833
R34649 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n84 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n83 29.4833
R34650 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n106 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n105 29.4833
R34651 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n113 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t7 27.6955
R34652 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n113 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t6 27.6955
R34653 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n120 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n119 15.4558
R34654 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n149 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n148 15.4558
R34655 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n32 15.4558
R34656 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n55 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n51 15.4558
R34657 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n74 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n71 15.4558
R34658 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n96 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n92 15.4558
R34659 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n42 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n41 13.5534
R34660 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n61 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n60 13.5534
R34661 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n81 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n80 13.5534
R34662 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n103 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n102 13.5534
R34663 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n113 9.67857
R34664 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n34 9.41227
R34665 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n55 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n54 9.41227
R34666 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n74 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n73 9.41227
R34667 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n96 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n95 9.41227
R34668 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n99 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n98 9.3037
R34669 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n117 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n121 9.3005
R34670 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n127 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n126 9.3005
R34671 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n146 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n150 9.3005
R34672 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n143 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n142 9.3005
R34673 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n41 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n40 9.3005
R34674 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n34 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n33 9.3005
R34675 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n30 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n28 9.3005
R34676 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n29 9.3005
R34677 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n45 9.3005
R34678 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n60 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n59 9.3005
R34679 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n54 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n53 9.3005
R34680 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n52 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n26 9.3005
R34681 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n66 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n65 9.3005
R34682 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n64 9.3005
R34683 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n80 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n79 9.3005
R34684 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n73 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n72 9.3005
R34685 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n69 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n25 9.3005
R34686 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n85 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n68 9.3005
R34687 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n85 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n84 9.3005
R34688 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n102 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n101 9.3005
R34689 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n95 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n94 9.3005
R34690 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n93 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n23 9.3005
R34691 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n108 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n107 9.3005
R34692 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n107 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n106 9.3005
R34693 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t2 8.2655
R34694 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t3 8.2655
R34695 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n11 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n10 7.26743
R34696 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n11 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n8 6.15568
R34697 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n127 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n123 5.64756
R34698 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n143 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n139 5.64756
R34699 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n31 5.64756
R34700 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n50 5.64756
R34701 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n85 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n70 5.64756
R34702 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n107 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n91 5.64756
R34703 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n135 5.29345
R34704 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n132 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n130 4.89462
R34705 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n153 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n151 4.89462
R34706 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n38 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n37 4.89462
R34707 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n58 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n57 4.89462
R34708 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n77 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n76 4.89462
R34709 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n100 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n99 4.89462
R34710 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n135 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n133 4.89462
R34711 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n129 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n127 4.51815
R34712 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n145 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n143 4.51815
R34713 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t11 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n7 35.3416
R34714 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n15 35.2708
R34715 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.t14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n14 35.2708
R34716 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n89 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n22 4.5005
R34717 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n110 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n22 4.5005
R34718 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n109 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n89 4.5005
R34719 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n110 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n109 4.5005
R34720 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n19 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n18 1.49962
R34721 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n88 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n17 4.5005
R34722 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n20 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n19 0.00981422
R34723 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n20 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n87 2.24659
R34724 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n1 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n2 1.12391
R34725 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n67 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n1 2.24659
R34726 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n4 1.12391
R34727 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n6 0.00725908
R34728 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n48 2.24659
R34729 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n34 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n30 4.14168
R34730 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n47 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n46 4.14168
R34731 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n54 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n52 4.14168
R34732 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n27 4.14168
R34733 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n73 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n69 4.14168
R34734 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n86 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n85 4.14168
R34735 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n95 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n93 4.14168
R34736 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n107 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n24 4.14168
R34737 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n125 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n124 3.93153
R34738 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n141 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n140 3.93153
R34739 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n43 3.93153
R34740 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n63 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n62 3.93153
R34741 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n83 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n82 3.93153
R34742 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n105 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n104 3.93153
R34743 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n116 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n132 3.07655
R34744 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n137 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n153 3.07514
R34745 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n100 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n22 3.03311
R34746 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n109 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n24 3.03311
R34747 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n77 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n17 3.03311
R34748 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n87 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n86 3.03311
R34749 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n58 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n5 3.03311
R34750 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n67 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n27 3.03311
R34751 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n38 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n6 3.03311
R34752 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n47 3.03311
R34753 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n136 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n145 3.03311
R34754 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n115 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n129 3.03311
R34755 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n112 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN 2.63881
R34756 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n12 2.28594
R34757 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n47 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n30 2.25932
R34758 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n52 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n27 2.25932
R34759 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n86 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n69 2.25932
R34760 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n93 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n24 2.25932
R34761 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n57 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n2 9.31071
R34762 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n98 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n21 2.25315
R34763 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n76 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n18 9.30786
R34764 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n129 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n128 1.88285
R34765 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n145 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n144 1.88285
R34766 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n132 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n131 1.50638
R34767 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n153 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n152 1.50638
R34768 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n41 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n38 1.50638
R34769 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n60 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n58 1.50638
R34770 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n80 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n77 1.50638
R34771 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n102 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n100 1.50638
R34772 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n135 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n134 1.50638
R34773 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n156 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n116 1.50133
R34774 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n33 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n32 1.4932
R34775 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n53 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n51 1.4932
R34776 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n94 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n92 1.4932
R34777 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n72 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n71 1.49258
R34778 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n78 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n19 1.4922
R34779 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n137 1.49213
R34780 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n117 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n120 1.49212
R34781 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n90 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n21 1.49182
R34782 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n49 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n1 1.49182
R34783 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n39 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n3 1.49182
R34784 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n146 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n149 1.49166
R34785 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n112 1.25694
R34786 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n123 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n122 0.753441
R34787 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n139 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n138 0.753441
R34788 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n42 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n31 0.753441
R34789 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n61 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n50 0.753441
R34790 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n81 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n70 0.753441
R34791 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n103 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n91 0.753441
R34792 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n111 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n110 0.55213
R34793 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n10 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n9 0.521921
R34794 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n157 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n114 0.29767
R34795 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n111 0.296016
R34796 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n157 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n156 0.196255
R34797 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n157 0.1855
R34798 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n89 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n88 0.1255
R34799 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n155 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n154 0.124821
R34800 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n11 0.0579027
R34801 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n40 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n39 0.0382131
R34802 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n59 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n49 0.0382131
R34803 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n101 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n90 0.0382131
R34804 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n79 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n78 0.0366935
R34805 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n116 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n115 0.0332098
R34806 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n137 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n136 0.0321501
R34807 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n15 0.269649
R34808 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n108 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n90 0.0216934
R34809 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n66 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n49 0.0216934
R34810 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n39 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n29 0.0216934
R34811 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n78 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n68 0.0208694
R34812 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n115 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n117 0.018819
R34813 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n136 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n146 0.0182083
R34814 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n154 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n16 0.018163
R34815 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n88 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n20 0.00981422
R34816 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n89 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n21 0.0134076
R34817 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n33 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n28 0.0123534
R34818 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n29 0.0123534
R34819 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n53 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n26 0.0123534
R34820 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n67 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n66 0.0123534
R34821 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n94 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n23 0.0123534
R34822 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n109 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n108 0.0123534
R34823 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n37 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n4 9.31071
R34824 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n2 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n5 0.00725908
R34825 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n98 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n22 0.0123089
R34826 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n72 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n25 0.0118636
R34827 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n87 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n68 0.0118636
R34828 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n18 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n17 0.00854565
R34829 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n15 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n7 0.254871
R34830 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n28 0.00696552
R34831 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n67 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n26 0.00696552
R34832 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n109 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n23 0.00696552
R34833 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n87 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n25 0.00669835
R34834 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n110 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n21 0.00525544
R34835 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n40 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n6 0.00481034
R34836 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n59 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n5 0.00481034
R34837 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n101 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n22 0.00481034
R34838 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n79 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n17 0.00463223
R34839 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n156 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n155 0.00457609
R34840 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n111 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n14 0.515676
R34841 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n1 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n3 0.251465
R34842 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n13 0.240989
R34843 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n114 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n0 0.180788
R34844 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n19 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN.n1 0.150243
R34845 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 356.022
R34846 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n64 292.5
R34847 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n28 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n23 152
R34848 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n33 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n22 152
R34849 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n38 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n21 152
R34850 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n43 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n20 152
R34851 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n19 152
R34852 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n53 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n18 152
R34853 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n58 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n17 152
R34854 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n60 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n59 152
R34855 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n55 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n54 152
R34856 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n50 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n49 152
R34857 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n45 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n44 152
R34858 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n40 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n39 152
R34859 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n34 152
R34860 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n30 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n29 152
R34861 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n64 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t0 147.756
R34862 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t1 105.415
R34863 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t5 84.8325
R34864 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t6 84.8325
R34865 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n13 60.1541
R34866 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n15 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 50.1642
R34867 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t3 48.6825
R34868 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t4 48.6825
R34869 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n62 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n61 45.1373
R34870 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 36.3683
R34871 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n1 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n60 33.7894
R34872 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n56 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n55 29.03
R34873 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n51 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n50 29.03
R34874 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n45 29.03
R34875 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n41 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n40 29.03
R34876 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n35 29.03
R34877 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n31 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n30 29.03
R34878 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n26 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n25 28.4823
R34879 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n25 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n24 26.4823
R34880 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n15 15.6972
R34881 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n59 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n11 16.3795
R34882 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n54 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n6 16.2631
R34883 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n49 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n8 16.1289
R34884 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n10 15.9761
R34885 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n65 10.4732
R34886 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n11 2.10258
R34887 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n6 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 2.08561
R34888 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n57 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n56 9.3005
R34889 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n8 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 2.07495
R34890 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n52 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n51 9.3005
R34891 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n10 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 2.07042
R34892 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n47 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n46 9.3005
R34893 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n9 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 2.07192
R34894 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n42 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n41 9.3005
R34895 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n7 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 2.0795
R34896 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n37 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n36 9.3005
R34897 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n32 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n5 2.77054
R34898 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n32 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n31 9.3005
R34899 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n5 2.09329
R34900 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n27 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n26 9.3005
R34901 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n2 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n1 18.3534
R34902 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n26 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n23 8.76414
R34903 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n31 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n22 7.66868
R34904 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n60 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n17 7.12095
R34905 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n63 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n62 6.98232
R34906 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n62 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 6.73734
R34907 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n21 6.57323
R34908 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n55 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n18 6.0255
R34909 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n28 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n27 6.02403
R34910 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n41 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n20 5.47777
R34911 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n33 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n32 5.27109
R34912 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n61 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 5.22977
R34913 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n63 5.04292
R34914 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n50 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n19 4.93005
R34915 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n59 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n58 4.89462
R34916 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 4.74124
R34917 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n2 4.55946
R34918 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n38 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n37 4.51815
R34919 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n37 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n7 2.64533
R34920 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n27 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n24 4.45253
R34921 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n46 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n19 4.38232
R34922 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n54 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n53 4.14168
R34923 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 3.87929
R34924 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n65 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 3.87929
R34925 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n45 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n20 3.83459
R34926 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n43 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n42 3.76521
R34927 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n42 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n9 2.50198
R34928 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n16 3.43953
R34929 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n49 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n48 3.38874
R34930 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n51 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n18 3.28686
R34931 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n47 3.01226
R34932 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n47 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n10 2.33997
R34933 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n40 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n21 2.73914
R34934 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n43 2.63579
R34935 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n39 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n9 15.804
R34936 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n53 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n52 2.25932
R34937 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n52 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n8 2.15681
R34938 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n56 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n17 2.19141
R34939 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n39 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n38 1.88285
R34940 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n34 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n7 15.6099
R34941 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n22 1.64368
R34942 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 1.52175
R34943 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n25 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.t2 1.50675
R34944 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n58 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n57 1.50638
R34945 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n57 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n6 1.95132
R34946 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 1.37511
R34947 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n15 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 1.1768
R34948 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n34 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n33 1.12991
R34949 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n29 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n5 15.3925
R34950 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n11 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n1 4.58496
R34951 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 0.679754
R34952 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n30 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n23 0.548227
R34953 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n61 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH 0.546841
R34954 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n24 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 0.471686
R34955 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 0.468612
R34956 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n29 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n28 0.376971
R34957 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n2 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 0.310701
R34958 a_10209_n9511.n10 a_10209_n9511.t2 120.01
R34959 a_10209_n9511.n3 a_10209_n9511.t4 92.9415
R34960 a_10209_n9511.n9 a_10209_n9511.n8 92.5005
R34961 a_10209_n9511.n3 a_10209_n9511.t3 92.4623
R34962 a_10209_n9511.n22 a_10209_n9511.t5 73.195
R34963 a_10209_n9511.n22 a_10209_n9511.t6 72.1651
R34964 a_10209_n9511.n17 a_10209_n9511.n16 29.4833
R34965 a_10209_n9511.n26 a_10209_n9511.t0 27.6955
R34966 a_10209_n9511.t1 a_10209_n9511.n41 27.6955
R34967 a_10209_n9511.n10 a_10209_n9511.n9 15.4607
R34968 a_10209_n9511.n0 a_10209_n9511.n12 9.3005
R34969 a_10209_n9511.n0 a_10209_n9511.n19 9.3005
R34970 a_10209_n9511.n0 a_10209_n9511.n18 9.3005
R34971 a_10209_n9511.n18 a_10209_n9511.n17 9.3005
R34972 a_10209_n9511.n0 a_10209_n9511.n11 9.3005
R34973 a_10209_n9511.n0 a_10209_n9511.n21 9.3005
R34974 a_10209_n9511.n0 a_10209_n9511.n20 9.3005
R34975 a_10209_n9511.n41 a_10209_n9511.n40 9.02061
R34976 a_10209_n9511.n41 a_10209_n9511.n7 9.02061
R34977 a_10209_n9511.n27 a_10209_n9511.n26 9.01961
R34978 a_10209_n9511.n25 a_10209_n9511.n23 8.28285
R34979 a_10209_n9511.n34 a_10209_n9511.n35 8.28285
R34980 a_10209_n9511.n18 a_10209_n9511.n14 5.64756
R34981 a_10209_n9511.n2 a_10209_n9511.n25 5.32161
R34982 a_10209_n9511.n2 a_10209_n9511.n29 5.31894
R34983 a_10209_n9511.n29 a_10209_n9511.n28 4.14168
R34984 a_10209_n9511.n39 a_10209_n9511.n38 4.14168
R34985 a_10209_n9511.n2 a_10209_n9511.n3 4.03426
R34986 a_10209_n9511.n16 a_10209_n9511.n15 3.93153
R34987 a_10209_n9511.n32 a_10209_n9511.n30 3.76521
R34988 a_10209_n9511.n6 a_10209_n9511.n5 3.76521
R34989 a_10209_n9511.n3 a_10209_n9511.n22 3.20519
R34990 a_10209_n9511.n1 a_10209_n9511.n34 3.11223
R34991 a_10209_n9511.n33 a_10209_n9511.n32 3.04478
R34992 a_10209_n9511.n39 a_10209_n9511.n1 3.03311
R34993 a_10209_n9511.n1 a_10209_n9511.n36 3.03311
R34994 a_10209_n9511.n25 a_10209_n9511.n24 3.01226
R34995 a_10209_n9511.n32 a_10209_n9511.n31 2.63579
R34996 a_10209_n9511.n7 a_10209_n9511.n6 2.63579
R34997 a_10209_n9511.n1 a_10209_n9511.n2 2.47579
R34998 a_10209_n9511.n2 a_10209_n9511.n33 2.27623
R34999 a_10209_n9511.n29 a_10209_n9511.n27 2.25932
R35000 a_10209_n9511.n40 a_10209_n9511.n39 2.25932
R35001 a_10209_n9511.n1 a_10209_n9511.n0 1.9858
R35002 a_10209_n9511.n5 a_10209_n9511.n4 1.88285
R35003 a_10209_n9511.n0 a_10209_n9511.n10 1.64258
R35004 a_10209_n9511.n14 a_10209_n9511.n13 0.753441
R35005 a_10209_n9511.n38 a_10209_n9511.n37 0.376971
R35006 a_3606_n3488.n3 a_3606_n3488.t6 136.804
R35007 a_3606_n3488.n3 a_3606_n3488.t3 136.325
R35008 a_3606_n3488.n10 a_3606_n3488.t2 119.999
R35009 a_3606_n3488.n26 a_3606_n3488.t4 93.9023
R35010 a_3606_n3488.n22 a_3606_n3488.t7 93.3044
R35011 a_3606_n3488.n22 a_3606_n3488.t5 93.0848
R35012 a_3606_n3488.n9 a_3606_n3488.n8 92.5005
R35013 a_3606_n3488.n27 a_3606_n3488.t8 92.4623
R35014 a_3606_n3488.n23 a_3606_n3488.t9 69.2281
R35015 a_3606_n3488.n17 a_3606_n3488.n16 29.4833
R35016 a_3606_n3488.n38 a_3606_n3488.t0 27.6955
R35017 a_3606_n3488.t1 a_3606_n3488.n49 27.6955
R35018 a_3606_n3488.n10 a_3606_n3488.n9 15.4626
R35019 a_3606_n3488.n0 a_3606_n3488.n20 9.3005
R35020 a_3606_n3488.n0 a_3606_n3488.n12 9.3005
R35021 a_3606_n3488.n0 a_3606_n3488.n11 9.3005
R35022 a_3606_n3488.n0 a_3606_n3488.n18 9.3005
R35023 a_3606_n3488.n18 a_3606_n3488.n17 9.3005
R35024 a_3606_n3488.n0 a_3606_n3488.n19 9.3005
R35025 a_3606_n3488.n0 a_3606_n3488.n21 9.3005
R35026 a_3606_n3488.n39 a_3606_n3488.n38 9.02061
R35027 a_3606_n3488.n49 a_3606_n3488.n48 9.02061
R35028 a_3606_n3488.n49 a_3606_n3488.n7 9.02061
R35029 a_3606_n3488.n30 a_3606_n3488.n29 8.28285
R35030 a_3606_n3488.n42 a_3606_n3488.n43 8.28285
R35031 a_3606_n3488.n18 a_3606_n3488.n14 5.64756
R35032 a_3606_n3488.n1 a_3606_n3488.n36 5.31864
R35033 a_3606_n3488.n40 a_3606_n3488.n37 4.14168
R35034 a_3606_n3488.n47 a_3606_n3488.n46 4.14168
R35035 a_3606_n3488.n1 a_3606_n3488.n27 4.06959
R35036 a_3606_n3488.n16 a_3606_n3488.n15 3.93153
R35037 a_3606_n3488.n36 a_3606_n3488.n35 3.76521
R35038 a_3606_n3488.n30 a_3606_n3488.n28 3.76521
R35039 a_3606_n3488.n6 a_3606_n3488.n5 3.76521
R35040 a_3606_n3488.n32 a_3606_n3488.n31 3.38874
R35041 a_3606_n3488.n2 a_3606_n3488.n42 3.11333
R35042 a_3606_n3488.n33 a_3606_n3488.n32 3.07249
R35043 a_3606_n3488.n33 a_3606_n3488.n30 3.07078
R35044 a_3606_n3488.n41 a_3606_n3488.n40 3.04338
R35045 a_3606_n3488.n47 a_3606_n3488.n2 3.03311
R35046 a_3606_n3488.n2 a_3606_n3488.n44 3.03311
R35047 a_3606_n3488.n36 a_3606_n3488.n34 2.63579
R35048 a_3606_n3488.n7 a_3606_n3488.n6 2.63579
R35049 a_3606_n3488.n1 a_3606_n3488.n41 2.27447
R35050 a_3606_n3488.n40 a_3606_n3488.n39 2.25932
R35051 a_3606_n3488.n48 a_3606_n3488.n47 2.25932
R35052 a_3606_n3488.n27 a_3606_n3488.n26 1.80772
R35053 a_3606_n3488.n3 a_3606_n3488.n25 1.61433
R35054 a_3606_n3488.n5 a_3606_n3488.n4 1.50638
R35055 a_3606_n3488.n0 a_3606_n3488.n10 1.45534
R35056 a_3606_n3488.n26 a_3606_n3488.n3 1.19419
R35057 a_3606_n3488.n24 a_3606_n3488.n23 0.944378
R35058 a_3606_n3488.n14 a_3606_n3488.n13 0.753441
R35059 a_3606_n3488.n46 a_3606_n3488.n45 0.753441
R35060 a_3606_n3488.n23 a_3606_n3488.n22 0.176176
R35061 a_3606_n3488.n2 a_3606_n3488.n1 2.36361
R35062 a_3606_n3488.n1 a_3606_n3488.n33 2.36353
R35063 a_3606_n3488.n24 a_3606_n3488.n0 1.14499
R35064 a_3606_n3488.n2 a_3606_n3488.n24 0.92021
R35065 SELA.n1 SELA.t3 186.374
R35066 SELA.n1 SELA.t4 170.308
R35067 SELA.n2 SELA.n1 139.876
R35068 SELA.n8 SELA.t0 84.8325
R35069 SELA.n9 SELA.t7 84.8325
R35070 SELA.n14 SELA.t8 84.8325
R35071 SELA.n22 SELA.t5 84.8325
R35072 SELA SELA.n10 84.6593
R35073 SELA.n11 SELA.n7 76.0005
R35074 SELA.n13 SELA.n12 76.0005
R35075 SELA.n16 SELA.n15 76.0005
R35076 SELA.n17 SELA.n6 76.0005
R35077 SELA.n21 SELA.n20 76.0005
R35078 SELA.n8 SELA.t6 48.6825
R35079 SELA.n9 SELA.t1 48.6825
R35080 SELA.n14 SELA.t2 48.6825
R35081 SELA.n22 SELA.t9 48.6825
R35082 SELA.n0 SELA 42.9181
R35083 SELA.n10 SELA.n8 34.8915
R35084 SELA.n13 SELA.n7 24.4602
R35085 SELA.n15 SELA.n13 24.4602
R35086 SELA.n21 SELA.n6 24.4602
R35087 SELA.n17 SELA 21.4593
R35088 SELA.n10 SELA.n9 21.2229
R35089 SELA.n14 SELA.n6 20.5035
R35090 SELA SELA.n11 19.2005
R35091 SELA.n20 SELA.n19 18.824
R35092 SELA.n11 SELA 16.9417
R35093 SELA SELA.n17 14.6829
R35094 SELA.n0 SELA 12.8005
R35095 SELA.n23 SELA.n22 12.2304
R35096 SELA.n22 SELA.n21 11.1512
R35097 SELA.n20 SELA 10.9181
R35098 SELA.n26 SELA.n25 9.3005
R35099 SELA.n30 SELA.n28 9.3005
R35100 SELA.n12 SELA 6.4005
R35101 SELA.n19 SELA 6.4005
R35102 SELA.n38 SELA 5.6255
R35103 SELA.n25 SELA.n24 5.20629
R35104 SELA.n3 SELA 4.98883
R35105 SELA.n37 SELA.n36 4.5005
R35106 SELA SELA.n16 4.14168
R35107 SELA.n15 SELA.n14 3.95722
R35108 SELA.n31 SELA 3.65919
R35109 SELA.n19 SELA.n18 3.42907
R35110 SELA.n9 SELA.n7 3.23781
R35111 SELA.n26 SELA.n5 3.2005
R35112 SELA.n32 SELA.n31 3.03171
R35113 SELA SELA.n30 2.51479
R35114 SELA.n27 SELA.n26 1.96244
R35115 SELA.n28 SELA.n27 1.83038
R35116 SELA SELA.n2 1.61978
R35117 SELA.n34 SELA 1.14315
R35118 SELA.n34 SELA.n33 1.10531
R35119 SELA.n36 SELA.n35 1.10429
R35120 SELA.n24 SELA.n23 1.0796
R35121 SELA.n30 SELA.n29 0.93044
R35122 SELA.n2 SELA.n0 0.925801
R35123 SELA.n33 SELA 0.592448
R35124 SELA.n18 SELA 0.457643
R35125 SELA.n3 SELA 0.232113
R35126 SELA SELA.n5 0.229071
R35127 SELA.n33 SELA.n32 0.128495
R35128 SELA.n31 SELA.n28 0.0395621
R35129 SELA.n4 SELA.n3 0.0278528
R35130 SELA.n37 SELA 0.0274737
R35131 SELA.n38 SELA.n37 0.0248421
R35132 SELA.n4 SELA 0.00479904
R35133 SELA.n35 SELA.n34 0.00434615
R35134 SELA SELA.n38 0.00181579
R35135 SELA.n36 SELA.n4 0.00100097
R35136 a_206_n3488.n5 a_206_n3488.t3 136.804
R35137 a_206_n3488.n5 a_206_n3488.t7 136.325
R35138 a_206_n3488.n20 a_206_n3488.t2 119.999
R35139 a_206_n3488.n11 a_206_n3488.t8 93.9023
R35140 a_206_n3488.n0 a_206_n3488.t5 93.3044
R35141 a_206_n3488.n0 a_206_n3488.t9 93.0848
R35142 a_206_n3488.n19 a_206_n3488.n18 92.5005
R35143 a_206_n3488.n12 a_206_n3488.t4 92.4623
R35144 a_206_n3488.n0 a_206_n3488.t6 69.2281
R35145 a_206_n3488.n27 a_206_n3488.n26 29.4833
R35146 a_206_n3488.n15 a_206_n3488.t0 27.6955
R35147 a_206_n3488.t1 a_206_n3488.n46 27.6955
R35148 a_206_n3488.n20 a_206_n3488.n19 15.4626
R35149 a_206_n3488.n2 a_206_n3488.n30 9.3005
R35150 a_206_n3488.n2 a_206_n3488.n22 9.3005
R35151 a_206_n3488.n2 a_206_n3488.n21 9.3005
R35152 a_206_n3488.n2 a_206_n3488.n28 9.3005
R35153 a_206_n3488.n28 a_206_n3488.n27 9.3005
R35154 a_206_n3488.n2 a_206_n3488.n29 9.3005
R35155 a_206_n3488.n2 a_206_n3488.n31 9.3005
R35156 a_206_n3488.n46 a_206_n3488.n45 9.02061
R35157 a_206_n3488.n46 a_206_n3488.n41 9.02061
R35158 a_206_n3488.n16 a_206_n3488.n15 9.01961
R35159 a_206_n3488.n35 a_206_n3488.n33 8.28285
R35160 a_206_n3488.n3 a_206_n3488.n8 8.28285
R35161 a_206_n3488.n28 a_206_n3488.n24 5.64756
R35162 a_206_n3488.n1 a_206_n3488.n35 5.32328
R35163 a_206_n3488.n13 a_206_n3488.n17 4.14168
R35164 a_206_n3488.n40 a_206_n3488.n7 4.14168
R35165 a_206_n3488.n1 a_206_n3488.n12 4.06959
R35166 a_206_n3488.n26 a_206_n3488.n25 3.93153
R35167 a_206_n3488.n38 a_206_n3488.n36 3.76521
R35168 a_206_n3488.n44 a_206_n3488.n43 3.76521
R35169 a_206_n3488.n35 a_206_n3488.n34 3.38874
R35170 a_206_n3488.n4 a_206_n3488.n3 3.11016
R35171 a_206_n3488.n14 a_206_n3488.n13 3.07321
R35172 a_206_n3488.n39 a_206_n3488.n38 3.04543
R35173 a_206_n3488.n40 a_206_n3488.n4 3.03311
R35174 a_206_n3488.n4 a_206_n3488.n9 3.03311
R35175 a_206_n3488.n38 a_206_n3488.n37 2.63579
R35176 a_206_n3488.n45 a_206_n3488.n44 2.63579
R35177 a_206_n3488.n4 a_206_n3488.n1 2.43716
R35178 a_206_n3488.n1 a_206_n3488.n14 2.36361
R35179 a_206_n3488.n1 a_206_n3488.n39 2.27338
R35180 a_206_n3488.n13 a_206_n3488.n16 2.25932
R35181 a_206_n3488.n41 a_206_n3488.n40 2.25932
R35182 a_206_n3488.n12 a_206_n3488.n11 1.80772
R35183 a_206_n3488.n5 a_206_n3488.n10 1.61433
R35184 a_206_n3488.n2 a_206_n3488.n20 1.45534
R35185 a_206_n3488.n11 a_206_n3488.n5 1.19419
R35186 a_206_n3488.n32 a_206_n3488.n2 1.14499
R35187 a_206_n3488.n43 a_206_n3488.n42 1.12991
R35188 a_206_n3488.n7 a_206_n3488.n6 1.12991
R35189 a_206_n3488.n32 a_206_n3488.n0 1.12005
R35190 a_206_n3488.n14 a_206_n3488.n32 0.839613
R35191 a_206_n3488.n24 a_206_n3488.n23 0.753441
R35192 a_3611_n9515.n10 a_3611_n9515.t2 120.01
R35193 a_3611_n9515.n3 a_3611_n9515.t6 92.9415
R35194 a_3611_n9515.n9 a_3611_n9515.n8 92.5005
R35195 a_3611_n9515.n3 a_3611_n9515.t5 92.4623
R35196 a_3611_n9515.n22 a_3611_n9515.t4 73.195
R35197 a_3611_n9515.n22 a_3611_n9515.t3 72.1651
R35198 a_3611_n9515.n17 a_3611_n9515.n16 29.4833
R35199 a_3611_n9515.n26 a_3611_n9515.t0 27.6955
R35200 a_3611_n9515.t1 a_3611_n9515.n41 27.6955
R35201 a_3611_n9515.n10 a_3611_n9515.n9 15.4607
R35202 a_3611_n9515.n0 a_3611_n9515.n12 9.3005
R35203 a_3611_n9515.n0 a_3611_n9515.n19 9.3005
R35204 a_3611_n9515.n0 a_3611_n9515.n18 9.3005
R35205 a_3611_n9515.n18 a_3611_n9515.n17 9.3005
R35206 a_3611_n9515.n0 a_3611_n9515.n11 9.3005
R35207 a_3611_n9515.n0 a_3611_n9515.n21 9.3005
R35208 a_3611_n9515.n0 a_3611_n9515.n20 9.3005
R35209 a_3611_n9515.n41 a_3611_n9515.n40 9.02061
R35210 a_3611_n9515.n41 a_3611_n9515.n7 9.02061
R35211 a_3611_n9515.n27 a_3611_n9515.n26 9.01961
R35212 a_3611_n9515.n25 a_3611_n9515.n23 8.28285
R35213 a_3611_n9515.n34 a_3611_n9515.n35 8.28285
R35214 a_3611_n9515.n18 a_3611_n9515.n14 5.64756
R35215 a_3611_n9515.n2 a_3611_n9515.n25 5.32161
R35216 a_3611_n9515.n2 a_3611_n9515.n29 5.31894
R35217 a_3611_n9515.n29 a_3611_n9515.n28 4.14168
R35218 a_3611_n9515.n39 a_3611_n9515.n38 4.14168
R35219 a_3611_n9515.n2 a_3611_n9515.n3 4.03426
R35220 a_3611_n9515.n16 a_3611_n9515.n15 3.93153
R35221 a_3611_n9515.n32 a_3611_n9515.n30 3.76521
R35222 a_3611_n9515.n6 a_3611_n9515.n5 3.76521
R35223 a_3611_n9515.n3 a_3611_n9515.n22 3.20519
R35224 a_3611_n9515.n1 a_3611_n9515.n34 3.11223
R35225 a_3611_n9515.n33 a_3611_n9515.n32 3.04478
R35226 a_3611_n9515.n39 a_3611_n9515.n1 3.03311
R35227 a_3611_n9515.n1 a_3611_n9515.n36 3.03311
R35228 a_3611_n9515.n25 a_3611_n9515.n24 3.01226
R35229 a_3611_n9515.n32 a_3611_n9515.n31 2.63579
R35230 a_3611_n9515.n7 a_3611_n9515.n6 2.63579
R35231 a_3611_n9515.n1 a_3611_n9515.n2 2.47579
R35232 a_3611_n9515.n2 a_3611_n9515.n33 2.27623
R35233 a_3611_n9515.n29 a_3611_n9515.n27 2.25932
R35234 a_3611_n9515.n40 a_3611_n9515.n39 2.25932
R35235 a_3611_n9515.n1 a_3611_n9515.n0 1.9858
R35236 a_3611_n9515.n5 a_3611_n9515.n4 1.88285
R35237 a_3611_n9515.n0 a_3611_n9515.n10 1.64258
R35238 a_3611_n9515.n14 a_3611_n9515.n13 0.753441
R35239 a_3611_n9515.n38 a_3611_n9515.n37 0.376971
R35240 a_206_n8490.n3 a_206_n8490.t6 136.804
R35241 a_206_n8490.n3 a_206_n8490.t4 136.325
R35242 a_206_n8490.n10 a_206_n8490.t2 119.999
R35243 a_206_n8490.n26 a_206_n8490.t3 93.9023
R35244 a_206_n8490.n22 a_206_n8490.t8 93.3044
R35245 a_206_n8490.n22 a_206_n8490.t5 93.0848
R35246 a_206_n8490.n9 a_206_n8490.n8 92.5005
R35247 a_206_n8490.n27 a_206_n8490.t7 92.4623
R35248 a_206_n8490.n23 a_206_n8490.t9 69.2281
R35249 a_206_n8490.n17 a_206_n8490.n16 29.4833
R35250 a_206_n8490.n38 a_206_n8490.t0 27.6955
R35251 a_206_n8490.t1 a_206_n8490.n49 27.6955
R35252 a_206_n8490.n10 a_206_n8490.n9 15.4626
R35253 a_206_n8490.n0 a_206_n8490.n20 9.3005
R35254 a_206_n8490.n0 a_206_n8490.n12 9.3005
R35255 a_206_n8490.n0 a_206_n8490.n11 9.3005
R35256 a_206_n8490.n0 a_206_n8490.n18 9.3005
R35257 a_206_n8490.n18 a_206_n8490.n17 9.3005
R35258 a_206_n8490.n0 a_206_n8490.n19 9.3005
R35259 a_206_n8490.n0 a_206_n8490.n21 9.3005
R35260 a_206_n8490.n39 a_206_n8490.n38 9.02061
R35261 a_206_n8490.n49 a_206_n8490.n48 9.02061
R35262 a_206_n8490.n49 a_206_n8490.n7 9.02061
R35263 a_206_n8490.n30 a_206_n8490.n29 8.28285
R35264 a_206_n8490.n42 a_206_n8490.n43 8.28285
R35265 a_206_n8490.n18 a_206_n8490.n14 5.64756
R35266 a_206_n8490.n1 a_206_n8490.n36 5.31864
R35267 a_206_n8490.n40 a_206_n8490.n37 4.14168
R35268 a_206_n8490.n47 a_206_n8490.n46 4.14168
R35269 a_206_n8490.n1 a_206_n8490.n27 4.06959
R35270 a_206_n8490.n16 a_206_n8490.n15 3.93153
R35271 a_206_n8490.n36 a_206_n8490.n35 3.76521
R35272 a_206_n8490.n30 a_206_n8490.n28 3.76521
R35273 a_206_n8490.n6 a_206_n8490.n5 3.76521
R35274 a_206_n8490.n32 a_206_n8490.n31 3.38874
R35275 a_206_n8490.n2 a_206_n8490.n42 3.11333
R35276 a_206_n8490.n33 a_206_n8490.n32 3.07249
R35277 a_206_n8490.n33 a_206_n8490.n30 3.07078
R35278 a_206_n8490.n41 a_206_n8490.n40 3.04338
R35279 a_206_n8490.n47 a_206_n8490.n2 3.03311
R35280 a_206_n8490.n2 a_206_n8490.n44 3.03311
R35281 a_206_n8490.n36 a_206_n8490.n34 2.63579
R35282 a_206_n8490.n7 a_206_n8490.n6 2.63579
R35283 a_206_n8490.n1 a_206_n8490.n41 2.27447
R35284 a_206_n8490.n40 a_206_n8490.n39 2.25932
R35285 a_206_n8490.n48 a_206_n8490.n47 2.25932
R35286 a_206_n8490.n27 a_206_n8490.n26 1.80772
R35287 a_206_n8490.n3 a_206_n8490.n25 1.61433
R35288 a_206_n8490.n5 a_206_n8490.n4 1.50638
R35289 a_206_n8490.n0 a_206_n8490.n10 1.45534
R35290 a_206_n8490.n26 a_206_n8490.n3 1.19419
R35291 a_206_n8490.n24 a_206_n8490.n23 0.944378
R35292 a_206_n8490.n14 a_206_n8490.n13 0.753441
R35293 a_206_n8490.n46 a_206_n8490.n45 0.753441
R35294 a_206_n8490.n23 a_206_n8490.n22 0.176176
R35295 a_206_n8490.n2 a_206_n8490.n1 2.36361
R35296 a_206_n8490.n1 a_206_n8490.n33 2.36353
R35297 a_206_n8490.n24 a_206_n8490.n0 1.14499
R35298 a_206_n8490.n2 a_206_n8490.n24 0.92021
R35299 B1.n66 B1.n65 185
R35300 B1.n64 B1.n57 185
R35301 B1.n24 B1.n15 185
R35302 B1.n23 B1.n22 185
R35303 B1.n69 B1.t1 120.037
R35304 B1.t2 B1.n14 120.037
R35305 B1.n59 B1.n57 112.831
R35306 B1.n22 B1.n21 112.831
R35307 B1.n68 B1.n67 104.172
R35308 B1.n27 B1.n26 104.172
R35309 B1.n68 B1.n56 92.5005
R35310 B1.n28 B1.n27 92.5005
R35311 B1.t1 B1.n68 66.8281
R35312 B1.n27 B1.t2 66.8281
R35313 B1.n6 B1.t6 35.2053
R35314 B1.n3 B1.t7 34.0571
R35315 B1.n67 B1.n66 29.4833
R35316 B1.n26 B1.n15 29.4833
R35317 B1.n1 B1.t3 27.6955
R35318 B1.n1 B1.t0 27.6955
R35319 B1.n45 B1.n44 19.0955
R35320 B1.n69 B1.n56 15.4558
R35321 B1.n28 B1.n14 15.4558
R35322 B1.n64 B1.n63 13.5534
R35323 B1.n23 B1.n18 13.5534
R35324 B1.n2 B1.n1 9.67857
R35325 B1.n41 B1.n34 9.30581
R35326 B1.n59 B1.n58 9.30424
R35327 B1.n21 B1.n20 9.30413
R35328 B1.n40 B1.n39 9.3005
R35329 B1.n46 B1.n45 9.3005
R35330 B1.n71 B1.n70 9.3005
R35331 B1.n55 B1.n52 9.3005
R35332 B1.n67 B1.n55 9.3005
R35333 B1.n63 B1.n62 9.3005
R35334 B1.n72 B1.n54 9.3005
R35335 B1.n29 B1.n13 9.3005
R35336 B1.n25 B1.n11 9.3005
R35337 B1.n26 B1.n25 9.3005
R35338 B1.n18 B1.n17 9.3005
R35339 B1.n31 B1.n30 9.3005
R35340 B1.n71 B1.n56 9.03579
R35341 B1.n29 B1.n28 9.03579
R35342 B1.n43 B1.n41 8.49366
R35343 B1.n43 B1.t4 8.2655
R35344 B1.n43 B1.t5 8.2655
R35345 B1.n44 B1.n43 7.97749
R35346 B1.n42 B1.n40 7.26743
R35347 B1.n43 B1.n42 6.15568
R35348 B1.n65 B1.n55 5.64756
R35349 B1.n25 B1.n24 5.64756
R35350 B1.n41 B1.n35 4.89462
R35351 B1.n60 B1.n59 4.89462
R35352 B1.n21 B1.n19 4.89462
R35353 B1.n73 B1.n55 4.51815
R35354 B1.n72 B1.n71 4.51815
R35355 B1.n25 B1.n12 4.51815
R35356 B1.n30 B1.n29 4.51815
R35357 B1.n5 B1.n4 4.5005
R35358 B1.n4 B1.n2 4.5005
R35359 B1.n51 B1.n9 4.5005
R35360 B1.n49 B1.n9 4.5005
R35361 B1.n51 B1.n50 4.5005
R35362 B1.n50 B1.n49 4.5005
R35363 B1.n74 B1.n53 4.5005
R35364 B1.n75 B1.n8 4.5005
R35365 B1.n53 B1.n8 4.5005
R35366 B1.n75 B1.n74 4.5005
R35367 B1.n48 B1.n32 4.5005
R35368 B1.n47 B1.n36 4.5005
R35369 B1.n48 B1.n47 4.5005
R35370 B1.n36 B1.n32 4.5005
R35371 B1.n38 B1.n33 4.5005
R35372 B1.n66 B1.n57 3.93153
R35373 B1.n22 B1.n15 3.93153
R35374 B1.n19 B1.n9 3.03311
R35375 B1.n50 B1.n12 3.03311
R35376 B1.n60 B1.n8 3.03311
R35377 B1.n74 B1.n73 3.03311
R35378 B1.n47 B1.n35 3.03311
R35379 B1.n3 B1.n0 2.2714
R35380 B1.n58 B1.n7 2.25261
R35381 B1.n20 B1.n10 2.25256
R35382 B1.n34 B1.n33 2.25127
R35383 B1.n37 B1.n33 2.24434
R35384 B1.n213 B1.n212 1.94045
R35385 B1.n86 B1.n85 1.94045
R35386 B1.n73 B1.n72 1.88285
R35387 B1.n30 B1.n12 1.88285
R35388 B1.n148 B1.n126 1.72426
R35389 B1.n131 B1.n130 1.7055
R35390 B1.n135 B1.n134 1.7055
R35391 B1.n139 B1.n138 1.7055
R35392 B1.n143 B1.n142 1.7055
R35393 B1.n147 B1.n146 1.7055
R35394 B1.n164 B1.n163 1.54412
R35395 B1.n45 B1.n35 1.50638
R35396 B1.n63 B1.n60 1.50638
R35397 B1.n19 B1.n18 1.50638
R35398 B1.n16 B1.n10 1.49213
R35399 B1.n70 B1.n69 1.49212
R35400 B1.n61 B1.n7 1.49182
R35401 B1.n14 B1.n13 1.49166
R35402 B1.n78 B1 1.05905
R35403 B1.n212 B1.n211 0.853
R35404 B1.n65 B1.n64 0.753441
R35405 B1.n24 B1.n23 0.753441
R35406 B1.n44 B1.n40 0.521921
R35407 B1.n181 B1.n180 0.513942
R35408 B1.n149 B1.n148 0.326891
R35409 B1.n77 B1.n6 0.29767
R35410 B1.n49 B1.n48 0.238951
R35411 B1.n77 B1.n76 0.196255
R35412 B1 B1.n77 0.1855
R35413 B1.n6 B1.n5 0.149538
R35414 B1.n75 B1.n51 0.124821
R35415 B1 B1.n216 0.0770766
R35416 B1.n126 B1 0.0686818
R35417 B1.n42 B1.n32 0.0579027
R35418 B1.n86 B1.n80 0.0511757
R35419 B1.n87 B1.n86 0.0511757
R35420 B1.n213 B1.n100 0.0511757
R35421 B1.n214 B1.n213 0.0511757
R35422 B1.n62 B1.n61 0.0396286
R35423 B1.n90 B1.n89 0.0387883
R35424 B1.n94 B1.n93 0.0387883
R35425 B1.n98 B1.n97 0.0387883
R35426 B1.n17 B1.n16 0.0383668
R35427 B1.n85 B1.n84 0.0323396
R35428 B1.n212 B1.n121 0.0323396
R35429 B1.n212 B1.n125 0.0323396
R35430 B1.n46 B1.n37 0.0314092
R35431 B1.n5 B1.n0 0.0281442
R35432 B1.n39 B1.n37 0.0271357
R35433 B1.n83 B1.n82 0.0229057
R35434 B1.n103 B1.n102 0.0229057
R35435 B1.n120 B1.n119 0.0229057
R35436 B1.n124 B1.n123 0.0229057
R35437 B1.n80 B1.n79 0.0218964
R35438 B1.n88 B1.n87 0.0218964
R35439 B1.n100 B1.n99 0.0218964
R35440 B1.n215 B1.n214 0.0218964
R35441 B1.n84 B1.n83 0.0217264
R35442 B1.n102 B1.n101 0.0217264
R35443 B1.n121 B1.n120 0.0217264
R35444 B1.n125 B1.n124 0.0217264
R35445 B1.n111 B1.n110 0.0205472
R35446 B1.n112 B1.n111 0.0205472
R35447 B1.n148 B1.n147 0.0203537
R35448 B1.n61 B1.n52 0.0202788
R35449 B1.n16 B1.n11 0.0196501
R35450 B1.n106 B1.n105 0.0193679
R35451 B1.n117 B1.n116 0.0193679
R35452 B1.n182 B1.n181 0.0189241
R35453 B1.n108 B1.n107 0.0181887
R35454 B1.n110 B1.n109 0.0181887
R35455 B1.n113 B1.n112 0.0181887
R35456 B1.n115 B1.n114 0.0181887
R35457 B1.n91 B1.n90 0.0173919
R35458 B1.n93 B1.n92 0.0173919
R35459 B1.n95 B1.n94 0.0173919
R35460 B1.n97 B1.n96 0.0173919
R35461 B1.n163 B1.n162 0.0169458
R35462 B1.n51 B1.n10 0.0168043
R35463 B1.n36 B1.n33 0.016125
R35464 B1.n128 B1.n127 0.0138019
R35465 B1.n131 B1.n129 0.0138019
R35466 B1.n132 B1.n131 0.0138019
R35467 B1.n135 B1.n133 0.0138019
R35468 B1.n136 B1.n135 0.0138019
R35469 B1.n139 B1.n137 0.0138019
R35470 B1.n140 B1.n139 0.0138019
R35471 B1.n143 B1.n141 0.0138019
R35472 B1.n144 B1.n143 0.0138019
R35473 B1.n147 B1.n145 0.0138019
R35474 B1.n180 B1.n179 0.0138019
R35475 B1.n178 B1.n177 0.0138019
R35476 B1.n177 B1.n176 0.0138019
R35477 B1.n175 B1.n174 0.0138019
R35478 B1.n174 B1.n173 0.0138019
R35479 B1.n172 B1.n171 0.0138019
R35480 B1.n171 B1.n170 0.0138019
R35481 B1.n169 B1.n168 0.0138019
R35482 B1.n168 B1.n167 0.0138019
R35483 B1.n166 B1.n165 0.0138019
R35484 B1.n165 B1.n164 0.0138019
R35485 B1.n161 B1.n160 0.0138019
R35486 B1.n160 B1.n159 0.0138019
R35487 B1.n158 B1.n157 0.0138019
R35488 B1.n157 B1.n156 0.0138019
R35489 B1.n155 B1.n154 0.0138019
R35490 B1.n154 B1.n153 0.0138019
R35491 B1.n152 B1.n151 0.0138019
R35492 B1.n151 B1.n150 0.0138019
R35493 B1.n74 B1.n52 0.013431
R35494 B1.n70 B1.n54 0.013431
R35495 B1.n50 B1.n11 0.013
R35496 B1.n31 B1.n13 0.013
R35497 B1.n183 B1.n182 0.0124717
R35498 B1.n184 B1.n183 0.0124717
R35499 B1.n211 B1.n204 0.0124717
R35500 B1.n211 B1.n210 0.0124717
R35501 B1.n38 B1.n32 0.0122521
R35502 B1.n58 B1.n8 0.0117689
R35503 B1.n20 B1.n9 0.0114102
R35504 B1.n105 B1.n104 0.0111132
R35505 B1.n107 B1.n106 0.0111132
R35506 B1.n116 B1.n115 0.0111132
R35507 B1.n118 B1.n117 0.0111132
R35508 B1.n47 B1.n34 0.0100704
R35509 B1.n76 B1.n7 0.0100109
R35510 B1.n109 B1.n108 0.00993396
R35511 B1.n114 B1.n113 0.00993396
R35512 B1.n187 B1.n186 0.00981132
R35513 B1.n202 B1.n201 0.00981132
R35514 B1.n208 B1.n207 0.00981132
R35515 B1.n92 B1.n91 0.00950901
R35516 B1.n96 B1.n95 0.00950901
R35517 B1.n129 B1.n128 0.00936793
R35518 B1.n133 B1.n132 0.00936793
R35519 B1.n137 B1.n136 0.00936793
R35520 B1.n141 B1.n140 0.00936793
R35521 B1.n145 B1.n144 0.00936793
R35522 B1.n186 B1.n185 0.00936793
R35523 B1.n192 B1.n191 0.00936793
R35524 B1.n197 B1.n196 0.00936793
R35525 B1.n203 B1.n202 0.00936793
R35526 B1.n209 B1.n208 0.00936793
R35527 B1.n179 B1.n178 0.00936793
R35528 B1.n176 B1.n175 0.00936793
R35529 B1.n173 B1.n172 0.00936793
R35530 B1.n170 B1.n169 0.00936793
R35531 B1.n167 B1.n166 0.00936793
R35532 B1.n162 B1.n161 0.00936793
R35533 B1.n159 B1.n158 0.00936793
R35534 B1.n156 B1.n155 0.00936793
R35535 B1.n153 B1.n152 0.00936793
R35536 B1.n150 B1.n149 0.00936793
R35537 B1.n82 B1.n81 0.00875472
R35538 B1.n104 B1.n103 0.00875472
R35539 B1.n119 B1.n118 0.00875472
R35540 B1.n123 B1.n122 0.00875472
R35541 B1.n79 B1.n78 0.00838288
R35542 B1.n89 B1.n88 0.00838288
R35543 B1.n99 B1.n98 0.00838288
R35544 B1.n216 B1.n215 0.00838288
R35545 B1.n194 B1.n193 0.00803774
R35546 B1.n195 B1.n194 0.00803774
R35547 B1.n189 B1.n188 0.00759434
R35548 B1.n200 B1.n199 0.00759434
R35549 B1.n193 B1.n192 0.00626415
R35550 B1.n196 B1.n195 0.00626415
R35551 B1.n74 B1.n54 0.00588793
R35552 B1.n50 B1.n31 0.00570833
R35553 B1.n206 B1.n205 0.00519331
R35554 B1.n62 B1.n8 0.00481034
R35555 B1.n47 B1.n46 0.0047735
R35556 B1.n17 B1.n9 0.00466667
R35557 B1.n53 B1.n7 0.00457609
R35558 B1.n76 B1.n75 0.00457609
R35559 B1.n188 B1.n187 0.00449057
R35560 B1.n190 B1.n189 0.00449057
R35561 B1.n199 B1.n198 0.00449057
R35562 B1.n201 B1.n200 0.00449057
R35563 B1.n207 B1.n206 0.00449057
R35564 B1.n2 B1.n0 0.00410577
R35565 B1.n39 B1.n38 0.00370513
R35566 B1.n191 B1.n190 0.00271698
R35567 B1.n198 B1.n197 0.00271698
R35568 B1.n48 B1.n33 0.00253804
R35569 B1.n4 B1.n3 0.00185919
R35570 B1.n49 B1.n10 0.0018587
R35571 B1.n185 B1.n184 0.00183019
R35572 B1.n204 B1.n203 0.00183019
R35573 B1.n210 B1.n209 0.00183019
R35574 a_10204_n3484.n5 a_10204_n3484.t3 136.804
R35575 a_10204_n3484.n5 a_10204_n3484.t9 136.325
R35576 a_10204_n3484.n20 a_10204_n3484.t2 119.999
R35577 a_10204_n3484.n11 a_10204_n3484.t7 93.9023
R35578 a_10204_n3484.n0 a_10204_n3484.t4 93.3044
R35579 a_10204_n3484.n0 a_10204_n3484.t8 93.0848
R35580 a_10204_n3484.n19 a_10204_n3484.n18 92.5005
R35581 a_10204_n3484.n12 a_10204_n3484.t5 92.4623
R35582 a_10204_n3484.n0 a_10204_n3484.t6 69.2281
R35583 a_10204_n3484.n27 a_10204_n3484.n26 29.4833
R35584 a_10204_n3484.n15 a_10204_n3484.t0 27.6955
R35585 a_10204_n3484.t1 a_10204_n3484.n46 27.6955
R35586 a_10204_n3484.n20 a_10204_n3484.n19 15.4626
R35587 a_10204_n3484.n2 a_10204_n3484.n30 9.3005
R35588 a_10204_n3484.n2 a_10204_n3484.n22 9.3005
R35589 a_10204_n3484.n2 a_10204_n3484.n21 9.3005
R35590 a_10204_n3484.n2 a_10204_n3484.n28 9.3005
R35591 a_10204_n3484.n28 a_10204_n3484.n27 9.3005
R35592 a_10204_n3484.n2 a_10204_n3484.n29 9.3005
R35593 a_10204_n3484.n2 a_10204_n3484.n31 9.3005
R35594 a_10204_n3484.n46 a_10204_n3484.n45 9.02061
R35595 a_10204_n3484.n46 a_10204_n3484.n41 9.02061
R35596 a_10204_n3484.n16 a_10204_n3484.n15 9.01961
R35597 a_10204_n3484.n35 a_10204_n3484.n33 8.28285
R35598 a_10204_n3484.n3 a_10204_n3484.n8 8.28285
R35599 a_10204_n3484.n28 a_10204_n3484.n24 5.64756
R35600 a_10204_n3484.n1 a_10204_n3484.n35 5.32328
R35601 a_10204_n3484.n13 a_10204_n3484.n17 4.14168
R35602 a_10204_n3484.n40 a_10204_n3484.n7 4.14168
R35603 a_10204_n3484.n1 a_10204_n3484.n12 4.06959
R35604 a_10204_n3484.n26 a_10204_n3484.n25 3.93153
R35605 a_10204_n3484.n38 a_10204_n3484.n36 3.76521
R35606 a_10204_n3484.n44 a_10204_n3484.n43 3.76521
R35607 a_10204_n3484.n35 a_10204_n3484.n34 3.38874
R35608 a_10204_n3484.n4 a_10204_n3484.n3 3.11016
R35609 a_10204_n3484.n14 a_10204_n3484.n13 3.07321
R35610 a_10204_n3484.n39 a_10204_n3484.n38 3.04543
R35611 a_10204_n3484.n40 a_10204_n3484.n4 3.03311
R35612 a_10204_n3484.n4 a_10204_n3484.n9 3.03311
R35613 a_10204_n3484.n38 a_10204_n3484.n37 2.63579
R35614 a_10204_n3484.n45 a_10204_n3484.n44 2.63579
R35615 a_10204_n3484.n4 a_10204_n3484.n1 2.43716
R35616 a_10204_n3484.n1 a_10204_n3484.n14 2.36361
R35617 a_10204_n3484.n1 a_10204_n3484.n39 2.27338
R35618 a_10204_n3484.n13 a_10204_n3484.n16 2.25932
R35619 a_10204_n3484.n41 a_10204_n3484.n40 2.25932
R35620 a_10204_n3484.n12 a_10204_n3484.n11 1.80772
R35621 a_10204_n3484.n5 a_10204_n3484.n10 1.61433
R35622 a_10204_n3484.n2 a_10204_n3484.n20 1.45534
R35623 a_10204_n3484.n11 a_10204_n3484.n5 1.19419
R35624 a_10204_n3484.n32 a_10204_n3484.n2 1.14499
R35625 a_10204_n3484.n43 a_10204_n3484.n42 1.12991
R35626 a_10204_n3484.n7 a_10204_n3484.n6 1.12991
R35627 a_10204_n3484.n32 a_10204_n3484.n0 1.12005
R35628 a_10204_n3484.n14 a_10204_n3484.n32 0.839613
R35629 a_10204_n3484.n24 a_10204_n3484.n23 0.753441
R35630 a_1425_9823.n79 a_1425_9823.t9 60.2505
R35631 a_1425_9823.n57 a_1425_9823.t6 60.2505
R35632 a_1425_9823.n43 a_1425_9823.t8 60.2505
R35633 a_1425_9823.n21 a_1425_9823.t7 60.2505
R35634 a_1425_9823.n0 a_1425_9823.n131 9.3005
R35635 a_1425_9823.n0 a_1425_9823.n129 9.3005
R35636 a_1425_9823.n4 a_1425_9823.n65 9.3005
R35637 a_1425_9823.n4 a_1425_9823.n66 9.3005
R35638 a_1425_9823.n4 a_1425_9823.n64 9.3005
R35639 a_1425_9823.n64 a_1425_9823.n63 9.3005
R35640 a_1425_9823.n5 a_1425_9823.n72 9.3005
R35641 a_1425_9823.n6 a_1425_9823.n89 9.3005
R35642 a_1425_9823.n5 a_1425_9823.n78 9.3005
R35643 a_1425_9823.n78 a_1425_9823.n77 9.3005
R35644 a_1425_9823.n5 a_1425_9823.n71 9.3005
R35645 a_1425_9823.n6 a_1425_9823.n87 9.3005
R35646 a_1425_9823.n87 a_1425_9823.n86 9.3005
R35647 a_1425_9823.n6 a_1425_9823.n88 9.3005
R35648 a_1425_9823.n3 a_1425_9823.n29 9.3005
R35649 a_1425_9823.n3 a_1425_9823.n30 9.3005
R35650 a_1425_9823.n3 a_1425_9823.n28 9.3005
R35651 a_1425_9823.n28 a_1425_9823.n27 9.3005
R35652 a_1425_9823.n2 a_1425_9823.n36 9.3005
R35653 a_1425_9823.n2 a_1425_9823.n42 9.3005
R35654 a_1425_9823.n42 a_1425_9823.n41 9.3005
R35655 a_1425_9823.n2 a_1425_9823.n35 9.3005
R35656 a_1425_9823.n1 a_1425_9823.n51 9.3005
R35657 a_1425_9823.n51 a_1425_9823.n50 9.3005
R35658 a_1425_9823.n1 a_1425_9823.n53 9.3005
R35659 a_1425_9823.n1 a_1425_9823.n52 9.3005
R35660 a_1425_9823.n8 a_1425_9823.n19 9.3005
R35661 a_1425_9823.n7 a_1425_9823.n14 9.3005
R35662 a_1425_9823.n162 a_1425_9823.n159 9.3005
R35663 a_1425_9823.n162 a_1425_9823.n160 9.3005
R35664 a_1425_9823.n80 a_1425_9823.n79 8.76429
R35665 a_1425_9823.n44 a_1425_9823.n43 8.76429
R35666 a_1425_9823.n85 a_1425_9823.n84 7.45411
R35667 a_1425_9823.n76 a_1425_9823.n75 7.45411
R35668 a_1425_9823.n62 a_1425_9823.n61 7.45411
R35669 a_1425_9823.n40 a_1425_9823.n39 7.45411
R35670 a_1425_9823.n49 a_1425_9823.n48 7.45411
R35671 a_1425_9823.n26 a_1425_9823.n25 7.45411
R35672 a_1425_9823.n58 a_1425_9823.n57 6.80105
R35673 a_1425_9823.n22 a_1425_9823.n21 6.80105
R35674 a_1425_9823.n83 a_1425_9823.n82 5.64756
R35675 a_1425_9823.n74 a_1425_9823.n73 5.64756
R35676 a_1425_9823.n60 a_1425_9823.n59 5.64756
R35677 a_1425_9823.n38 a_1425_9823.n37 5.64756
R35678 a_1425_9823.n47 a_1425_9823.n46 5.64756
R35679 a_1425_9823.n24 a_1425_9823.n23 5.64756
R35680 a_1425_9823.n112 a_1425_9823.t3 5.5395
R35681 a_1425_9823.n112 a_1425_9823.t2 5.5395
R35682 a_1425_9823.n162 a_1425_9823.t1 5.5395
R35683 a_1425_9823.t4 a_1425_9823.n162 5.5395
R35684 a_1425_9823.n70 a_1425_9823.n69 4.73575
R35685 a_1425_9823.n68 a_1425_9823.n67 4.73575
R35686 a_1425_9823.n34 a_1425_9823.n33 4.73575
R35687 a_1425_9823.n32 a_1425_9823.n31 4.73575
R35688 a_1425_9823.n81 a_1425_9823.n80 4.6505
R35689 a_1425_9823.n45 a_1425_9823.n44 4.6505
R35690 a_1425_9823.n135 a_1425_9823.n134 4.51815
R35691 a_1425_9823.n17 a_1425_9823.n16 4.51815
R35692 a_1425_9823.n155 a_1425_9823.n154 4.51815
R35693 a_1425_9823.n0 a_1425_9823.n128 4.5005
R35694 a_1425_9823.n124 a_1425_9823.n133 4.5005
R35695 a_1425_9823.n125 a_1425_9823.n123 4.5005
R35696 a_1425_9823.n118 a_1425_9823.n116 4.5005
R35697 a_1425_9823.n8 a_1425_9823.n12 4.5005
R35698 a_1425_9823.n7 a_1425_9823.n17 4.5005
R35699 a_1425_9823.n102 a_1425_9823.n107 4.5005
R35700 a_1425_9823.n139 a_1425_9823.n147 4.5005
R35701 a_1425_9823.n152 a_1425_9823.n151 4.5005
R35702 a_1425_9823.n138 a_1425_9823.n141 4.5005
R35703 a_1425_9823.n162 a_1425_9823.n161 4.35791
R35704 a_1425_9823.n91 a_1425_9823.n93 4.24504
R35705 a_1425_9823.n54 a_1425_9823.n56 4.24504
R35706 a_1425_9823.n12 a_1425_9823.n11 3.76521
R35707 a_1425_9823.n4 a_1425_9823.n58 3.42768
R35708 a_1425_9823.n3 a_1425_9823.n22 3.42768
R35709 a_1425_9823.n123 a_1425_9823.n119 3.38874
R35710 a_1425_9823.n147 a_1425_9823.n144 3.38874
R35711 a_1425_9823.n131 a_1425_9823.n130 3.38537
R35712 a_1425_9823.n158 a_1425_9823.n157 3.38537
R35713 a_1425_9823.n97 a_1425_9823.t0 3.3065
R35714 a_1425_9823.n97 a_1425_9823.t5 3.3065
R35715 a_1425_9823.n107 a_1425_9823.n105 3.28194
R35716 a_1425_9823.n99 a_1425_9823.n98 3.15821
R35717 a_1425_9823.n117 a_1425_9823.n135 3.03311
R35718 a_1425_9823.n153 a_1425_9823.n155 3.03311
R35719 a_1425_9823.n107 a_1425_9823.n106 3.01226
R35720 a_1425_9823.n12 a_1425_9823.n10 2.63579
R35721 a_1425_9823.n14 a_1425_9823.n13 2.61733
R35722 a_1425_9823.n0 a_1425_9823.n126 2.57914
R35723 a_1425_9823.n122 a_1425_9823.n121 2.25932
R35724 a_1425_9823.n146 a_1425_9823.n145 2.25932
R35725 a_1425_9823.n19 a_1425_9823.n18 2.24766
R35726 a_1425_9823.n116 a_1425_9823.n114 2.22452
R35727 a_1425_9823.n151 a_1425_9823.n149 2.22452
R35728 a_1425_9823.n162 a_1425_9823.n148 1.99078
R35729 a_1425_9823.n17 a_1425_9823.n15 1.88285
R35730 a_1425_9823.n113 a_1425_9823.n112 1.72048
R35731 a_1425_9823.n99 a_1425_9823.n97 1.61799
R35732 a_1425_9823.n108 a_1425_9823.n96 1.51434
R35733 a_1425_9823.n96 a_1425_9823.n8 1.51334
R35734 a_1425_9823.n128 a_1425_9823.n127 1.50638
R35735 a_1425_9823.n159 a_1425_9823.n158 1.50638
R35736 a_1425_9823.n142 a_1425_9823.n143 1.50638
R35737 a_1425_9823.n101 a_1425_9823.n100 1.12991
R35738 a_1425_9823.n95 a_1425_9823.n94 3.28829
R35739 a_1425_9823.n86 a_1425_9823.n85 0.994314
R35740 a_1425_9823.n77 a_1425_9823.n76 0.994314
R35741 a_1425_9823.n63 a_1425_9823.n62 0.994314
R35742 a_1425_9823.n41 a_1425_9823.n40 0.994314
R35743 a_1425_9823.n50 a_1425_9823.n49 0.994314
R35744 a_1425_9823.n27 a_1425_9823.n26 0.994314
R35745 a_1425_9823.n111 a_1425_9823.n156 0.829361
R35746 a_1425_9823.n133 a_1425_9823.n132 0.753441
R35747 a_1425_9823.n87 a_1425_9823.n83 0.753441
R35748 a_1425_9823.n78 a_1425_9823.n74 0.753441
R35749 a_1425_9823.n64 a_1425_9823.n60 0.753441
R35750 a_1425_9823.n42 a_1425_9823.n38 0.753441
R35751 a_1425_9823.n51 a_1425_9823.n47 0.753441
R35752 a_1425_9823.n28 a_1425_9823.n24 0.753441
R35753 a_1425_9823.n141 a_1425_9823.n140 0.753441
R35754 a_1425_9823.n137 a_1425_9823.n136 0.754708
R35755 a_1425_9823.n93 a_1425_9823.n92 0.709906
R35756 a_1425_9823.n56 a_1425_9823.n55 0.709906
R35757 a_1425_9823.n109 a_1425_9823.n137 0.678625
R35758 a_1425_9823.n70 a_1425_9823.n68 0.458354
R35759 a_1425_9823.n34 a_1425_9823.n32 0.458354
R35760 a_1425_9823.n123 a_1425_9823.n122 0.376971
R35761 a_1425_9823.n121 a_1425_9823.n120 0.376971
R35762 a_1425_9823.n104 a_1425_9823.n103 0.376971
R35763 a_1425_9823.n147 a_1425_9823.n146 0.376971
R35764 a_1425_9823.n95 a_1425_9823.n20 0.242354
R35765 a_1425_9823.n136 a_1425_9823.n113 0.225683
R35766 a_1425_9823.n108 a_1425_9823.n99 0.224119
R35767 a_1425_9823.n6 a_1425_9823.n81 0.190717
R35768 a_1425_9823.n81 a_1425_9823.n5 0.190717
R35769 a_1425_9823.n45 a_1425_9823.n2 0.190717
R35770 a_1425_9823.n1 a_1425_9823.n45 0.190717
R35771 a_1425_9823.n94 a_1425_9823.n54 0.159981
R35772 a_1425_9823.n94 a_1425_9823.n91 0.159717
R35773 a_1425_9823.n138 a_1425_9823.n142 4.63429
R35774 a_1425_9823.n105 a_1425_9823.n104 0.0902327
R35775 a_1425_9823.n117 a_1425_9823.n125 0.0900802
R35776 a_1425_9823.n136 a_1425_9823.n118 0.0608541
R35777 a_1425_9823.n111 a_1425_9823.n110 0.0528649
R35778 a_1425_9823.n156 a_1425_9823.n153 0.0511262
R35779 a_1425_9823.n156 a_1425_9823.n139 0.040511
R35780 a_1425_9823.n114 a_1425_9823.n115 0.0303633
R35781 a_1425_9823.n149 a_1425_9823.n150 0.0303633
R35782 a_1425_9823.n102 a_1425_9823.n101 4.54542
R35783 a_1425_9823.n152 a_1425_9823.n148 0.0122188
R35784 a_1425_9823.n153 a_1425_9823.n152 0.0454219
R35785 a_1425_9823.n139 a_1425_9823.n138 0.0454219
R35786 a_1425_9823.n118 a_1425_9823.n117 0.0454219
R35787 a_1425_9823.n125 a_1425_9823.n124 0.0454219
R35788 a_1425_9823.n111 a_1425_9823.n109 0.022561
R35789 a_1425_9823.n111 a_1425_9823.n20 0.847626
R35790 a_1425_9823.n108 a_1425_9823.n102 0.0883906
R35791 a_1425_9823.n96 a_1425_9823.n95 0.905839
R35792 a_1425_9823.n91 a_1425_9823.n90 0.0410417
R35793 a_1425_9823.n8 a_1425_9823.n9 2.77239
R35794 a_1425_9823.n5 a_1425_9823.n70 0.205546
R35795 a_1425_9823.n68 a_1425_9823.n4 0.205546
R35796 a_1425_9823.n32 a_1425_9823.n3 0.205546
R35797 a_1425_9823.n2 a_1425_9823.n34 0.205546
R35798 a_1425_9823.n54 a_1425_9823.n1 0.177485
R35799 a_1425_9823.n124 a_1425_9823.n0 0.171838
R35800 a_1425_9823.n8 a_1425_9823.n7 0.167464
R35801 a_1425_9823.n90 a_1425_9823.n6 0.137941
R35802 B2.n101 B2.n100 185
R35803 B2.n99 B2.n92 185
R35804 B2.n59 B2.n50 185
R35805 B2.n58 B2.n57 185
R35806 B2.n104 B2.t4 120.037
R35807 B2.t5 B2.n49 120.037
R35808 B2.n94 B2.n92 112.831
R35809 B2.n57 B2.n56 112.831
R35810 B2.n103 B2.n102 104.172
R35811 B2.n62 B2.n61 104.172
R35812 B2.n103 B2.n91 92.5005
R35813 B2.n63 B2.n62 92.5005
R35814 B2.t4 B2.n103 66.8281
R35815 B2.n62 B2.t5 66.8281
R35816 B2.n41 B2.t0 35.2053
R35817 B2.n38 B2.t1 34.0571
R35818 B2.n102 B2.n101 29.4833
R35819 B2.n61 B2.n50 29.4833
R35820 B2.n36 B2.t6 27.6955
R35821 B2.n36 B2.t7 27.6955
R35822 B2.n80 B2.n79 19.0955
R35823 B2.n104 B2.n91 15.4558
R35824 B2.n63 B2.n49 15.4558
R35825 B2.n99 B2.n98 13.5534
R35826 B2.n58 B2.n53 13.5534
R35827 B2.n37 B2.n36 9.67857
R35828 B2.n76 B2.n69 9.30581
R35829 B2.n94 B2.n93 9.30424
R35830 B2.n56 B2.n55 9.30413
R35831 B2.n75 B2.n74 9.3005
R35832 B2.n81 B2.n80 9.3005
R35833 B2.n106 B2.n105 9.3005
R35834 B2.n90 B2.n87 9.3005
R35835 B2.n102 B2.n90 9.3005
R35836 B2.n98 B2.n97 9.3005
R35837 B2.n107 B2.n89 9.3005
R35838 B2.n64 B2.n48 9.3005
R35839 B2.n60 B2.n46 9.3005
R35840 B2.n61 B2.n60 9.3005
R35841 B2.n53 B2.n52 9.3005
R35842 B2.n66 B2.n65 9.3005
R35843 B2.n106 B2.n91 9.03579
R35844 B2.n64 B2.n63 9.03579
R35845 B2.n78 B2.n76 8.49366
R35846 B2.n78 B2.t2 8.2655
R35847 B2.n78 B2.t3 8.2655
R35848 B2.n79 B2.n78 7.97749
R35849 B2.n77 B2.n75 7.26743
R35850 B2.n78 B2.n77 6.15568
R35851 B2.n100 B2.n90 5.64756
R35852 B2.n60 B2.n59 5.64756
R35853 B2.n76 B2.n70 4.89462
R35854 B2.n95 B2.n94 4.89462
R35855 B2.n56 B2.n54 4.89462
R35856 B2.n108 B2.n90 4.51815
R35857 B2.n107 B2.n106 4.51815
R35858 B2.n60 B2.n47 4.51815
R35859 B2.n65 B2.n64 4.51815
R35860 B2.n40 B2.n39 4.5005
R35861 B2.n39 B2.n37 4.5005
R35862 B2.n86 B2.n44 4.5005
R35863 B2.n84 B2.n44 4.5005
R35864 B2.n86 B2.n85 4.5005
R35865 B2.n85 B2.n84 4.5005
R35866 B2.n109 B2.n88 4.5005
R35867 B2.n110 B2.n43 4.5005
R35868 B2.n88 B2.n43 4.5005
R35869 B2.n110 B2.n109 4.5005
R35870 B2.n83 B2.n67 4.5005
R35871 B2.n82 B2.n71 4.5005
R35872 B2.n83 B2.n82 4.5005
R35873 B2.n71 B2.n67 4.5005
R35874 B2.n73 B2.n68 4.5005
R35875 B2.n114 B2.n34 4.5005
R35876 B2.n127 B2.n28 4.5005
R35877 B2.n139 B2.n138 4.5005
R35878 B2.n141 B2.n20 4.5005
R35879 B2.n8 B2.n7 4.5005
R35880 B2.n167 B2.n166 4.5005
R35881 B2.n164 B2.n163 4.5005
R35882 B2.n137 B2.n21 4.5005
R35883 B2.n126 B2.n125 4.5005
R35884 B2.n116 B2.n115 4.5005
R35885 B2.n15 B2.n14 4.5005
R35886 B2.n1 B2.n0 4.5005
R35887 B2.n101 B2.n92 3.93153
R35888 B2.n57 B2.n50 3.93153
R35889 B2.n211 B2.n2 3.4201
R35890 B2.n152 B2.n151 3.4105
R35891 B2.n154 B2.n153 3.4105
R35892 B2.n24 B2.n22 3.4105
R35893 B2.n136 B2.n23 3.4105
R35894 B2.n124 B2.n123 3.4105
R35895 B2.n113 B2.n33 3.4105
R35896 B2.n118 B2.n117 3.4105
R35897 B2.n129 B2.n128 3.4105
R35898 B2.n140 B2.n19 3.4105
R35899 B2.n143 B2.n142 3.4105
R35900 B2.n13 B2.n11 3.4105
R35901 B2.n162 B2.n161 3.4105
R35902 B2.n169 B2.n168 3.4105
R35903 B2.n216 B2.n215 3.4105
R35904 B2.n172 B2.n3 3.4105
R35905 B2.n122 B2.n121 3.4105
R35906 B2.n32 B2.n26 3.4105
R35907 B2.n134 B2.n133 3.4105
R35908 B2.n25 B2.n17 3.4105
R35909 B2.n148 B2.n147 3.4105
R35910 B2.n149 B2.n10 3.4105
R35911 B2.n158 B2.n9 3.4105
R35912 B2.n160 B2.n159 3.4105
R35913 B2.n171 B2.n170 3.4105
R35914 B2.n131 B2.n130 3.4105
R35915 B2.n156 B2.n155 3.4105
R35916 B2.n190 B2.n185 3.4105
R35917 B2.n208 B2.n173 3.4105
R35918 B2.n207 B2.n206 3.4105
R35919 B2.n204 B2.n203 3.4105
R35920 B2.n202 B2.n176 3.4105
R35921 B2.n182 B2.n177 3.4105
R35922 B2.n183 B2.n180 3.4105
R35923 B2.n196 B2.n181 3.4105
R35924 B2.n195 B2.n194 3.4105
R35925 B2.n192 B2.n191 3.4105
R35926 B2.n54 B2.n44 3.03311
R35927 B2.n85 B2.n47 3.03311
R35928 B2.n95 B2.n43 3.03311
R35929 B2.n109 B2.n108 3.03311
R35930 B2.n82 B2.n70 3.03311
R35931 B2.n38 B2.n35 2.2714
R35932 B2.n93 B2.n42 2.25261
R35933 B2.n55 B2.n45 2.25256
R35934 B2.n69 B2.n68 2.25127
R35935 B2.n72 B2.n68 2.24434
R35936 B2.n165 B2.n6 1.94045
R35937 B2.n30 B2.n29 1.94045
R35938 B2.n108 B2.n107 1.88285
R35939 B2.n65 B2.n47 1.88285
R35940 B2.n209 B2.n174 1.79984
R35941 B2.n189 B2.n186 1.72491
R35942 B2.n215 B2.n2 1.72009
R35943 B2.n145 B2.n144 1.7055
R35944 B2.n175 B2.n174 1.7055
R35945 B2.n201 B2.n200 1.7055
R35946 B2.n199 B2.n198 1.7055
R35947 B2.n193 B2.n179 1.7055
R35948 B2.n188 B2.n187 1.7055
R35949 B2.n217 B2 1.563
R35950 B2.n217 B2 1.563
R35951 B2.n211 B2.n210 1.54227
R35952 B2.n80 B2.n70 1.50638
R35953 B2.n98 B2.n95 1.50638
R35954 B2.n54 B2.n53 1.50638
R35955 B2.n51 B2.n45 1.49213
R35956 B2.n105 B2.n104 1.49212
R35957 B2.n96 B2.n42 1.49182
R35958 B2.n49 B2.n48 1.49166
R35959 B2.n215 B2.n214 1.13717
R35960 B2.n151 B2.n150 1.13717
R35961 B2.n154 B2.n12 1.13717
R35962 B2.n129 B2.n27 1.13717
R35963 B2.n136 B2.n135 1.13717
R35964 B2.n19 B2.n18 1.13717
R35965 B2.n143 B2.n16 1.13717
R35966 B2.n113 B2 1.06286
R35967 B2.n120 B2.n31 0.853
R35968 B2.n31 B2.n30 0.853
R35969 B2.n132 B2.n131 0.853
R35970 B2.n146 B2.n145 0.853
R35971 B2.n157 B2.n156 0.853
R35972 B2.n6 B2.n5 0.853
R35973 B2.n5 B2.n4 0.853
R35974 B2.n213 B2.n212 0.853
R35975 B2.n205 B2.n175 0.853
R35976 B2.n201 B2.n178 0.853
R35977 B2.n198 B2.n197 0.853
R35978 B2.n193 B2.n184 0.853
R35979 B2.n100 B2.n99 0.753441
R35980 B2.n59 B2.n58 0.753441
R35981 B2.n119 B2.n33 0.690775
R35982 B2.n210 B2.n209 0.681308
R35983 B2.n79 B2.n75 0.521921
R35984 B2.n120 B2.n119 0.513942
R35985 B2.n190 B2.n189 0.32799
R35986 B2.n112 B2.n41 0.29767
R35987 B2.n84 B2.n83 0.238951
R35988 B2.n112 B2.n111 0.196255
R35989 B2 B2.n112 0.1855
R35990 B2.n41 B2.n40 0.149538
R35991 B2.n110 B2.n86 0.124821
R35992 B2.n200 B2.n174 0.0948396
R35993 B2.n200 B2.n199 0.0948396
R35994 B2.n199 B2.n179 0.0948396
R35995 B2.n187 B2.n179 0.0948396
R35996 B2.n187 B2.n186 0.0948396
R35997 B2.n217 B2.n216 0.0784817
R35998 B2.n186 B2 0.0783302
R35999 B2.n77 B2.n67 0.0579027
R36000 B2.n115 B2.n29 0.0521055
R36001 B2.n126 B2.n29 0.0521055
R36002 B2.n165 B2.n164 0.0521055
R36003 B2.n166 B2.n165 0.0521055
R36004 B2.n97 B2.n96 0.0396286
R36005 B2.n128 B2.n23 0.0394908
R36006 B2.n142 B2.n140 0.0394908
R36007 B2.n153 B2.n152 0.0394908
R36008 B2.n52 B2.n51 0.0383668
R36009 B2.n117 B2.n30 0.0323396
R36010 B2.n124 B2.n30 0.0323396
R36011 B2.n162 B2.n6 0.0323396
R36012 B2.n168 B2.n6 0.0323396
R36013 B2.n81 B2.n72 0.0314092
R36014 B2.n40 B2.n35 0.0281442
R36015 B2.n74 B2.n72 0.0271357
R36016 B2.n116 B2.n34 0.0229057
R36017 B2.n125 B2.n28 0.0229057
R36018 B2.n163 B2.n8 0.0229057
R36019 B2.n167 B2.n1 0.0229057
R36020 B2.n115 B2.n114 0.022289
R36021 B2.n127 B2.n126 0.022289
R36022 B2.n164 B2.n7 0.022289
R36023 B2.n166 B2.n0 0.022289
R36024 B2.n117 B2.n116 0.0217264
R36025 B2.n125 B2.n124 0.0217264
R36026 B2.n163 B2.n162 0.0217264
R36027 B2.n168 B2.n167 0.0217264
R36028 B2.n189 B2.n188 0.0210321
R36029 B2.n144 B2.n19 0.0205472
R36030 B2.n144 B2.n143 0.0205472
R36031 B2.n96 B2.n87 0.0202788
R36032 B2.n51 B2.n46 0.0196501
R36033 B2.n130 B2.n22 0.0193679
R36034 B2.n155 B2.n13 0.0193679
R36035 B2.n119 B2.n118 0.0189241
R36036 B2.n137 B2.n136 0.0181887
R36037 B2.n138 B2.n19 0.0181887
R36038 B2.n143 B2.n20 0.0181887
R36039 B2.n151 B2.n15 0.0181887
R36040 B2.n210 B2.n173 0.0179016
R36041 B2.n23 B2.n21 0.0177018
R36042 B2.n140 B2.n139 0.0177018
R36043 B2.n142 B2.n141 0.0177018
R36044 B2.n152 B2.n14 0.0177018
R36045 B2.n86 B2.n45 0.0168043
R36046 B2.n71 B2.n68 0.016125
R36047 B2.n206 B2.n205 0.0146
R36048 B2.n205 B2.n204 0.0146
R36049 B2.n178 B2.n176 0.0146
R36050 B2.n182 B2.n178 0.0146
R36051 B2.n197 B2.n183 0.0146
R36052 B2.n197 B2.n196 0.0146
R36053 B2.n195 B2.n184 0.0146
R36054 B2.n191 B2.n184 0.0146
R36055 B2.n209 B2.n208 0.0143235
R36056 B2.n207 B2.n175 0.0143235
R36057 B2.n203 B2.n175 0.0143235
R36058 B2.n202 B2.n201 0.0143235
R36059 B2.n201 B2.n177 0.0143235
R36060 B2.n198 B2.n180 0.0143235
R36061 B2.n198 B2.n181 0.0143235
R36062 B2.n194 B2.n193 0.0143235
R36063 B2.n193 B2.n192 0.0143235
R36064 B2.n188 B2.n185 0.0143235
R36065 B2.n121 B2.n120 0.0138019
R36066 B2.n132 B2.n26 0.0138019
R36067 B2.n133 B2.n132 0.0138019
R36068 B2.n146 B2.n17 0.0138019
R36069 B2.n147 B2.n146 0.0138019
R36070 B2.n157 B2.n10 0.0138019
R36071 B2.n158 B2.n157 0.0138019
R36072 B2.n159 B2.n4 0.0138019
R36073 B2.n171 B2.n4 0.0138019
R36074 B2.n212 B2.n172 0.0138019
R36075 B2.n212 B2.n211 0.0138019
R36076 B2.n109 B2.n87 0.013431
R36077 B2.n105 B2.n89 0.013431
R36078 B2.n85 B2.n46 0.013
R36079 B2.n66 B2.n48 0.013
R36080 B2.n118 B2.n31 0.0124717
R36081 B2.n123 B2.n31 0.0124717
R36082 B2.n161 B2.n5 0.0124717
R36083 B2.n169 B2.n5 0.0124717
R36084 B2.n73 B2.n67 0.0122521
R36085 B2.n93 B2.n43 0.0117689
R36086 B2.n55 B2.n44 0.0114102
R36087 B2.n130 B2.n129 0.0111132
R36088 B2.n136 B2.n22 0.0111132
R36089 B2.n151 B2.n13 0.0111132
R36090 B2.n155 B2.n154 0.0111132
R36091 B2.n82 B2.n69 0.0100704
R36092 B2.n111 B2.n42 0.0100109
R36093 B2.n138 B2.n137 0.00993396
R36094 B2.n20 B2.n15 0.00993396
R36095 B2.n206 B2.n173 0.0099
R36096 B2.n204 B2.n176 0.0099
R36097 B2.n183 B2.n182 0.0099
R36098 B2.n196 B2.n195 0.0099
R36099 B2.n191 B2.n190 0.0099
R36100 B2.n32 B2.n27 0.00981132
R36101 B2.n12 B2.n9 0.00981132
R36102 B2.n214 B2.n3 0.00981132
R36103 B2.n208 B2.n207 0.00971569
R36104 B2.n203 B2.n202 0.00971569
R36105 B2.n180 B2.n177 0.00971569
R36106 B2.n194 B2.n181 0.00971569
R36107 B2.n192 B2.n185 0.00971569
R36108 B2.n139 B2.n21 0.00967431
R36109 B2.n141 B2.n14 0.00967431
R36110 B2.n122 B2.n32 0.00936793
R36111 B2.n134 B2.n25 0.00936793
R36112 B2.n149 B2.n148 0.00936793
R36113 B2.n160 B2.n9 0.00936793
R36114 B2.n170 B2.n3 0.00936793
R36115 B2.n121 B2.n26 0.00936793
R36116 B2.n133 B2.n17 0.00936793
R36117 B2.n147 B2.n10 0.00936793
R36118 B2.n159 B2.n158 0.00936793
R36119 B2.n172 B2.n171 0.00936793
R36120 B2.n34 B2.n33 0.00875472
R36121 B2.n129 B2.n28 0.00875472
R36122 B2.n154 B2.n8 0.00875472
R36123 B2.n215 B2.n1 0.00875472
R36124 B2.n114 B2.n113 0.00852752
R36125 B2.n128 B2.n127 0.00852752
R36126 B2.n153 B2.n7 0.00852752
R36127 B2.n216 B2.n0 0.00852752
R36128 B2.n145 B2.n18 0.00803774
R36129 B2.n145 B2.n16 0.00803774
R36130 B2.n131 B2.n24 0.00759434
R36131 B2.n156 B2.n11 0.00759434
R36132 B2.n25 B2.n18 0.00626415
R36133 B2.n148 B2.n16 0.00626415
R36134 B2.n109 B2.n89 0.00588793
R36135 B2.n85 B2.n66 0.00570833
R36136 B2.n213 B2.n2 0.00519331
R36137 B2 B2.n217 0.00508716
R36138 B2.n97 B2.n43 0.00481034
R36139 B2.n82 B2.n81 0.0047735
R36140 B2.n52 B2.n44 0.00466667
R36141 B2.n88 B2.n42 0.00457609
R36142 B2.n111 B2.n110 0.00457609
R36143 B2.n131 B2.n27 0.00449057
R36144 B2.n135 B2.n24 0.00449057
R36145 B2.n150 B2.n11 0.00449057
R36146 B2.n156 B2.n12 0.00449057
R36147 B2.n214 B2.n213 0.00449057
R36148 B2.n37 B2.n35 0.00410577
R36149 B2.n74 B2.n73 0.00370513
R36150 B2.n135 B2.n134 0.00271698
R36151 B2.n150 B2.n149 0.00271698
R36152 B2.n83 B2.n68 0.00253804
R36153 B2.n39 B2.n38 0.00185919
R36154 B2.n84 B2.n45 0.0018587
R36155 B2.n123 B2.n122 0.00183019
R36156 B2.n161 B2.n160 0.00183019
R36157 B2.n170 B2.n169 0.00183019
R36158 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 356.022
R36159 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n65 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n64 292.5
R36160 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n28 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n23 152
R36161 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n33 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n22 152
R36162 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n38 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n21 152
R36163 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n43 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n20 152
R36164 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n48 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n19 152
R36165 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n53 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n18 152
R36166 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n58 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n17 152
R36167 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n60 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n59 152
R36168 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n55 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n54 152
R36169 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n50 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n49 152
R36170 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n45 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n44 152
R36171 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n40 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n39 152
R36172 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n35 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n34 152
R36173 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n30 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n29 152
R36174 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n64 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t0 147.756
R36175 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t1 105.415
R36176 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n13 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t5 84.8325
R36177 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t6 84.8325
R36178 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n13 60.1541
R36179 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n15 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 50.1642
R36180 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n13 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t3 48.6825
R36181 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n14 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t4 48.6825
R36182 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n62 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n61 45.1373
R36183 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 36.3683
R36184 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n1 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n60 33.7894
R36185 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n56 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n55 29.03
R36186 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n51 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n50 29.03
R36187 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n46 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n45 29.03
R36188 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n41 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n40 29.03
R36189 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n36 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n35 29.03
R36190 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n31 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n30 29.03
R36191 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n26 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n25 28.4823
R36192 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n25 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n24 26.4823
R36193 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n16 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n15 15.6972
R36194 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n59 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n11 16.3795
R36195 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n54 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n6 16.2631
R36196 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n49 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n8 16.1289
R36197 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n44 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n10 15.9761
R36198 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n65 10.4732
R36199 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n11 2.10258
R36200 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n6 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 2.08561
R36201 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n57 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n56 9.3005
R36202 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n8 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 2.07495
R36203 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n52 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n51 9.3005
R36204 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n10 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 2.07042
R36205 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n47 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n46 9.3005
R36206 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n9 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 2.07192
R36207 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n42 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n41 9.3005
R36208 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n7 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 2.0795
R36209 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n37 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n36 9.3005
R36210 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n32 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n5 2.77054
R36211 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n32 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n31 9.3005
R36212 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n5 2.09329
R36213 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n27 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n26 9.3005
R36214 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n2 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n1 18.3534
R36215 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n26 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n23 8.76414
R36216 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n31 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n22 7.66868
R36217 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n60 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n17 7.12095
R36218 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n63 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n62 6.98232
R36219 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n62 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 6.73734
R36220 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n36 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n21 6.57323
R36221 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n55 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n18 6.0255
R36222 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n28 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n27 6.02403
R36223 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n41 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n20 5.47777
R36224 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n33 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n32 5.27109
R36225 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n61 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 5.22977
R36226 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n63 5.04292
R36227 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n50 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n19 4.93005
R36228 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n59 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n58 4.89462
R36229 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 4.74124
R36230 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n2 4.55946
R36231 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n38 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n37 4.51815
R36232 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n37 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n7 2.64533
R36233 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n27 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n24 4.45253
R36234 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n46 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n19 4.38232
R36235 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n54 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n53 4.14168
R36236 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n12 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 3.87929
R36237 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n65 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 3.87929
R36238 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n45 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n20 3.83459
R36239 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n43 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n42 3.76521
R36240 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n42 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n9 2.50198
R36241 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n16 3.43953
R36242 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n49 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n48 3.38874
R36243 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n51 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n18 3.28686
R36244 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n48 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n47 3.01226
R36245 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n47 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n10 2.33997
R36246 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n40 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n21 2.73914
R36247 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n44 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n43 2.63579
R36248 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n39 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n9 15.804
R36249 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n53 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n52 2.25932
R36250 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n52 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n8 2.15681
R36251 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n56 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n17 2.19141
R36252 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n39 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n38 1.88285
R36253 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n34 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n7 15.6099
R36254 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n35 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n22 1.64368
R36255 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n16 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 1.52175
R36256 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n25 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.t2 1.50675
R36257 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n58 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n57 1.50638
R36258 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n57 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n6 1.95132
R36259 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 1.37511
R36260 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n15 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 1.1768
R36261 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n34 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n33 1.12991
R36262 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n29 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n5 15.3925
R36263 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n11 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n1 4.58496
R36264 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n4 0.679754
R36265 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n30 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n23 0.548227
R36266 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n61 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH 0.546841
R36267 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n24 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 0.471686
R36268 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 0.468612
R36269 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n29 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n28 0.376971
R36270 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n2 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOH.n0 0.310701
R36271 a_8085_2982.n109 a_8085_2982.t3 120.501
R36272 a_8085_2982.n21 a_8085_2982.t1 69.2068
R36273 a_8085_2982.n59 a_8085_2982.t2 60.2505
R36274 a_8085_2982.n46 a_8085_2982.n45 31.4488
R36275 a_8085_2982.n24 a_8085_2982.n23 27.5177
R36276 a_8085_2982.n7 a_8085_2982.n3 26.107
R36277 a_8085_2982.n35 a_8085_2982.n34 23.5867
R36278 a_8085_2982.n13 a_8085_2982.n12 19.6557
R36279 a_8085_2982.n3 a_8085_2982.n2 15.7246
R36280 a_8085_2982.n14 a_8085_2982.n13 13.7591
R36281 a_8085_2982.n36 a_8085_2982.n35 9.82809
R36282 a_8085_2982.n86 a_8085_2982.n85 9.3005
R36283 a_8085_2982.n69 a_8085_2982.n68 9.3005
R36284 a_8085_2982.n123 a_8085_2982.n122 9.3005
R36285 a_8085_2982.n104 a_8085_2982.n103 9.3005
R36286 a_8085_2982.n50 a_8085_2982.n52 9.3005
R36287 a_8085_2982.n15 a_8085_2982.n14 9.3005
R36288 a_8085_2982.n37 a_8085_2982.n36 9.3005
R36289 a_8085_2982.n28 a_8085_2982.n38 9.3005
R36290 a_8085_2982.n26 a_8085_2982.n25 9.3005
R36291 a_8085_2982.n39 a_8085_2982.n41 9.3005
R36292 a_8085_2982.n48 a_8085_2982.n47 9.3005
R36293 a_8085_2982.n1 a_8085_2982.n139 9.3005
R36294 a_8085_2982.n131 a_8085_2982.n146 9.3005
R36295 a_8085_2982.n1 a_8085_2982.n138 9.3005
R36296 a_8085_2982.n0 a_8085_2982.n134 9.3005
R36297 a_8085_2982.n131 a_8085_2982.n145 9.3005
R36298 a_8085_2982.n60 a_8085_2982.n59 8.76429
R36299 a_8085_2982.n110 a_8085_2982.n109 8.76429
R36300 a_8085_2982.n67 a_8085_2982.n66 8.21641
R36301 a_8085_2982.n84 a_8085_2982.n83 8.21641
R36302 a_8085_2982.n102 a_8085_2982.n101 7.45411
R36303 a_8085_2982.n121 a_8085_2982.n120 7.45411
R36304 a_8085_2982.n25 a_8085_2982.n24 5.89705
R36305 a_8085_2982.n150 a_8085_2982.n149 5.38095
R36306 a_8085_2982.n8 a_8085_2982.n7 5.20544
R36307 a_8085_2982.n56 a_8085_2982.n54 4.87224
R36308 a_8085_2982.n89 a_8085_2982.n74 4.86623
R36309 a_8085_2982.n92 a_8085_2982.n90 4.84151
R36310 a_8085_2982.n126 a_8085_2982.n108 4.83995
R36311 a_8085_2982.n111 a_8085_2982.n110 4.6505
R36312 a_8085_2982.n0 a_8085_2982.n133 4.5298
R36313 a_8085_2982.n30 a_8085_2982.n31 4.51815
R36314 a_8085_2982.n33 a_8085_2982.n32 4.51815
R36315 a_8085_2982.n55 a_8085_2982.n70 4.5005
R36316 a_8085_2982.n57 a_8085_2982.n63 4.5005
R36317 a_8085_2982.n77 a_8085_2982.n81 4.5005
R36318 a_8085_2982.n82 a_8085_2982.n88 4.5005
R36319 a_8085_2982.n91 a_8085_2982.n105 4.5005
R36320 a_8085_2982.n93 a_8085_2982.n98 4.5005
R36321 a_8085_2982.n114 a_8085_2982.n118 4.5005
R36322 a_8085_2982.n119 a_8085_2982.n125 4.5005
R36323 a_8085_2982.n8 a_8085_2982.n16 4.5005
R36324 a_8085_2982.n42 a_8085_2982.n49 4.5005
R36325 a_8085_2982.n29 a_8085_2982.n27 4.5005
R36326 a_8085_2982.n94 a_8085_2982.n95 4.5005
R36327 a_8085_2982.n113 a_8085_2982.n112 4.5005
R36328 a_8085_2982.n1 a_8085_2982.n137 4.5005
R36329 a_8085_2982.n130 a_8085_2982.n144 4.5005
R36330 a_8085_2982.n58 a_8085_2982.n60 4.14168
R36331 a_8085_2982.n76 a_8085_2982.n75 4.14168
R36332 a_8085_2982.n49 a_8085_2982.n43 4.14168
R36333 a_8085_2982.n88 a_8085_2982.n86 3.76521
R36334 a_8085_2982.n125 a_8085_2982.n123 3.76521
R36335 a_8085_2982.n16 a_8085_2982.n9 3.76521
R36336 a_8085_2982.n11 a_8085_2982.n10 3.76521
R36337 a_8085_2982.n70 a_8085_2982.n69 3.38874
R36338 a_8085_2982.n105 a_8085_2982.n104 3.38874
R36339 a_8085_2982.n6 a_8085_2982.n5 3.38874
R36340 a_8085_2982.n130 a_8085_2982.n141 3.17178
R36341 a_8085_2982.n70 a_8085_2982.n64 3.01226
R36342 a_8085_2982.n81 a_8085_2982.n80 3.01226
R36343 a_8085_2982.n105 a_8085_2982.n99 3.01226
R36344 a_8085_2982.n98 a_8085_2982.n96 3.01226
R36345 a_8085_2982.n5 a_8085_2982.n4 3.01226
R36346 a_8085_2982.t0 a_8085_2982.n151 2.77
R36347 a_8085_2982.n63 a_8085_2982.n61 2.63579
R36348 a_8085_2982.n88 a_8085_2982.n87 2.63579
R36349 a_8085_2982.n118 a_8085_2982.n117 2.63579
R36350 a_8085_2982.n125 a_8085_2982.n124 2.63579
R36351 a_8085_2982.n16 a_8085_2982.n15 2.63579
R36352 a_8085_2982.n15 a_8085_2982.n11 2.63579
R36353 a_8085_2982.n53 a_8085_2982.n21 2.41452
R36354 a_8085_2982.n107 a_8085_2982.n127 2.28493
R36355 a_8085_2982.n49 a_8085_2982.n48 2.25932
R36356 a_8085_2982.n52 a_8085_2982.n51 2.25932
R36357 a_8085_2982.n47 a_8085_2982.n46 1.96602
R36358 a_8085_2982.n30 a_8085_2982.n37 1.88285
R36359 a_8085_2982.n37 a_8085_2982.n33 1.88285
R36360 a_8085_2982.n151 a_8085_2982.n150 1.84417
R36361 a_8085_2982.n81 a_8085_2982.n78 1.50638
R36362 a_8085_2982.n118 a_8085_2982.n115 1.50638
R36363 a_8085_2982.n117 a_8085_2982.n116 1.50638
R36364 a_8085_2982.n27 a_8085_2982.n26 1.50638
R36365 a_8085_2982.n41 a_8085_2982.n40 1.50638
R36366 a_8085_2982.n151 a_8085_2982.n140 1.32032
R36367 a_8085_2982.n151 a_8085_2982.n148 1.29978
R36368 a_8085_2982.n18 a_8085_2982.n129 1.24675
R36369 a_8085_2982.n107 a_8085_2982.n92 1.21366
R36370 a_8085_2982.n71 a_8085_2982.n89 1.15702
R36371 a_8085_2982.n73 a_8085_2982.n56 1.21147
R36372 a_8085_2982.n106 a_8085_2982.n126 1.15482
R36373 a_8085_2982.n63 a_8085_2982.n62 1.12991
R36374 a_8085_2982.n80 a_8085_2982.n79 1.12991
R36375 a_8085_2982.n98 a_8085_2982.n97 1.12991
R36376 a_8085_2982.n26 a_8085_2982.n22 1.12991
R36377 a_8085_2982.n68 a_8085_2982.n67 1.09595
R36378 a_8085_2982.n85 a_8085_2982.n84 1.09595
R36379 a_8085_2982.n1 a_8085_2982.n132 1.04835
R36380 a_8085_2982.n147 a_8085_2982.n127 0.996877
R36381 a_8085_2982.n103 a_8085_2982.n102 0.994314
R36382 a_8085_2982.n122 a_8085_2982.n121 0.994314
R36383 a_8085_2982.n17 a_8085_2982.n53 0.994096
R36384 a_8085_2982.n72 a_8085_2982.n128 0.963
R36385 a_8085_2982.n69 a_8085_2982.n65 0.753441
R36386 a_8085_2982.n104 a_8085_2982.n100 0.753441
R36387 a_8085_2982.n137 a_8085_2982.n135 0.753441
R36388 a_8085_2982.n140 a_8085_2982.n1 0.418831
R36389 a_8085_2982.n148 a_8085_2982.n147 0.386668
R36390 a_8085_2982.n48 a_8085_2982.n44 0.376971
R36391 a_8085_2982.n144 a_8085_2982.n142 0.376971
R36392 a_8085_2982.n7 a_8085_2982.n6 0.319725
R36393 a_8085_2982.n135 a_8085_2982.n136 0.121922
R36394 a_8085_2982.n142 a_8085_2982.n143 0.110027
R36395 a_8085_2982.n147 a_8085_2982.n131 0.0843535
R36396 a_8085_2982.n53 a_8085_2982.n50 0.0827519
R36397 a_8085_2982.n107 a_8085_2982.n106 0.0590938
R36398 a_8085_2982.n42 a_8085_2982.n39 0.100109
R36399 a_8085_2982.n126 a_8085_2982.n119 0.0371012
R36400 a_8085_2982.n131 a_8085_2982.n130 0.0337031
R36401 a_8085_2982.n20 a_8085_2982.n18 0.0287031
R36402 a_8085_2982.n20 a_8085_2982.n19 0.028
R36403 a_8085_2982.n128 a_8085_2982.n107 0.028
R36404 a_8085_2982.n129 a_8085_2982.n73 0.028
R36405 a_8085_2982.n73 a_8085_2982.n72 0.0276737
R36406 a_8085_2982.n113 a_8085_2982.n111 0.0239375
R36407 a_8085_2982.n77 a_8085_2982.n76 4.5892
R36408 a_8085_2982.n114 a_8085_2982.n113 0.0892218
R36409 a_8085_2982.n93 a_8085_2982.n94 0.0883906
R36410 a_8085_2982.n57 a_8085_2982.n58 4.58839
R36411 a_8085_2982.n20 a_8085_2982.n17 0.119641
R36412 a_8085_2982.n28 a_8085_2982.n30 4.61452
R36413 a_8085_2982.n73 a_8085_2982.n71 0.0590938
R36414 a_8085_2982.n82 a_8085_2982.n77 0.0454219
R36415 a_8085_2982.n119 a_8085_2982.n114 0.0454219
R36416 a_8085_2982.n91 a_8085_2982.n93 0.0454219
R36417 a_8085_2982.n55 a_8085_2982.n57 0.0454219
R36418 a_8085_2982.n92 a_8085_2982.n91 0.0388205
R36419 a_8085_2982.n89 a_8085_2982.n82 0.0385721
R36420 a_8085_2982.n56 a_8085_2982.n55 0.0373496
R36421 a_8085_2982.n50 a_8085_2982.n42 0.0337031
R36422 a_8085_2982.n39 a_8085_2982.n29 0.0337031
R36423 a_8085_2982.n29 a_8085_2982.n28 0.0268395
R36424 a_8085_2982.n20 a_8085_2982.n8 1.5962
R36425 a_8085_2982.n1 a_8085_2982.n0 0.225375
R36426 EF_R2RVCE_0.comparator_0.VBP.n29 EF_R2RVCE_0.comparator_0.VBP.t3 116.841
R36427 EF_R2RVCE_0.comparator_0.VBP.n56 EF_R2RVCE_0.comparator_0.VBP.t2 60.2505
R36428 EF_R2RVCE_0.comparator_0.VBP.n98 EF_R2RVCE_0.comparator_0.VBP.t4 60.2505
R36429 EF_R2RVCE_0.comparator_0.VBP.n110 EF_R2RVCE_0.comparator_0.VBP.t5 60.2505
R36430 EF_R2RVCE_0.comparator_0.VBP.n33 EF_R2RVCE_0.comparator_0.VBP.n32 52.6902
R36431 EF_R2RVCE_0.comparator_0.VBP.n41 EF_R2RVCE_0.comparator_0.VBP.n40 46.104
R36432 EF_R2RVCE_0.comparator_0.VBP.n89 EF_R2RVCE_0.comparator_0.VBP.n88 39.5177
R36433 EF_R2RVCE_0.comparator_0.VBP.n81 EF_R2RVCE_0.comparator_0.VBP.n80 32.9315
R36434 EF_R2RVCE_0.comparator_0.VBP.n72 EF_R2RVCE_0.comparator_0.VBP.n71 29.6384
R36435 EF_R2RVCE_0.comparator_0.VBP.n71 EF_R2RVCE_0.comparator_0.VBP.n70 26.3453
R36436 EF_R2RVCE_0.comparator_0.VBP.n82 EF_R2RVCE_0.comparator_0.VBP.n81 23.0522
R36437 EF_R2RVCE_0.comparator_0.VBP.n90 EF_R2RVCE_0.comparator_0.VBP.n89 16.466
R36438 EF_R2RVCE_0.comparator_0.VBP.n42 EF_R2RVCE_0.comparator_0.VBP.n41 9.87981
R36439 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n36 9.3005
R36440 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n44 9.3005
R36441 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n43 9.3005
R36442 EF_R2RVCE_0.comparator_0.VBP.n43 EF_R2RVCE_0.comparator_0.VBP.n42 9.3005
R36443 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n37 9.3005
R36444 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n35 9.3005
R36445 EF_R2RVCE_0.comparator_0.VBP.n35 EF_R2RVCE_0.comparator_0.VBP.n34 9.3005
R36446 EF_R2RVCE_0.comparator_0.VBP.n8 EF_R2RVCE_0.comparator_0.VBP.n76 9.3005
R36447 EF_R2RVCE_0.comparator_0.VBP.n83 EF_R2RVCE_0.comparator_0.VBP.n82 9.3005
R36448 EF_R2RVCE_0.comparator_0.VBP.n91 EF_R2RVCE_0.comparator_0.VBP.n90 9.3005
R36449 EF_R2RVCE_0.comparator_0.VBP.n8 EF_R2RVCE_0.comparator_0.VBP.n73 9.3005
R36450 EF_R2RVCE_0.comparator_0.VBP.n73 EF_R2RVCE_0.comparator_0.VBP.n72 9.3005
R36451 EF_R2RVCE_0.comparator_0.VBP.n65 EF_R2RVCE_0.comparator_0.VBP.n64 9.3005
R36452 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n59 9.3005
R36453 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n48 9.3005
R36454 EF_R2RVCE_0.comparator_0.VBP.n54 EF_R2RVCE_0.comparator_0.VBP.n53 9.3005
R36455 EF_R2RVCE_0.comparator_0.VBP.n4 EF_R2RVCE_0.comparator_0.VBP.n107 9.3005
R36456 EF_R2RVCE_0.comparator_0.VBP.n4 EF_R2RVCE_0.comparator_0.VBP.n105 9.3005
R36457 EF_R2RVCE_0.comparator_0.VBP.n105 EF_R2RVCE_0.comparator_0.VBP.n104 9.3005
R36458 EF_R2RVCE_0.comparator_0.VBP.n4 EF_R2RVCE_0.comparator_0.VBP.n106 9.3005
R36459 EF_R2RVCE_0.comparator_0.VBP.n5 EF_R2RVCE_0.comparator_0.VBP.n117 9.3005
R36460 EF_R2RVCE_0.comparator_0.VBP.n117 EF_R2RVCE_0.comparator_0.VBP.n116 9.3005
R36461 EF_R2RVCE_0.comparator_0.VBP.n5 EF_R2RVCE_0.comparator_0.VBP.n119 9.3005
R36462 EF_R2RVCE_0.comparator_0.VBP.n5 EF_R2RVCE_0.comparator_0.VBP.n118 9.3005
R36463 EF_R2RVCE_0.comparator_0.VBP.n6 EF_R2RVCE_0.comparator_0.VBP.n18 9.3005
R36464 EF_R2RVCE_0.comparator_0.VBP.n6 EF_R2RVCE_0.comparator_0.VBP.n13 9.3005
R36465 EF_R2RVCE_0.comparator_0.VBP.n57 EF_R2RVCE_0.comparator_0.VBP.n56 8.76429
R36466 EF_R2RVCE_0.comparator_0.VBP.n52 EF_R2RVCE_0.comparator_0.VBP.n51 7.45411
R36467 EF_R2RVCE_0.comparator_0.VBP.n63 EF_R2RVCE_0.comparator_0.VBP.n62 7.45411
R36468 EF_R2RVCE_0.comparator_0.VBP.n103 EF_R2RVCE_0.comparator_0.VBP.n102 7.45411
R36469 EF_R2RVCE_0.comparator_0.VBP.n115 EF_R2RVCE_0.comparator_0.VBP.n114 7.45411
R36470 EF_R2RVCE_0.comparator_0.VBP.n99 EF_R2RVCE_0.comparator_0.VBP.n98 6.80105
R36471 EF_R2RVCE_0.comparator_0.VBP.n111 EF_R2RVCE_0.comparator_0.VBP.n110 6.801
R36472 EF_R2RVCE_0.comparator_0.VBP.n31 EF_R2RVCE_0.comparator_0.VBP.n30 6.02403
R36473 EF_R2RVCE_0.comparator_0.VBP.n2 EF_R2RVCE_0.comparator_0.VBP.n93 6.0005
R36474 EF_R2RVCE_0.comparator_0.VBP.n2 EF_R2RVCE_0.comparator_0.VBP.n86 6.0005
R36475 EF_R2RVCE_0.comparator_0.VBP.n50 EF_R2RVCE_0.comparator_0.VBP.n49 5.64756
R36476 EF_R2RVCE_0.comparator_0.VBP.n61 EF_R2RVCE_0.comparator_0.VBP.n60 5.64756
R36477 EF_R2RVCE_0.comparator_0.VBP.n101 EF_R2RVCE_0.comparator_0.VBP.n100 5.64756
R36478 EF_R2RVCE_0.comparator_0.VBP.n113 EF_R2RVCE_0.comparator_0.VBP.n112 5.64756
R36479 EF_R2RVCE_0.comparator_0.VBP.n39 EF_R2RVCE_0.comparator_0.VBP.n38 5.27109
R36480 EF_R2RVCE_0.comparator_0.VBP.n10 EF_R2RVCE_0.comparator_0.VBP.n69 5.25098
R36481 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n47 4.88281
R36482 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n58 4.88086
R36483 EF_R2RVCE_0.comparator_0.VBP.n1 EF_R2RVCE_0.comparator_0.VBP.n9 4.54542
R36484 EF_R2RVCE_0.comparator_0.VBP.n16 EF_R2RVCE_0.comparator_0.VBP.n15 4.51815
R36485 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n55 4.5005
R36486 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n66 4.5005
R36487 EF_R2RVCE_0.comparator_0.VBP.n8 EF_R2RVCE_0.comparator_0.VBP.n78 4.5005
R36488 EF_R2RVCE_0.comparator_0.VBP.n10 EF_R2RVCE_0.comparator_0.VBP.n68 4.5005
R36489 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n46 4.5005
R36490 EF_R2RVCE_0.comparator_0.VBP.n6 EF_R2RVCE_0.comparator_0.VBP.n16 4.5005
R36491 EF_R2RVCE_0.comparator_0.VBP.n6 EF_R2RVCE_0.comparator_0.VBP.n21 4.5005
R36492 EF_R2RVCE_0.comparator_0.VBP.n1 EF_R2RVCE_0.comparator_0.VBP.n26 4.5005
R36493 EF_R2RVCE_0.comparator_0.VBP.n4 EF_R2RVCE_0.comparator_0.VBP.n97 4.24504
R36494 EF_R2RVCE_0.comparator_0.VBP.n5 EF_R2RVCE_0.comparator_0.VBP.n109 4.24504
R36495 EF_R2RVCE_0.comparator_0.VBP.n3 EF_R2RVCE_0.comparator_0.VBP.n29 4.23684
R36496 EF_R2RVCE_0.comparator_0.VBP.n93 EF_R2RVCE_0.comparator_0.VBP.n87 4.14168
R36497 EF_R2RVCE_0.comparator_0.VBP.n21 EF_R2RVCE_0.comparator_0.VBP.n20 3.76521
R36498 EF_R2RVCE_0.comparator_0.VBP.n5 EF_R2RVCE_0.comparator_0.VBP.n111 3.42853
R36499 EF_R2RVCE_0.comparator_0.VBP.n4 EF_R2RVCE_0.comparator_0.VBP.n99 3.42768
R36500 EF_R2RVCE_0.comparator_0.VBP.n86 EF_R2RVCE_0.comparator_0.VBP.n79 3.38874
R36501 EF_R2RVCE_0.comparator_0.VBP.n27 EF_R2RVCE_0.comparator_0.VBP.t0 3.3065
R36502 EF_R2RVCE_0.comparator_0.VBP.n27 EF_R2RVCE_0.comparator_0.VBP.t1 3.3065
R36503 EF_R2RVCE_0.comparator_0.VBP.n34 EF_R2RVCE_0.comparator_0.VBP.n33 3.2936
R36504 EF_R2RVCE_0.comparator_0.VBP.n26 EF_R2RVCE_0.comparator_0.VBP.n24 3.74814
R36505 EF_R2RVCE_0.comparator_0.VBP EF_R2RVCE_0.comparator_0.VBP.n95 3.26842
R36506 EF_R2RVCE_0.comparator_0.VBP.n1 EF_R2RVCE_0.comparator_0.VBP.n28 3.15814
R36507 EF_R2RVCE_0.comparator_0.VBP.n0 EF_R2RVCE_0.comparator_0.VBP.n57 3.03311
R36508 EF_R2RVCE_0.comparator_0.VBP.n75 EF_R2RVCE_0.comparator_0.VBP.n74 3.01226
R36509 EF_R2RVCE_0.comparator_0.VBP.n26 EF_R2RVCE_0.comparator_0.VBP.n25 3.01226
R36510 EF_R2RVCE_0.comparator_0.VBP.n6 EF_R2RVCE_0.comparator_0.VBP.n11 2.77255
R36511 EF_R2RVCE_0.comparator_0.VBP.n21 EF_R2RVCE_0.comparator_0.VBP.n19 2.63579
R36512 EF_R2RVCE_0.comparator_0.VBP.n13 EF_R2RVCE_0.comparator_0.VBP.n12 2.61733
R36513 EF_R2RVCE_0.comparator_0.VBP.n85 EF_R2RVCE_0.comparator_0.VBP.n84 2.25932
R36514 EF_R2RVCE_0.comparator_0.VBP.n18 EF_R2RVCE_0.comparator_0.VBP.n17 2.24766
R36515 EF_R2RVCE_0.comparator_0.VBP.n92 EF_R2RVCE_0.comparator_0.VBP.n91 1.88285
R36516 EF_R2RVCE_0.comparator_0.VBP.n76 EF_R2RVCE_0.comparator_0.VBP.n75 1.88285
R36517 EF_R2RVCE_0.comparator_0.VBP.n16 EF_R2RVCE_0.comparator_0.VBP.n14 1.88285
R36518 EF_R2RVCE_0.comparator_0.VBP.n7 EF_R2RVCE_0.comparator_0.VBP.n0 1.85011
R36519 EF_R2RVCE_0.comparator_0.VBP.n22 EF_R2RVCE_0.comparator_0.VBP.n1 1.82596
R36520 EF_R2RVCE_0.comparator_0.VBP.n120 EF_R2RVCE_0.comparator_0.VBP.n5 1.75631
R36521 EF_R2RVCE_0.comparator_0.VBP.n2 EF_R2RVCE_0.comparator_0.VBP.n3 1.74716
R36522 EF_R2RVCE_0.comparator_0.VBP.n22 EF_R2RVCE_0.comparator_0.VBP.n6 1.6803
R36523 EF_R2RVCE_0.comparator_0.VBP.n1 EF_R2RVCE_0.comparator_0.VBP.n27 1.61775
R36524 EF_R2RVCE_0.comparator_0.VBP.n2 EF_R2RVCE_0.comparator_0.VBP.n8 1.60792
R36525 EF_R2RVCE_0.comparator_0.VBP.n2 EF_R2RVCE_0.comparator_0.VBP.n10 1.55128
R36526 EF_R2RVCE_0.comparator_0.VBP.n68 EF_R2RVCE_0.comparator_0.VBP.n67 1.50638
R36527 EF_R2RVCE_0.comparator_0.VBP EF_R2RVCE_0.comparator_0.VBP.n120 1.3155
R36528 EF_R2RVCE_0.comparator_0.VBP.n43 EF_R2RVCE_0.comparator_0.VBP.n39 1.12991
R36529 EF_R2RVCE_0.comparator_0.VBP.n9 EF_R2RVCE_0.comparator_0.VBP.n23 1.12991
R36530 EF_R2RVCE_0.comparator_0.VBP.n95 EF_R2RVCE_0.comparator_0.VBP.n22 1.04295
R36531 EF_R2RVCE_0.comparator_0.VBP.n53 EF_R2RVCE_0.comparator_0.VBP.n52 0.994314
R36532 EF_R2RVCE_0.comparator_0.VBP.n64 EF_R2RVCE_0.comparator_0.VBP.n63 0.994314
R36533 EF_R2RVCE_0.comparator_0.VBP.n104 EF_R2RVCE_0.comparator_0.VBP.n103 0.994314
R36534 EF_R2RVCE_0.comparator_0.VBP.n116 EF_R2RVCE_0.comparator_0.VBP.n115 0.994314
R36535 EF_R2RVCE_0.comparator_0.VBP.n94 EF_R2RVCE_0.comparator_0.VBP.n2 0.794925
R36536 EF_R2RVCE_0.comparator_0.VBP.n46 EF_R2RVCE_0.comparator_0.VBP.n45 0.753441
R36537 EF_R2RVCE_0.comparator_0.VBP.n78 EF_R2RVCE_0.comparator_0.VBP.n77 0.753441
R36538 EF_R2RVCE_0.comparator_0.VBP.n55 EF_R2RVCE_0.comparator_0.VBP.n54 0.753441
R36539 EF_R2RVCE_0.comparator_0.VBP.n54 EF_R2RVCE_0.comparator_0.VBP.n50 0.753441
R36540 EF_R2RVCE_0.comparator_0.VBP.n65 EF_R2RVCE_0.comparator_0.VBP.n61 0.753441
R36541 EF_R2RVCE_0.comparator_0.VBP.n66 EF_R2RVCE_0.comparator_0.VBP.n65 0.753441
R36542 EF_R2RVCE_0.comparator_0.VBP.n105 EF_R2RVCE_0.comparator_0.VBP.n101 0.753441
R36543 EF_R2RVCE_0.comparator_0.VBP.n117 EF_R2RVCE_0.comparator_0.VBP.n113 0.753441
R36544 EF_R2RVCE_0.comparator_0.VBP.n2 EF_R2RVCE_0.comparator_0.VBP.n7 0.748981
R36545 EF_R2RVCE_0.comparator_0.VBP.n97 EF_R2RVCE_0.comparator_0.VBP.n96 0.709906
R36546 EF_R2RVCE_0.comparator_0.VBP.n109 EF_R2RVCE_0.comparator_0.VBP.n108 0.709906
R36547 EF_R2RVCE_0.comparator_0.VBP.n5 EF_R2RVCE_0.comparator_0.VBP.n4 0.673704
R36548 EF_R2RVCE_0.comparator_0.VBP.n95 EF_R2RVCE_0.comparator_0.VBP.n94 0.577213
R36549 EF_R2RVCE_0.comparator_0.VBP.n7 EF_R2RVCE_0.comparator_0.VBP 0.538902
R36550 EF_R2RVCE_0.comparator_0.VBP.n35 EF_R2RVCE_0.comparator_0.VBP.n31 0.376971
R36551 EF_R2RVCE_0.comparator_0.VBP.n93 EF_R2RVCE_0.comparator_0.VBP.n92 0.376971
R36552 EF_R2RVCE_0.comparator_0.VBP.n86 EF_R2RVCE_0.comparator_0.VBP.n85 0.376971
R36553 EF_R2RVCE_0.comparator_0.VBP.n84 EF_R2RVCE_0.comparator_0.VBP.n83 0.376971
R36554 A1.n66 A1.n65 185
R36555 A1.n64 A1.n57 185
R36556 A1.n24 A1.n15 185
R36557 A1.n23 A1.n22 185
R36558 A1.n69 A1.t5 120.037
R36559 A1.t6 A1.n14 120.037
R36560 A1.n59 A1.n57 112.831
R36561 A1.n22 A1.n21 112.831
R36562 A1.n68 A1.n67 104.172
R36563 A1.n27 A1.n26 104.172
R36564 A1.n68 A1.n56 92.5005
R36565 A1.n28 A1.n27 92.5005
R36566 A1.t5 A1.n68 66.8281
R36567 A1.n27 A1.t6 66.8281
R36568 A1.n6 A1.t0 35.2053
R36569 A1.n3 A1.t1 34.0571
R36570 A1.n67 A1.n66 29.4833
R36571 A1.n26 A1.n15 29.4833
R36572 A1.n1 A1.t7 27.6955
R36573 A1.n1 A1.t4 27.6955
R36574 A1.n45 A1.n44 19.0955
R36575 A1.n69 A1.n56 15.4558
R36576 A1.n28 A1.n14 15.4558
R36577 A1.n64 A1.n63 13.5534
R36578 A1.n23 A1.n18 13.5534
R36579 A1.n2 A1.n1 9.67857
R36580 A1.n41 A1.n34 9.30581
R36581 A1.n59 A1.n58 9.30424
R36582 A1.n21 A1.n20 9.30413
R36583 A1.n40 A1.n39 9.3005
R36584 A1.n46 A1.n45 9.3005
R36585 A1.n71 A1.n70 9.3005
R36586 A1.n55 A1.n52 9.3005
R36587 A1.n67 A1.n55 9.3005
R36588 A1.n63 A1.n62 9.3005
R36589 A1.n72 A1.n54 9.3005
R36590 A1.n29 A1.n13 9.3005
R36591 A1.n25 A1.n11 9.3005
R36592 A1.n26 A1.n25 9.3005
R36593 A1.n18 A1.n17 9.3005
R36594 A1.n31 A1.n30 9.3005
R36595 A1.n71 A1.n56 9.03579
R36596 A1.n29 A1.n28 9.03579
R36597 A1.n43 A1.n41 8.49366
R36598 A1.n43 A1.t2 8.2655
R36599 A1.n43 A1.t3 8.2655
R36600 A1.n44 A1.n43 7.97749
R36601 A1.n42 A1.n40 7.26743
R36602 A1.n43 A1.n42 6.15568
R36603 A1.n65 A1.n55 5.64756
R36604 A1.n25 A1.n24 5.64756
R36605 A1.n41 A1.n35 4.89462
R36606 A1.n60 A1.n59 4.89462
R36607 A1.n21 A1.n19 4.89462
R36608 A1.n73 A1.n55 4.51815
R36609 A1.n72 A1.n71 4.51815
R36610 A1.n25 A1.n12 4.51815
R36611 A1.n30 A1.n29 4.51815
R36612 A1.n5 A1.n4 4.5005
R36613 A1.n4 A1.n2 4.5005
R36614 A1.n51 A1.n9 4.5005
R36615 A1.n49 A1.n9 4.5005
R36616 A1.n51 A1.n50 4.5005
R36617 A1.n50 A1.n49 4.5005
R36618 A1.n74 A1.n53 4.5005
R36619 A1.n75 A1.n8 4.5005
R36620 A1.n53 A1.n8 4.5005
R36621 A1.n75 A1.n74 4.5005
R36622 A1.n48 A1.n32 4.5005
R36623 A1.n47 A1.n36 4.5005
R36624 A1.n48 A1.n47 4.5005
R36625 A1.n36 A1.n32 4.5005
R36626 A1.n38 A1.n33 4.5005
R36627 A1.n66 A1.n57 3.93153
R36628 A1.n22 A1.n15 3.93153
R36629 A1.n19 A1.n9 3.03311
R36630 A1.n50 A1.n12 3.03311
R36631 A1.n60 A1.n8 3.03311
R36632 A1.n74 A1.n73 3.03311
R36633 A1.n47 A1.n35 3.03311
R36634 A1.n3 A1.n0 2.2714
R36635 A1.n58 A1.n7 2.25261
R36636 A1.n20 A1.n10 2.25256
R36637 A1.n34 A1.n33 2.25127
R36638 A1.n37 A1.n33 2.24434
R36639 A1.n213 A1.n212 1.94045
R36640 A1.n73 A1.n72 1.88285
R36641 A1.n30 A1.n12 1.88285
R36642 A1.n148 A1.n126 1.72424
R36643 A1.n131 A1.n130 1.7055
R36644 A1.n135 A1.n134 1.7055
R36645 A1.n139 A1.n138 1.7055
R36646 A1.n143 A1.n142 1.7055
R36647 A1.n147 A1.n146 1.7055
R36648 A1.n164 A1.n163 1.51869
R36649 A1.n45 A1.n35 1.50638
R36650 A1.n63 A1.n60 1.50638
R36651 A1.n19 A1.n18 1.50638
R36652 A1.n16 A1.n10 1.49213
R36653 A1.n70 A1.n69 1.49212
R36654 A1.n61 A1.n7 1.49182
R36655 A1.n14 A1.n13 1.49166
R36656 A1.n217 A1 1.09946
R36657 A1.n78 A1 1.04529
R36658 A1.n212 A1.n211 0.853
R36659 A1.n217 A1 0.797375
R36660 A1.n65 A1.n64 0.753441
R36661 A1.n24 A1.n23 0.753441
R36662 A1.n44 A1.n40 0.521921
R36663 A1.n181 A1.n180 0.513942
R36664 A1.n149 A1.n148 0.326031
R36665 A1.n77 A1.n6 0.29767
R36666 A1.n49 A1.n48 0.238951
R36667 A1.n77 A1.n76 0.196255
R36668 A1 A1.n77 0.1855
R36669 A1.n6 A1.n5 0.149538
R36670 A1.n75 A1.n51 0.124821
R36671 A1.n217 A1.n216 0.0869486
R36672 A1.n126 A1 0.0741607
R36673 A1.n42 A1.n32 0.0579027
R36674 A1.n81 A1.n80 0.0530701
R36675 A1.n82 A1.n81 0.0530701
R36676 A1.n213 A1.n95 0.0530701
R36677 A1.n214 A1.n213 0.0530701
R36678 A1.n85 A1.n84 0.0402196
R36679 A1.n89 A1.n88 0.0402196
R36680 A1.n93 A1.n92 0.0402196
R36681 A1.n62 A1.n61 0.0396286
R36682 A1.n17 A1.n16 0.0383668
R36683 A1.n100 A1.n99 0.0323396
R36684 A1.n101 A1.n100 0.0323396
R36685 A1.n212 A1.n121 0.0323396
R36686 A1.n212 A1.n125 0.0323396
R36687 A1.n46 A1.n37 0.0314092
R36688 A1.n5 A1.n0 0.0281442
R36689 A1.n39 A1.n37 0.0271357
R36690 A1.n98 A1.n97 0.0229057
R36691 A1.n103 A1.n102 0.0229057
R36692 A1.n120 A1.n119 0.0229057
R36693 A1.n124 A1.n123 0.0229057
R36694 A1.n80 A1.n79 0.0226963
R36695 A1.n83 A1.n82 0.0226963
R36696 A1.n95 A1.n94 0.0226963
R36697 A1.n215 A1.n214 0.0226963
R36698 A1.n99 A1.n98 0.0217264
R36699 A1.n102 A1.n101 0.0217264
R36700 A1.n121 A1.n120 0.0217264
R36701 A1.n125 A1.n124 0.0217264
R36702 A1.n111 A1.n110 0.0205472
R36703 A1.n112 A1.n111 0.0205472
R36704 A1.n148 A1.n147 0.0203694
R36705 A1.n61 A1.n52 0.0202788
R36706 A1.n16 A1.n11 0.0196501
R36707 A1.n106 A1.n105 0.0193679
R36708 A1.n117 A1.n116 0.0193679
R36709 A1.n182 A1.n181 0.0189241
R36710 A1.n108 A1.n107 0.0181887
R36711 A1.n110 A1.n109 0.0181887
R36712 A1.n113 A1.n112 0.0181887
R36713 A1.n115 A1.n114 0.0181887
R36714 A1.n86 A1.n85 0.0180234
R36715 A1.n88 A1.n87 0.0180234
R36716 A1.n90 A1.n89 0.0180234
R36717 A1.n92 A1.n91 0.0180234
R36718 A1.n51 A1.n10 0.0168043
R36719 A1.n163 A1.n162 0.0163662
R36720 A1.n36 A1.n33 0.016125
R36721 A1.n128 A1.n127 0.0138019
R36722 A1.n131 A1.n129 0.0138019
R36723 A1.n132 A1.n131 0.0138019
R36724 A1.n135 A1.n133 0.0138019
R36725 A1.n136 A1.n135 0.0138019
R36726 A1.n139 A1.n137 0.0138019
R36727 A1.n140 A1.n139 0.0138019
R36728 A1.n143 A1.n141 0.0138019
R36729 A1.n144 A1.n143 0.0138019
R36730 A1.n147 A1.n145 0.0138019
R36731 A1.n180 A1.n179 0.0138019
R36732 A1.n178 A1.n177 0.0138019
R36733 A1.n177 A1.n176 0.0138019
R36734 A1.n175 A1.n174 0.0138019
R36735 A1.n174 A1.n173 0.0138019
R36736 A1.n172 A1.n171 0.0138019
R36737 A1.n171 A1.n170 0.0138019
R36738 A1.n169 A1.n168 0.0138019
R36739 A1.n168 A1.n167 0.0138019
R36740 A1.n166 A1.n165 0.0138019
R36741 A1.n165 A1.n164 0.0138019
R36742 A1.n74 A1.n52 0.013431
R36743 A1.n70 A1.n54 0.013431
R36744 A1.n161 A1.n160 0.0133182
R36745 A1.n160 A1.n159 0.0133182
R36746 A1.n158 A1.n157 0.0133182
R36747 A1.n157 A1.n156 0.0133182
R36748 A1.n155 A1.n154 0.0133182
R36749 A1.n154 A1.n153 0.0133182
R36750 A1.n152 A1.n151 0.0133182
R36751 A1.n151 A1.n150 0.0133182
R36752 A1.n50 A1.n11 0.013
R36753 A1.n31 A1.n13 0.013
R36754 A1.n183 A1.n182 0.0124717
R36755 A1.n184 A1.n183 0.0124717
R36756 A1.n211 A1.n204 0.0124717
R36757 A1.n211 A1.n210 0.0124717
R36758 A1.n38 A1.n32 0.0122521
R36759 A1.n58 A1.n8 0.0117689
R36760 A1.n20 A1.n9 0.0114102
R36761 A1.n105 A1.n104 0.0111132
R36762 A1.n107 A1.n106 0.0111132
R36763 A1.n116 A1.n115 0.0111132
R36764 A1.n118 A1.n117 0.0111132
R36765 A1.n47 A1.n34 0.0100704
R36766 A1.n76 A1.n7 0.0100109
R36767 A1.n109 A1.n108 0.00993396
R36768 A1.n114 A1.n113 0.00993396
R36769 A1.n87 A1.n86 0.0098458
R36770 A1.n91 A1.n90 0.0098458
R36771 A1 A1.n217 0.0098458
R36772 A1.n187 A1.n186 0.00981132
R36773 A1.n202 A1.n201 0.00981132
R36774 A1.n208 A1.n207 0.00981132
R36775 A1.n129 A1.n128 0.00936793
R36776 A1.n133 A1.n132 0.00936793
R36777 A1.n137 A1.n136 0.00936793
R36778 A1.n141 A1.n140 0.00936793
R36779 A1.n145 A1.n144 0.00936793
R36780 A1.n186 A1.n185 0.00936793
R36781 A1.n192 A1.n191 0.00936793
R36782 A1.n197 A1.n196 0.00936793
R36783 A1.n203 A1.n202 0.00936793
R36784 A1.n209 A1.n208 0.00936793
R36785 A1.n179 A1.n178 0.00936793
R36786 A1.n176 A1.n175 0.00936793
R36787 A1.n173 A1.n172 0.00936793
R36788 A1.n170 A1.n169 0.00936793
R36789 A1.n167 A1.n166 0.00936793
R36790 A1.n162 A1.n161 0.00904545
R36791 A1.n159 A1.n158 0.00904545
R36792 A1.n156 A1.n155 0.00904545
R36793 A1.n153 A1.n152 0.00904545
R36794 A1.n150 A1.n149 0.00904545
R36795 A1.n97 A1.n96 0.00875472
R36796 A1.n104 A1.n103 0.00875472
R36797 A1.n119 A1.n118 0.00875472
R36798 A1.n123 A1.n122 0.00875472
R36799 A1.n79 A1.n78 0.00867757
R36800 A1.n84 A1.n83 0.00867757
R36801 A1.n94 A1.n93 0.00867757
R36802 A1.n216 A1.n215 0.00867757
R36803 A1.n194 A1.n193 0.00803774
R36804 A1.n195 A1.n194 0.00803774
R36805 A1.n189 A1.n188 0.00759434
R36806 A1.n200 A1.n199 0.00759434
R36807 A1.n193 A1.n192 0.00626415
R36808 A1.n196 A1.n195 0.00626415
R36809 A1.n74 A1.n54 0.00588793
R36810 A1.n50 A1.n31 0.00570833
R36811 A1.n206 A1.n205 0.00519331
R36812 A1.n62 A1.n8 0.00481034
R36813 A1.n47 A1.n46 0.0047735
R36814 A1.n17 A1.n9 0.00466667
R36815 A1.n53 A1.n7 0.00457609
R36816 A1.n76 A1.n75 0.00457609
R36817 A1.n188 A1.n187 0.00449057
R36818 A1.n190 A1.n189 0.00449057
R36819 A1.n199 A1.n198 0.00449057
R36820 A1.n201 A1.n200 0.00449057
R36821 A1.n207 A1.n206 0.00449057
R36822 A1.n2 A1.n0 0.00410577
R36823 A1.n39 A1.n38 0.00370513
R36824 A1.n191 A1.n190 0.00271698
R36825 A1.n198 A1.n197 0.00271698
R36826 A1.n48 A1.n33 0.00253804
R36827 A1.n4 A1.n3 0.00185919
R36828 A1.n49 A1.n10 0.0018587
R36829 A1.n185 A1.n184 0.00183019
R36830 A1.n204 A1.n203 0.00183019
R36831 A1.n210 A1.n209 0.00183019
R36832 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 356.022
R36833 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n65 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n64 292.5
R36834 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n28 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n23 152
R36835 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n33 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n22 152
R36836 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n38 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n21 152
R36837 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n43 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n20 152
R36838 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n48 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n19 152
R36839 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n53 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n18 152
R36840 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n58 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n17 152
R36841 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n60 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n59 152
R36842 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n55 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n54 152
R36843 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n50 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n49 152
R36844 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n45 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n44 152
R36845 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n40 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n39 152
R36846 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n35 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n34 152
R36847 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n30 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n29 152
R36848 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n64 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t0 147.756
R36849 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t1 105.415
R36850 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n13 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t5 84.8325
R36851 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t6 84.8325
R36852 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n13 60.1541
R36853 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n15 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 50.1642
R36854 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n13 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t2 48.6825
R36855 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n14 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t4 48.6825
R36856 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n62 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n61 45.1373
R36857 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 36.3683
R36858 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n1 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n60 33.7894
R36859 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n56 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n55 29.03
R36860 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n51 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n50 29.03
R36861 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n46 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n45 29.03
R36862 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n41 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n40 29.03
R36863 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n36 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n35 29.03
R36864 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n31 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n30 29.03
R36865 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n26 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n25 28.4823
R36866 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n25 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n24 26.4823
R36867 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n16 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n15 15.6972
R36868 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n59 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n11 16.3795
R36869 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n54 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n6 16.2631
R36870 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n49 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n8 16.1289
R36871 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n44 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n10 15.9761
R36872 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n65 10.4732
R36873 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n11 2.10258
R36874 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n6 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 2.08561
R36875 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n57 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n56 9.3005
R36876 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n8 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 2.07495
R36877 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n52 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n51 9.3005
R36878 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n10 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 2.07042
R36879 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n47 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n46 9.3005
R36880 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n9 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 2.07192
R36881 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n42 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n41 9.3005
R36882 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n7 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 2.0795
R36883 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n37 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n36 9.3005
R36884 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n32 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n5 2.77054
R36885 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n32 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n31 9.3005
R36886 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n5 2.09329
R36887 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n27 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n26 9.3005
R36888 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n2 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n1 18.3534
R36889 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n26 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n23 8.76414
R36890 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n31 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n22 7.66868
R36891 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n60 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n17 7.12095
R36892 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n63 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n62 6.98232
R36893 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n62 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 6.73734
R36894 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n36 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n21 6.57323
R36895 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n55 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n18 6.0255
R36896 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n28 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n27 6.02403
R36897 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n41 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n20 5.47777
R36898 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n33 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n32 5.27109
R36899 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n61 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 5.22977
R36900 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n63 5.04292
R36901 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n50 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n19 4.93005
R36902 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n59 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n58 4.89462
R36903 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 4.74124
R36904 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n2 4.55946
R36905 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n38 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n37 4.51815
R36906 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n37 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n7 2.64533
R36907 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n27 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n24 4.45253
R36908 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n46 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n19 4.38232
R36909 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n54 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n53 4.14168
R36910 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n12 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 3.87929
R36911 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n65 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 3.87929
R36912 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n45 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n20 3.83459
R36913 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n43 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n42 3.76521
R36914 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n42 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n9 2.50198
R36915 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n16 3.43953
R36916 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n49 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n48 3.38874
R36917 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n51 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n18 3.28686
R36918 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n48 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n47 3.01226
R36919 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n47 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n10 2.33997
R36920 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n40 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n21 2.73914
R36921 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n44 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n43 2.63579
R36922 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n39 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n9 15.804
R36923 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n53 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n52 2.25932
R36924 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n52 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n8 2.15681
R36925 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n56 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n17 2.19141
R36926 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n39 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n38 1.88285
R36927 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n34 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n7 15.6099
R36928 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n35 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n22 1.64368
R36929 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n16 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 1.52175
R36930 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n25 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.t3 1.50675
R36931 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n58 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n57 1.50638
R36932 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n57 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n6 1.95132
R36933 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 1.37511
R36934 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n15 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 1.1768
R36935 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n34 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n33 1.12991
R36936 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n29 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n5 15.3925
R36937 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n11 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n1 4.58496
R36938 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n4 0.679754
R36939 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n30 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n23 0.548227
R36940 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n61 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH 0.546841
R36941 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n24 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 0.471686
R36942 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 0.468612
R36943 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n29 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n28 0.376971
R36944 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n2 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOH.n0 0.310701
R36945 EF_R2RVCE_0.comparator_0.VOUTANALOG.n49 EF_R2RVCE_0.comparator_0.VOUTANALOG.t9 129.037
R36946 EF_R2RVCE_0.comparator_0.VOUTANALOG.n49 EF_R2RVCE_0.comparator_0.VOUTANALOG.t10 68.9672
R36947 EF_R2RVCE_0.comparator_0.VOUTANALOG.n69 EF_R2RVCE_0.comparator_0.VOUTANALOG.t0 35.3798
R36948 EF_R2RVCE_0.comparator_0.VOUTANALOG.n64 EF_R2RVCE_0.comparator_0.VOUTANALOG.n63 31.4488
R36949 EF_R2RVCE_0.comparator_0.VOUTANALOG.n70 EF_R2RVCE_0.comparator_0.VOUTANALOG.n69 31.4488
R36950 EF_R2RVCE_0.comparator_0.VOUTANALOG.n56 EF_R2RVCE_0.comparator_0.VOUTANALOG.n55 27.5177
R36951 EF_R2RVCE_0.comparator_0.VOUTANALOG.n78 EF_R2RVCE_0.comparator_0.VOUTANALOG.n77 27.5177
R36952 EF_R2RVCE_0.comparator_0.VOUTANALOG.n14 EF_R2RVCE_0.comparator_0.VOUTANALOG.n13 23.5867
R36953 EF_R2RVCE_0.comparator_0.VOUTANALOG.n86 EF_R2RVCE_0.comparator_0.VOUTANALOG.n85 23.5867
R36954 EF_R2RVCE_0.comparator_0.VOUTANALOG.n26 EF_R2RVCE_0.comparator_0.VOUTANALOG.n25 21.6212
R36955 EF_R2RVCE_0.comparator_0.VOUTANALOG.n115 EF_R2RVCE_0.comparator_0.VOUTANALOG.n114 21.6212
R36956 EF_R2RVCE_0.comparator_0.VOUTANALOG.n8 EF_R2RVCE_0.comparator_0.VOUTANALOG.n7 19.6557
R36957 EF_R2RVCE_0.comparator_0.VOUTANALOG.n94 EF_R2RVCE_0.comparator_0.VOUTANALOG.n93 19.6557
R36958 EF_R2RVCE_0.comparator_0.VOUTANALOG.n34 EF_R2RVCE_0.comparator_0.VOUTANALOG.n33 17.6902
R36959 EF_R2RVCE_0.comparator_0.VOUTANALOG.n104 EF_R2RVCE_0.comparator_0.VOUTANALOG.n103 17.6902
R36960 EF_R2RVCE_0.comparator_0.VOUTANALOG.n33 EF_R2RVCE_0.comparator_0.VOUTANALOG.n32 15.7246
R36961 EF_R2RVCE_0.comparator_0.VOUTANALOG.n103 EF_R2RVCE_0.comparator_0.VOUTANALOG.n102 15.7246
R36962 EF_R2RVCE_0.comparator_0.VOUTANALOG.n9 EF_R2RVCE_0.comparator_0.VOUTANALOG.n8 13.7591
R36963 EF_R2RVCE_0.comparator_0.VOUTANALOG.n95 EF_R2RVCE_0.comparator_0.VOUTANALOG.n94 13.7591
R36964 EF_R2RVCE_0.comparator_0.VOUTANALOG.n25 EF_R2RVCE_0.comparator_0.VOUTANALOG.n24 11.7936
R36965 EF_R2RVCE_0.comparator_0.VOUTANALOG.n114 EF_R2RVCE_0.comparator_0.VOUTANALOG.n113 11.7936
R36966 EF_R2RVCE_0.comparator_0.VOUTANALOG.n15 EF_R2RVCE_0.comparator_0.VOUTANALOG.n14 9.82809
R36967 EF_R2RVCE_0.comparator_0.VOUTANALOG.n87 EF_R2RVCE_0.comparator_0.VOUTANALOG.n86 9.82809
R36968 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n51 9.31585
R36969 EF_R2RVCE_0.comparator_0.VOUTANALOG.n117 EF_R2RVCE_0.comparator_0.VOUTANALOG.n118 9.3005
R36970 EF_R2RVCE_0.comparator_0.VOUTANALOG.n107 EF_R2RVCE_0.comparator_0.VOUTANALOG.n106 9.3005
R36971 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n97 9.3005
R36972 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n89 9.3005
R36973 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n81 9.3005
R36974 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n73 9.3005
R36975 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n60 9.3005
R36976 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n52 9.3005
R36977 EF_R2RVCE_0.comparator_0.VOUTANALOG.n3 EF_R2RVCE_0.comparator_0.VOUTANALOG.n16 9.3005
R36978 EF_R2RVCE_0.comparator_0.VOUTANALOG.n3 EF_R2RVCE_0.comparator_0.VOUTANALOG.n37 9.3005
R36979 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n29 9.3005
R36980 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n21 9.3005
R36981 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n20 9.3005
R36982 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n27 9.3005
R36983 EF_R2RVCE_0.comparator_0.VOUTANALOG.n27 EF_R2RVCE_0.comparator_0.VOUTANALOG.n26 9.3005
R36984 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n28 9.3005
R36985 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n35 9.3005
R36986 EF_R2RVCE_0.comparator_0.VOUTANALOG.n35 EF_R2RVCE_0.comparator_0.VOUTANALOG.n34 9.3005
R36987 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n36 9.3005
R36988 EF_R2RVCE_0.comparator_0.VOUTANALOG.n3 EF_R2RVCE_0.comparator_0.VOUTANALOG.n10 9.3005
R36989 EF_R2RVCE_0.comparator_0.VOUTANALOG.n10 EF_R2RVCE_0.comparator_0.VOUTANALOG.n9 9.3005
R36990 EF_R2RVCE_0.comparator_0.VOUTANALOG.n3 EF_R2RVCE_0.comparator_0.VOUTANALOG.n17 9.3005
R36991 EF_R2RVCE_0.comparator_0.VOUTANALOG.n4 EF_R2RVCE_0.comparator_0.VOUTANALOG.n15 9.3005
R36992 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n58 9.3005
R36993 EF_R2RVCE_0.comparator_0.VOUTANALOG.n58 EF_R2RVCE_0.comparator_0.VOUTANALOG.n57 9.3005
R36994 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n59 9.3005
R36995 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n66 9.3005
R36996 EF_R2RVCE_0.comparator_0.VOUTANALOG.n66 EF_R2RVCE_0.comparator_0.VOUTANALOG.n65 9.3005
R36997 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n72 9.3005
R36998 EF_R2RVCE_0.comparator_0.VOUTANALOG.n72 EF_R2RVCE_0.comparator_0.VOUTANALOG.n71 9.3005
R36999 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 EF_R2RVCE_0.comparator_0.VOUTANALOG.n74 9.3005
R37000 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n80 9.3005
R37001 EF_R2RVCE_0.comparator_0.VOUTANALOG.n80 EF_R2RVCE_0.comparator_0.VOUTANALOG.n79 9.3005
R37002 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n82 9.3005
R37003 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n88 9.3005
R37004 EF_R2RVCE_0.comparator_0.VOUTANALOG.n88 EF_R2RVCE_0.comparator_0.VOUTANALOG.n87 9.3005
R37005 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n90 9.3005
R37006 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n96 9.3005
R37007 EF_R2RVCE_0.comparator_0.VOUTANALOG.n96 EF_R2RVCE_0.comparator_0.VOUTANALOG.n95 9.3005
R37008 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n98 9.3005
R37009 EF_R2RVCE_0.comparator_0.VOUTANALOG.n99 EF_R2RVCE_0.comparator_0.VOUTANALOG.n105 9.3005
R37010 EF_R2RVCE_0.comparator_0.VOUTANALOG.n105 EF_R2RVCE_0.comparator_0.VOUTANALOG.n104 9.3005
R37011 EF_R2RVCE_0.comparator_0.VOUTANALOG.n108 EF_R2RVCE_0.comparator_0.VOUTANALOG.n109 9.3005
R37012 EF_R2RVCE_0.comparator_0.VOUTANALOG.n110 EF_R2RVCE_0.comparator_0.VOUTANALOG.n116 9.3005
R37013 EF_R2RVCE_0.comparator_0.VOUTANALOG.n116 EF_R2RVCE_0.comparator_0.VOUTANALOG.n115 9.3005
R37014 EF_R2RVCE_0.comparator_0.VOUTANALOG.n120 EF_R2RVCE_0.comparator_0.VOUTANALOG.n119 9.3005
R37015 EF_R2RVCE_0.comparator_0.VOUTANALOG.n139 EF_R2RVCE_0.comparator_0.VOUTANALOG.n137 8.0439
R37016 EF_R2RVCE_0.comparator_0.VOUTANALOG.n173 EF_R2RVCE_0.comparator_0.VOUTANALOG.n172 7.45281
R37017 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n19 6.4629
R37018 EF_R2RVCE_0.comparator_0.VOUTANALOG.n121 EF_R2RVCE_0.comparator_0.VOUTANALOG.n50 6.44763
R37019 EF_R2RVCE_0.comparator_0.VOUTANALOG.n62 EF_R2RVCE_0.comparator_0.VOUTANALOG.n61 6.02403
R37020 EF_R2RVCE_0.comparator_0.VOUTANALOG.n68 EF_R2RVCE_0.comparator_0.VOUTANALOG.n67 6.02403
R37021 EF_R2RVCE_0.comparator_0.VOUTANALOG.n57 EF_R2RVCE_0.comparator_0.VOUTANALOG.n56 5.89705
R37022 EF_R2RVCE_0.comparator_0.VOUTANALOG.n79 EF_R2RVCE_0.comparator_0.VOUTANALOG.n78 5.89705
R37023 EF_R2RVCE_0.comparator_0.VOUTANALOG.n130 EF_R2RVCE_0.comparator_0.VOUTANALOG.n128 5.63
R37024 EF_R2RVCE_0.comparator_0.VOUTANALOG.n131 EF_R2RVCE_0.comparator_0.VOUTANALOG.t8 5.5395
R37025 EF_R2RVCE_0.comparator_0.VOUTANALOG.n131 EF_R2RVCE_0.comparator_0.VOUTANALOG.t7 5.5395
R37026 EF_R2RVCE_0.comparator_0.VOUTANALOG.n179 EF_R2RVCE_0.comparator_0.VOUTANALOG.t1 5.5395
R37027 EF_R2RVCE_0.comparator_0.VOUTANALOG.n179 EF_R2RVCE_0.comparator_0.VOUTANALOG.t2 5.5395
R37028 EF_R2RVCE_0.comparator_0.VOUTANALOG.n54 EF_R2RVCE_0.comparator_0.VOUTANALOG.n53 5.27109
R37029 EF_R2RVCE_0.comparator_0.VOUTANALOG.n76 EF_R2RVCE_0.comparator_0.VOUTANALOG.n75 5.27109
R37030 EF_R2RVCE_0.comparator_0.VOUTANALOG.n48 EF_R2RVCE_0.comparator_0.VOUTANALOG.n178 4.7471
R37031 EF_R2RVCE_0.comparator_0.VOUTANALOG.n12 EF_R2RVCE_0.comparator_0.VOUTANALOG.n11 4.51815
R37032 EF_R2RVCE_0.comparator_0.VOUTANALOG.n84 EF_R2RVCE_0.comparator_0.VOUTANALOG.n83 4.51815
R37033 EF_R2RVCE_0.comparator_0.VOUTANALOG.n47 EF_R2RVCE_0.comparator_0.VOUTANALOG.n134 4.5005
R37034 EF_R2RVCE_0.comparator_0.VOUTANALOG.n46 EF_R2RVCE_0.comparator_0.VOUTANALOG.n126 4.5005
R37035 EF_R2RVCE_0.comparator_0.VOUTANALOG.n140 EF_R2RVCE_0.comparator_0.VOUTANALOG.n145 4.5005
R37036 EF_R2RVCE_0.comparator_0.VOUTANALOG.n141 EF_R2RVCE_0.comparator_0.VOUTANALOG.n139 4.5005
R37037 EF_R2RVCE_0.comparator_0.VOUTANALOG.n155 EF_R2RVCE_0.comparator_0.VOUTANALOG.n157 4.5005
R37038 EF_R2RVCE_0.comparator_0.VOUTANALOG.n150 EF_R2RVCE_0.comparator_0.VOUTANALOG.n154 4.5005
R37039 EF_R2RVCE_0.comparator_0.VOUTANALOG.n164 EF_R2RVCE_0.comparator_0.VOUTANALOG.n162 4.5005
R37040 EF_R2RVCE_0.comparator_0.VOUTANALOG.n163 EF_R2RVCE_0.comparator_0.VOUTANALOG.n173 4.5005
R37041 EF_R2RVCE_0.comparator_0.VOUTANALOG.n174 EF_R2RVCE_0.comparator_0.VOUTANALOG.n177 4.5005
R37042 EF_R2RVCE_0.comparator_0.VOUTANALOG.n166 EF_R2RVCE_0.comparator_0.VOUTANALOG.n170 4.5005
R37043 EF_R2RVCE_0.comparator_0.VOUTANALOG.n159 EF_R2RVCE_0.comparator_0.VOUTANALOG.n158 4.3695
R37044 EF_R2RVCE_0.comparator_0.VOUTANALOG.n154 EF_R2RVCE_0.comparator_0.VOUTANALOG.n152 4.14168
R37045 EF_R2RVCE_0.comparator_0.VOUTANALOG.n27 EF_R2RVCE_0.comparator_0.VOUTANALOG.n23 4.14168
R37046 EF_R2RVCE_0.comparator_0.VOUTANALOG.n116 EF_R2RVCE_0.comparator_0.VOUTANALOG.n112 4.14168
R37047 EF_R2RVCE_0.comparator_0.VOUTANALOG.n177 EF_R2RVCE_0.comparator_0.VOUTANALOG.n175 4.14168
R37048 EF_R2RVCE_0.comparator_0.VOUTANALOG.n134 EF_R2RVCE_0.comparator_0.VOUTANALOG.n133 3.76521
R37049 EF_R2RVCE_0.comparator_0.VOUTANALOG.n157 EF_R2RVCE_0.comparator_0.VOUTANALOG.n156 3.76521
R37050 EF_R2RVCE_0.comparator_0.VOUTANALOG.n145 EF_R2RVCE_0.comparator_0.VOUTANALOG.n142 3.76521
R37051 EF_R2RVCE_0.comparator_0.VOUTANALOG.n6 EF_R2RVCE_0.comparator_0.VOUTANALOG.n5 3.76521
R37052 EF_R2RVCE_0.comparator_0.VOUTANALOG.n92 EF_R2RVCE_0.comparator_0.VOUTANALOG.n91 3.76521
R37053 EF_R2RVCE_0.comparator_0.VOUTANALOG.n162 EF_R2RVCE_0.comparator_0.VOUTANALOG.n160 3.75958
R37054 EF_R2RVCE_0.comparator_0.VOUTANALOG.n126 EF_R2RVCE_0.comparator_0.VOUTANALOG.n123 3.38874
R37055 EF_R2RVCE_0.comparator_0.VOUTANALOG.n139 EF_R2RVCE_0.comparator_0.VOUTANALOG.n138 3.38874
R37056 EF_R2RVCE_0.comparator_0.VOUTANALOG.n35 EF_R2RVCE_0.comparator_0.VOUTANALOG.n31 3.38874
R37057 EF_R2RVCE_0.comparator_0.VOUTANALOG.n105 EF_R2RVCE_0.comparator_0.VOUTANALOG.n101 3.38874
R37058 EF_R2RVCE_0.comparator_0.VOUTANALOG.n170 EF_R2RVCE_0.comparator_0.VOUTANALOG.n167 3.38874
R37059 EF_R2RVCE_0.comparator_0.VOUTANALOG.n45 EF_R2RVCE_0.comparator_0.VOUTANALOG.n44 3.38238
R37060 EF_R2RVCE_0.comparator_0.VOUTANALOG.n148 EF_R2RVCE_0.comparator_0.VOUTANALOG.t3 3.3065
R37061 EF_R2RVCE_0.comparator_0.VOUTANALOG.n148 EF_R2RVCE_0.comparator_0.VOUTANALOG.t6 3.3065
R37062 EF_R2RVCE_0.comparator_0.VOUTANALOG.n181 EF_R2RVCE_0.comparator_0.VOUTANALOG.t4 3.3065
R37063 EF_R2RVCE_0.comparator_0.VOUTANALOG.n181 EF_R2RVCE_0.comparator_0.VOUTANALOG.t5 3.3065
R37064 EF_R2RVCE_0.comparator_0.VOUTANALOG.n39 EF_R2RVCE_0.comparator_0.VOUTANALOG.n181 3.21133
R37065 EF_R2RVCE_0.comparator_0.VOUTANALOG.n126 EF_R2RVCE_0.comparator_0.VOUTANALOG.n125 3.01226
R37066 EF_R2RVCE_0.comparator_0.VOUTANALOG.n31 EF_R2RVCE_0.comparator_0.VOUTANALOG.n30 3.01226
R37067 EF_R2RVCE_0.comparator_0.VOUTANALOG.n101 EF_R2RVCE_0.comparator_0.VOUTANALOG.n100 3.01226
R37068 EF_R2RVCE_0.comparator_0.VOUTANALOG.n170 EF_R2RVCE_0.comparator_0.VOUTANALOG.n168 3.01226
R37069 EF_R2RVCE_0.comparator_0.VOUTANALOG.n134 EF_R2RVCE_0.comparator_0.VOUTANALOG.n132 2.63579
R37070 EF_R2RVCE_0.comparator_0.VOUTANALOG.n145 EF_R2RVCE_0.comparator_0.VOUTANALOG.n144 2.63579
R37071 EF_R2RVCE_0.comparator_0.VOUTANALOG.n10 EF_R2RVCE_0.comparator_0.VOUTANALOG.n6 2.63579
R37072 EF_R2RVCE_0.comparator_0.VOUTANALOG.n96 EF_R2RVCE_0.comparator_0.VOUTANALOG.n92 2.63579
R37073 EF_R2RVCE_0.comparator_0.VOUTANALOG.n173 EF_R2RVCE_0.comparator_0.VOUTANALOG.n171 2.63579
R37074 EF_R2RVCE_0.comparator_0.VOUTANALOG.n122 EF_R2RVCE_0.comparator_0.VOUTANALOG.n18 2.48927
R37075 EF_R2RVCE_0.comparator_0.VOUTANALOG.n154 EF_R2RVCE_0.comparator_0.VOUTANALOG.n151 2.25932
R37076 EF_R2RVCE_0.comparator_0.VOUTANALOG.n23 EF_R2RVCE_0.comparator_0.VOUTANALOG.n22 2.25932
R37077 EF_R2RVCE_0.comparator_0.VOUTANALOG.n112 EF_R2RVCE_0.comparator_0.VOUTANALOG.n111 2.25932
R37078 EF_R2RVCE_0.comparator_0.VOUTANALOG.n18 EF_R2RVCE_0.comparator_0.VOUTANALOG.n121 2.22642
R37079 EF_R2RVCE_0.comparator_0.VOUTANALOG.n180 EF_R2RVCE_0.comparator_0.VOUTANALOG.n179 2.1242
R37080 EF_R2RVCE_0.comparator_0.VOUTANALOG.n65 EF_R2RVCE_0.comparator_0.VOUTANALOG.n64 1.96602
R37081 EF_R2RVCE_0.comparator_0.VOUTANALOG.n71 EF_R2RVCE_0.comparator_0.VOUTANALOG.n70 1.96602
R37082 EF_R2RVCE_0.comparator_0.VOUTANALOG.n159 EF_R2RVCE_0.comparator_0.VOUTANALOG.n136 1.95996
R37083 EF_R2RVCE_0.comparator_0.VOUTANALOG.n47 EF_R2RVCE_0.comparator_0.VOUTANALOG.n131 1.90815
R37084 EF_R2RVCE_0.comparator_0.VOUTANALOG.n4 EF_R2RVCE_0.comparator_0.VOUTANALOG.n12 1.88285
R37085 EF_R2RVCE_0.comparator_0.VOUTANALOG.n88 EF_R2RVCE_0.comparator_0.VOUTANALOG.n84 1.88285
R37086 EF_R2RVCE_0.comparator_0.VOUTANALOG.n45 EF_R2RVCE_0.comparator_0.VOUTANALOG.n43 1.88285
R37087 EF_R2RVCE_0.comparator_0.VOUTANALOG EF_R2RVCE_0.comparator_0.VOUTANALOG.n48 1.8055
R37088 EF_R2RVCE_0.comparator_0.VOUTANALOG.n149 EF_R2RVCE_0.comparator_0.VOUTANALOG.n148 1.52639
R37089 EF_R2RVCE_0.comparator_0.VOUTANALOG.n177 EF_R2RVCE_0.comparator_0.VOUTANALOG.n176 1.50638
R37090 EF_R2RVCE_0.comparator_0.VOUTANALOG.n38 EF_R2RVCE_0.comparator_0.VOUTANALOG.n41 6.0005
R37091 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 EF_R2RVCE_0.comparator_0.VOUTANALOG.n18 2.51704
R37092 EF_R2RVCE_0.comparator_0.VOUTANALOG.n135 EF_R2RVCE_0.comparator_0.VOUTANALOG.n47 1.13289
R37093 EF_R2RVCE_0.comparator_0.VOUTANALOG.n58 EF_R2RVCE_0.comparator_0.VOUTANALOG.n54 1.12991
R37094 EF_R2RVCE_0.comparator_0.VOUTANALOG.n80 EF_R2RVCE_0.comparator_0.VOUTANALOG.n76 1.12991
R37095 EF_R2RVCE_0.comparator_0.VOUTANALOG.n41 EF_R2RVCE_0.comparator_0.VOUTANALOG.n40 1.12991
R37096 EF_R2RVCE_0.comparator_0.VOUTANALOG.n150 EF_R2RVCE_0.comparator_0.VOUTANALOG.n149 0.978783
R37097 EF_R2RVCE_0.comparator_0.VOUTANALOG.n166 EF_R2RVCE_0.comparator_0.VOUTANALOG.n165 0.944917
R37098 EF_R2RVCE_0.comparator_0.VOUTANALOG.n146 EF_R2RVCE_0.comparator_0.VOUTANALOG.n147 0.938895
R37099 EF_R2RVCE_0.comparator_0.VOUTANALOG.n48 EF_R2RVCE_0.comparator_0.VOUTANALOG.n182 0.824928
R37100 EF_R2RVCE_0.comparator_0.VOUTANALOG.n43 EF_R2RVCE_0.comparator_0.VOUTANALOG.n42 0.753441
R37101 EF_R2RVCE_0.comparator_0.VOUTANALOG.n182 EF_R2RVCE_0.comparator_0.VOUTANALOG.n39 0.699656
R37102 EF_R2RVCE_0.comparator_0.VOUTANALOG.n48 EF_R2RVCE_0.comparator_0.VOUTANALOG.n159 0.504252
R37103 EF_R2RVCE_0.comparator_0.VOUTANALOG.n66 EF_R2RVCE_0.comparator_0.VOUTANALOG.n62 0.376971
R37104 EF_R2RVCE_0.comparator_0.VOUTANALOG.n72 EF_R2RVCE_0.comparator_0.VOUTANALOG.n68 0.376971
R37105 EF_R2RVCE_0.comparator_0.VOUTANALOG.n178 EF_R2RVCE_0.comparator_0.VOUTANALOG.n180 0.350345
R37106 EF_R2RVCE_0.comparator_0.VOUTANALOG EF_R2RVCE_0.comparator_0.VOUTANALOG.n122 0.327011
R37107 EF_R2RVCE_0.comparator_0.VOUTANALOG.n122 EF_R2RVCE_0.comparator_0.VOUTANALOG.n49 0.289671
R37108 EF_R2RVCE_0.comparator_0.VOUTANALOG.n127 EF_R2RVCE_0.comparator_0.VOUTANALOG.n130 0.278788
R37109 EF_R2RVCE_0.comparator_0.VOUTANALOG.n128 EF_R2RVCE_0.comparator_0.VOUTANALOG.n129 0.161367
R37110 EF_R2RVCE_0.comparator_0.VOUTANALOG.n123 EF_R2RVCE_0.comparator_0.VOUTANALOG.n124 0.150167
R37111 EF_R2RVCE_0.comparator_0.VOUTANALOG.n47 EF_R2RVCE_0.comparator_0.VOUTANALOG.n46 0.143833
R37112 EF_R2RVCE_0.comparator_0.VOUTANALOG.n46 EF_R2RVCE_0.comparator_0.VOUTANALOG.n127 0.1366
R37113 EF_R2RVCE_0.comparator_0.VOUTANALOG.n38 EF_R2RVCE_0.comparator_0.VOUTANALOG.n39 0.0960207
R37114 EF_R2RVCE_0.comparator_0.VOUTANALOG.n164 EF_R2RVCE_0.comparator_0.VOUTANALOG.n163 0.0905088
R37115 EF_R2RVCE_0.comparator_0.VOUTANALOG.n45 EF_R2RVCE_0.comparator_0.VOUTANALOG.n38 6.07651
R37116 EF_R2RVCE_0.comparator_0.VOUTANALOG.n178 EF_R2RVCE_0.comparator_0.VOUTANALOG.n174 0.0722992
R37117 EF_R2RVCE_0.comparator_0.VOUTANALOG.n121 EF_R2RVCE_0.comparator_0.VOUTANALOG.n120 0.061862
R37118 EF_R2RVCE_0.comparator_0.VOUTANALOG.n110 EF_R2RVCE_0.comparator_0.VOUTANALOG.n108 0.058614
R37119 EF_R2RVCE_0.comparator_0.VOUTANALOG.n158 EF_R2RVCE_0.comparator_0.VOUTANALOG.n141 0.0456361
R37120 EF_R2RVCE_0.comparator_0.VOUTANALOG.n141 EF_R2RVCE_0.comparator_0.VOUTANALOG.n140 0.0454219
R37121 EF_R2RVCE_0.comparator_0.VOUTANALOG.n155 EF_R2RVCE_0.comparator_0.VOUTANALOG.n150 0.0454219
R37122 EF_R2RVCE_0.comparator_0.VOUTANALOG.n163 EF_R2RVCE_0.comparator_0.VOUTANALOG.n166 0.0454219
R37123 EF_R2RVCE_0.comparator_0.VOUTANALOG.n174 EF_R2RVCE_0.comparator_0.VOUTANALOG.n164 0.0454219
R37124 EF_R2RVCE_0.comparator_0.VOUTANALOG.n158 EF_R2RVCE_0.comparator_0.VOUTANALOG.n155 0.045375
R37125 EF_R2RVCE_0.comparator_0.VOUTANALOG.n140 EF_R2RVCE_0.comparator_0.VOUTANALOG.n146 0.0439417
R37126 EF_R2RVCE_0.comparator_0.VOUTANALOG.n136 EF_R2RVCE_0.comparator_0.VOUTANALOG.n135 0.028
R37127 EF_R2RVCE_0.comparator_0.VOUTANALOG.n152 EF_R2RVCE_0.comparator_0.VOUTANALOG.n153 0.0189846
R37128 EF_R2RVCE_0.comparator_0.VOUTANALOG.n142 EF_R2RVCE_0.comparator_0.VOUTANALOG.n143 0.0189846
R37129 EF_R2RVCE_0.comparator_0.VOUTANALOG.n117 EF_R2RVCE_0.comparator_0.VOUTANALOG.n110 0.0125614
R37130 EF_R2RVCE_0.comparator_0.VOUTANALOG.n107 EF_R2RVCE_0.comparator_0.VOUTANALOG.n99 0.0103684
R37131 EF_R2RVCE_0.comparator_0.VOUTANALOG.n108 EF_R2RVCE_0.comparator_0.VOUTANALOG.n107 0.00927193
R37132 EF_R2RVCE_0.comparator_0.VOUTANALOG.n120 EF_R2RVCE_0.comparator_0.VOUTANALOG.n117 0.00707895
R37133 EF_R2RVCE_0.comparator_0.VOUTANALOG.n168 EF_R2RVCE_0.comparator_0.VOUTANALOG.n169 0.00688753
R37134 EF_R2RVCE_0.comparator_0.VOUTANALOG.n160 EF_R2RVCE_0.comparator_0.VOUTANALOG.n161 0.00688753
R37135 EF_R2RVCE_0.comparator_0.VOUTANALOG.n3 EF_R2RVCE_0.comparator_0.VOUTANALOG.n4 9.30598
R37136 EF_R2RVCE_0.comparator_0.VOUTANALOG.n3 EF_R2RVCE_0.comparator_0.VOUTANALOG.n2 0.29046
R37137 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 EF_R2RVCE_0.comparator_0.VOUTANALOG.n0 0.234053
R37138 EF_R2RVCE_0.comparator_0.VOUTANALOG.n99 EF_R2RVCE_0.comparator_0.VOUTANALOG.n1 0.230763
R37139 a_4503_2982.n20 a_4503_2982.t9 60.2505
R37140 a_4503_2982.n41 a_4503_2982.t8 60.2505
R37141 a_4503_2982.n63 a_4503_2982.t6 60.2505
R37142 a_4503_2982.n75 a_4503_2982.t4 60.2505
R37143 a_4503_2982.n1 a_4503_2982.n83 9.3005
R37144 a_4503_2982.n1 a_4503_2982.n84 9.3005
R37145 a_4503_2982.n1 a_4503_2982.n82 9.3005
R37146 a_4503_2982.n82 a_4503_2982.n81 9.3005
R37147 a_4503_2982.n2 a_4503_2982.n72 9.3005
R37148 a_4503_2982.n3 a_4503_2982.n56 9.3005
R37149 a_4503_2982.n3 a_4503_2982.n55 9.3005
R37150 a_4503_2982.n3 a_4503_2982.n62 9.3005
R37151 a_4503_2982.n62 a_4503_2982.n61 9.3005
R37152 a_4503_2982.n2 a_4503_2982.n71 9.3005
R37153 a_4503_2982.n71 a_4503_2982.n70 9.3005
R37154 a_4503_2982.n2 a_4503_2982.n73 9.3005
R37155 a_4503_2982.n4 a_4503_2982.n50 9.3005
R37156 a_4503_2982.n5 a_4503_2982.n34 9.3005
R37157 a_4503_2982.n5 a_4503_2982.n33 9.3005
R37158 a_4503_2982.n5 a_4503_2982.n40 9.3005
R37159 a_4503_2982.n40 a_4503_2982.n39 9.3005
R37160 a_4503_2982.n4 a_4503_2982.n49 9.3005
R37161 a_4503_2982.n49 a_4503_2982.n48 9.3005
R37162 a_4503_2982.n4 a_4503_2982.n51 9.3005
R37163 a_4503_2982.n6 a_4503_2982.n28 9.3005
R37164 a_4503_2982.n6 a_4503_2982.n27 9.3005
R37165 a_4503_2982.n27 a_4503_2982.n26 9.3005
R37166 a_4503_2982.n6 a_4503_2982.n29 9.3005
R37167 a_4503_2982.n0 a_4503_2982.n90 9.3005
R37168 a_4503_2982.n120 a_4503_2982.n99 10.743
R37169 a_4503_2982.n64 a_4503_2982.n63 8.76429
R37170 a_4503_2982.n42 a_4503_2982.n41 8.76429
R37171 a_4503_2982.n25 a_4503_2982.n24 7.45411
R37172 a_4503_2982.n38 a_4503_2982.n37 7.45411
R37173 a_4503_2982.n47 a_4503_2982.n46 7.45411
R37174 a_4503_2982.n60 a_4503_2982.n59 7.45411
R37175 a_4503_2982.n69 a_4503_2982.n68 7.45411
R37176 a_4503_2982.n80 a_4503_2982.n79 7.45411
R37177 a_4503_2982.n21 a_4503_2982.n20 6.80105
R37178 a_4503_2982.n76 a_4503_2982.n75 6.80105
R37179 a_4503_2982.n23 a_4503_2982.n22 5.64756
R37180 a_4503_2982.n36 a_4503_2982.n35 5.64756
R37181 a_4503_2982.n45 a_4503_2982.n44 5.64756
R37182 a_4503_2982.n58 a_4503_2982.n57 5.64756
R37183 a_4503_2982.n67 a_4503_2982.n66 5.64756
R37184 a_4503_2982.n78 a_4503_2982.n77 5.64756
R37185 a_4503_2982.n95 a_4503_2982.t7 5.5395
R37186 a_4503_2982.n95 a_4503_2982.t5 5.5395
R37187 a_4503_2982.n89 a_4503_2982.n88 4.95584
R37188 a_4503_2982.n30 a_4503_2982.n19 4.73575
R37189 a_4503_2982.n32 a_4503_2982.n31 4.73575
R37190 a_4503_2982.n52 a_4503_2982.n18 4.73575
R37191 a_4503_2982.n54 a_4503_2982.n53 4.73575
R37192 a_4503_2982.n74 a_4503_2982.n17 4.73575
R37193 a_4503_2982.n86 a_4503_2982.n85 4.73575
R37194 a_4503_2982.n109 a_4503_2982.n12 4.66695
R37195 a_4503_2982.n65 a_4503_2982.n64 4.6505
R37196 a_4503_2982.n43 a_4503_2982.n42 4.6505
R37197 a_4503_2982.n9 a_4503_2982.n104 4.5005
R37198 a_4503_2982.n10 a_4503_2982.n108 4.5005
R37199 a_4503_2982.n0 a_4503_2982.n16 4.5005
R37200 a_4503_2982.n12 a_4503_2982.n98 4.5005
R37201 a_4503_2982.n11 a_4503_2982.n94 4.5005
R37202 a_4503_2982.n7 a_4503_2982.n111 4.5005
R37203 a_4503_2982.n7 a_4503_2982.n113 4.5005
R37204 a_4503_2982.n8 a_4503_2982.n116 4.5005
R37205 a_4503_2982.n108 a_4503_2982.n107 4.14168
R37206 a_4503_2982.n98 a_4503_2982.n97 3.76521
R37207 a_4503_2982.n113 a_4503_2982.n112 3.76521
R37208 a_4503_2982.n6 a_4503_2982.n21 3.42768
R37209 a_4503_2982.n1 a_4503_2982.n76 3.42768
R37210 a_4503_2982.n94 a_4503_2982.n92 3.38874
R37211 a_4503_2982.n16 a_4503_2982.n15 3.38874
R37212 a_4503_2982.n105 a_4503_2982.t2 3.3065
R37213 a_4503_2982.n105 a_4503_2982.t1 3.3065
R37214 a_4503_2982.n120 a_4503_2982.t0 3.3065
R37215 a_4503_2982.t3 a_4503_2982.n120 3.3065
R37216 a_4503_2982.n94 a_4503_2982.n93 3.01226
R37217 a_4503_2982.n16 a_4503_2982.n14 3.01226
R37218 a_4503_2982.n120 a_4503_2982.n119 2.66355
R37219 a_4503_2982.n98 a_4503_2982.n96 2.63579
R37220 a_4503_2982.n103 a_4503_2982.n102 2.25932
R37221 a_4503_2982.n115 a_4503_2982.n114 2.25932
R37222 a_4503_2982.n109 a_4503_2982.n101 1.62138
R37223 a_4503_2982.n120 a_4503_2982.n118 1.46878
R37224 a_4503_2982.n26 a_4503_2982.n25 0.994314
R37225 a_4503_2982.n39 a_4503_2982.n38 0.994314
R37226 a_4503_2982.n48 a_4503_2982.n47 0.994314
R37227 a_4503_2982.n61 a_4503_2982.n60 0.994314
R37228 a_4503_2982.n70 a_4503_2982.n69 0.994314
R37229 a_4503_2982.n81 a_4503_2982.n80 0.994314
R37230 a_4503_2982.n7 a_4503_2982.n109 0.763998
R37231 a_4503_2982.n27 a_4503_2982.n23 0.753441
R37232 a_4503_2982.n40 a_4503_2982.n36 0.753441
R37233 a_4503_2982.n49 a_4503_2982.n45 0.753441
R37234 a_4503_2982.n62 a_4503_2982.n58 0.753441
R37235 a_4503_2982.n71 a_4503_2982.n67 0.753441
R37236 a_4503_2982.n82 a_4503_2982.n78 0.753441
R37237 a_4503_2982.n101 a_4503_2982.n100 0.594417
R37238 a_4503_2982.n9 a_4503_2982.n105 2.11614
R37239 a_4503_2982.n118 a_4503_2982.n117 0.555026
R37240 a_4503_2982.n32 a_4503_2982.n30 0.458354
R37241 a_4503_2982.n54 a_4503_2982.n52 0.458354
R37242 a_4503_2982.n12 a_4503_2982.n95 1.90913
R37243 a_4503_2982.n108 a_4503_2982.n106 0.376971
R37244 a_4503_2982.n104 a_4503_2982.n103 0.376971
R37245 a_4503_2982.n111 a_4503_2982.n110 0.376971
R37246 a_4503_2982.n116 a_4503_2982.n115 0.376971
R37247 a_4503_2982.n87 a_4503_2982.n74 0.229427
R37248 a_4503_2982.n87 a_4503_2982.n86 0.229427
R37249 a_4503_2982.n89 a_4503_2982.n87 0.215848
R37250 a_4503_2982.n30 a_4503_2982.n6 0.205546
R37251 a_4503_2982.n5 a_4503_2982.n32 0.205546
R37252 a_4503_2982.n52 a_4503_2982.n4 0.205546
R37253 a_4503_2982.n3 a_4503_2982.n54 0.205546
R37254 a_4503_2982.n74 a_4503_2982.n2 0.205546
R37255 a_4503_2982.n86 a_4503_2982.n1 0.205546
R37256 a_4503_2982.n43 a_4503_2982.n5 0.190717
R37257 a_4503_2982.n4 a_4503_2982.n43 0.190717
R37258 a_4503_2982.n65 a_4503_2982.n3 0.190717
R37259 a_4503_2982.n2 a_4503_2982.n65 0.190717
R37260 a_4503_2982.n11 a_4503_2982.n0 0.169804
R37261 a_4503_2982.n14 a_4503_2982.n13 0.161367
R37262 a_4503_2982.n92 a_4503_2982.n91 0.150167
R37263 a_4503_2982.n0 a_4503_2982.n89 0.140745
R37264 a_4503_2982.n12 a_4503_2982.n11 0.14187
R37265 a_4503_2982.n8 a_4503_2982.n7 0.135023
R37266 a_4503_2982.n101 a_4503_2982.n10 0.116464
R37267 a_4503_2982.n117 a_4503_2982.n8 0.094364
R37268 a_4503_2982.n10 a_4503_2982.n9 0.0905048
R37269 EN.n0 EN.t1 186.374
R37270 EN.n0 EN.t0 170.308
R37271 EN.n1 EN 101.761
R37272 EN.n2 EN.n1 101.561
R37273 EN.n1 EN.n0 77.4126
R37274 EN.n4 EN.n3 6.39139
R37275 EN.n3 EN.n2 3.02951
R37276 EN.n2 EN 2.24783
R37277 EN.n3 EN 1.9547
R37278 EN EN.n4 0.878376
R37279 EN.n4 EN 0.0508071
R37280 a_6809_n9511.n10 a_6809_n9511.t2 120.01
R37281 a_6809_n9511.n3 a_6809_n9511.t5 92.9415
R37282 a_6809_n9511.n9 a_6809_n9511.n8 92.5005
R37283 a_6809_n9511.n3 a_6809_n9511.t4 92.4623
R37284 a_6809_n9511.n22 a_6809_n9511.t6 73.195
R37285 a_6809_n9511.n22 a_6809_n9511.t3 72.1651
R37286 a_6809_n9511.n17 a_6809_n9511.n16 29.4833
R37287 a_6809_n9511.n26 a_6809_n9511.t0 27.6955
R37288 a_6809_n9511.t1 a_6809_n9511.n41 27.6955
R37289 a_6809_n9511.n10 a_6809_n9511.n9 15.4607
R37290 a_6809_n9511.n0 a_6809_n9511.n12 9.3005
R37291 a_6809_n9511.n0 a_6809_n9511.n19 9.3005
R37292 a_6809_n9511.n0 a_6809_n9511.n18 9.3005
R37293 a_6809_n9511.n18 a_6809_n9511.n17 9.3005
R37294 a_6809_n9511.n0 a_6809_n9511.n11 9.3005
R37295 a_6809_n9511.n0 a_6809_n9511.n21 9.3005
R37296 a_6809_n9511.n0 a_6809_n9511.n20 9.3005
R37297 a_6809_n9511.n41 a_6809_n9511.n40 9.02061
R37298 a_6809_n9511.n41 a_6809_n9511.n7 9.02061
R37299 a_6809_n9511.n27 a_6809_n9511.n26 9.01961
R37300 a_6809_n9511.n25 a_6809_n9511.n23 8.28285
R37301 a_6809_n9511.n34 a_6809_n9511.n35 8.28285
R37302 a_6809_n9511.n18 a_6809_n9511.n14 5.64756
R37303 a_6809_n9511.n2 a_6809_n9511.n25 5.32161
R37304 a_6809_n9511.n2 a_6809_n9511.n29 5.31894
R37305 a_6809_n9511.n29 a_6809_n9511.n28 4.14168
R37306 a_6809_n9511.n39 a_6809_n9511.n38 4.14168
R37307 a_6809_n9511.n2 a_6809_n9511.n3 4.03426
R37308 a_6809_n9511.n16 a_6809_n9511.n15 3.93153
R37309 a_6809_n9511.n32 a_6809_n9511.n30 3.76521
R37310 a_6809_n9511.n6 a_6809_n9511.n5 3.76521
R37311 a_6809_n9511.n3 a_6809_n9511.n22 3.20519
R37312 a_6809_n9511.n1 a_6809_n9511.n34 3.11223
R37313 a_6809_n9511.n33 a_6809_n9511.n32 3.04478
R37314 a_6809_n9511.n39 a_6809_n9511.n1 3.03311
R37315 a_6809_n9511.n1 a_6809_n9511.n36 3.03311
R37316 a_6809_n9511.n25 a_6809_n9511.n24 3.01226
R37317 a_6809_n9511.n32 a_6809_n9511.n31 2.63579
R37318 a_6809_n9511.n7 a_6809_n9511.n6 2.63579
R37319 a_6809_n9511.n1 a_6809_n9511.n2 2.47579
R37320 a_6809_n9511.n2 a_6809_n9511.n33 2.27623
R37321 a_6809_n9511.n29 a_6809_n9511.n27 2.25932
R37322 a_6809_n9511.n40 a_6809_n9511.n39 2.25932
R37323 a_6809_n9511.n1 a_6809_n9511.n0 1.9858
R37324 a_6809_n9511.n5 a_6809_n9511.n4 1.88285
R37325 a_6809_n9511.n0 a_6809_n9511.n10 1.64258
R37326 a_6809_n9511.n14 a_6809_n9511.n13 0.753441
R37327 a_6809_n9511.n38 a_6809_n9511.n37 0.376971
R37328 a_211_n9515.n19 a_211_n9515.t2 120.01
R37329 a_211_n9515.n3 a_211_n9515.t4 92.9415
R37330 a_211_n9515.n18 a_211_n9515.n17 92.5005
R37331 a_211_n9515.n3 a_211_n9515.t3 92.4623
R37332 a_211_n9515.n10 a_211_n9515.t6 73.195
R37333 a_211_n9515.n10 a_211_n9515.t5 72.1651
R37334 a_211_n9515.n26 a_211_n9515.n25 29.4833
R37335 a_211_n9515.n14 a_211_n9515.t0 27.6955
R37336 a_211_n9515.t1 a_211_n9515.n43 27.6955
R37337 a_211_n9515.n19 a_211_n9515.n18 15.4607
R37338 a_211_n9515.n0 a_211_n9515.n21 9.3005
R37339 a_211_n9515.n0 a_211_n9515.n28 9.3005
R37340 a_211_n9515.n0 a_211_n9515.n27 9.3005
R37341 a_211_n9515.n27 a_211_n9515.n26 9.3005
R37342 a_211_n9515.n0 a_211_n9515.n20 9.3005
R37343 a_211_n9515.n0 a_211_n9515.n30 9.3005
R37344 a_211_n9515.n0 a_211_n9515.n29 9.3005
R37345 a_211_n9515.n43 a_211_n9515.n42 9.02061
R37346 a_211_n9515.n43 a_211_n9515.n7 9.02061
R37347 a_211_n9515.n15 a_211_n9515.n14 9.01961
R37348 a_211_n9515.n33 a_211_n9515.n31 8.28285
R37349 a_211_n9515.n38 a_211_n9515.n39 8.28285
R37350 a_211_n9515.n27 a_211_n9515.n23 5.64756
R37351 a_211_n9515.n11 a_211_n9515.n33 5.32317
R37352 a_211_n9515.n12 a_211_n9515.n16 4.14168
R37353 a_211_n9515.n41 a_211_n9515.n9 4.14168
R37354 a_211_n9515.n2 a_211_n9515.n3 4.03426
R37355 a_211_n9515.n25 a_211_n9515.n24 3.93153
R37356 a_211_n9515.n36 a_211_n9515.n34 3.76521
R37357 a_211_n9515.n6 a_211_n9515.n5 3.76521
R37358 a_211_n9515.n3 a_211_n9515.n10 3.20519
R37359 a_211_n9515.n1 a_211_n9515.n38 3.10911
R37360 a_211_n9515.n13 a_211_n9515.n12 3.07353
R37361 a_211_n9515.n37 a_211_n9515.n36 3.04526
R37362 a_211_n9515.n1 a_211_n9515.n40 3.03311
R37363 a_211_n9515.n41 a_211_n9515.n1 3.03311
R37364 a_211_n9515.n33 a_211_n9515.n32 3.01226
R37365 a_211_n9515.n36 a_211_n9515.n35 2.63579
R37366 a_211_n9515.n7 a_211_n9515.n6 2.63579
R37367 a_211_n9515.n1 a_211_n9515.n2 2.32466
R37368 a_211_n9515.n11 a_211_n9515.n37 2.27176
R37369 a_211_n9515.n12 a_211_n9515.n15 2.25932
R37370 a_211_n9515.n42 a_211_n9515.n41 2.25932
R37371 a_211_n9515.n11 a_211_n9515.n13 2.2484
R37372 a_211_n9515.n13 a_211_n9515.n0 1.90545
R37373 a_211_n9515.n5 a_211_n9515.n4 1.88285
R37374 a_211_n9515.n0 a_211_n9515.n19 1.64258
R37375 a_211_n9515.n23 a_211_n9515.n22 0.753441
R37376 a_211_n9515.n9 a_211_n9515.n8 0.376971
R37377 a_211_n9515.n2 a_211_n9515.n11 0.227894
R37378 a_1355_5983.n34 a_1355_5983.t9 60.2505
R37379 a_1355_5983.n56 a_1355_5983.t8 60.2505
R37380 a_1355_5983.n79 a_1355_5983.t2 60.2505
R37381 a_1355_5983.n22 a_1355_5983.t0 60.2505
R37382 a_1355_5983.n1 a_1355_5983.n43 9.3005
R37383 a_1355_5983.n2 a_1355_5983.n48 9.3005
R37384 a_1355_5983.n3 a_1355_5983.n66 9.3005
R37385 a_1355_5983.n4 a_1355_5983.n71 9.3005
R37386 a_1355_5983.n5 a_1355_5983.n89 9.3005
R37387 a_1355_5983.n6 a_1355_5983.n31 9.3005
R37388 a_1355_5983.n6 a_1355_5983.n30 9.3005
R37389 a_1355_5983.n6 a_1355_5983.n29 9.3005
R37390 a_1355_5983.n29 a_1355_5983.n28 9.3005
R37391 a_1355_5983.n5 a_1355_5983.n88 9.3005
R37392 a_1355_5983.n5 a_1355_5983.n87 9.3005
R37393 a_1355_5983.n87 a_1355_5983.n86 9.3005
R37394 a_1355_5983.n4 a_1355_5983.n72 9.3005
R37395 a_1355_5983.n4 a_1355_5983.n78 9.3005
R37396 a_1355_5983.n78 a_1355_5983.n77 9.3005
R37397 a_1355_5983.n3 a_1355_5983.n65 9.3005
R37398 a_1355_5983.n3 a_1355_5983.n64 9.3005
R37399 a_1355_5983.n64 a_1355_5983.n63 9.3005
R37400 a_1355_5983.n2 a_1355_5983.n49 9.3005
R37401 a_1355_5983.n2 a_1355_5983.n55 9.3005
R37402 a_1355_5983.n55 a_1355_5983.n54 9.3005
R37403 a_1355_5983.n1 a_1355_5983.n41 9.3005
R37404 a_1355_5983.n41 a_1355_5983.n40 9.3005
R37405 a_1355_5983.n1 a_1355_5983.n42 9.3005
R37406 a_1355_5983.n0 a_1355_5983.n95 9.3005
R37407 a_1355_5983.n121 a_1355_5983.n100 10.743
R37408 a_1355_5983.n80 a_1355_5983.n79 8.76429
R37409 a_1355_5983.n57 a_1355_5983.n56 8.76429
R37410 a_1355_5983.n27 a_1355_5983.n26 7.45411
R37411 a_1355_5983.n85 a_1355_5983.n84 7.45411
R37412 a_1355_5983.n76 a_1355_5983.n75 7.45411
R37413 a_1355_5983.n62 a_1355_5983.n61 7.45411
R37414 a_1355_5983.n53 a_1355_5983.n52 7.45411
R37415 a_1355_5983.n39 a_1355_5983.n38 7.45411
R37416 a_1355_5983.n23 a_1355_5983.n22 6.80334
R37417 a_1355_5983.n35 a_1355_5983.n34 6.80105
R37418 a_1355_5983.n25 a_1355_5983.n24 5.64756
R37419 a_1355_5983.n83 a_1355_5983.n82 5.64756
R37420 a_1355_5983.n74 a_1355_5983.n73 5.64756
R37421 a_1355_5983.n60 a_1355_5983.n59 5.64756
R37422 a_1355_5983.n51 a_1355_5983.n50 5.64756
R37423 a_1355_5983.n37 a_1355_5983.n36 5.64756
R37424 a_1355_5983.n96 a_1355_5983.t1 5.5395
R37425 a_1355_5983.n96 a_1355_5983.t3 5.5395
R37426 a_1355_5983.n94 a_1355_5983.n93 4.95584
R37427 a_1355_5983.n33 a_1355_5983.n32 4.73575
R37428 a_1355_5983.n91 a_1355_5983.n90 4.73575
R37429 a_1355_5983.n70 a_1355_5983.n69 4.73575
R37430 a_1355_5983.n68 a_1355_5983.n67 4.73575
R37431 a_1355_5983.n47 a_1355_5983.n46 4.73575
R37432 a_1355_5983.n45 a_1355_5983.n44 4.73575
R37433 a_1355_5983.n11 a_1355_5983.n13 4.66506
R37434 a_1355_5983.n81 a_1355_5983.n80 4.6505
R37435 a_1355_5983.n58 a_1355_5983.n57 4.6505
R37436 a_1355_5983.n7 a_1355_5983.n108 4.5005
R37437 a_1355_5983.n8 a_1355_5983.n105 4.5005
R37438 a_1355_5983.n0 a_1355_5983.n21 4.5005
R37439 a_1355_5983.n13 a_1355_5983.n99 4.5005
R37440 a_1355_5983.n12 a_1355_5983.n17 4.5005
R37441 a_1355_5983.n10 a_1355_5983.n118 4.5005
R37442 a_1355_5983.n9 a_1355_5983.n113 4.5005
R37443 a_1355_5983.n9 a_1355_5983.n115 4.5005
R37444 a_1355_5983.n105 a_1355_5983.n104 4.14168
R37445 a_1355_5983.n99 a_1355_5983.n98 3.76521
R37446 a_1355_5983.n115 a_1355_5983.n114 3.76521
R37447 a_1355_5983.n1 a_1355_5983.n35 3.42768
R37448 a_1355_5983.n6 a_1355_5983.n23 3.42683
R37449 a_1355_5983.n17 a_1355_5983.n15 3.38874
R37450 a_1355_5983.n21 a_1355_5983.n20 3.38874
R37451 a_1355_5983.n109 a_1355_5983.t5 3.3065
R37452 a_1355_5983.n109 a_1355_5983.t6 3.3065
R37453 a_1355_5983.t7 a_1355_5983.n121 3.3065
R37454 a_1355_5983.n121 a_1355_5983.t4 3.3065
R37455 a_1355_5983.n17 a_1355_5983.n16 3.01226
R37456 a_1355_5983.n21 a_1355_5983.n19 3.01226
R37457 a_1355_5983.n121 a_1355_5983.n101 2.66355
R37458 a_1355_5983.n99 a_1355_5983.n97 2.63579
R37459 a_1355_5983.n107 a_1355_5983.n106 2.25932
R37460 a_1355_5983.n117 a_1355_5983.n116 2.25932
R37461 a_1355_5983.n121 a_1355_5983.n120 1.4688
R37462 a_1355_5983.n13 a_1355_5983.n96 1.90914
R37463 a_1355_5983.n28 a_1355_5983.n27 0.994314
R37464 a_1355_5983.n86 a_1355_5983.n85 0.994314
R37465 a_1355_5983.n77 a_1355_5983.n76 0.994314
R37466 a_1355_5983.n63 a_1355_5983.n62 0.994314
R37467 a_1355_5983.n54 a_1355_5983.n53 0.994314
R37468 a_1355_5983.n40 a_1355_5983.n39 0.994314
R37469 a_1355_5983.n111 a_1355_5983.n102 0.920917
R37470 a_1355_5983.n9 a_1355_5983.n11 0.764358
R37471 a_1355_5983.n29 a_1355_5983.n25 0.753441
R37472 a_1355_5983.n87 a_1355_5983.n83 0.753441
R37473 a_1355_5983.n78 a_1355_5983.n74 0.753441
R37474 a_1355_5983.n64 a_1355_5983.n60 0.753441
R37475 a_1355_5983.n55 a_1355_5983.n51 0.753441
R37476 a_1355_5983.n41 a_1355_5983.n37 0.753441
R37477 a_1355_5983.n11 a_1355_5983.n111 0.700686
R37478 a_1355_5983.n102 a_1355_5983.n110 0.594011
R37479 a_1355_5983.n7 a_1355_5983.n109 2.11687
R37480 a_1355_5983.n120 a_1355_5983.n119 0.555
R37481 a_1355_5983.n70 a_1355_5983.n68 0.458354
R37482 a_1355_5983.n47 a_1355_5983.n45 0.458354
R37483 a_1355_5983.n105 a_1355_5983.n103 0.376971
R37484 a_1355_5983.n108 a_1355_5983.n107 0.376971
R37485 a_1355_5983.n113 a_1355_5983.n112 0.376971
R37486 a_1355_5983.n118 a_1355_5983.n117 0.376971
R37487 a_1355_5983.n92 a_1355_5983.n33 0.229427
R37488 a_1355_5983.n92 a_1355_5983.n91 0.229427
R37489 a_1355_5983.n94 a_1355_5983.n92 0.215848
R37490 a_1355_5983.n33 a_1355_5983.n6 0.205546
R37491 a_1355_5983.n91 a_1355_5983.n5 0.205546
R37492 a_1355_5983.n4 a_1355_5983.n70 0.205546
R37493 a_1355_5983.n68 a_1355_5983.n3 0.205546
R37494 a_1355_5983.n2 a_1355_5983.n47 0.205546
R37495 a_1355_5983.n45 a_1355_5983.n1 0.205546
R37496 a_1355_5983.n5 a_1355_5983.n81 0.190717
R37497 a_1355_5983.n81 a_1355_5983.n4 0.190717
R37498 a_1355_5983.n3 a_1355_5983.n58 0.190717
R37499 a_1355_5983.n58 a_1355_5983.n2 0.190717
R37500 a_1355_5983.n12 a_1355_5983.n0 0.169805
R37501 a_1355_5983.n19 a_1355_5983.n18 0.161367
R37502 a_1355_5983.n15 a_1355_5983.n14 0.150167
R37503 a_1355_5983.n0 a_1355_5983.n94 0.140745
R37504 a_1355_5983.n13 a_1355_5983.n12 0.142842
R37505 a_1355_5983.n10 a_1355_5983.n9 0.135433
R37506 a_1355_5983.n102 a_1355_5983.n8 0.116866
R37507 a_1355_5983.n119 a_1355_5983.n10 0.0933679
R37508 a_1355_5983.n8 a_1355_5983.n7 0.0905048
R37509 a_1755_6080.n76 a_1755_6080.t0 60.2505
R37510 a_1755_6080.n53 a_1755_6080.t7 60.2505
R37511 a_1755_6080.n30 a_1755_6080.t6 60.2505
R37512 a_1755_6080.n90 a_1755_6080.t2 60.2505
R37513 a_1755_6080.n140 a_1755_6080.n10 10.3264
R37514 a_1755_6080.n140 a_1755_6080.n11 9.57347
R37515 a_1755_6080.n7 a_1755_6080.n98 9.3005
R37516 a_1755_6080.n100 a_1755_6080.n99 9.3005
R37517 a_1755_6080.n7 a_1755_6080.n97 9.3005
R37518 a_1755_6080.n97 a_1755_6080.n96 9.3005
R37519 a_1755_6080.n64 a_1755_6080.n63 9.3005
R37520 a_1755_6080.n1 a_1755_6080.n45 9.3005
R37521 a_1755_6080.n40 a_1755_6080.n39 9.3005
R37522 a_1755_6080.n0 a_1755_6080.n38 9.3005
R37523 a_1755_6080.n0 a_1755_6080.n37 9.3005
R37524 a_1755_6080.n37 a_1755_6080.n36 9.3005
R37525 a_1755_6080.n2 a_1755_6080.n46 9.3005
R37526 a_1755_6080.n2 a_1755_6080.n52 9.3005
R37527 a_1755_6080.n52 a_1755_6080.n51 9.3005
R37528 a_1755_6080.n3 a_1755_6080.n62 9.3005
R37529 a_1755_6080.n3 a_1755_6080.n61 9.3005
R37530 a_1755_6080.n61 a_1755_6080.n60 9.3005
R37531 a_1755_6080.n4 a_1755_6080.n68 9.3005
R37532 a_1755_6080.n5 a_1755_6080.n75 9.3005
R37533 a_1755_6080.n75 a_1755_6080.n74 9.3005
R37534 a_1755_6080.n5 a_1755_6080.n69 9.3005
R37535 a_1755_6080.n6 a_1755_6080.n84 9.3005
R37536 a_1755_6080.n84 a_1755_6080.n83 9.3005
R37537 a_1755_6080.n87 a_1755_6080.n86 9.3005
R37538 a_1755_6080.n6 a_1755_6080.n85 9.3005
R37539 a_1755_6080.n112 a_1755_6080.n113 9.3005
R37540 a_1755_6080.n110 a_1755_6080.n111 9.3005
R37541 a_1755_6080.n108 a_1755_6080.n109 9.3005
R37542 a_1755_6080.n106 a_1755_6080.n107 9.3005
R37543 a_1755_6080.n105 a_1755_6080.n104 9.3005
R37544 a_1755_6080.n54 a_1755_6080.n53 8.76429
R37545 a_1755_6080.n77 a_1755_6080.n76 8.76429
R37546 a_1755_6080.n35 a_1755_6080.n34 8.21641
R37547 a_1755_6080.n50 a_1755_6080.n49 8.21641
R37548 a_1755_6080.n59 a_1755_6080.n58 8.21641
R37549 a_1755_6080.n95 a_1755_6080.n94 8.21641
R37550 a_1755_6080.n73 a_1755_6080.n72 8.21641
R37551 a_1755_6080.n82 a_1755_6080.n81 8.21641
R37552 a_1755_6080.n140 a_1755_6080.n27 8.139
R37553 a_1755_6080.n140 a_1755_6080.n24 8.11104
R37554 a_1755_6080.n140 a_1755_6080.n21 8.08351
R37555 a_1755_6080.n140 a_1755_6080.n18 8.05639
R37556 a_1755_6080.n133 a_1755_6080.n132 8.0439
R37557 a_1755_6080.n140 a_1755_6080.n15 8.02969
R37558 a_1755_6080.n140 a_1755_6080.n12 8.00339
R37559 a_1755_6080.n31 a_1755_6080.n30 6.92242
R37560 a_1755_6080.n91 a_1755_6080.n90 6.92012
R37561 a_1755_6080.n33 a_1755_6080.n32 5.64756
R37562 a_1755_6080.n48 a_1755_6080.n47 5.64756
R37563 a_1755_6080.n57 a_1755_6080.n56 5.64756
R37564 a_1755_6080.n93 a_1755_6080.n92 5.64756
R37565 a_1755_6080.n71 a_1755_6080.n70 5.64756
R37566 a_1755_6080.n80 a_1755_6080.n79 5.64756
R37567 a_1755_6080.n122 a_1755_6080.n120 5.62996
R37568 a_1755_6080.n127 a_1755_6080.t5 5.5395
R37569 a_1755_6080.n127 a_1755_6080.t4 5.5395
R37570 a_1755_6080.n42 a_1755_6080.n41 4.76425
R37571 a_1755_6080.n44 a_1755_6080.n43 4.76425
R37572 a_1755_6080.n66 a_1755_6080.n65 4.76425
R37573 a_1755_6080.n101 a_1755_6080.n89 4.76425
R37574 a_1755_6080.n67 a_1755_6080.n29 4.76425
R37575 a_1755_6080.n88 a_1755_6080.n28 4.76425
R37576 a_1755_6080.n55 a_1755_6080.n54 4.6505
R37577 a_1755_6080.n78 a_1755_6080.n77 4.6505
R37578 a_1755_6080.n9 a_1755_6080.n130 4.5005
R37579 a_1755_6080.n8 a_1755_6080.n126 4.5005
R37580 a_1755_6080.n135 a_1755_6080.n137 4.5005
R37581 a_1755_6080.n134 a_1755_6080.n133 4.5005
R37582 a_1755_6080.n117 a_1755_6080.n118 4.5005
R37583 a_1755_6080.n114 a_1755_6080.n116 4.5005
R37584 a_1755_6080.n14 a_1755_6080.n13 4.14168
R37585 a_1755_6080.n130 a_1755_6080.n129 3.76521
R37586 a_1755_6080.n7 a_1755_6080.n91 3.47756
R37587 a_1755_6080.n0 a_1755_6080.n31 3.4767
R37588 a_1755_6080.n126 a_1755_6080.n123 3.38874
R37589 a_1755_6080.n17 a_1755_6080.n16 3.38874
R37590 a_1755_6080.n140 a_1755_6080.t1 3.3065
R37591 a_1755_6080.t3 a_1755_6080.n140 3.3065
R37592 a_1755_6080.n126 a_1755_6080.n125 3.01226
R37593 a_1755_6080.n130 a_1755_6080.n128 2.63579
R37594 a_1755_6080.n20 a_1755_6080.n19 2.63579
R37595 a_1755_6080.n137 a_1755_6080.n136 2.63579
R37596 a_1755_6080.n116 a_1755_6080.n115 2.25932
R37597 a_1755_6080.n9 a_1755_6080.n127 1.90814
R37598 a_1755_6080.n23 a_1755_6080.n22 1.88285
R37599 a_1755_6080.n140 a_1755_6080.n139 1.52638
R37600 a_1755_6080.n26 a_1755_6080.n25 1.12991
R37601 a_1755_6080.n36 a_1755_6080.n35 1.09595
R37602 a_1755_6080.n51 a_1755_6080.n50 1.09595
R37603 a_1755_6080.n60 a_1755_6080.n59 1.09595
R37604 a_1755_6080.n96 a_1755_6080.n95 1.09595
R37605 a_1755_6080.n74 a_1755_6080.n73 1.09595
R37606 a_1755_6080.n83 a_1755_6080.n82 1.09595
R37607 a_1755_6080.n139 a_1755_6080.n138 0.93881
R37608 a_1755_6080.n37 a_1755_6080.n33 0.753441
R37609 a_1755_6080.n52 a_1755_6080.n48 0.753441
R37610 a_1755_6080.n61 a_1755_6080.n57 0.753441
R37611 a_1755_6080.n97 a_1755_6080.n93 0.753441
R37612 a_1755_6080.n75 a_1755_6080.n71 0.753441
R37613 a_1755_6080.n84 a_1755_6080.n80 0.753441
R37614 a_1755_6080.n15 a_1755_6080.n14 0.461175
R37615 a_1755_6080.n44 a_1755_6080.n42 0.458354
R37616 a_1755_6080.n67 a_1755_6080.n66 0.458354
R37617 a_1755_6080.n18 a_1755_6080.n17 0.430121
R37618 a_1755_6080.n21 a_1755_6080.n20 0.398603
R37619 a_1755_6080.n24 a_1755_6080.n23 0.366615
R37620 a_1755_6080.n27 a_1755_6080.n26 0.334147
R37621 a_1755_6080.n119 a_1755_6080.n122 0.27883
R37622 a_1755_6080.n102 a_1755_6080.n88 0.229427
R37623 a_1755_6080.n102 a_1755_6080.n101 0.229427
R37624 a_1755_6080.n103 a_1755_6080.n102 0.191391
R37625 a_1755_6080.n106 a_1755_6080.n105 0.190717
R37626 a_1755_6080.n108 a_1755_6080.n106 0.190717
R37627 a_1755_6080.n110 a_1755_6080.n108 0.190717
R37628 a_1755_6080.n112 a_1755_6080.n110 0.190717
R37629 a_1755_6080.n55 a_1755_6080.n2 0.190717
R37630 a_1755_6080.n3 a_1755_6080.n55 0.190717
R37631 a_1755_6080.n78 a_1755_6080.n5 0.190717
R37632 a_1755_6080.n6 a_1755_6080.n78 0.190717
R37633 a_1755_6080.n114 a_1755_6080.n112 0.169023
R37634 a_1755_6080.n105 a_1755_6080.n103 0.164777
R37635 a_1755_6080.n120 a_1755_6080.n121 0.161367
R37636 a_1755_6080.n42 a_1755_6080.n40 0.15935
R37637 a_1755_6080.n1 a_1755_6080.n44 0.15935
R37638 a_1755_6080.n66 a_1755_6080.n64 0.15935
R37639 a_1755_6080.n4 a_1755_6080.n67 0.15935
R37640 a_1755_6080.n88 a_1755_6080.n87 0.15935
R37641 a_1755_6080.n101 a_1755_6080.n100 0.15935
R37642 a_1755_6080.n123 a_1755_6080.n124 0.150167
R37643 a_1755_6080.n9 a_1755_6080.n8 0.143833
R37644 a_1755_6080.n8 a_1755_6080.n119 0.1366
R37645 a_1755_6080.n100 a_1755_6080.n7 0.0466957
R37646 a_1755_6080.n87 a_1755_6080.n6 0.0466957
R37647 a_1755_6080.n5 a_1755_6080.n4 0.0466957
R37648 a_1755_6080.n64 a_1755_6080.n3 0.0466957
R37649 a_1755_6080.n2 a_1755_6080.n1 0.0466957
R37650 a_1755_6080.n40 a_1755_6080.n0 0.0466957
R37651 a_1755_6080.n134 a_1755_6080.n131 0.0456361
R37652 a_1755_6080.n117 a_1755_6080.n114 0.0454219
R37653 a_1755_6080.n135 a_1755_6080.n134 0.0454219
R37654 a_1755_6080.n131 a_1755_6080.n117 0.045375
R37655 a_1755_6080.n138 a_1755_6080.n135 0.0439417
R37656 a_1755_6080.n131 a_1755_6080.n9 7.51529
R37657 A2.n107 A2.n106 185
R37658 A2.n105 A2.n98 185
R37659 A2.n65 A2.n56 185
R37660 A2.n64 A2.n63 185
R37661 A2.n110 A2.t6 120.037
R37662 A2.t7 A2.n55 120.037
R37663 A2.n100 A2.n98 112.831
R37664 A2.n63 A2.n62 112.831
R37665 A2.n109 A2.n108 104.172
R37666 A2.n68 A2.n67 104.172
R37667 A2.n109 A2.n97 92.5005
R37668 A2.n69 A2.n68 92.5005
R37669 A2.t6 A2.n109 66.8281
R37670 A2.n68 A2.t7 66.8281
R37671 A2.n47 A2.t2 35.2053
R37672 A2.n44 A2.t3 34.0571
R37673 A2.n108 A2.n107 29.4833
R37674 A2.n67 A2.n56 29.4833
R37675 A2.n42 A2.t4 27.6955
R37676 A2.n42 A2.t5 27.6955
R37677 A2.n86 A2.n85 19.0955
R37678 A2.n110 A2.n97 15.4558
R37679 A2.n69 A2.n55 15.4558
R37680 A2.n105 A2.n104 13.5534
R37681 A2.n64 A2.n59 13.5534
R37682 A2.n43 A2.n42 9.67857
R37683 A2.n82 A2.n75 9.30581
R37684 A2.n100 A2.n99 9.30424
R37685 A2.n62 A2.n61 9.30413
R37686 A2.n81 A2.n80 9.3005
R37687 A2.n87 A2.n86 9.3005
R37688 A2.n112 A2.n111 9.3005
R37689 A2.n96 A2.n93 9.3005
R37690 A2.n108 A2.n96 9.3005
R37691 A2.n104 A2.n103 9.3005
R37692 A2.n113 A2.n95 9.3005
R37693 A2.n70 A2.n54 9.3005
R37694 A2.n66 A2.n52 9.3005
R37695 A2.n67 A2.n66 9.3005
R37696 A2.n59 A2.n58 9.3005
R37697 A2.n72 A2.n71 9.3005
R37698 A2.n112 A2.n97 9.03579
R37699 A2.n70 A2.n69 9.03579
R37700 A2.n84 A2.n82 8.49366
R37701 A2.n84 A2.t0 8.2655
R37702 A2.n84 A2.t1 8.2655
R37703 A2.n85 A2.n84 7.97749
R37704 A2.n83 A2.n81 7.26743
R37705 A2.n84 A2.n83 6.15568
R37706 A2.n106 A2.n96 5.64756
R37707 A2.n66 A2.n65 5.64756
R37708 A2.n82 A2.n76 4.89462
R37709 A2.n101 A2.n100 4.89462
R37710 A2.n62 A2.n60 4.89462
R37711 A2.n114 A2.n96 4.51815
R37712 A2.n113 A2.n112 4.51815
R37713 A2.n66 A2.n53 4.51815
R37714 A2.n71 A2.n70 4.51815
R37715 A2.n46 A2.n45 4.5005
R37716 A2.n45 A2.n43 4.5005
R37717 A2.n92 A2.n50 4.5005
R37718 A2.n90 A2.n50 4.5005
R37719 A2.n92 A2.n91 4.5005
R37720 A2.n91 A2.n90 4.5005
R37721 A2.n115 A2.n94 4.5005
R37722 A2.n116 A2.n49 4.5005
R37723 A2.n94 A2.n49 4.5005
R37724 A2.n116 A2.n115 4.5005
R37725 A2.n89 A2.n73 4.5005
R37726 A2.n88 A2.n77 4.5005
R37727 A2.n89 A2.n88 4.5005
R37728 A2.n77 A2.n73 4.5005
R37729 A2.n79 A2.n74 4.5005
R37730 A2.n107 A2.n98 3.93153
R37731 A2.n63 A2.n56 3.93153
R37732 A2.n219 A2 3.5005
R37733 A2.n148 A2 3.1255
R37734 A2.n60 A2.n50 3.03311
R37735 A2.n91 A2.n53 3.03311
R37736 A2.n101 A2.n49 3.03311
R37737 A2.n115 A2.n114 3.03311
R37738 A2.n88 A2.n76 3.03311
R37739 A2.n44 A2.n41 2.2714
R37740 A2.n99 A2.n48 2.25261
R37741 A2.n61 A2.n51 2.25256
R37742 A2.n75 A2.n74 2.25127
R37743 A2.n78 A2.n74 2.24434
R37744 A2.n153 A2.n152 1.94045
R37745 A2.n136 A2.n135 1.94045
R37746 A2.n114 A2.n113 1.88285
R37747 A2.n71 A2.n53 1.88285
R37748 A2.n218 A2.n217 1.72425
R37749 A2.n148 A2 1.563
R37750 A2.n202 A2.n201 1.54186
R37751 A2.n86 A2.n76 1.50638
R37752 A2.n104 A2.n101 1.50638
R37753 A2.n60 A2.n59 1.50638
R37754 A2.n57 A2.n51 1.49213
R37755 A2.n111 A2.n110 1.49212
R37756 A2.n102 A2.n48 1.49182
R37757 A2.n55 A2.n54 1.49166
R37758 A2.n119 A2 1.06297
R37759 A2.n157 A2.n153 0.853
R37760 A2.n200 A2.n199 0.853
R37761 A2.n106 A2.n105 0.753441
R37762 A2.n65 A2.n64 0.753441
R37763 A2.n0 A2 0.744783
R37764 A2.n181 A2.n140 0.690775
R37765 A2.n85 A2.n81 0.521921
R37766 A2.n182 A2.n181 0.513942
R37767 A2.n217 A2.n216 0.326453
R37768 A2.n118 A2.n47 0.29767
R37769 A2.n90 A2.n89 0.238951
R37770 A2.n118 A2.n117 0.196255
R37771 A2 A2.n118 0.1855
R37772 A2.n47 A2.n46 0.149538
R37773 A2.n116 A2.n92 0.124821
R37774 A2.n1 A2.n0 0.0882193
R37775 A2.n2 A2.n1 0.0882193
R37776 A2.n3 A2.n2 0.0882193
R37777 A2.n4 A2.n3 0.0882193
R37778 A2.n5 A2.n4 0.0882193
R37779 A2.n218 A2.n5 0.0882193
R37780 A2.n149 A2.n148 0.0807752
R37781 A2.n219 A2.n218 0.0640965
R37782 A2.n83 A2.n73 0.0579027
R37783 A2.n135 A2.n121 0.0521055
R37784 A2.n135 A2.n134 0.0521055
R37785 A2.n152 A2.n147 0.0521055
R37786 A2.n152 A2.n151 0.0521055
R37787 A2.n103 A2.n102 0.0396286
R37788 A2.n132 A2.n131 0.0394908
R37789 A2.n128 A2.n127 0.0394908
R37790 A2.n124 A2.n123 0.0394908
R37791 A2.n58 A2.n57 0.0383668
R37792 A2.n137 A2.n136 0.0323396
R37793 A2.n136 A2.n40 0.0323396
R37794 A2.n153 A2.n142 0.0323396
R37795 A2.n153 A2.n146 0.0323396
R37796 A2.n87 A2.n78 0.0314092
R37797 A2.n46 A2.n41 0.0281442
R37798 A2.n80 A2.n78 0.0271357
R37799 A2.n139 A2.n138 0.0229057
R37800 A2.n39 A2.n38 0.0229057
R37801 A2.n145 A2.n144 0.0229057
R37802 A2.n121 A2.n120 0.022289
R37803 A2.n134 A2.n133 0.022289
R37804 A2.n151 A2.n150 0.022289
R37805 A2.n138 A2.n137 0.0217264
R37806 A2.n40 A2.n39 0.0217264
R37807 A2.n142 A2.n141 0.0217264
R37808 A2.n146 A2.n145 0.0217264
R37809 A2.n31 A2.n30 0.0205472
R37810 A2.n30 A2.n29 0.0205472
R37811 A2.n217 A2.n21 0.0203617
R37812 A2.n102 A2.n93 0.0202788
R37813 A2.n57 A2.n52 0.0196501
R37814 A2.n36 A2.n35 0.0193679
R37815 A2.n25 A2.n24 0.0193679
R37816 A2.n181 A2.n180 0.0189241
R37817 A2.n34 A2.n33 0.0181887
R37818 A2.n32 A2.n31 0.0181887
R37819 A2.n29 A2.n28 0.0181887
R37820 A2.n27 A2.n26 0.0181887
R37821 A2.n131 A2.n130 0.0177018
R37822 A2.n129 A2.n128 0.0177018
R37823 A2.n127 A2.n126 0.0177018
R37824 A2.n125 A2.n124 0.0177018
R37825 A2.n92 A2.n51 0.0168043
R37826 A2.n203 A2.n202 0.0166506
R37827 A2.n77 A2.n74 0.016125
R37828 A2.n7 A2.n6 0.0138019
R37829 A2.n9 A2.n8 0.0138019
R37830 A2.n10 A2.n9 0.0138019
R37831 A2.n12 A2.n11 0.0138019
R37832 A2.n13 A2.n12 0.0138019
R37833 A2.n15 A2.n14 0.0138019
R37834 A2.n16 A2.n15 0.0138019
R37835 A2.n18 A2.n17 0.0138019
R37836 A2.n19 A2.n18 0.0138019
R37837 A2.n21 A2.n20 0.0138019
R37838 A2.n183 A2.n182 0.0138019
R37839 A2.n185 A2.n184 0.0138019
R37840 A2.n186 A2.n185 0.0138019
R37841 A2.n188 A2.n187 0.0138019
R37842 A2.n189 A2.n188 0.0138019
R37843 A2.n191 A2.n190 0.0138019
R37844 A2.n192 A2.n191 0.0138019
R37845 A2.n194 A2.n193 0.0138019
R37846 A2.n195 A2.n194 0.0138019
R37847 A2.n200 A2.n196 0.0138019
R37848 A2.n201 A2.n200 0.0136459
R37849 A2.n205 A2.n204 0.0135556
R37850 A2.n206 A2.n205 0.0135556
R37851 A2.n208 A2.n207 0.0135556
R37852 A2.n209 A2.n208 0.0135556
R37853 A2.n211 A2.n210 0.0135556
R37854 A2.n212 A2.n211 0.0135556
R37855 A2.n214 A2.n213 0.0135556
R37856 A2.n215 A2.n214 0.0135556
R37857 A2.n115 A2.n93 0.013431
R37858 A2.n111 A2.n95 0.013431
R37859 A2.n91 A2.n52 0.013
R37860 A2.n72 A2.n54 0.013
R37861 A2.n180 A2.n179 0.0124717
R37862 A2.n179 A2.n178 0.0124717
R37863 A2.n158 A2.n157 0.0124717
R37864 A2.n157 A2.n156 0.0124717
R37865 A2.n79 A2.n73 0.0122521
R37866 A2.n99 A2.n49 0.0117689
R37867 A2.n61 A2.n50 0.0114102
R37868 A2.n37 A2.n36 0.0111132
R37869 A2.n35 A2.n34 0.0111132
R37870 A2.n26 A2.n25 0.0111132
R37871 A2.n24 A2.n23 0.0111132
R37872 A2.n88 A2.n75 0.0100704
R37873 A2.n117 A2.n48 0.0100109
R37874 A2.n33 A2.n32 0.00993396
R37875 A2.n28 A2.n27 0.00993396
R37876 A2.n176 A2.n175 0.00981132
R37877 A2.n161 A2.n160 0.00981132
R37878 A2.n130 A2.n129 0.00967431
R37879 A2.n126 A2.n125 0.00967431
R37880 A2.n8 A2.n7 0.00936793
R37881 A2.n11 A2.n10 0.00936793
R37882 A2.n14 A2.n13 0.00936793
R37883 A2.n17 A2.n16 0.00936793
R37884 A2.n20 A2.n19 0.00936793
R37885 A2.n177 A2.n176 0.00936793
R37886 A2.n171 A2.n170 0.00936793
R37887 A2.n166 A2.n165 0.00936793
R37888 A2.n160 A2.n159 0.00936793
R37889 A2.n155 A2.n154 0.00936793
R37890 A2.n184 A2.n183 0.00936793
R37891 A2.n187 A2.n186 0.00936793
R37892 A2.n190 A2.n189 0.00936793
R37893 A2.n193 A2.n192 0.00936793
R37894 A2.n196 A2.n195 0.00936793
R37895 A2.n204 A2.n203 0.0092037
R37896 A2.n207 A2.n206 0.0092037
R37897 A2.n210 A2.n209 0.0092037
R37898 A2.n213 A2.n212 0.0092037
R37899 A2.n216 A2.n215 0.0092037
R37900 A2.n140 A2.n139 0.00875472
R37901 A2.n38 A2.n37 0.00875472
R37902 A2.n23 A2.n22 0.00875472
R37903 A2.n144 A2.n143 0.00875472
R37904 A2.n120 A2.n119 0.00852752
R37905 A2.n133 A2.n132 0.00852752
R37906 A2.n123 A2.n122 0.00852752
R37907 A2.n150 A2.n149 0.00852752
R37908 A2.n169 A2.n168 0.00803774
R37909 A2.n168 A2.n167 0.00803774
R37910 A2.n174 A2.n173 0.00759434
R37911 A2.n163 A2.n162 0.00759434
R37912 A2.n170 A2.n169 0.00626415
R37913 A2.n167 A2.n166 0.00626415
R37914 A2.n115 A2.n95 0.00588793
R37915 A2.n91 A2.n72 0.00570833
R37916 A2.n199 A2.n198 0.00519331
R37917 A2.n103 A2.n49 0.00481034
R37918 A2.n88 A2.n87 0.0047735
R37919 A2.n58 A2.n50 0.00466667
R37920 A2.n94 A2.n48 0.00457609
R37921 A2.n117 A2.n116 0.00457609
R37922 A2.n175 A2.n174 0.00449057
R37923 A2.n173 A2.n172 0.00449057
R37924 A2.n164 A2.n163 0.00449057
R37925 A2.n162 A2.n161 0.00449057
R37926 A2.n199 A2.n197 0.00449057
R37927 A2.n43 A2.n41 0.00410577
R37928 A2.n80 A2.n79 0.00370513
R37929 A2.n148 A2 0.00279358
R37930 A2.n172 A2.n171 0.00271698
R37931 A2.n165 A2.n164 0.00271698
R37932 A2 A2.n219 0.00269298
R37933 A2.n89 A2.n74 0.00253804
R37934 A2.n45 A2.n44 0.00185919
R37935 A2.n90 A2.n51 0.0018587
R37936 A2.n178 A2.n177 0.00183019
R37937 A2.n159 A2.n158 0.00183019
R37938 A2.n156 A2.n155 0.00183019
C0 a_10180_3343# a_10136_2294# 0.139f
C1 EF_R2RVCE_0.comparator_0.VOUTANALOG EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.00128f
C2 a_10475_5424# DVDD 0.449f
C3 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN m3_n495_n10736# 1.49e-19
C4 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL a_3441_n11595# 0.0195f
C5 a_n227_n10525# SELA 0.00242f
C6 a_211_n4513# VDD 1.98f
C7 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3611_n4513# 0.124f
C8 a_6371_n10521# m3_6103_n10732# 0.0049f
C9 a_9771_n10521# a_10039_n11591# 0.0272f
C10 a_3073_n10613# a_3173_n10525# 0.405f
C11 a_7578_n10857# VDD 0.484f
C12 a_10015_9447# a_10015_8387# 0.14f
C13 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_7578_n10857# 9.6e-19
C14 a_6809_n4509# VDD 1.98f
C15 a_3441_n11595# DVDD 0.261f
C16 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6809_n4509# 0.124f
C17 a_10015_9447# VSS 0.00938f
C18 a_10162_2241# EN 0.00364f
C19 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN VSS 0.061f
C20 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL SELA 0.746f
C21 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10209_n4509# 0.124f
C22 VDD B1 1.47f
C23 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN 0.181f
C24 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB B1 0.925f
C25 B1 SELB 0.0415f
C26 a_6371_n10521# a_7064_n11635# 0.265f
C27 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN m3_2905_n10736# 1.49e-19
C28 DVDD SELA 1.01f
C29 a_3073_n10613# a_3441_n11595# 0.139f
C30 a_10180_3343# VSS 9.56e-19
C31 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD 5.01f
C32 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN 0.238f
C33 a_6271_n10609# DVDD 0.417f
C34 VDD EN 0.258f
C35 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN 0.181f
C36 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN VDD 4.87f
C37 a_10618_2709# a_10162_2241# 0.265f
C38 a_10180_3343# a_10914_2086# 3.88e-20
C39 a_10235_4600# DVDD 0.0708f
C40 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB A2 1.2e-19
C41 a_5555_8917# VDD 0.522f
C42 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_n327_n10613# 0.00112f
C43 a_3173_n10525# a_4380_n10861# 0.289f
C44 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN m3_6103_n10732# 1.49e-19
C45 VDD A2 1.49f
C46 a_5555_8917# a_5555_7857# 0.14f
C47 a_9771_n10521# VDD 1.08f
C48 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_9771_n10521# 9.91e-19
C49 A2 SELB 0.083f
C50 a_466_n11639# A1 0.00648f
C51 a_6639_n11591# DVDD 0.261f
C52 DVDD VO 0.997f
C53 EF_R2RVCE_0.comparator_0.VBP EF_AMUX2to1ISO_1.VO 0.015f
C54 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A EN 2.07e-19
C55 DVDD B2 0.165f
C56 a_10618_2709# VDD 0.844f
C57 m3_9503_n10732# B1 0.00123f
C58 a_10475_5424# a_10179_5308# 0.136f
C59 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10475_5424# 0.00606f
C60 a_10136_2294# VSS 0.00922f
C61 a_4380_n10861# a_3441_n11595# 6.24e-19
C62 EF_AMUX2to1ISO_0.VO VSS 5.82f
C63 EF_R2RVCE_0.comparator_0.VBN EF_AMUX2to1ISO_1.VO 0.507f
C64 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB A1 0.931f
C65 a_7578_n10857# DVDD 0.0117f
C66 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN m3_9503_n10732# 1.49e-19
C67 a_10039_n11591# VDD 0.15f
C68 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10978_n10857# 9.6e-19
C69 m3_2905_n10736# A1 0.00124f
C70 EF_AMUX2to1ISO_0.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB 0.0349f
C71 VDD A1 1.47f
C72 a_10618_2709# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.018f
C73 a_10136_2294# a_10914_2086# 6.7e-19
C74 EF_R2RVCE_0.comparator_bias_0.down a_5553_10507# 0.028f
C75 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_466_n11639# 3.13e-19
C76 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_980_n10861# 0.00261f
C77 m3_n495_n10736# VSS 0.00203f
C78 DVDD B1 0.484f
C79 a_9771_n10521# m3_9503_n10732# 0.0049f
C80 a_4380_n10861# a_6271_n10609# 6.31e-19
C81 a_466_n11639# VDD 0.609f
C82 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_5553_10507# 5.39e-19
C83 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10475_5424# 0.00564f
C84 a_41_n11595# A1 0.00532f
C85 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_AMUX2to1ISO_1.VO 0.0445f
C86 DVDD EN 0.362f
C87 a_10162_2241# VDD 0.592f
C88 EF_R2RVCE_0.comparator_bias_0.up a_5553_10507# 0.0709f
C89 a_10475_5424# a_10169_4802# 7.97e-19
C90 a_10179_5308# a_10235_4600# 0.166f
C91 a_466_n11639# a_41_n11595# 0.461f
C92 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10235_4600# 0.00852f
C93 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB m3_2905_n10736# 9.58e-19
C94 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.comparator_0.VOUTANALOG 0.542f
C95 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3866_n11639# 3.13e-19
C96 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3073_n10613# 0.00112f
C97 a_10914_2086# VSS 7.15e-21
C98 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD 3.5f
C99 a_n327_n10613# m3_n495_n10736# 0.00773f
C100 DVDD A2 0.165f
C101 a_9771_n10521# DVDD 0.118f
C102 m3_2905_n10736# VDD 0.237f
C103 a_10179_5308# VO 0.169f
C104 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB VDD 3.5f
C105 a_n227_n10525# A1 0.00597f
C106 VDD SELB 0.0598f
C107 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB SELB 3.18e-19
C108 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y VO 0.0203f
C109 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.comparator_0.VOUTANALOG 0.00123f
C110 a_10162_2241# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.0172f
C111 a_10618_2709# DVDD 0.0862f
C112 a_5555_7857# VDD 0.684f
C113 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_41_n11595# 1.09e-19
C114 a_n327_n10613# VSS 0.0102f
C115 a_3073_n10613# A2 7.86e-19
C116 a_n227_n10525# a_466_n11639# 0.265f
C117 a_6271_n10609# a_6371_n10521# 0.405f
C118 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB m3_6103_n10732# 0.00159f
C119 a_41_n11595# VDD 0.153f
C120 a_10464_n11635# B2 0.00646f
C121 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL A1 0.0308f
C122 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10235_4600# 0.224f
C123 EF_R2RVCE_0.comparator_0.VOUTANALOG EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A 0.266f
C124 a_10039_n11591# DVDD 0.261f
C125 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A VDD 1.4f
C126 DVDD A1 0.49f
C127 EF_AMUX2to1ISO_1.VO a_3611_n4513# 6.66e-19
C128 a_10235_4600# a_10169_4802# 0.17f
C129 a_10475_5424# a_10180_3343# 4.85e-19
C130 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A VO 0.043f
C131 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_4380_n10861# 0.00261f
C132 a_6371_n10521# a_6639_n11591# 0.0272f
C133 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_n227_n10525# 5.11e-19
C134 EF_AMUX2to1ISO_1.VO a_10209_n4509# 1.07f
C135 a_466_n11639# DVDD 0.157f
C136 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB m3_9503_n10732# 9.58e-19
C137 m3_9503_n10732# VDD 0.237f
C138 a_n227_n10525# VDD 1.07f
C139 a_10169_4802# VO 0.0178f
C140 a_3073_n10613# A1 0.00572f
C141 EF_R2RVCE_0.comparator_bias_0.down a_5555_8917# 0.0111f
C142 a_10179_5308# EN 3.53e-19
C143 a_10162_2241# DVDD 0.104f
C144 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EN 0.0155f
C145 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL 4.83e-20
C146 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN 2.82f
C147 a_n227_n10525# a_41_n11595# 0.0272f
C148 a_4380_n10861# A2 0.00601f
C149 a_6371_n10521# a_7578_n10857# 0.289f
C150 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL VDD 0.0593f
C151 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN a_6271_n10609# 0.00112f
C152 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB DVDD 0.0846f
C153 m3_2905_n10736# DVDD 0.0559f
C154 VDD DVDD 11.9f
C155 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB DVDD 0.0843f
C156 a_6371_n10521# B1 0.00598f
C157 DVDD SELB 1.09f
C158 EF_R2RVCE_0.comparator_bias_0.up a_5555_8917# 0.096f
C159 a_10235_4600# a_10180_3343# 0.00306f
C160 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10618_2709# 0.0104f
C161 a_9771_n10521# a_10464_n11635# 0.265f
C162 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_3073_n10613# 0.00651f
C163 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A EN 0.0784f
C164 a_3073_n10613# m3_2905_n10736# 0.00773f
C165 a_9671_n10609# B2 8.08e-19
C166 a_41_n11595# DVDD 0.25f
C167 a_n327_n10613# a_980_n10861# 3.88e-20
C168 a_3073_n10613# VDD 0.34f
C169 a_211_n4513# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN 1.5f
C170 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL B1 0.0306f
C171 a_10169_4802# EN 0.00512f
C172 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A DVDD 0.0104f
C173 EF_R2RVCE_0.comparator_0.VBP VDD 10.8f
C174 a_3611_n4513# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN 1.5f
C175 a_6371_n10521# A2 0.00374f
C176 a_3173_n10525# a_3866_n11639# 0.265f
C177 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN a_7578_n10857# 0.00261f
C178 a_10464_n11635# a_10039_n11591# 0.461f
C179 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10618_2709# 2.44e-19
C180 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3173_n10525# 5.11e-19
C181 a_6809_n4509# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN 1.5f
C182 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_0.VO 5.55f
C183 m3_9503_n10732# DVDD 0.0554f
C184 a_n227_n10525# DVDD 0.113f
C185 EF_R2RVCE_0.comparator_0.VBN VDD 9.94f
C186 a_10209_n4509# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN 1.5f
C187 a_9671_n10609# B1 0.00567f
C188 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN B1 2.82f
C189 a_10235_4600# a_10136_2294# 6.27e-20
C190 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10162_2241# 0.0148f
C191 EF_R2RVCE_0.comparator_0.VOUTANALOG EF_AMUX2to1ISO_0.VO 0.359f
C192 m3_n495_n10736# SELA 0.00585f
C193 a_10013_10507# VDD 0.697f
C194 a_9771_n10521# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL 0.00242f
C195 a_3866_n11639# a_3441_n11595# 0.461f
C196 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_3441_n11595# 1.09e-19
C197 a_10978_n10857# B2 0.00602f
C198 EF_R2RVCE_0.comparator_bias_0.down VDD 11.6f
C199 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL DVDD 1.16f
C200 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_9671_n10609# 0.00112f
C201 a_4380_n10861# VDD 0.484f
C202 a_5553_10507# VSS 0.0239f
C203 a_10180_3343# EN 0.229f
C204 VSS SELA 0.0339f
C205 EF_AMUX2to1ISO_1.VO VSS 4.27f
C206 a_10179_5308# VDD 0.251f
C207 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y VDD 4.91f
C208 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB 0.153f
C209 a_3073_n10613# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL 0.231f
C210 a_9671_n10609# a_9771_n10521# 0.405f
C211 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN A2 5.23e-19
C212 EF_AMUX2to1ISO_0.VO a_211_n4513# 1.07f
C213 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_6271_n10609# 0.00876f
C214 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL a_10039_n11591# 0.0195f
C215 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10162_2241# 2.14e-19
C216 EF_R2RVCE_0.comparator_0.VOUTANALOG VSS 13.5f
C217 a_10464_n11635# VDD 0.608f
C218 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB 0.0349f
C219 EF_R2RVCE_0.comparator_bias_0.up VDD 5.51f
C220 a_3073_n10613# DVDD 0.422f
C221 EF_R2RVCE_0.comparator_bias_0.up a_5555_7857# 0.222f
C222 a_10180_3343# a_10618_2709# 0.405f
C223 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.823f
C224 a_n327_n10613# SELA 0.232f
C225 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A VDD 3.17f
C226 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_6639_n11591# 1.55e-20
C227 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN A1 2.82f
C228 a_6271_n10609# m3_6103_n10732# 0.00773f
C229 a_9671_n10609# a_10039_n11591# 0.139f
C230 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_10978_n10857# 0.00261f
C231 a_6371_n10521# VDD 1.08f
C232 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6371_n10521# 5.11e-19
C233 EF_AMUX2to1ISO_0.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN 2.82f
C234 a_6371_n10521# SELB 0.00242f
C235 a_10136_2294# EN 0.0106f
C236 a_211_n4513# VSS 0.00149f
C237 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB B2 0.93f
C238 a_10169_4802# VDD 0.0956f
C239 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_3611_n4513# 0.00474f
C240 a_9771_n10521# a_10978_n10857# 0.289f
C241 a_6271_n10609# a_7064_n11635# 8.36e-19
C242 a_3611_n4513# VDD 1.98f
C243 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_6809_n4509# 0.00631f
C244 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL 4.83e-20
C245 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL VDD 0.0593f
C246 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL SELB 0.746f
C247 a_4380_n10861# DVDD 0.0117f
C248 a_10209_n4509# VDD 1.98f
C249 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_10209_n4509# 0.00474f
C250 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN 1.28f
C251 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB B1 1.67e-19
C252 a_10618_2709# a_10136_2294# 0.0246f
C253 a_10180_3343# a_10162_2241# 8.36e-19
C254 a_10179_5308# DVDD 0.467f
C255 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y DVDD 0.0702f
C256 EF_R2RVCE_0.comparator_0.VBN EF_R2RVCE_0.comparator_0.VBP 1.78f
C257 a_10015_9447# VDD 0.508f
C258 a_7064_n11635# a_6639_n11591# 0.461f
C259 VSS EN 0.00384f
C260 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN VDD 5.02f
C261 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN 1.28f
C262 a_10978_n10857# a_10039_n11591# 6.24e-19
C263 a_3073_n10613# a_4380_n10861# 3.88e-20
C264 a_9671_n10609# VDD 0.34f
C265 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_9671_n10609# 0.00651f
C266 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN VDD 5.01f
C267 a_10464_n11635# DVDD 0.155f
C268 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN 1.28f
C269 a_5555_8917# VSS 0.00163f
C270 a_10914_2086# EN 7.57e-19
C271 EF_R2RVCE_0.comparator_bias_0.down EF_R2RVCE_0.comparator_0.VBP 0.175f
C272 a_10180_3343# VDD 0.192f
C273 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN 1.28f
C274 a_3866_n11639# A2 0.00645f
C275 a_7578_n10857# a_7064_n11635# 2.63e-19
C276 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB A2 0.93f
C277 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.comparator_0.VBP 5.81e-20
C278 a_3173_n10525# a_3441_n11595# 0.0272f
C279 a_10618_2709# VSS 3.07e-21
C280 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A DVDD 0.0901f
C281 EF_R2RVCE_0.comparator_bias_0.down EF_R2RVCE_0.comparator_0.VBN 3.35f
C282 a_6371_n10521# DVDD 0.118f
C283 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_9771_n10521# 5.11e-19
C284 a_7064_n11635# B1 0.00649f
C285 a_10136_2294# a_10162_2241# 0.461f
C286 a_10618_2709# a_10914_2086# 0.289f
C287 a_10180_3343# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.00283f
C288 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.comparator_0.VBP 1.63e-19
C289 a_10169_4802# DVDD 0.0333f
C290 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_n227_n10525# 0.00263f
C291 m3_6103_n10732# A2 0.00196f
C292 a_9671_n10609# m3_9503_n10732# 0.00773f
C293 VSS A1 0.00275f
C294 a_10978_n10857# VDD 0.484f
C295 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10013_10507# 0.0374f
C296 EF_AMUX2to1ISO_0.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB 0.175f
C297 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL DVDD 1.16f
C298 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.comparator_0.VBN 0.0447f
C299 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.comparator_bias_0.down 1.53f
C300 a_10136_2294# VDD 0.147f
C301 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10039_n11591# 1.09e-19
C302 EF_AMUX2to1ISO_0.VO VDD 10.9f
C303 a_10209_n4509# DVDD 2.27e-19
C304 a_10475_5424# a_10235_4600# 0.25f
C305 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10179_5308# 0.00834f
C306 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.comparator_bias_0.down 1.18f
C307 a_10162_2241# VSS 1.27e-19
C308 a_9671_n10609# DVDD 0.422f
C309 m3_n495_n10736# VDD 0.235f
C310 a_10475_5424# VO 0.0695f
C311 a_n327_n10613# A1 8.51e-19
C312 a_10162_2241# a_10914_2086# 2.63e-19
C313 a_10136_2294# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.00919f
C314 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y 2.12f
C315 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB VSS 0.00208f
C316 a_10180_3343# DVDD 0.381f
C317 a_10015_8387# VDD 0.512f
C318 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB 1.07e-19
C319 VDD VSS 0.191p
C320 a_n327_n10613# a_466_n11639# 8.36e-19
C321 a_3866_n11639# VDD 0.609f
C322 a_3866_n11639# SELB 0.00104f
C323 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10179_5308# 0.0131f
C324 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB 2.19e-19
C325 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD 3.56f
C326 EF_R2RVCE_0.comparator_0.VOUTANALOG EF_AMUX2to1ISO_1.VO 0.0398f
C327 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A 0.179f
C328 a_5555_7857# VSS 0.0236f
C329 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB SELB 8.51e-20
C330 a_10914_2086# VDD 0.421f
C331 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB 1.07e-19
C332 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB VDD 3.31f
C333 a_41_n11595# VSS 0.0025f
C334 a_10179_5308# a_10169_4802# 0.249f
C335 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10169_4802# 0.00899f
C336 EF_R2RVCE_0.comparator_bias_0.up EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A 1.44e-19
C337 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_3173_n10525# 0.00263f
C338 a_6271_n10609# a_6639_n11591# 0.139f
C339 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A VSS 0.00644f
C340 a_n227_n10525# m3_n495_n10736# 0.0049f
C341 a_10978_n10857# DVDD 0.012f
C342 m3_6103_n10732# VDD 0.238f
C343 a_n327_n10613# VDD 0.338f
C344 a_10013_10507# a_10015_9447# 0.139f
C345 a_10235_4600# VO 0.0204f
C346 a_980_n10861# A1 0.00605f
C347 a_10914_2086# EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.A 0.145f
C348 a_10475_5424# EN 0.00163f
C349 a_10136_2294# DVDD 0.169f
C350 a_n227_n10525# VSS 0.00321f
C351 EF_AMUX2to1ISO_1.VO a_6809_n4509# 1.07f
C352 a_10464_n11635# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL 0.0044f
C353 a_3173_n10525# A2 0.00591f
C354 a_n327_n10613# a_41_n11595# 0.139f
C355 a_980_n10861# a_466_n11639# 2.63e-19
C356 a_6271_n10609# a_7578_n10857# 3.88e-20
C357 a_7064_n11635# VDD 0.609f
C358 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_7064_n11635# 3.13e-19
C359 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10015_9447# 0.0424f
C360 a_7064_n11635# SELB 0.00457f
C361 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10169_4802# 0.0308f
C362 m3_n495_n10736# DVDD 0.00403f
C363 a_6271_n10609# B1 8.72e-19
C364 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN 0.00175f
C365 EF_R2RVCE_0.comparator_bias_0.up a_10015_9447# 0.00243f
C366 a_10179_5308# a_10180_3343# 2.43e-19
C367 a_3866_n11639# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL 0.0044f
C368 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10180_3343# 0.00999f
C369 EF_R2RVCE_0.comparator_0.VBP EF_AMUX2to1ISO_0.VO 0.385f
C370 a_3441_n11595# A2 0.00528f
C371 a_9671_n10609# a_10464_n11635# 8.36e-19
C372 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_980_n10861# 9.6e-19
C373 a_7578_n10857# a_6639_n11591# 6.24e-19
C374 VSS DVDD 0.00695f
C375 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN 2.82f
C376 a_3866_n11639# DVDD 0.155f
C377 a_n327_n10613# a_n227_n10525# 0.405f
C378 a_5553_10507# a_5555_8917# 0.14f
C379 a_980_n10861# VDD 0.484f
C380 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB DVDD 0.077f
C381 a_3173_n10525# A1 0.00228f
C382 a_6639_n11591# B1 0.00533f
C383 a_10235_4600# EN 0.00732f
C384 a_10914_2086# DVDD 9.52e-19
C385 EF_R2RVCE_0.comparator_0.VBN EF_AMUX2to1ISO_0.VO 0.091f
C386 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB DVDD 0.152f
C387 a_3073_n10613# a_3866_n11639# 8.36e-19
C388 a_6271_n10609# A2 0.00788f
C389 a_980_n10861# a_41_n11595# 6.24e-19
C390 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN a_6371_n10521# 0.00263f
C391 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10180_3343# 0.00654f
C392 VO EN 0.00366f
C393 EF_R2RVCE_0.comparator_0.VBP VSS 2.22f
C394 a_3441_n11595# A1 0.00153f
C395 m3_6103_n10732# DVDD 0.0554f
C396 a_n327_n10613# DVDD 0.389f
C397 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN B2 2.82f
C398 a_7578_n10857# B1 0.00605f
C399 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN a_3611_n4513# 2.44e-20
C400 a_10169_4802# a_10180_3343# 0.00246f
C401 a_10235_4600# a_10618_2709# 9.75e-19
C402 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10136_2294# 0.0177f
C403 a_6639_n11591# A2 0.0029f
C404 a_10978_n10857# a_10464_n11635# 2.63e-19
C405 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_3173_n10525# 9.91e-19
C406 a_9671_n10609# EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.DINL 0.231f
C407 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN a_6809_n4509# 1.05e-19
C408 EF_R2RVCE_0.comparator_0.VBN VSS 11.1f
C409 A1 SELA 0.0418f
C410 a_9771_n10521# B2 0.00595f
C411 a_3173_n10525# m3_2905_n10736# 0.0049f
C412 a_7064_n11635# DVDD 0.157f
C413 a_n227_n10525# a_980_n10861# 0.289f
C414 a_10013_10507# a_10015_8387# 4.42e-21
C415 a_3173_n10525# VDD 1.08f
C416 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_tg_0.VIN a_10209_n4509# 2.44e-20
C417 a_10013_10507# VSS 0.0638f
C418 a_10475_5424# VDD 0.17f
C419 EF_R2RVCE_0.comparator_bias_0.down VSS 1.27f
C420 a_466_n11639# SELA 0.00457f
C421 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN B1 3.48e-19
C422 a_4380_n10861# a_3866_n11639# 2.63e-19
C423 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10015_8387# 0.0424f
C424 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A a_10136_2294# 0.00121f
C425 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_4380_n10861# 9.6e-19
C426 a_3441_n11595# VDD 0.151f
C427 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y VSS 2.64f
C428 a_10039_n11591# B2 0.00529f
C429 a_980_n10861# DVDD 0.0117f
C430 a_9771_n10521# B1 0.00226f
C431 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB SELA 3.18e-19
C432 EF_R2RVCE_0.comparator_bias_0.up a_10015_8387# 0.176f
C433 a_10169_4802# a_10136_2294# 1.11e-20
C434 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB 2.03e-19
C435 EF_R2RVCE_0.sky130_fd_sc_hvl__inv_4_0.Y a_10914_2086# 0.00403f
C436 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN A2 2.82f
C437 EF_R2RVCE_0.comparator_bias_0.up VSS 1.22f
C438 a_5553_10507# VDD 0.701f
C439 VDD SELA 0.0685f
C440 EF_AMUX2to1ISO_1.VO VDD 12f
C441 EF_AMUX2to1ISO_1.VO EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB 0.171f
C442 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_tg_0.VIN a_9771_n10521# 0.00263f
C443 a_6271_n10609# VDD 0.343f
C444 EF_AMUX2to1ISO_0.VO a_3611_n4513# 1.07f
C445 a_6271_n10609# SELB 0.232f
C446 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_10464_n11635# 3.13e-19
C447 a_10618_2709# EN 0.0207f
C448 EF_R2RVCE_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.A VSS 0.825f
C449 a_10235_4600# VDD 0.517f
C450 EF_R2RVCE_0.comparator_0.VOUTANALOG VDD 5.14f
C451 a_41_n11595# SELA 0.021f
C452 a_10039_n11591# B1 0.00152f
C453 a_3173_n10525# EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.DINL 0.00242f
C454 a_9671_n10609# a_10978_n10857# 3.88e-20
C455 a_5555_7857# EF_R2RVCE_0.comparator_0.VOUTANALOG 2.82e-19
C456 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_ls_0.DOHB a_6371_n10521# 0.00182f
C457 EF_AMUX2to1ISO_0.VO EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_tg_0.VIN 2.82f
C458 VDD VO 0.294f
C459 a_6639_n11591# VDD 0.15f
C460 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_6639_n11591# 1.09e-19
C461 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_0.single_tg_0.VIN A1 4.34e-19
C462 a_6639_n11591# SELB 0.021f
C463 a_3173_n10525# DVDD 0.118f
C464 VDD B2 1.4f
C465 EF_AMUX2to1ISO_1.single_ls_2tgwd_sw_1.single_ls_0.DOHB B2 1.2e-19
C466 EF_AMUX2to1ISO_0.single_ls_2tgwd_sw_1.single_ls_0.DOHB a_211_n4513# 0.124f
.ends

