VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_R2RVC02
  CLASS BLOCK ;
  FOREIGN EF_R2RVC02 ;
  ORIGIN 8.090 42.230 ;
  SIZE 78.410 BY 98.600 ;
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 263.488281 ;
    PORT
      LAYER met3 ;
        RECT -7.590 52.790 -7.070 53.570 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 433.882782 ;
    PORT
      LAYER met4 ;
        RECT -7.630 55.380 -7.250 55.750 ;
    END
  END VDD
  PIN DVSS
    ANTENNADIFFAREA 107.239799 ;
    PORT
      LAYER met3 ;
        RECT 69.790 1.410 70.060 2.170 ;
    END
  END DVSS
  PIN DVDD
    ANTENNADIFFAREA 7.633700 ;
    PORT
      LAYER met3 ;
        RECT 69.680 26.580 69.940 27.310 ;
    END
  END DVDD
  PIN SELB
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met2 ;
        RECT 35.210 -41.680 35.560 -40.960 ;
    END
  END SELB
  PIN SELA
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met2 ;
        RECT 2.030 -41.680 2.320 -41.020 ;
    END
  END SELA
  PIN VO
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 69.820 22.220 69.970 22.460 ;
    END
  END VO
  PIN B2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met4 ;
        RECT 63.320 -41.610 63.560 -41.190 ;
    END
  END B2
  PIN B1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met4 ;
        RECT 46.530 -41.270 46.760 -41.010 ;
    END
  END B1
  PIN A2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met4 ;
        RECT 30.000 -41.660 30.420 -41.120 ;
    END
  END A2
  PIN A1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met4 ;
        RECT 13.120 -42.000 13.930 -39.280 ;
    END
  END A1
  OBS
      LAYER li1 ;
        RECT 0.330 -39.890 64.300 52.065 ;
      LAYER met1 ;
        RECT -0.130 -40.050 67.280 51.750 ;
      LAYER met2 ;
        RECT -1.080 -40.680 70.210 51.750 ;
        RECT -1.080 -40.740 34.930 -40.680 ;
        RECT -1.080 -41.960 1.750 -40.740 ;
        RECT 2.600 -41.960 34.930 -40.740 ;
        RECT 35.840 -41.960 70.210 -40.680 ;
        RECT -1.080 -42.230 70.210 -41.960 ;
      LAYER met3 ;
        RECT -8.090 53.970 70.320 56.360 ;
        RECT -8.090 52.390 -7.990 53.970 ;
        RECT -6.670 52.390 70.320 53.970 ;
        RECT -8.090 27.710 70.320 52.390 ;
        RECT -8.090 26.180 69.280 27.710 ;
        RECT -8.090 22.860 70.320 26.180 ;
        RECT -8.090 21.820 69.420 22.860 ;
        RECT -8.090 2.570 70.320 21.820 ;
        RECT -8.090 1.010 69.390 2.570 ;
        RECT -8.090 -42.230 70.320 1.010 ;
      LAYER met4 ;
        RECT -8.060 56.150 69.760 56.370 ;
        RECT -8.060 54.980 -8.030 56.150 ;
        RECT -6.850 54.980 69.760 56.150 ;
        RECT -8.060 -38.880 69.760 54.980 ;
        RECT -8.060 -42.210 12.720 -38.880 ;
        RECT 14.330 -40.610 69.760 -38.880 ;
        RECT 14.330 -40.720 46.130 -40.610 ;
        RECT 14.330 -42.060 29.600 -40.720 ;
        RECT 30.820 -41.670 46.130 -40.720 ;
        RECT 47.160 -40.790 69.760 -40.610 ;
        RECT 47.160 -41.670 62.920 -40.790 ;
        RECT 30.820 -42.010 62.920 -41.670 ;
        RECT 63.960 -42.010 69.760 -40.790 ;
        RECT 30.820 -42.060 69.760 -42.010 ;
        RECT 14.330 -42.210 69.760 -42.060 ;
  END
END EF_R2RVC02
END LIBRARY

