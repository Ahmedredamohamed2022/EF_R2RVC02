magic
tech sky130A
magscale 1 2
timestamp 1694943448
<< nwell >>
rect 507806 647830 518378 649916
rect 507806 646042 513113 647830
<< pwell >>
rect 513380 646078 518338 647724
<< mvnmos >>
rect 514514 646368 514914 647368
rect 514972 646368 515372 647368
rect 515430 646368 515830 647368
rect 515888 646368 516288 647368
rect 516346 646368 516746 647368
rect 516804 646368 517204 647368
<< mvpmos >>
rect 514355 649378 517355 649578
rect 513709 648213 514109 649213
rect 514167 648213 514567 649213
rect 514625 648213 515025 649213
rect 515083 648213 515483 649213
rect 515659 648213 516059 649213
rect 516117 648213 516517 649213
rect 516575 648213 516975 649213
rect 517033 648213 517433 649213
rect 517609 648213 518009 649213
<< mvndiff >>
rect 514456 647327 514514 647368
rect 514456 647293 514468 647327
rect 514502 647293 514514 647327
rect 514456 647259 514514 647293
rect 514456 647225 514468 647259
rect 514502 647225 514514 647259
rect 514456 647191 514514 647225
rect 514456 647157 514468 647191
rect 514502 647157 514514 647191
rect 514456 647123 514514 647157
rect 514456 647089 514468 647123
rect 514502 647089 514514 647123
rect 514456 647055 514514 647089
rect 514456 647021 514468 647055
rect 514502 647021 514514 647055
rect 514456 646987 514514 647021
rect 514456 646953 514468 646987
rect 514502 646953 514514 646987
rect 514456 646919 514514 646953
rect 514456 646885 514468 646919
rect 514502 646885 514514 646919
rect 514456 646851 514514 646885
rect 514456 646817 514468 646851
rect 514502 646817 514514 646851
rect 514456 646783 514514 646817
rect 514456 646749 514468 646783
rect 514502 646749 514514 646783
rect 514456 646715 514514 646749
rect 514456 646681 514468 646715
rect 514502 646681 514514 646715
rect 514456 646647 514514 646681
rect 514456 646613 514468 646647
rect 514502 646613 514514 646647
rect 514456 646579 514514 646613
rect 514456 646545 514468 646579
rect 514502 646545 514514 646579
rect 514456 646511 514514 646545
rect 514456 646477 514468 646511
rect 514502 646477 514514 646511
rect 514456 646443 514514 646477
rect 514456 646409 514468 646443
rect 514502 646409 514514 646443
rect 514456 646368 514514 646409
rect 514914 647327 514972 647368
rect 514914 647293 514926 647327
rect 514960 647293 514972 647327
rect 514914 647259 514972 647293
rect 514914 647225 514926 647259
rect 514960 647225 514972 647259
rect 514914 647191 514972 647225
rect 514914 647157 514926 647191
rect 514960 647157 514972 647191
rect 514914 647123 514972 647157
rect 514914 647089 514926 647123
rect 514960 647089 514972 647123
rect 514914 647055 514972 647089
rect 514914 647021 514926 647055
rect 514960 647021 514972 647055
rect 514914 646987 514972 647021
rect 514914 646953 514926 646987
rect 514960 646953 514972 646987
rect 514914 646919 514972 646953
rect 514914 646885 514926 646919
rect 514960 646885 514972 646919
rect 514914 646851 514972 646885
rect 514914 646817 514926 646851
rect 514960 646817 514972 646851
rect 514914 646783 514972 646817
rect 514914 646749 514926 646783
rect 514960 646749 514972 646783
rect 514914 646715 514972 646749
rect 514914 646681 514926 646715
rect 514960 646681 514972 646715
rect 514914 646647 514972 646681
rect 514914 646613 514926 646647
rect 514960 646613 514972 646647
rect 514914 646579 514972 646613
rect 514914 646545 514926 646579
rect 514960 646545 514972 646579
rect 514914 646511 514972 646545
rect 514914 646477 514926 646511
rect 514960 646477 514972 646511
rect 514914 646443 514972 646477
rect 514914 646409 514926 646443
rect 514960 646409 514972 646443
rect 514914 646368 514972 646409
rect 515372 647327 515430 647368
rect 515372 647293 515384 647327
rect 515418 647293 515430 647327
rect 515372 647259 515430 647293
rect 515372 647225 515384 647259
rect 515418 647225 515430 647259
rect 515372 647191 515430 647225
rect 515372 647157 515384 647191
rect 515418 647157 515430 647191
rect 515372 647123 515430 647157
rect 515372 647089 515384 647123
rect 515418 647089 515430 647123
rect 515372 647055 515430 647089
rect 515372 647021 515384 647055
rect 515418 647021 515430 647055
rect 515372 646987 515430 647021
rect 515372 646953 515384 646987
rect 515418 646953 515430 646987
rect 515372 646919 515430 646953
rect 515372 646885 515384 646919
rect 515418 646885 515430 646919
rect 515372 646851 515430 646885
rect 515372 646817 515384 646851
rect 515418 646817 515430 646851
rect 515372 646783 515430 646817
rect 515372 646749 515384 646783
rect 515418 646749 515430 646783
rect 515372 646715 515430 646749
rect 515372 646681 515384 646715
rect 515418 646681 515430 646715
rect 515372 646647 515430 646681
rect 515372 646613 515384 646647
rect 515418 646613 515430 646647
rect 515372 646579 515430 646613
rect 515372 646545 515384 646579
rect 515418 646545 515430 646579
rect 515372 646511 515430 646545
rect 515372 646477 515384 646511
rect 515418 646477 515430 646511
rect 515372 646443 515430 646477
rect 515372 646409 515384 646443
rect 515418 646409 515430 646443
rect 515372 646368 515430 646409
rect 515830 647327 515888 647368
rect 515830 647293 515842 647327
rect 515876 647293 515888 647327
rect 515830 647259 515888 647293
rect 515830 647225 515842 647259
rect 515876 647225 515888 647259
rect 515830 647191 515888 647225
rect 515830 647157 515842 647191
rect 515876 647157 515888 647191
rect 515830 647123 515888 647157
rect 515830 647089 515842 647123
rect 515876 647089 515888 647123
rect 515830 647055 515888 647089
rect 515830 647021 515842 647055
rect 515876 647021 515888 647055
rect 515830 646987 515888 647021
rect 515830 646953 515842 646987
rect 515876 646953 515888 646987
rect 515830 646919 515888 646953
rect 515830 646885 515842 646919
rect 515876 646885 515888 646919
rect 515830 646851 515888 646885
rect 515830 646817 515842 646851
rect 515876 646817 515888 646851
rect 515830 646783 515888 646817
rect 515830 646749 515842 646783
rect 515876 646749 515888 646783
rect 515830 646715 515888 646749
rect 515830 646681 515842 646715
rect 515876 646681 515888 646715
rect 515830 646647 515888 646681
rect 515830 646613 515842 646647
rect 515876 646613 515888 646647
rect 515830 646579 515888 646613
rect 515830 646545 515842 646579
rect 515876 646545 515888 646579
rect 515830 646511 515888 646545
rect 515830 646477 515842 646511
rect 515876 646477 515888 646511
rect 515830 646443 515888 646477
rect 515830 646409 515842 646443
rect 515876 646409 515888 646443
rect 515830 646368 515888 646409
rect 516288 647327 516346 647368
rect 516288 647293 516300 647327
rect 516334 647293 516346 647327
rect 516288 647259 516346 647293
rect 516288 647225 516300 647259
rect 516334 647225 516346 647259
rect 516288 647191 516346 647225
rect 516288 647157 516300 647191
rect 516334 647157 516346 647191
rect 516288 647123 516346 647157
rect 516288 647089 516300 647123
rect 516334 647089 516346 647123
rect 516288 647055 516346 647089
rect 516288 647021 516300 647055
rect 516334 647021 516346 647055
rect 516288 646987 516346 647021
rect 516288 646953 516300 646987
rect 516334 646953 516346 646987
rect 516288 646919 516346 646953
rect 516288 646885 516300 646919
rect 516334 646885 516346 646919
rect 516288 646851 516346 646885
rect 516288 646817 516300 646851
rect 516334 646817 516346 646851
rect 516288 646783 516346 646817
rect 516288 646749 516300 646783
rect 516334 646749 516346 646783
rect 516288 646715 516346 646749
rect 516288 646681 516300 646715
rect 516334 646681 516346 646715
rect 516288 646647 516346 646681
rect 516288 646613 516300 646647
rect 516334 646613 516346 646647
rect 516288 646579 516346 646613
rect 516288 646545 516300 646579
rect 516334 646545 516346 646579
rect 516288 646511 516346 646545
rect 516288 646477 516300 646511
rect 516334 646477 516346 646511
rect 516288 646443 516346 646477
rect 516288 646409 516300 646443
rect 516334 646409 516346 646443
rect 516288 646368 516346 646409
rect 516746 647327 516804 647368
rect 516746 647293 516758 647327
rect 516792 647293 516804 647327
rect 516746 647259 516804 647293
rect 516746 647225 516758 647259
rect 516792 647225 516804 647259
rect 516746 647191 516804 647225
rect 516746 647157 516758 647191
rect 516792 647157 516804 647191
rect 516746 647123 516804 647157
rect 516746 647089 516758 647123
rect 516792 647089 516804 647123
rect 516746 647055 516804 647089
rect 516746 647021 516758 647055
rect 516792 647021 516804 647055
rect 516746 646987 516804 647021
rect 516746 646953 516758 646987
rect 516792 646953 516804 646987
rect 516746 646919 516804 646953
rect 516746 646885 516758 646919
rect 516792 646885 516804 646919
rect 516746 646851 516804 646885
rect 516746 646817 516758 646851
rect 516792 646817 516804 646851
rect 516746 646783 516804 646817
rect 516746 646749 516758 646783
rect 516792 646749 516804 646783
rect 516746 646715 516804 646749
rect 516746 646681 516758 646715
rect 516792 646681 516804 646715
rect 516746 646647 516804 646681
rect 516746 646613 516758 646647
rect 516792 646613 516804 646647
rect 516746 646579 516804 646613
rect 516746 646545 516758 646579
rect 516792 646545 516804 646579
rect 516746 646511 516804 646545
rect 516746 646477 516758 646511
rect 516792 646477 516804 646511
rect 516746 646443 516804 646477
rect 516746 646409 516758 646443
rect 516792 646409 516804 646443
rect 516746 646368 516804 646409
rect 517204 647327 517262 647368
rect 517204 647293 517216 647327
rect 517250 647293 517262 647327
rect 517204 647259 517262 647293
rect 517204 647225 517216 647259
rect 517250 647225 517262 647259
rect 517204 647191 517262 647225
rect 517204 647157 517216 647191
rect 517250 647157 517262 647191
rect 517204 647123 517262 647157
rect 517204 647089 517216 647123
rect 517250 647089 517262 647123
rect 517204 647055 517262 647089
rect 517204 647021 517216 647055
rect 517250 647021 517262 647055
rect 517204 646987 517262 647021
rect 517204 646953 517216 646987
rect 517250 646953 517262 646987
rect 517204 646919 517262 646953
rect 517204 646885 517216 646919
rect 517250 646885 517262 646919
rect 517204 646851 517262 646885
rect 517204 646817 517216 646851
rect 517250 646817 517262 646851
rect 517204 646783 517262 646817
rect 517204 646749 517216 646783
rect 517250 646749 517262 646783
rect 517204 646715 517262 646749
rect 517204 646681 517216 646715
rect 517250 646681 517262 646715
rect 517204 646647 517262 646681
rect 517204 646613 517216 646647
rect 517250 646613 517262 646647
rect 517204 646579 517262 646613
rect 517204 646545 517216 646579
rect 517250 646545 517262 646579
rect 517204 646511 517262 646545
rect 517204 646477 517216 646511
rect 517250 646477 517262 646511
rect 517204 646443 517262 646477
rect 517204 646409 517216 646443
rect 517250 646409 517262 646443
rect 517204 646368 517262 646409
<< mvpdiff >>
rect 514297 649563 514355 649578
rect 514297 649529 514309 649563
rect 514343 649529 514355 649563
rect 514297 649495 514355 649529
rect 514297 649461 514309 649495
rect 514343 649461 514355 649495
rect 514297 649427 514355 649461
rect 514297 649393 514309 649427
rect 514343 649393 514355 649427
rect 514297 649378 514355 649393
rect 517355 649563 517413 649578
rect 517355 649529 517367 649563
rect 517401 649529 517413 649563
rect 517355 649495 517413 649529
rect 517355 649461 517367 649495
rect 517401 649461 517413 649495
rect 517355 649427 517413 649461
rect 517355 649393 517367 649427
rect 517401 649393 517413 649427
rect 517355 649378 517413 649393
rect 513651 649172 513709 649213
rect 513651 649138 513663 649172
rect 513697 649138 513709 649172
rect 513651 649104 513709 649138
rect 513651 649070 513663 649104
rect 513697 649070 513709 649104
rect 513651 649036 513709 649070
rect 513651 649002 513663 649036
rect 513697 649002 513709 649036
rect 513651 648968 513709 649002
rect 513651 648934 513663 648968
rect 513697 648934 513709 648968
rect 513651 648900 513709 648934
rect 513651 648866 513663 648900
rect 513697 648866 513709 648900
rect 513651 648832 513709 648866
rect 513651 648798 513663 648832
rect 513697 648798 513709 648832
rect 513651 648764 513709 648798
rect 513651 648730 513663 648764
rect 513697 648730 513709 648764
rect 513651 648696 513709 648730
rect 513651 648662 513663 648696
rect 513697 648662 513709 648696
rect 513651 648628 513709 648662
rect 513651 648594 513663 648628
rect 513697 648594 513709 648628
rect 513651 648560 513709 648594
rect 513651 648526 513663 648560
rect 513697 648526 513709 648560
rect 513651 648492 513709 648526
rect 513651 648458 513663 648492
rect 513697 648458 513709 648492
rect 513651 648424 513709 648458
rect 513651 648390 513663 648424
rect 513697 648390 513709 648424
rect 513651 648356 513709 648390
rect 513651 648322 513663 648356
rect 513697 648322 513709 648356
rect 513651 648288 513709 648322
rect 513651 648254 513663 648288
rect 513697 648254 513709 648288
rect 513651 648213 513709 648254
rect 514109 649172 514167 649213
rect 514109 649138 514121 649172
rect 514155 649138 514167 649172
rect 514109 649104 514167 649138
rect 514109 649070 514121 649104
rect 514155 649070 514167 649104
rect 514109 649036 514167 649070
rect 514109 649002 514121 649036
rect 514155 649002 514167 649036
rect 514109 648968 514167 649002
rect 514109 648934 514121 648968
rect 514155 648934 514167 648968
rect 514109 648900 514167 648934
rect 514109 648866 514121 648900
rect 514155 648866 514167 648900
rect 514109 648832 514167 648866
rect 514109 648798 514121 648832
rect 514155 648798 514167 648832
rect 514109 648764 514167 648798
rect 514109 648730 514121 648764
rect 514155 648730 514167 648764
rect 514109 648696 514167 648730
rect 514109 648662 514121 648696
rect 514155 648662 514167 648696
rect 514109 648628 514167 648662
rect 514109 648594 514121 648628
rect 514155 648594 514167 648628
rect 514109 648560 514167 648594
rect 514109 648526 514121 648560
rect 514155 648526 514167 648560
rect 514109 648492 514167 648526
rect 514109 648458 514121 648492
rect 514155 648458 514167 648492
rect 514109 648424 514167 648458
rect 514109 648390 514121 648424
rect 514155 648390 514167 648424
rect 514109 648356 514167 648390
rect 514109 648322 514121 648356
rect 514155 648322 514167 648356
rect 514109 648288 514167 648322
rect 514109 648254 514121 648288
rect 514155 648254 514167 648288
rect 514109 648213 514167 648254
rect 514567 649172 514625 649213
rect 514567 649138 514579 649172
rect 514613 649138 514625 649172
rect 514567 649104 514625 649138
rect 514567 649070 514579 649104
rect 514613 649070 514625 649104
rect 514567 649036 514625 649070
rect 514567 649002 514579 649036
rect 514613 649002 514625 649036
rect 514567 648968 514625 649002
rect 514567 648934 514579 648968
rect 514613 648934 514625 648968
rect 514567 648900 514625 648934
rect 514567 648866 514579 648900
rect 514613 648866 514625 648900
rect 514567 648832 514625 648866
rect 514567 648798 514579 648832
rect 514613 648798 514625 648832
rect 514567 648764 514625 648798
rect 514567 648730 514579 648764
rect 514613 648730 514625 648764
rect 514567 648696 514625 648730
rect 514567 648662 514579 648696
rect 514613 648662 514625 648696
rect 514567 648628 514625 648662
rect 514567 648594 514579 648628
rect 514613 648594 514625 648628
rect 514567 648560 514625 648594
rect 514567 648526 514579 648560
rect 514613 648526 514625 648560
rect 514567 648492 514625 648526
rect 514567 648458 514579 648492
rect 514613 648458 514625 648492
rect 514567 648424 514625 648458
rect 514567 648390 514579 648424
rect 514613 648390 514625 648424
rect 514567 648356 514625 648390
rect 514567 648322 514579 648356
rect 514613 648322 514625 648356
rect 514567 648288 514625 648322
rect 514567 648254 514579 648288
rect 514613 648254 514625 648288
rect 514567 648213 514625 648254
rect 515025 649172 515083 649213
rect 515025 649138 515037 649172
rect 515071 649138 515083 649172
rect 515025 649104 515083 649138
rect 515025 649070 515037 649104
rect 515071 649070 515083 649104
rect 515025 649036 515083 649070
rect 515025 649002 515037 649036
rect 515071 649002 515083 649036
rect 515025 648968 515083 649002
rect 515025 648934 515037 648968
rect 515071 648934 515083 648968
rect 515025 648900 515083 648934
rect 515025 648866 515037 648900
rect 515071 648866 515083 648900
rect 515025 648832 515083 648866
rect 515025 648798 515037 648832
rect 515071 648798 515083 648832
rect 515025 648764 515083 648798
rect 515025 648730 515037 648764
rect 515071 648730 515083 648764
rect 515025 648696 515083 648730
rect 515025 648662 515037 648696
rect 515071 648662 515083 648696
rect 515025 648628 515083 648662
rect 515025 648594 515037 648628
rect 515071 648594 515083 648628
rect 515025 648560 515083 648594
rect 515025 648526 515037 648560
rect 515071 648526 515083 648560
rect 515025 648492 515083 648526
rect 515025 648458 515037 648492
rect 515071 648458 515083 648492
rect 515025 648424 515083 648458
rect 515025 648390 515037 648424
rect 515071 648390 515083 648424
rect 515025 648356 515083 648390
rect 515025 648322 515037 648356
rect 515071 648322 515083 648356
rect 515025 648288 515083 648322
rect 515025 648254 515037 648288
rect 515071 648254 515083 648288
rect 515025 648213 515083 648254
rect 515483 649172 515541 649213
rect 515483 649138 515495 649172
rect 515529 649138 515541 649172
rect 515483 649104 515541 649138
rect 515483 649070 515495 649104
rect 515529 649070 515541 649104
rect 515483 649036 515541 649070
rect 515483 649002 515495 649036
rect 515529 649002 515541 649036
rect 515483 648968 515541 649002
rect 515483 648934 515495 648968
rect 515529 648934 515541 648968
rect 515483 648900 515541 648934
rect 515483 648866 515495 648900
rect 515529 648866 515541 648900
rect 515483 648832 515541 648866
rect 515483 648798 515495 648832
rect 515529 648798 515541 648832
rect 515483 648764 515541 648798
rect 515483 648730 515495 648764
rect 515529 648730 515541 648764
rect 515483 648696 515541 648730
rect 515483 648662 515495 648696
rect 515529 648662 515541 648696
rect 515483 648628 515541 648662
rect 515483 648594 515495 648628
rect 515529 648594 515541 648628
rect 515483 648560 515541 648594
rect 515483 648526 515495 648560
rect 515529 648526 515541 648560
rect 515483 648492 515541 648526
rect 515483 648458 515495 648492
rect 515529 648458 515541 648492
rect 515483 648424 515541 648458
rect 515483 648390 515495 648424
rect 515529 648390 515541 648424
rect 515483 648356 515541 648390
rect 515483 648322 515495 648356
rect 515529 648322 515541 648356
rect 515483 648288 515541 648322
rect 515483 648254 515495 648288
rect 515529 648254 515541 648288
rect 515483 648213 515541 648254
rect 515601 649172 515659 649213
rect 515601 649138 515613 649172
rect 515647 649138 515659 649172
rect 515601 649104 515659 649138
rect 515601 649070 515613 649104
rect 515647 649070 515659 649104
rect 515601 649036 515659 649070
rect 515601 649002 515613 649036
rect 515647 649002 515659 649036
rect 515601 648968 515659 649002
rect 515601 648934 515613 648968
rect 515647 648934 515659 648968
rect 515601 648900 515659 648934
rect 515601 648866 515613 648900
rect 515647 648866 515659 648900
rect 515601 648832 515659 648866
rect 515601 648798 515613 648832
rect 515647 648798 515659 648832
rect 515601 648764 515659 648798
rect 515601 648730 515613 648764
rect 515647 648730 515659 648764
rect 515601 648696 515659 648730
rect 515601 648662 515613 648696
rect 515647 648662 515659 648696
rect 515601 648628 515659 648662
rect 515601 648594 515613 648628
rect 515647 648594 515659 648628
rect 515601 648560 515659 648594
rect 515601 648526 515613 648560
rect 515647 648526 515659 648560
rect 515601 648492 515659 648526
rect 515601 648458 515613 648492
rect 515647 648458 515659 648492
rect 515601 648424 515659 648458
rect 515601 648390 515613 648424
rect 515647 648390 515659 648424
rect 515601 648356 515659 648390
rect 515601 648322 515613 648356
rect 515647 648322 515659 648356
rect 515601 648288 515659 648322
rect 515601 648254 515613 648288
rect 515647 648254 515659 648288
rect 515601 648213 515659 648254
rect 516059 649172 516117 649213
rect 516059 649138 516071 649172
rect 516105 649138 516117 649172
rect 516059 649104 516117 649138
rect 516059 649070 516071 649104
rect 516105 649070 516117 649104
rect 516059 649036 516117 649070
rect 516059 649002 516071 649036
rect 516105 649002 516117 649036
rect 516059 648968 516117 649002
rect 516059 648934 516071 648968
rect 516105 648934 516117 648968
rect 516059 648900 516117 648934
rect 516059 648866 516071 648900
rect 516105 648866 516117 648900
rect 516059 648832 516117 648866
rect 516059 648798 516071 648832
rect 516105 648798 516117 648832
rect 516059 648764 516117 648798
rect 516059 648730 516071 648764
rect 516105 648730 516117 648764
rect 516059 648696 516117 648730
rect 516059 648662 516071 648696
rect 516105 648662 516117 648696
rect 516059 648628 516117 648662
rect 516059 648594 516071 648628
rect 516105 648594 516117 648628
rect 516059 648560 516117 648594
rect 516059 648526 516071 648560
rect 516105 648526 516117 648560
rect 516059 648492 516117 648526
rect 516059 648458 516071 648492
rect 516105 648458 516117 648492
rect 516059 648424 516117 648458
rect 516059 648390 516071 648424
rect 516105 648390 516117 648424
rect 516059 648356 516117 648390
rect 516059 648322 516071 648356
rect 516105 648322 516117 648356
rect 516059 648288 516117 648322
rect 516059 648254 516071 648288
rect 516105 648254 516117 648288
rect 516059 648213 516117 648254
rect 516517 649172 516575 649213
rect 516517 649138 516529 649172
rect 516563 649138 516575 649172
rect 516517 649104 516575 649138
rect 516517 649070 516529 649104
rect 516563 649070 516575 649104
rect 516517 649036 516575 649070
rect 516517 649002 516529 649036
rect 516563 649002 516575 649036
rect 516517 648968 516575 649002
rect 516517 648934 516529 648968
rect 516563 648934 516575 648968
rect 516517 648900 516575 648934
rect 516517 648866 516529 648900
rect 516563 648866 516575 648900
rect 516517 648832 516575 648866
rect 516517 648798 516529 648832
rect 516563 648798 516575 648832
rect 516517 648764 516575 648798
rect 516517 648730 516529 648764
rect 516563 648730 516575 648764
rect 516517 648696 516575 648730
rect 516517 648662 516529 648696
rect 516563 648662 516575 648696
rect 516517 648628 516575 648662
rect 516517 648594 516529 648628
rect 516563 648594 516575 648628
rect 516517 648560 516575 648594
rect 516517 648526 516529 648560
rect 516563 648526 516575 648560
rect 516517 648492 516575 648526
rect 516517 648458 516529 648492
rect 516563 648458 516575 648492
rect 516517 648424 516575 648458
rect 516517 648390 516529 648424
rect 516563 648390 516575 648424
rect 516517 648356 516575 648390
rect 516517 648322 516529 648356
rect 516563 648322 516575 648356
rect 516517 648288 516575 648322
rect 516517 648254 516529 648288
rect 516563 648254 516575 648288
rect 516517 648213 516575 648254
rect 516975 649172 517033 649213
rect 516975 649138 516987 649172
rect 517021 649138 517033 649172
rect 516975 649104 517033 649138
rect 516975 649070 516987 649104
rect 517021 649070 517033 649104
rect 516975 649036 517033 649070
rect 516975 649002 516987 649036
rect 517021 649002 517033 649036
rect 516975 648968 517033 649002
rect 516975 648934 516987 648968
rect 517021 648934 517033 648968
rect 516975 648900 517033 648934
rect 516975 648866 516987 648900
rect 517021 648866 517033 648900
rect 516975 648832 517033 648866
rect 516975 648798 516987 648832
rect 517021 648798 517033 648832
rect 516975 648764 517033 648798
rect 516975 648730 516987 648764
rect 517021 648730 517033 648764
rect 516975 648696 517033 648730
rect 516975 648662 516987 648696
rect 517021 648662 517033 648696
rect 516975 648628 517033 648662
rect 516975 648594 516987 648628
rect 517021 648594 517033 648628
rect 516975 648560 517033 648594
rect 516975 648526 516987 648560
rect 517021 648526 517033 648560
rect 516975 648492 517033 648526
rect 516975 648458 516987 648492
rect 517021 648458 517033 648492
rect 516975 648424 517033 648458
rect 516975 648390 516987 648424
rect 517021 648390 517033 648424
rect 516975 648356 517033 648390
rect 516975 648322 516987 648356
rect 517021 648322 517033 648356
rect 516975 648288 517033 648322
rect 516975 648254 516987 648288
rect 517021 648254 517033 648288
rect 516975 648213 517033 648254
rect 517433 649172 517491 649213
rect 517433 649138 517445 649172
rect 517479 649138 517491 649172
rect 517433 649104 517491 649138
rect 517433 649070 517445 649104
rect 517479 649070 517491 649104
rect 517433 649036 517491 649070
rect 517433 649002 517445 649036
rect 517479 649002 517491 649036
rect 517433 648968 517491 649002
rect 517433 648934 517445 648968
rect 517479 648934 517491 648968
rect 517433 648900 517491 648934
rect 517433 648866 517445 648900
rect 517479 648866 517491 648900
rect 517433 648832 517491 648866
rect 517433 648798 517445 648832
rect 517479 648798 517491 648832
rect 517433 648764 517491 648798
rect 517433 648730 517445 648764
rect 517479 648730 517491 648764
rect 517433 648696 517491 648730
rect 517433 648662 517445 648696
rect 517479 648662 517491 648696
rect 517433 648628 517491 648662
rect 517433 648594 517445 648628
rect 517479 648594 517491 648628
rect 517433 648560 517491 648594
rect 517433 648526 517445 648560
rect 517479 648526 517491 648560
rect 517433 648492 517491 648526
rect 517433 648458 517445 648492
rect 517479 648458 517491 648492
rect 517433 648424 517491 648458
rect 517433 648390 517445 648424
rect 517479 648390 517491 648424
rect 517433 648356 517491 648390
rect 517433 648322 517445 648356
rect 517479 648322 517491 648356
rect 517433 648288 517491 648322
rect 517433 648254 517445 648288
rect 517479 648254 517491 648288
rect 517433 648213 517491 648254
rect 517551 649172 517609 649213
rect 517551 649138 517563 649172
rect 517597 649138 517609 649172
rect 517551 649104 517609 649138
rect 517551 649070 517563 649104
rect 517597 649070 517609 649104
rect 517551 649036 517609 649070
rect 517551 649002 517563 649036
rect 517597 649002 517609 649036
rect 517551 648968 517609 649002
rect 517551 648934 517563 648968
rect 517597 648934 517609 648968
rect 517551 648900 517609 648934
rect 517551 648866 517563 648900
rect 517597 648866 517609 648900
rect 517551 648832 517609 648866
rect 517551 648798 517563 648832
rect 517597 648798 517609 648832
rect 517551 648764 517609 648798
rect 517551 648730 517563 648764
rect 517597 648730 517609 648764
rect 517551 648696 517609 648730
rect 517551 648662 517563 648696
rect 517597 648662 517609 648696
rect 517551 648628 517609 648662
rect 517551 648594 517563 648628
rect 517597 648594 517609 648628
rect 517551 648560 517609 648594
rect 517551 648526 517563 648560
rect 517597 648526 517609 648560
rect 517551 648492 517609 648526
rect 517551 648458 517563 648492
rect 517597 648458 517609 648492
rect 517551 648424 517609 648458
rect 517551 648390 517563 648424
rect 517597 648390 517609 648424
rect 517551 648356 517609 648390
rect 517551 648322 517563 648356
rect 517597 648322 517609 648356
rect 517551 648288 517609 648322
rect 517551 648254 517563 648288
rect 517597 648254 517609 648288
rect 517551 648213 517609 648254
rect 518009 649172 518067 649213
rect 518009 649138 518021 649172
rect 518055 649138 518067 649172
rect 518009 649104 518067 649138
rect 518009 649070 518021 649104
rect 518055 649070 518067 649104
rect 518009 649036 518067 649070
rect 518009 649002 518021 649036
rect 518055 649002 518067 649036
rect 518009 648968 518067 649002
rect 518009 648934 518021 648968
rect 518055 648934 518067 648968
rect 518009 648900 518067 648934
rect 518009 648866 518021 648900
rect 518055 648866 518067 648900
rect 518009 648832 518067 648866
rect 518009 648798 518021 648832
rect 518055 648798 518067 648832
rect 518009 648764 518067 648798
rect 518009 648730 518021 648764
rect 518055 648730 518067 648764
rect 518009 648696 518067 648730
rect 518009 648662 518021 648696
rect 518055 648662 518067 648696
rect 518009 648628 518067 648662
rect 518009 648594 518021 648628
rect 518055 648594 518067 648628
rect 518009 648560 518067 648594
rect 518009 648526 518021 648560
rect 518055 648526 518067 648560
rect 518009 648492 518067 648526
rect 518009 648458 518021 648492
rect 518055 648458 518067 648492
rect 518009 648424 518067 648458
rect 518009 648390 518021 648424
rect 518055 648390 518067 648424
rect 518009 648356 518067 648390
rect 518009 648322 518021 648356
rect 518055 648322 518067 648356
rect 518009 648288 518067 648322
rect 518009 648254 518021 648288
rect 518055 648254 518067 648288
rect 518009 648213 518067 648254
<< mvndiffc >>
rect 514468 647293 514502 647327
rect 514468 647225 514502 647259
rect 514468 647157 514502 647191
rect 514468 647089 514502 647123
rect 514468 647021 514502 647055
rect 514468 646953 514502 646987
rect 514468 646885 514502 646919
rect 514468 646817 514502 646851
rect 514468 646749 514502 646783
rect 514468 646681 514502 646715
rect 514468 646613 514502 646647
rect 514468 646545 514502 646579
rect 514468 646477 514502 646511
rect 514468 646409 514502 646443
rect 514926 647293 514960 647327
rect 514926 647225 514960 647259
rect 514926 647157 514960 647191
rect 514926 647089 514960 647123
rect 514926 647021 514960 647055
rect 514926 646953 514960 646987
rect 514926 646885 514960 646919
rect 514926 646817 514960 646851
rect 514926 646749 514960 646783
rect 514926 646681 514960 646715
rect 514926 646613 514960 646647
rect 514926 646545 514960 646579
rect 514926 646477 514960 646511
rect 514926 646409 514960 646443
rect 515384 647293 515418 647327
rect 515384 647225 515418 647259
rect 515384 647157 515418 647191
rect 515384 647089 515418 647123
rect 515384 647021 515418 647055
rect 515384 646953 515418 646987
rect 515384 646885 515418 646919
rect 515384 646817 515418 646851
rect 515384 646749 515418 646783
rect 515384 646681 515418 646715
rect 515384 646613 515418 646647
rect 515384 646545 515418 646579
rect 515384 646477 515418 646511
rect 515384 646409 515418 646443
rect 515842 647293 515876 647327
rect 515842 647225 515876 647259
rect 515842 647157 515876 647191
rect 515842 647089 515876 647123
rect 515842 647021 515876 647055
rect 515842 646953 515876 646987
rect 515842 646885 515876 646919
rect 515842 646817 515876 646851
rect 515842 646749 515876 646783
rect 515842 646681 515876 646715
rect 515842 646613 515876 646647
rect 515842 646545 515876 646579
rect 515842 646477 515876 646511
rect 515842 646409 515876 646443
rect 516300 647293 516334 647327
rect 516300 647225 516334 647259
rect 516300 647157 516334 647191
rect 516300 647089 516334 647123
rect 516300 647021 516334 647055
rect 516300 646953 516334 646987
rect 516300 646885 516334 646919
rect 516300 646817 516334 646851
rect 516300 646749 516334 646783
rect 516300 646681 516334 646715
rect 516300 646613 516334 646647
rect 516300 646545 516334 646579
rect 516300 646477 516334 646511
rect 516300 646409 516334 646443
rect 516758 647293 516792 647327
rect 516758 647225 516792 647259
rect 516758 647157 516792 647191
rect 516758 647089 516792 647123
rect 516758 647021 516792 647055
rect 516758 646953 516792 646987
rect 516758 646885 516792 646919
rect 516758 646817 516792 646851
rect 516758 646749 516792 646783
rect 516758 646681 516792 646715
rect 516758 646613 516792 646647
rect 516758 646545 516792 646579
rect 516758 646477 516792 646511
rect 516758 646409 516792 646443
rect 517216 647293 517250 647327
rect 517216 647225 517250 647259
rect 517216 647157 517250 647191
rect 517216 647089 517250 647123
rect 517216 647021 517250 647055
rect 517216 646953 517250 646987
rect 517216 646885 517250 646919
rect 517216 646817 517250 646851
rect 517216 646749 517250 646783
rect 517216 646681 517250 646715
rect 517216 646613 517250 646647
rect 517216 646545 517250 646579
rect 517216 646477 517250 646511
rect 517216 646409 517250 646443
<< mvpdiffc >>
rect 514309 649529 514343 649563
rect 514309 649461 514343 649495
rect 514309 649393 514343 649427
rect 517367 649529 517401 649563
rect 517367 649461 517401 649495
rect 517367 649393 517401 649427
rect 513663 649138 513697 649172
rect 513663 649070 513697 649104
rect 513663 649002 513697 649036
rect 513663 648934 513697 648968
rect 513663 648866 513697 648900
rect 513663 648798 513697 648832
rect 513663 648730 513697 648764
rect 513663 648662 513697 648696
rect 513663 648594 513697 648628
rect 513663 648526 513697 648560
rect 513663 648458 513697 648492
rect 513663 648390 513697 648424
rect 513663 648322 513697 648356
rect 513663 648254 513697 648288
rect 514121 649138 514155 649172
rect 514121 649070 514155 649104
rect 514121 649002 514155 649036
rect 514121 648934 514155 648968
rect 514121 648866 514155 648900
rect 514121 648798 514155 648832
rect 514121 648730 514155 648764
rect 514121 648662 514155 648696
rect 514121 648594 514155 648628
rect 514121 648526 514155 648560
rect 514121 648458 514155 648492
rect 514121 648390 514155 648424
rect 514121 648322 514155 648356
rect 514121 648254 514155 648288
rect 514579 649138 514613 649172
rect 514579 649070 514613 649104
rect 514579 649002 514613 649036
rect 514579 648934 514613 648968
rect 514579 648866 514613 648900
rect 514579 648798 514613 648832
rect 514579 648730 514613 648764
rect 514579 648662 514613 648696
rect 514579 648594 514613 648628
rect 514579 648526 514613 648560
rect 514579 648458 514613 648492
rect 514579 648390 514613 648424
rect 514579 648322 514613 648356
rect 514579 648254 514613 648288
rect 515037 649138 515071 649172
rect 515037 649070 515071 649104
rect 515037 649002 515071 649036
rect 515037 648934 515071 648968
rect 515037 648866 515071 648900
rect 515037 648798 515071 648832
rect 515037 648730 515071 648764
rect 515037 648662 515071 648696
rect 515037 648594 515071 648628
rect 515037 648526 515071 648560
rect 515037 648458 515071 648492
rect 515037 648390 515071 648424
rect 515037 648322 515071 648356
rect 515037 648254 515071 648288
rect 515495 649138 515529 649172
rect 515495 649070 515529 649104
rect 515495 649002 515529 649036
rect 515495 648934 515529 648968
rect 515495 648866 515529 648900
rect 515495 648798 515529 648832
rect 515495 648730 515529 648764
rect 515495 648662 515529 648696
rect 515495 648594 515529 648628
rect 515495 648526 515529 648560
rect 515495 648458 515529 648492
rect 515495 648390 515529 648424
rect 515495 648322 515529 648356
rect 515495 648254 515529 648288
rect 515613 649138 515647 649172
rect 515613 649070 515647 649104
rect 515613 649002 515647 649036
rect 515613 648934 515647 648968
rect 515613 648866 515647 648900
rect 515613 648798 515647 648832
rect 515613 648730 515647 648764
rect 515613 648662 515647 648696
rect 515613 648594 515647 648628
rect 515613 648526 515647 648560
rect 515613 648458 515647 648492
rect 515613 648390 515647 648424
rect 515613 648322 515647 648356
rect 515613 648254 515647 648288
rect 516071 649138 516105 649172
rect 516071 649070 516105 649104
rect 516071 649002 516105 649036
rect 516071 648934 516105 648968
rect 516071 648866 516105 648900
rect 516071 648798 516105 648832
rect 516071 648730 516105 648764
rect 516071 648662 516105 648696
rect 516071 648594 516105 648628
rect 516071 648526 516105 648560
rect 516071 648458 516105 648492
rect 516071 648390 516105 648424
rect 516071 648322 516105 648356
rect 516071 648254 516105 648288
rect 516529 649138 516563 649172
rect 516529 649070 516563 649104
rect 516529 649002 516563 649036
rect 516529 648934 516563 648968
rect 516529 648866 516563 648900
rect 516529 648798 516563 648832
rect 516529 648730 516563 648764
rect 516529 648662 516563 648696
rect 516529 648594 516563 648628
rect 516529 648526 516563 648560
rect 516529 648458 516563 648492
rect 516529 648390 516563 648424
rect 516529 648322 516563 648356
rect 516529 648254 516563 648288
rect 516987 649138 517021 649172
rect 516987 649070 517021 649104
rect 516987 649002 517021 649036
rect 516987 648934 517021 648968
rect 516987 648866 517021 648900
rect 516987 648798 517021 648832
rect 516987 648730 517021 648764
rect 516987 648662 517021 648696
rect 516987 648594 517021 648628
rect 516987 648526 517021 648560
rect 516987 648458 517021 648492
rect 516987 648390 517021 648424
rect 516987 648322 517021 648356
rect 516987 648254 517021 648288
rect 517445 649138 517479 649172
rect 517445 649070 517479 649104
rect 517445 649002 517479 649036
rect 517445 648934 517479 648968
rect 517445 648866 517479 648900
rect 517445 648798 517479 648832
rect 517445 648730 517479 648764
rect 517445 648662 517479 648696
rect 517445 648594 517479 648628
rect 517445 648526 517479 648560
rect 517445 648458 517479 648492
rect 517445 648390 517479 648424
rect 517445 648322 517479 648356
rect 517445 648254 517479 648288
rect 517563 649138 517597 649172
rect 517563 649070 517597 649104
rect 517563 649002 517597 649036
rect 517563 648934 517597 648968
rect 517563 648866 517597 648900
rect 517563 648798 517597 648832
rect 517563 648730 517597 648764
rect 517563 648662 517597 648696
rect 517563 648594 517597 648628
rect 517563 648526 517597 648560
rect 517563 648458 517597 648492
rect 517563 648390 517597 648424
rect 517563 648322 517597 648356
rect 517563 648254 517597 648288
rect 518021 649138 518055 649172
rect 518021 649070 518055 649104
rect 518021 649002 518055 649036
rect 518021 648934 518055 648968
rect 518021 648866 518055 648900
rect 518021 648798 518055 648832
rect 518021 648730 518055 648764
rect 518021 648662 518055 648696
rect 518021 648594 518055 648628
rect 518021 648526 518055 648560
rect 518021 648458 518055 648492
rect 518021 648390 518055 648424
rect 518021 648322 518055 648356
rect 518021 648254 518055 648288
<< mvpsubdiff >>
rect 513406 647672 518312 647698
rect 513406 647666 514380 647672
rect 513406 646136 513454 647666
rect 514304 647570 514380 647666
rect 517338 647666 518312 647672
rect 517338 647570 517414 647666
rect 514304 647544 517414 647570
rect 514304 646258 514352 647544
rect 517366 646258 517414 647544
rect 514304 646232 517414 646258
rect 514304 646136 514380 646232
rect 513406 646130 514380 646136
rect 517338 646136 517414 646232
rect 518264 646136 518312 647666
rect 517338 646130 518312 646136
rect 513406 646104 518312 646130
<< mvnsubdiff >>
rect 507872 649814 507992 649848
rect 508026 649814 508060 649848
rect 508094 649814 508128 649848
rect 508162 649814 508196 649848
rect 508230 649814 508264 649848
rect 508298 649814 508332 649848
rect 508366 649814 508400 649848
rect 508434 649814 508468 649848
rect 508502 649814 508536 649848
rect 508570 649814 508604 649848
rect 508638 649814 508672 649848
rect 508706 649814 508740 649848
rect 508774 649814 508808 649848
rect 508842 649814 508876 649848
rect 508910 649814 508944 649848
rect 508978 649814 509012 649848
rect 509046 649814 509080 649848
rect 509114 649814 509148 649848
rect 509182 649814 509216 649848
rect 509250 649814 509284 649848
rect 509318 649814 509352 649848
rect 509386 649814 509420 649848
rect 509454 649814 509488 649848
rect 509522 649814 509556 649848
rect 509590 649814 509624 649848
rect 509658 649814 509692 649848
rect 509726 649814 509760 649848
rect 509794 649814 509828 649848
rect 509862 649814 509896 649848
rect 509930 649814 509964 649848
rect 509998 649814 510032 649848
rect 510066 649814 510100 649848
rect 510134 649814 510168 649848
rect 510202 649814 510236 649848
rect 510270 649814 510304 649848
rect 510338 649814 510372 649848
rect 510406 649814 510440 649848
rect 510474 649814 510508 649848
rect 510542 649814 510576 649848
rect 510610 649814 510644 649848
rect 510678 649814 510712 649848
rect 510746 649814 510780 649848
rect 510814 649814 510848 649848
rect 510882 649814 510916 649848
rect 510950 649814 510984 649848
rect 511018 649814 511052 649848
rect 511086 649814 511120 649848
rect 511154 649814 511188 649848
rect 511222 649814 511256 649848
rect 511290 649814 511324 649848
rect 511358 649814 511392 649848
rect 511426 649814 511460 649848
rect 511494 649814 511528 649848
rect 511562 649814 511596 649848
rect 511630 649814 511664 649848
rect 511698 649814 511732 649848
rect 511766 649814 511800 649848
rect 511834 649814 511868 649848
rect 511902 649814 511936 649848
rect 511970 649814 512004 649848
rect 512038 649814 512072 649848
rect 512106 649814 512140 649848
rect 512174 649814 512208 649848
rect 512242 649814 512276 649848
rect 512310 649814 512344 649848
rect 512378 649814 512412 649848
rect 512446 649814 512480 649848
rect 512514 649814 512548 649848
rect 512582 649814 512616 649848
rect 512650 649814 512684 649848
rect 512718 649814 512752 649848
rect 512786 649814 512820 649848
rect 512854 649814 512888 649848
rect 512922 649814 513047 649848
rect 507872 649736 507906 649814
rect 513013 649736 513047 649814
rect 507872 649668 507906 649702
rect 507872 649600 507906 649634
rect 507872 649532 507906 649566
rect 507872 649464 507906 649498
rect 507872 649396 507906 649430
rect 513013 649668 513047 649702
rect 513013 649600 513047 649634
rect 513013 649532 513047 649566
rect 513013 649464 513047 649498
rect 507872 649328 507906 649362
rect 507872 649260 507906 649294
rect 507872 649192 507906 649226
rect 513013 649396 513047 649430
rect 513013 649328 513047 649362
rect 513013 649260 513047 649294
rect 513013 649192 513047 649226
rect 507872 649124 507906 649158
rect 507872 649056 507906 649090
rect 507872 648988 507906 649022
rect 507872 648920 507906 648954
rect 513013 649124 513047 649158
rect 513013 649056 513047 649090
rect 513013 648988 513047 649022
rect 513013 648920 513047 648954
rect 507872 648852 507906 648886
rect 507872 648784 507906 648818
rect 507872 648716 507906 648750
rect 507872 648648 507906 648682
rect 513013 648852 513047 648886
rect 513013 648784 513047 648818
rect 513013 648716 513047 648750
rect 507872 648580 507906 648614
rect 507872 648512 507906 648546
rect 507872 648444 507906 648478
rect 507872 648376 507906 648410
rect 513013 648648 513047 648682
rect 513013 648580 513047 648614
rect 513013 648512 513047 648546
rect 513013 648444 513047 648478
rect 513013 648376 513047 648410
rect 507872 648308 507906 648342
rect 507872 648240 507906 648274
rect 507872 648172 507906 648206
rect 507872 648104 507906 648138
rect 513013 648308 513047 648342
rect 513013 648240 513047 648274
rect 513013 648172 513047 648206
rect 507872 648036 507906 648070
rect 507872 647968 507906 648002
rect 507872 647900 507906 647934
rect 507872 647832 507906 647866
rect 513013 648104 513047 648138
rect 513013 648036 513047 648070
rect 513013 647968 513047 648002
rect 513013 647900 513047 647934
rect 513406 649824 518312 649850
rect 513406 649722 513432 649824
rect 513534 649722 513598 649824
rect 518120 649722 518184 649824
rect 518286 649722 518312 649824
rect 513406 649696 518312 649722
rect 513406 649672 513560 649696
rect 513406 648074 513432 649672
rect 513534 648074 513560 649672
rect 518158 649672 518312 649696
rect 513406 648050 513560 648074
rect 518158 648074 518184 649672
rect 518286 648074 518312 649672
rect 518158 648050 518312 648074
rect 513406 648024 518312 648050
rect 513406 647922 513432 648024
rect 513534 647922 513598 648024
rect 518120 647922 518184 648024
rect 518286 647922 518312 648024
rect 513406 647896 518312 647922
rect 507872 647764 507906 647798
rect 507872 647696 507906 647730
rect 507872 647628 507906 647662
rect 507872 647560 507906 647594
rect 513013 647832 513047 647866
rect 513013 647764 513047 647798
rect 513013 647696 513047 647730
rect 513013 647628 513047 647662
rect 507872 647492 507906 647526
rect 507872 647424 507906 647458
rect 507872 647356 507906 647390
rect 507872 647288 507906 647322
rect 513013 647560 513047 647594
rect 513013 647492 513047 647526
rect 513013 647424 513047 647458
rect 513013 647356 513047 647390
rect 507872 647220 507906 647254
rect 507872 647152 507906 647186
rect 507872 647084 507906 647118
rect 513013 647288 513047 647322
rect 513013 647220 513047 647254
rect 513013 647152 513047 647186
rect 513013 647084 513047 647118
rect 507872 647016 507906 647050
rect 507872 646948 507906 646982
rect 507872 646880 507906 646914
rect 507872 646812 507906 646846
rect 507872 646744 507906 646778
rect 513013 647016 513047 647050
rect 513013 646948 513047 646982
rect 513013 646880 513047 646914
rect 513013 646812 513047 646846
rect 507872 646676 507906 646710
rect 507872 646608 507906 646642
rect 507872 646540 507906 646574
rect 513013 646744 513047 646778
rect 513013 646676 513047 646710
rect 513013 646608 513047 646642
rect 513013 646540 513047 646574
rect 507872 646472 507906 646506
rect 507872 646404 507906 646438
rect 507872 646336 507906 646370
rect 507872 646268 507906 646302
rect 513013 646472 513047 646506
rect 513013 646404 513047 646438
rect 513013 646336 513047 646370
rect 513013 646268 513047 646302
rect 507872 646142 507906 646234
rect 513013 646142 513047 646234
rect 507872 646108 507992 646142
rect 508026 646108 508060 646142
rect 508094 646108 508128 646142
rect 508162 646108 508196 646142
rect 508230 646108 508264 646142
rect 508298 646108 508332 646142
rect 508366 646108 508400 646142
rect 508434 646108 508468 646142
rect 508502 646108 508536 646142
rect 508570 646108 508604 646142
rect 508638 646108 508672 646142
rect 508706 646108 508740 646142
rect 508774 646108 508808 646142
rect 508842 646108 508876 646142
rect 508910 646108 508944 646142
rect 508978 646108 509012 646142
rect 509046 646108 509080 646142
rect 509114 646108 509148 646142
rect 509182 646108 509216 646142
rect 509250 646108 509284 646142
rect 509318 646108 509352 646142
rect 509386 646108 509420 646142
rect 509454 646108 509488 646142
rect 509522 646108 509556 646142
rect 509590 646108 509624 646142
rect 509658 646108 509692 646142
rect 509726 646108 509760 646142
rect 509794 646108 509828 646142
rect 509862 646108 509896 646142
rect 509930 646108 509964 646142
rect 509998 646108 510032 646142
rect 510066 646108 510100 646142
rect 510134 646108 510168 646142
rect 510202 646108 510236 646142
rect 510270 646108 510304 646142
rect 510338 646108 510372 646142
rect 510406 646108 510440 646142
rect 510474 646108 510508 646142
rect 510542 646108 510576 646142
rect 510610 646108 510644 646142
rect 510678 646108 510712 646142
rect 510746 646108 510780 646142
rect 510814 646108 510848 646142
rect 510882 646108 510916 646142
rect 510950 646108 510984 646142
rect 511018 646108 511052 646142
rect 511086 646108 511120 646142
rect 511154 646108 511188 646142
rect 511222 646108 511256 646142
rect 511290 646108 511324 646142
rect 511358 646108 511392 646142
rect 511426 646108 511460 646142
rect 511494 646108 511528 646142
rect 511562 646108 511596 646142
rect 511630 646108 511664 646142
rect 511698 646108 511732 646142
rect 511766 646108 511800 646142
rect 511834 646108 511868 646142
rect 511902 646108 511936 646142
rect 511970 646108 512004 646142
rect 512038 646108 512072 646142
rect 512106 646108 512140 646142
rect 512174 646108 512208 646142
rect 512242 646108 512276 646142
rect 512310 646108 512344 646142
rect 512378 646108 512412 646142
rect 512446 646108 512480 646142
rect 512514 646108 512548 646142
rect 512582 646108 512616 646142
rect 512650 646108 512684 646142
rect 512718 646108 512752 646142
rect 512786 646108 512820 646142
rect 512854 646108 512888 646142
rect 512922 646108 513047 646142
<< mvpsubdiffcont >>
rect 513454 646136 514304 647666
rect 514380 647570 517338 647672
rect 514380 646130 517338 646232
rect 517414 646136 518264 647666
<< mvnsubdiffcont >>
rect 507992 649814 508026 649848
rect 508060 649814 508094 649848
rect 508128 649814 508162 649848
rect 508196 649814 508230 649848
rect 508264 649814 508298 649848
rect 508332 649814 508366 649848
rect 508400 649814 508434 649848
rect 508468 649814 508502 649848
rect 508536 649814 508570 649848
rect 508604 649814 508638 649848
rect 508672 649814 508706 649848
rect 508740 649814 508774 649848
rect 508808 649814 508842 649848
rect 508876 649814 508910 649848
rect 508944 649814 508978 649848
rect 509012 649814 509046 649848
rect 509080 649814 509114 649848
rect 509148 649814 509182 649848
rect 509216 649814 509250 649848
rect 509284 649814 509318 649848
rect 509352 649814 509386 649848
rect 509420 649814 509454 649848
rect 509488 649814 509522 649848
rect 509556 649814 509590 649848
rect 509624 649814 509658 649848
rect 509692 649814 509726 649848
rect 509760 649814 509794 649848
rect 509828 649814 509862 649848
rect 509896 649814 509930 649848
rect 509964 649814 509998 649848
rect 510032 649814 510066 649848
rect 510100 649814 510134 649848
rect 510168 649814 510202 649848
rect 510236 649814 510270 649848
rect 510304 649814 510338 649848
rect 510372 649814 510406 649848
rect 510440 649814 510474 649848
rect 510508 649814 510542 649848
rect 510576 649814 510610 649848
rect 510644 649814 510678 649848
rect 510712 649814 510746 649848
rect 510780 649814 510814 649848
rect 510848 649814 510882 649848
rect 510916 649814 510950 649848
rect 510984 649814 511018 649848
rect 511052 649814 511086 649848
rect 511120 649814 511154 649848
rect 511188 649814 511222 649848
rect 511256 649814 511290 649848
rect 511324 649814 511358 649848
rect 511392 649814 511426 649848
rect 511460 649814 511494 649848
rect 511528 649814 511562 649848
rect 511596 649814 511630 649848
rect 511664 649814 511698 649848
rect 511732 649814 511766 649848
rect 511800 649814 511834 649848
rect 511868 649814 511902 649848
rect 511936 649814 511970 649848
rect 512004 649814 512038 649848
rect 512072 649814 512106 649848
rect 512140 649814 512174 649848
rect 512208 649814 512242 649848
rect 512276 649814 512310 649848
rect 512344 649814 512378 649848
rect 512412 649814 512446 649848
rect 512480 649814 512514 649848
rect 512548 649814 512582 649848
rect 512616 649814 512650 649848
rect 512684 649814 512718 649848
rect 512752 649814 512786 649848
rect 512820 649814 512854 649848
rect 512888 649814 512922 649848
rect 507872 649702 507906 649736
rect 507872 649634 507906 649668
rect 507872 649566 507906 649600
rect 507872 649498 507906 649532
rect 507872 649430 507906 649464
rect 513013 649702 513047 649736
rect 513013 649634 513047 649668
rect 513013 649566 513047 649600
rect 513013 649498 513047 649532
rect 513013 649430 513047 649464
rect 507872 649362 507906 649396
rect 507872 649294 507906 649328
rect 507872 649226 507906 649260
rect 507872 649158 507906 649192
rect 513013 649362 513047 649396
rect 513013 649294 513047 649328
rect 513013 649226 513047 649260
rect 507872 649090 507906 649124
rect 507872 649022 507906 649056
rect 507872 648954 507906 648988
rect 507872 648886 507906 648920
rect 513013 649158 513047 649192
rect 513013 649090 513047 649124
rect 513013 649022 513047 649056
rect 513013 648954 513047 648988
rect 507872 648818 507906 648852
rect 507872 648750 507906 648784
rect 507872 648682 507906 648716
rect 513013 648886 513047 648920
rect 513013 648818 513047 648852
rect 513013 648750 513047 648784
rect 513013 648682 513047 648716
rect 507872 648614 507906 648648
rect 507872 648546 507906 648580
rect 507872 648478 507906 648512
rect 507872 648410 507906 648444
rect 507872 648342 507906 648376
rect 513013 648614 513047 648648
rect 513013 648546 513047 648580
rect 513013 648478 513047 648512
rect 513013 648410 513047 648444
rect 507872 648274 507906 648308
rect 507872 648206 507906 648240
rect 507872 648138 507906 648172
rect 513013 648342 513047 648376
rect 513013 648274 513047 648308
rect 513013 648206 513047 648240
rect 513013 648138 513047 648172
rect 507872 648070 507906 648104
rect 507872 648002 507906 648036
rect 507872 647934 507906 647968
rect 507872 647866 507906 647900
rect 513013 648070 513047 648104
rect 513013 648002 513047 648036
rect 513013 647934 513047 647968
rect 513013 647866 513047 647900
rect 513432 649722 513534 649824
rect 513598 649722 518120 649824
rect 518184 649722 518286 649824
rect 513432 648074 513534 649672
rect 518184 648074 518286 649672
rect 513432 647922 513534 648024
rect 513598 647922 518120 648024
rect 518184 647922 518286 648024
rect 507872 647798 507906 647832
rect 507872 647730 507906 647764
rect 507872 647662 507906 647696
rect 507872 647594 507906 647628
rect 513013 647798 513047 647832
rect 513013 647730 513047 647764
rect 513013 647662 513047 647696
rect 513013 647594 513047 647628
rect 507872 647526 507906 647560
rect 507872 647458 507906 647492
rect 507872 647390 507906 647424
rect 507872 647322 507906 647356
rect 513013 647526 513047 647560
rect 513013 647458 513047 647492
rect 513013 647390 513047 647424
rect 513013 647322 513047 647356
rect 507872 647254 507906 647288
rect 507872 647186 507906 647220
rect 507872 647118 507906 647152
rect 507872 647050 507906 647084
rect 513013 647254 513047 647288
rect 513013 647186 513047 647220
rect 513013 647118 513047 647152
rect 507872 646982 507906 647016
rect 507872 646914 507906 646948
rect 507872 646846 507906 646880
rect 507872 646778 507906 646812
rect 513013 647050 513047 647084
rect 513013 646982 513047 647016
rect 513013 646914 513047 646948
rect 513013 646846 513047 646880
rect 513013 646778 513047 646812
rect 507872 646710 507906 646744
rect 507872 646642 507906 646676
rect 507872 646574 507906 646608
rect 507872 646506 507906 646540
rect 513013 646710 513047 646744
rect 513013 646642 513047 646676
rect 513013 646574 513047 646608
rect 507872 646438 507906 646472
rect 507872 646370 507906 646404
rect 507872 646302 507906 646336
rect 507872 646234 507906 646268
rect 513013 646506 513047 646540
rect 513013 646438 513047 646472
rect 513013 646370 513047 646404
rect 513013 646302 513047 646336
rect 513013 646234 513047 646268
rect 507992 646108 508026 646142
rect 508060 646108 508094 646142
rect 508128 646108 508162 646142
rect 508196 646108 508230 646142
rect 508264 646108 508298 646142
rect 508332 646108 508366 646142
rect 508400 646108 508434 646142
rect 508468 646108 508502 646142
rect 508536 646108 508570 646142
rect 508604 646108 508638 646142
rect 508672 646108 508706 646142
rect 508740 646108 508774 646142
rect 508808 646108 508842 646142
rect 508876 646108 508910 646142
rect 508944 646108 508978 646142
rect 509012 646108 509046 646142
rect 509080 646108 509114 646142
rect 509148 646108 509182 646142
rect 509216 646108 509250 646142
rect 509284 646108 509318 646142
rect 509352 646108 509386 646142
rect 509420 646108 509454 646142
rect 509488 646108 509522 646142
rect 509556 646108 509590 646142
rect 509624 646108 509658 646142
rect 509692 646108 509726 646142
rect 509760 646108 509794 646142
rect 509828 646108 509862 646142
rect 509896 646108 509930 646142
rect 509964 646108 509998 646142
rect 510032 646108 510066 646142
rect 510100 646108 510134 646142
rect 510168 646108 510202 646142
rect 510236 646108 510270 646142
rect 510304 646108 510338 646142
rect 510372 646108 510406 646142
rect 510440 646108 510474 646142
rect 510508 646108 510542 646142
rect 510576 646108 510610 646142
rect 510644 646108 510678 646142
rect 510712 646108 510746 646142
rect 510780 646108 510814 646142
rect 510848 646108 510882 646142
rect 510916 646108 510950 646142
rect 510984 646108 511018 646142
rect 511052 646108 511086 646142
rect 511120 646108 511154 646142
rect 511188 646108 511222 646142
rect 511256 646108 511290 646142
rect 511324 646108 511358 646142
rect 511392 646108 511426 646142
rect 511460 646108 511494 646142
rect 511528 646108 511562 646142
rect 511596 646108 511630 646142
rect 511664 646108 511698 646142
rect 511732 646108 511766 646142
rect 511800 646108 511834 646142
rect 511868 646108 511902 646142
rect 511936 646108 511970 646142
rect 512004 646108 512038 646142
rect 512072 646108 512106 646142
rect 512140 646108 512174 646142
rect 512208 646108 512242 646142
rect 512276 646108 512310 646142
rect 512344 646108 512378 646142
rect 512412 646108 512446 646142
rect 512480 646108 512514 646142
rect 512548 646108 512582 646142
rect 512616 646108 512650 646142
rect 512684 646108 512718 646142
rect 512752 646108 512786 646142
rect 512820 646108 512854 646142
rect 512888 646108 512922 646142
<< poly >>
rect 514355 649578 517355 649604
rect 514355 649331 517355 649378
rect 514355 649297 514376 649331
rect 514410 649297 514444 649331
rect 514478 649297 514512 649331
rect 514546 649297 514580 649331
rect 514614 649297 514648 649331
rect 514682 649297 514716 649331
rect 514750 649297 514784 649331
rect 514818 649297 514852 649331
rect 514886 649297 514920 649331
rect 514954 649297 514988 649331
rect 515022 649297 515056 649331
rect 515090 649297 515124 649331
rect 515158 649297 515192 649331
rect 515226 649297 515260 649331
rect 515294 649297 515328 649331
rect 515362 649297 515396 649331
rect 515430 649297 515464 649331
rect 515498 649297 515532 649331
rect 515566 649297 515600 649331
rect 515634 649297 515668 649331
rect 515702 649297 515736 649331
rect 515770 649297 515804 649331
rect 515838 649297 515872 649331
rect 515906 649297 515940 649331
rect 515974 649297 516008 649331
rect 516042 649297 516076 649331
rect 516110 649297 516144 649331
rect 516178 649297 516212 649331
rect 516246 649297 516280 649331
rect 516314 649297 516348 649331
rect 516382 649297 516416 649331
rect 516450 649297 516484 649331
rect 516518 649297 516552 649331
rect 516586 649297 516620 649331
rect 516654 649297 516688 649331
rect 516722 649297 516756 649331
rect 516790 649297 516824 649331
rect 516858 649297 516892 649331
rect 516926 649297 516960 649331
rect 516994 649297 517028 649331
rect 517062 649297 517096 649331
rect 517130 649297 517164 649331
rect 517198 649297 517232 649331
rect 517266 649297 517300 649331
rect 517334 649297 517355 649331
rect 514355 649281 517355 649297
rect 513709 649213 514109 649239
rect 514167 649213 514567 649239
rect 514625 649213 515025 649239
rect 515083 649213 515483 649239
rect 515659 649213 516059 649239
rect 516117 649213 516517 649239
rect 516575 649213 516975 649239
rect 517033 649213 517433 649239
rect 517609 649213 518009 649239
rect 513709 648166 514109 648213
rect 513709 648132 513756 648166
rect 513790 648132 513824 648166
rect 513858 648132 513892 648166
rect 513926 648132 513960 648166
rect 513994 648132 514028 648166
rect 514062 648132 514109 648166
rect 513709 648116 514109 648132
rect 514167 648166 514567 648213
rect 514167 648132 514214 648166
rect 514248 648132 514282 648166
rect 514316 648132 514350 648166
rect 514384 648132 514418 648166
rect 514452 648132 514486 648166
rect 514520 648132 514567 648166
rect 514167 648116 514567 648132
rect 514625 648166 515025 648213
rect 514625 648132 514672 648166
rect 514706 648132 514740 648166
rect 514774 648132 514808 648166
rect 514842 648132 514876 648166
rect 514910 648132 514944 648166
rect 514978 648132 515025 648166
rect 514625 648116 515025 648132
rect 515083 648166 515483 648213
rect 515083 648132 515130 648166
rect 515164 648132 515198 648166
rect 515232 648132 515266 648166
rect 515300 648132 515334 648166
rect 515368 648132 515402 648166
rect 515436 648132 515483 648166
rect 515083 648116 515483 648132
rect 515659 648166 516059 648213
rect 515659 648132 515706 648166
rect 515740 648132 515774 648166
rect 515808 648132 515842 648166
rect 515876 648132 515910 648166
rect 515944 648132 515978 648166
rect 516012 648132 516059 648166
rect 515659 648116 516059 648132
rect 516117 648166 516517 648213
rect 516117 648132 516164 648166
rect 516198 648132 516232 648166
rect 516266 648132 516300 648166
rect 516334 648132 516368 648166
rect 516402 648132 516436 648166
rect 516470 648132 516517 648166
rect 516117 648116 516517 648132
rect 516575 648166 516975 648213
rect 516575 648132 516622 648166
rect 516656 648132 516690 648166
rect 516724 648132 516758 648166
rect 516792 648132 516826 648166
rect 516860 648132 516894 648166
rect 516928 648132 516975 648166
rect 516575 648116 516975 648132
rect 517033 648166 517433 648213
rect 517033 648132 517080 648166
rect 517114 648132 517148 648166
rect 517182 648132 517216 648166
rect 517250 648132 517284 648166
rect 517318 648132 517352 648166
rect 517386 648132 517433 648166
rect 517033 648116 517433 648132
rect 517609 648166 518009 648213
rect 517609 648132 517656 648166
rect 517690 648132 517724 648166
rect 517758 648132 517792 648166
rect 517826 648132 517860 648166
rect 517894 648132 517928 648166
rect 517962 648132 518009 648166
rect 517609 648116 518009 648132
rect 514514 647440 514914 647456
rect 514514 647406 514561 647440
rect 514595 647406 514629 647440
rect 514663 647406 514697 647440
rect 514731 647406 514765 647440
rect 514799 647406 514833 647440
rect 514867 647406 514914 647440
rect 514514 647368 514914 647406
rect 514972 647440 515372 647456
rect 514972 647406 515019 647440
rect 515053 647406 515087 647440
rect 515121 647406 515155 647440
rect 515189 647406 515223 647440
rect 515257 647406 515291 647440
rect 515325 647406 515372 647440
rect 514972 647368 515372 647406
rect 515430 647440 515830 647456
rect 515430 647406 515477 647440
rect 515511 647406 515545 647440
rect 515579 647406 515613 647440
rect 515647 647406 515681 647440
rect 515715 647406 515749 647440
rect 515783 647406 515830 647440
rect 515430 647368 515830 647406
rect 515888 647440 516288 647456
rect 515888 647406 515935 647440
rect 515969 647406 516003 647440
rect 516037 647406 516071 647440
rect 516105 647406 516139 647440
rect 516173 647406 516207 647440
rect 516241 647406 516288 647440
rect 515888 647368 516288 647406
rect 516346 647440 516746 647456
rect 516346 647406 516393 647440
rect 516427 647406 516461 647440
rect 516495 647406 516529 647440
rect 516563 647406 516597 647440
rect 516631 647406 516665 647440
rect 516699 647406 516746 647440
rect 516346 647368 516746 647406
rect 516804 647440 517204 647456
rect 516804 647406 516851 647440
rect 516885 647406 516919 647440
rect 516953 647406 516987 647440
rect 517021 647406 517055 647440
rect 517089 647406 517123 647440
rect 517157 647406 517204 647440
rect 516804 647368 517204 647406
rect 514514 646342 514914 646368
rect 514972 646342 515372 646368
rect 515430 646342 515830 646368
rect 515888 646342 516288 646368
rect 516346 646342 516746 646368
rect 516804 646342 517204 646368
<< polycont >>
rect 514376 649297 514410 649331
rect 514444 649297 514478 649331
rect 514512 649297 514546 649331
rect 514580 649297 514614 649331
rect 514648 649297 514682 649331
rect 514716 649297 514750 649331
rect 514784 649297 514818 649331
rect 514852 649297 514886 649331
rect 514920 649297 514954 649331
rect 514988 649297 515022 649331
rect 515056 649297 515090 649331
rect 515124 649297 515158 649331
rect 515192 649297 515226 649331
rect 515260 649297 515294 649331
rect 515328 649297 515362 649331
rect 515396 649297 515430 649331
rect 515464 649297 515498 649331
rect 515532 649297 515566 649331
rect 515600 649297 515634 649331
rect 515668 649297 515702 649331
rect 515736 649297 515770 649331
rect 515804 649297 515838 649331
rect 515872 649297 515906 649331
rect 515940 649297 515974 649331
rect 516008 649297 516042 649331
rect 516076 649297 516110 649331
rect 516144 649297 516178 649331
rect 516212 649297 516246 649331
rect 516280 649297 516314 649331
rect 516348 649297 516382 649331
rect 516416 649297 516450 649331
rect 516484 649297 516518 649331
rect 516552 649297 516586 649331
rect 516620 649297 516654 649331
rect 516688 649297 516722 649331
rect 516756 649297 516790 649331
rect 516824 649297 516858 649331
rect 516892 649297 516926 649331
rect 516960 649297 516994 649331
rect 517028 649297 517062 649331
rect 517096 649297 517130 649331
rect 517164 649297 517198 649331
rect 517232 649297 517266 649331
rect 517300 649297 517334 649331
rect 513756 648132 513790 648166
rect 513824 648132 513858 648166
rect 513892 648132 513926 648166
rect 513960 648132 513994 648166
rect 514028 648132 514062 648166
rect 514214 648132 514248 648166
rect 514282 648132 514316 648166
rect 514350 648132 514384 648166
rect 514418 648132 514452 648166
rect 514486 648132 514520 648166
rect 514672 648132 514706 648166
rect 514740 648132 514774 648166
rect 514808 648132 514842 648166
rect 514876 648132 514910 648166
rect 514944 648132 514978 648166
rect 515130 648132 515164 648166
rect 515198 648132 515232 648166
rect 515266 648132 515300 648166
rect 515334 648132 515368 648166
rect 515402 648132 515436 648166
rect 515706 648132 515740 648166
rect 515774 648132 515808 648166
rect 515842 648132 515876 648166
rect 515910 648132 515944 648166
rect 515978 648132 516012 648166
rect 516164 648132 516198 648166
rect 516232 648132 516266 648166
rect 516300 648132 516334 648166
rect 516368 648132 516402 648166
rect 516436 648132 516470 648166
rect 516622 648132 516656 648166
rect 516690 648132 516724 648166
rect 516758 648132 516792 648166
rect 516826 648132 516860 648166
rect 516894 648132 516928 648166
rect 517080 648132 517114 648166
rect 517148 648132 517182 648166
rect 517216 648132 517250 648166
rect 517284 648132 517318 648166
rect 517352 648132 517386 648166
rect 517656 648132 517690 648166
rect 517724 648132 517758 648166
rect 517792 648132 517826 648166
rect 517860 648132 517894 648166
rect 517928 648132 517962 648166
rect 514561 647406 514595 647440
rect 514629 647406 514663 647440
rect 514697 647406 514731 647440
rect 514765 647406 514799 647440
rect 514833 647406 514867 647440
rect 515019 647406 515053 647440
rect 515087 647406 515121 647440
rect 515155 647406 515189 647440
rect 515223 647406 515257 647440
rect 515291 647406 515325 647440
rect 515477 647406 515511 647440
rect 515545 647406 515579 647440
rect 515613 647406 515647 647440
rect 515681 647406 515715 647440
rect 515749 647406 515783 647440
rect 515935 647406 515969 647440
rect 516003 647406 516037 647440
rect 516071 647406 516105 647440
rect 516139 647406 516173 647440
rect 516207 647406 516241 647440
rect 516393 647406 516427 647440
rect 516461 647406 516495 647440
rect 516529 647406 516563 647440
rect 516597 647406 516631 647440
rect 516665 647406 516699 647440
rect 516851 647406 516885 647440
rect 516919 647406 516953 647440
rect 516987 647406 517021 647440
rect 517055 647406 517089 647440
rect 517123 647406 517157 647440
<< xpolycontact >>
rect 508013 649427 508445 649709
rect 512473 649427 512905 649709
rect 508013 648897 508445 649179
rect 512473 648897 512905 649179
rect 508011 648367 508443 648649
rect 512471 648367 512903 648649
rect 508011 647837 508443 648119
rect 512471 647837 512903 648119
rect 508011 647307 508443 647589
rect 512471 647307 512903 647589
rect 508011 646777 508443 647059
rect 512471 646777 512903 647059
rect 508011 646247 508443 646529
rect 512471 646247 512903 646529
<< ppolyres >>
rect 508445 649427 512473 649709
rect 508445 648897 512473 649179
rect 508443 648367 512471 648649
rect 508443 647837 512471 648119
rect 508443 647307 512471 647589
rect 508443 646777 512471 647059
rect 508443 646247 512471 646529
<< locali >>
rect 507872 649814 507992 649848
rect 508026 649814 508060 649848
rect 508094 649814 508128 649848
rect 508162 649814 508196 649848
rect 508230 649814 508264 649848
rect 508298 649814 508332 649848
rect 508366 649814 508400 649848
rect 508434 649814 508468 649848
rect 508502 649814 508536 649848
rect 508570 649814 508604 649848
rect 508638 649814 508672 649848
rect 508706 649814 508740 649848
rect 508774 649814 508808 649848
rect 508842 649814 508876 649848
rect 508910 649814 508944 649848
rect 508978 649814 509012 649848
rect 509046 649814 509080 649848
rect 509114 649814 509148 649848
rect 509182 649814 509216 649848
rect 509250 649814 509284 649848
rect 509318 649814 509352 649848
rect 509386 649814 509420 649848
rect 509454 649814 509488 649848
rect 509522 649814 509556 649848
rect 509590 649814 509624 649848
rect 509658 649814 509692 649848
rect 509726 649814 509760 649848
rect 509794 649814 509828 649848
rect 509862 649814 509896 649848
rect 509930 649814 509964 649848
rect 509998 649814 510032 649848
rect 510066 649814 510100 649848
rect 510134 649814 510168 649848
rect 510202 649814 510236 649848
rect 510270 649814 510304 649848
rect 510338 649814 510372 649848
rect 510406 649814 510440 649848
rect 510474 649814 510508 649848
rect 510542 649814 510576 649848
rect 510610 649814 510644 649848
rect 510678 649814 510712 649848
rect 510746 649814 510780 649848
rect 510814 649814 510848 649848
rect 510882 649814 510916 649848
rect 510950 649814 510984 649848
rect 511018 649814 511052 649848
rect 511086 649814 511120 649848
rect 511154 649814 511188 649848
rect 511222 649814 511256 649848
rect 511290 649814 511324 649848
rect 511358 649814 511392 649848
rect 511426 649814 511460 649848
rect 511494 649814 511528 649848
rect 511562 649814 511596 649848
rect 511630 649814 511664 649848
rect 511698 649814 511732 649848
rect 511766 649814 511800 649848
rect 511834 649814 511868 649848
rect 511902 649814 511936 649848
rect 511970 649814 512004 649848
rect 512038 649814 512072 649848
rect 512106 649814 512140 649848
rect 512174 649814 512208 649848
rect 512242 649814 512276 649848
rect 512310 649814 512344 649848
rect 512378 649814 512412 649848
rect 512446 649814 512480 649848
rect 512514 649814 512548 649848
rect 512582 649814 512616 649848
rect 512650 649814 512684 649848
rect 512718 649814 512752 649848
rect 512786 649814 512820 649848
rect 512854 649814 512888 649848
rect 512922 649842 513047 649848
rect 512922 649824 518304 649842
rect 512922 649814 513432 649824
rect 507872 649736 507906 649814
rect 513013 649793 513432 649814
rect 513013 649736 513147 649793
rect 507872 649668 507906 649702
rect 507872 649600 507906 649634
rect 507872 649532 507906 649566
rect 507872 649464 507906 649498
rect 507872 649396 507906 649430
rect 513047 649702 513147 649736
rect 513013 649668 513147 649702
rect 513047 649634 513147 649668
rect 513013 649600 513147 649634
rect 513047 649566 513147 649600
rect 513013 649532 513147 649566
rect 513047 649498 513147 649532
rect 513013 649464 513147 649498
rect 513047 649430 513147 649464
rect 507872 649328 507906 649362
rect 507872 649260 507906 649294
rect 507872 649192 507906 649226
rect 513013 649396 513147 649430
rect 513047 649362 513147 649396
rect 513013 649328 513147 649362
rect 513047 649294 513147 649328
rect 513013 649260 513147 649294
rect 513047 649226 513147 649260
rect 513013 649192 513147 649226
rect 507872 649124 507906 649158
rect 507872 649056 507906 649090
rect 507872 648988 507906 649022
rect 507872 648920 507906 648954
rect 513047 649158 513147 649192
rect 513013 649124 513147 649158
rect 513047 649090 513147 649124
rect 513013 649056 513147 649090
rect 513047 649022 513147 649056
rect 513013 648988 513147 649022
rect 513047 648954 513147 648988
rect 513013 648920 513147 648954
rect 507872 648852 507906 648886
rect 507872 648784 507906 648818
rect 507872 648716 507906 648750
rect 507872 648648 507906 648682
rect 513047 648886 513147 648920
rect 513013 648852 513147 648886
rect 513047 648818 513147 648852
rect 513013 648784 513147 648818
rect 513047 648750 513147 648784
rect 513013 648716 513147 648750
rect 513047 648682 513147 648716
rect 507872 648580 507906 648614
rect 507872 648512 507906 648546
rect 507872 648444 507906 648478
rect 507872 648376 507906 648410
rect 513013 648648 513147 648682
rect 513047 648614 513147 648648
rect 513013 648580 513147 648614
rect 513047 648546 513147 648580
rect 513013 648512 513147 648546
rect 513047 648478 513147 648512
rect 513013 648444 513147 648478
rect 513047 648410 513147 648444
rect 513013 648376 513147 648410
rect 507872 648308 507906 648342
rect 507872 648240 507906 648274
rect 507872 648172 507906 648206
rect 507872 648104 507906 648138
rect 513047 648342 513147 648376
rect 513013 648308 513147 648342
rect 513047 648274 513147 648308
rect 513013 648240 513147 648274
rect 513047 648206 513147 648240
rect 513013 648172 513147 648206
rect 513047 648138 513147 648172
rect 507872 648036 507906 648070
rect 507872 647968 507906 648002
rect 507872 647900 507906 647934
rect 507872 647832 507906 647866
rect 513013 648104 513147 648138
rect 513047 648070 513147 648104
rect 513013 648036 513147 648070
rect 513047 648002 513147 648036
rect 513013 647968 513147 648002
rect 513047 647934 513147 647968
rect 513013 647900 513147 647934
rect 513047 647866 513147 647900
rect 507872 647764 507906 647798
rect 507872 647696 507906 647730
rect 507872 647628 507906 647662
rect 507872 647560 507906 647594
rect 513013 647832 513147 647866
rect 513047 647798 513147 647832
rect 513013 647764 513147 647798
rect 513047 647730 513147 647764
rect 513013 647696 513147 647730
rect 513047 647662 513147 647696
rect 513013 647628 513147 647662
rect 513047 647594 513147 647628
rect 507872 647492 507906 647526
rect 507872 647424 507906 647458
rect 507872 647356 507906 647390
rect 507872 647288 507906 647322
rect 513013 647560 513147 647594
rect 513047 647526 513147 647560
rect 513013 647492 513147 647526
rect 513047 647458 513147 647492
rect 513013 647424 513147 647458
rect 513047 647390 513147 647424
rect 513013 647356 513147 647390
rect 513047 647322 513147 647356
rect 507872 647220 507906 647254
rect 507872 647152 507906 647186
rect 507872 647084 507906 647118
rect 513013 647288 513147 647322
rect 513047 647254 513147 647288
rect 513013 647220 513147 647254
rect 513047 647186 513147 647220
rect 513013 647152 513147 647186
rect 513047 647118 513147 647152
rect 513013 647084 513147 647118
rect 507872 647016 507906 647050
rect 507872 646948 507906 646982
rect 507872 646880 507906 646914
rect 507872 646812 507906 646846
rect 507872 646744 507906 646778
rect 513047 647050 513147 647084
rect 513013 647016 513147 647050
rect 513047 646982 513147 647016
rect 513013 646948 513147 646982
rect 513047 646914 513147 646948
rect 513013 646880 513147 646914
rect 513047 646846 513147 646880
rect 513013 646812 513147 646846
rect 513047 646778 513147 646812
rect 507872 646676 507906 646710
rect 507872 646608 507906 646642
rect 507872 646540 507906 646574
rect 513013 646744 513147 646778
rect 513047 646710 513147 646744
rect 513013 646676 513147 646710
rect 513047 646642 513147 646676
rect 513013 646608 513147 646642
rect 513047 646574 513147 646608
rect 513013 646540 513147 646574
rect 507872 646472 507906 646506
rect 507872 646404 507906 646438
rect 507872 646336 507906 646370
rect 507872 646268 507906 646302
rect 513047 646506 513147 646540
rect 513013 646472 513147 646506
rect 513047 646438 513147 646472
rect 513013 646404 513147 646438
rect 513047 646370 513147 646404
rect 513013 646336 513147 646370
rect 513047 646302 513147 646336
rect 513013 646268 513147 646302
rect 507872 646142 507906 646234
rect 513047 646234 513147 646268
rect 513013 646159 513147 646234
rect 513253 649722 513432 649793
rect 513534 649722 513598 649824
rect 518120 649722 518184 649824
rect 518286 649722 518304 649824
rect 513253 649704 518304 649722
rect 513253 649672 513552 649704
rect 513253 648074 513432 649672
rect 513534 648074 513552 649672
rect 518166 649672 518304 649704
rect 514309 649563 514343 649582
rect 514309 649495 514343 649497
rect 514309 649459 514343 649461
rect 514309 649374 514343 649393
rect 517367 649563 517401 649582
rect 517367 649495 517401 649497
rect 517367 649459 517401 649461
rect 517367 649374 517401 649393
rect 514355 649297 514376 649331
rect 514432 649297 514444 649331
rect 514504 649297 514512 649331
rect 514576 649297 514580 649331
rect 514682 649297 514686 649331
rect 514750 649297 514758 649331
rect 514818 649297 514830 649331
rect 514886 649297 514902 649331
rect 514954 649297 514974 649331
rect 515022 649297 515046 649331
rect 515090 649297 515118 649331
rect 515158 649297 515190 649331
rect 515226 649297 515260 649331
rect 515296 649297 515328 649331
rect 515368 649297 515396 649331
rect 515440 649297 515464 649331
rect 515512 649297 515532 649331
rect 515584 649297 515600 649331
rect 515656 649297 515668 649331
rect 515728 649297 515736 649331
rect 515800 649297 515804 649331
rect 515906 649297 515910 649331
rect 515974 649297 515982 649331
rect 516042 649297 516054 649331
rect 516110 649297 516126 649331
rect 516178 649297 516198 649331
rect 516246 649297 516270 649331
rect 516314 649297 516342 649331
rect 516382 649297 516414 649331
rect 516450 649297 516484 649331
rect 516520 649297 516552 649331
rect 516592 649297 516620 649331
rect 516664 649297 516688 649331
rect 516736 649297 516756 649331
rect 516808 649297 516824 649331
rect 516880 649297 516892 649331
rect 516952 649297 516960 649331
rect 517024 649297 517028 649331
rect 517130 649297 517134 649331
rect 517198 649297 517206 649331
rect 517266 649297 517278 649331
rect 517334 649297 517355 649331
rect 513663 649198 513697 649217
rect 513663 649126 513697 649138
rect 513663 649054 513697 649070
rect 513663 648982 513697 649002
rect 513663 648910 513697 648934
rect 513663 648838 513697 648866
rect 513663 648766 513697 648798
rect 513663 648696 513697 648730
rect 513663 648628 513697 648660
rect 513663 648560 513697 648588
rect 513663 648492 513697 648516
rect 513663 648424 513697 648444
rect 513663 648356 513697 648372
rect 513663 648288 513697 648300
rect 513663 648209 513697 648228
rect 514121 649198 514155 649217
rect 514121 649126 514155 649138
rect 514121 649054 514155 649070
rect 514121 648982 514155 649002
rect 514121 648910 514155 648934
rect 514121 648838 514155 648866
rect 514121 648766 514155 648798
rect 514121 648696 514155 648730
rect 514121 648628 514155 648660
rect 514121 648560 514155 648588
rect 514121 648492 514155 648516
rect 514121 648424 514155 648444
rect 514121 648356 514155 648372
rect 514121 648288 514155 648300
rect 514121 648209 514155 648228
rect 514579 649198 514613 649217
rect 514579 649126 514613 649138
rect 514579 649054 514613 649070
rect 514579 648982 514613 649002
rect 514579 648910 514613 648934
rect 514579 648838 514613 648866
rect 514579 648766 514613 648798
rect 514579 648696 514613 648730
rect 514579 648628 514613 648660
rect 514579 648560 514613 648588
rect 514579 648492 514613 648516
rect 514579 648424 514613 648444
rect 514579 648356 514613 648372
rect 514579 648288 514613 648300
rect 514579 648209 514613 648228
rect 515037 649198 515071 649217
rect 515037 649126 515071 649138
rect 515037 649054 515071 649070
rect 515037 648982 515071 649002
rect 515037 648910 515071 648934
rect 515037 648838 515071 648866
rect 515037 648766 515071 648798
rect 515037 648696 515071 648730
rect 515037 648628 515071 648660
rect 515037 648560 515071 648588
rect 515037 648492 515071 648516
rect 515037 648424 515071 648444
rect 515037 648356 515071 648372
rect 515037 648288 515071 648300
rect 515037 648209 515071 648228
rect 515495 649198 515529 649217
rect 515495 649126 515529 649138
rect 515495 649054 515529 649070
rect 515495 648982 515529 649002
rect 515495 648910 515529 648934
rect 515495 648838 515529 648866
rect 515495 648766 515529 648798
rect 515495 648696 515529 648730
rect 515495 648628 515529 648660
rect 515495 648560 515529 648588
rect 515495 648492 515529 648516
rect 515495 648424 515529 648444
rect 515495 648356 515529 648372
rect 515495 648288 515529 648300
rect 515495 648209 515529 648228
rect 515613 649198 515647 649217
rect 515613 649126 515647 649138
rect 515613 649054 515647 649070
rect 515613 648982 515647 649002
rect 515613 648910 515647 648934
rect 515613 648838 515647 648866
rect 515613 648766 515647 648798
rect 515613 648696 515647 648730
rect 515613 648628 515647 648660
rect 515613 648560 515647 648588
rect 515613 648492 515647 648516
rect 515613 648424 515647 648444
rect 515613 648356 515647 648372
rect 515613 648288 515647 648300
rect 515613 648209 515647 648228
rect 516071 649198 516105 649217
rect 516071 649126 516105 649138
rect 516071 649054 516105 649070
rect 516071 648982 516105 649002
rect 516071 648910 516105 648934
rect 516071 648838 516105 648866
rect 516071 648766 516105 648798
rect 516071 648696 516105 648730
rect 516071 648628 516105 648660
rect 516071 648560 516105 648588
rect 516071 648492 516105 648516
rect 516071 648424 516105 648444
rect 516071 648356 516105 648372
rect 516071 648288 516105 648300
rect 516071 648209 516105 648228
rect 516529 649198 516563 649217
rect 516529 649126 516563 649138
rect 516529 649054 516563 649070
rect 516529 648982 516563 649002
rect 516529 648910 516563 648934
rect 516529 648838 516563 648866
rect 516529 648766 516563 648798
rect 516529 648696 516563 648730
rect 516529 648628 516563 648660
rect 516529 648560 516563 648588
rect 516529 648492 516563 648516
rect 516529 648424 516563 648444
rect 516529 648356 516563 648372
rect 516529 648288 516563 648300
rect 516529 648209 516563 648228
rect 516987 649198 517021 649217
rect 516987 649126 517021 649138
rect 516987 649054 517021 649070
rect 516987 648982 517021 649002
rect 516987 648910 517021 648934
rect 516987 648838 517021 648866
rect 516987 648766 517021 648798
rect 516987 648696 517021 648730
rect 516987 648628 517021 648660
rect 516987 648560 517021 648588
rect 516987 648492 517021 648516
rect 516987 648424 517021 648444
rect 516987 648356 517021 648372
rect 516987 648288 517021 648300
rect 516987 648209 517021 648228
rect 517445 649198 517479 649217
rect 517445 649126 517479 649138
rect 517445 649054 517479 649070
rect 517445 648982 517479 649002
rect 517445 648910 517479 648934
rect 517445 648838 517479 648866
rect 517445 648766 517479 648798
rect 517445 648696 517479 648730
rect 517445 648628 517479 648660
rect 517445 648560 517479 648588
rect 517445 648492 517479 648516
rect 517445 648424 517479 648444
rect 517445 648356 517479 648372
rect 517445 648288 517479 648300
rect 517445 648209 517479 648228
rect 517563 649198 517597 649217
rect 517563 649126 517597 649138
rect 517563 649054 517597 649070
rect 517563 648982 517597 649002
rect 517563 648910 517597 648934
rect 517563 648838 517597 648866
rect 517563 648766 517597 648798
rect 517563 648696 517597 648730
rect 517563 648628 517597 648660
rect 517563 648560 517597 648588
rect 517563 648492 517597 648516
rect 517563 648424 517597 648444
rect 517563 648356 517597 648372
rect 517563 648288 517597 648300
rect 517563 648209 517597 648228
rect 518021 649198 518055 649217
rect 518021 649126 518055 649138
rect 518021 649054 518055 649070
rect 518021 648982 518055 649002
rect 518021 648910 518055 648934
rect 518021 648838 518055 648866
rect 518021 648766 518055 648798
rect 518021 648696 518055 648730
rect 518021 648628 518055 648660
rect 518021 648560 518055 648588
rect 518021 648492 518055 648516
rect 518021 648424 518055 648444
rect 518021 648356 518055 648372
rect 518021 648288 518055 648300
rect 518021 648209 518055 648228
rect 513709 648132 513748 648166
rect 513790 648132 513820 648166
rect 513858 648132 513892 648166
rect 513926 648132 513960 648166
rect 513998 648132 514028 648166
rect 514070 648132 514109 648166
rect 514167 648132 514206 648166
rect 514248 648132 514278 648166
rect 514316 648132 514350 648166
rect 514384 648132 514418 648166
rect 514456 648132 514486 648166
rect 514528 648132 514567 648166
rect 514625 648132 514664 648166
rect 514706 648132 514736 648166
rect 514774 648132 514808 648166
rect 514842 648132 514876 648166
rect 514914 648132 514944 648166
rect 514986 648132 515025 648166
rect 515083 648132 515122 648166
rect 515164 648132 515194 648166
rect 515232 648132 515266 648166
rect 515300 648132 515334 648166
rect 515372 648132 515402 648166
rect 515444 648132 515483 648166
rect 515659 648132 515698 648166
rect 515740 648132 515770 648166
rect 515808 648132 515842 648166
rect 515876 648132 515910 648166
rect 515948 648132 515978 648166
rect 516020 648132 516059 648166
rect 516117 648132 516156 648166
rect 516198 648132 516228 648166
rect 516266 648132 516300 648166
rect 516334 648132 516368 648166
rect 516406 648132 516436 648166
rect 516478 648132 516517 648166
rect 516575 648132 516614 648166
rect 516656 648132 516686 648166
rect 516724 648132 516758 648166
rect 516792 648132 516826 648166
rect 516864 648132 516894 648166
rect 516936 648132 516975 648166
rect 517033 648132 517072 648166
rect 517114 648132 517144 648166
rect 517182 648132 517216 648166
rect 517250 648132 517284 648166
rect 517322 648132 517352 648166
rect 517394 648132 517433 648166
rect 517609 648132 517648 648166
rect 517690 648132 517720 648166
rect 517758 648132 517792 648166
rect 517826 648132 517860 648166
rect 517898 648132 517928 648166
rect 517970 648132 518009 648166
rect 513253 648042 513552 648074
rect 518166 648074 518184 649672
rect 518286 648074 518304 649672
rect 518166 648042 518304 648074
rect 513253 648024 518304 648042
rect 513253 647922 513432 648024
rect 513534 647922 513598 648024
rect 518120 647922 518184 648024
rect 518286 647922 518304 648024
rect 513253 647904 518304 647922
rect 513253 646159 513293 647904
rect 513013 646142 513293 646159
rect 507872 646108 507992 646142
rect 508026 646108 508060 646142
rect 508094 646108 508128 646142
rect 508162 646108 508196 646142
rect 508230 646108 508264 646142
rect 508298 646108 508332 646142
rect 508366 646108 508400 646142
rect 508434 646108 508468 646142
rect 508502 646108 508536 646142
rect 508570 646108 508604 646142
rect 508638 646108 508672 646142
rect 508706 646108 508740 646142
rect 508774 646108 508808 646142
rect 508842 646108 508876 646142
rect 508910 646108 508944 646142
rect 508978 646108 509012 646142
rect 509046 646108 509080 646142
rect 509114 646108 509148 646142
rect 509182 646108 509216 646142
rect 509250 646108 509284 646142
rect 509318 646108 509352 646142
rect 509386 646108 509420 646142
rect 509454 646108 509488 646142
rect 509522 646108 509556 646142
rect 509590 646108 509624 646142
rect 509658 646108 509692 646142
rect 509726 646108 509760 646142
rect 509794 646108 509828 646142
rect 509862 646108 509896 646142
rect 509930 646108 509964 646142
rect 509998 646108 510032 646142
rect 510066 646108 510100 646142
rect 510134 646108 510168 646142
rect 510202 646108 510236 646142
rect 510270 646108 510304 646142
rect 510338 646108 510372 646142
rect 510406 646108 510440 646142
rect 510474 646108 510508 646142
rect 510542 646108 510576 646142
rect 510610 646108 510644 646142
rect 510678 646108 510712 646142
rect 510746 646108 510780 646142
rect 510814 646108 510848 646142
rect 510882 646108 510916 646142
rect 510950 646108 510984 646142
rect 511018 646108 511052 646142
rect 511086 646108 511120 646142
rect 511154 646108 511188 646142
rect 511222 646108 511256 646142
rect 511290 646108 511324 646142
rect 511358 646108 511392 646142
rect 511426 646108 511460 646142
rect 511494 646108 511528 646142
rect 511562 646108 511596 646142
rect 511630 646108 511664 646142
rect 511698 646108 511732 646142
rect 511766 646108 511800 646142
rect 511834 646108 511868 646142
rect 511902 646108 511936 646142
rect 511970 646108 512004 646142
rect 512038 646108 512072 646142
rect 512106 646108 512140 646142
rect 512174 646108 512208 646142
rect 512242 646108 512276 646142
rect 512310 646108 512344 646142
rect 512378 646108 512412 646142
rect 512446 646108 512480 646142
rect 512514 646108 512548 646142
rect 512582 646108 512616 646142
rect 512650 646108 512684 646142
rect 512718 646108 512752 646142
rect 512786 646108 512820 646142
rect 512854 646108 512888 646142
rect 512922 646108 513293 646142
rect 513414 647672 518304 647690
rect 513414 647666 514380 647672
rect 513414 646136 513454 647666
rect 514304 647570 514380 647666
rect 517338 647666 518304 647672
rect 517338 647570 517414 647666
rect 514304 647552 517414 647570
rect 514304 646250 514344 647552
rect 514514 647406 514553 647440
rect 514595 647406 514625 647440
rect 514663 647406 514697 647440
rect 514731 647406 514765 647440
rect 514803 647406 514833 647440
rect 514875 647406 514914 647440
rect 514972 647406 515011 647440
rect 515053 647406 515083 647440
rect 515121 647406 515155 647440
rect 515189 647406 515223 647440
rect 515261 647406 515291 647440
rect 515333 647406 515372 647440
rect 515430 647406 515469 647440
rect 515511 647406 515541 647440
rect 515579 647406 515613 647440
rect 515647 647406 515681 647440
rect 515719 647406 515749 647440
rect 515791 647406 515830 647440
rect 515888 647406 515927 647440
rect 515969 647406 515999 647440
rect 516037 647406 516071 647440
rect 516105 647406 516139 647440
rect 516177 647406 516207 647440
rect 516249 647406 516288 647440
rect 516346 647406 516385 647440
rect 516427 647406 516457 647440
rect 516495 647406 516529 647440
rect 516563 647406 516597 647440
rect 516635 647406 516665 647440
rect 516707 647406 516746 647440
rect 516804 647406 516843 647440
rect 516885 647406 516915 647440
rect 516953 647406 516987 647440
rect 517021 647406 517055 647440
rect 517093 647406 517123 647440
rect 517165 647406 517204 647440
rect 514468 647353 514502 647372
rect 514468 647281 514502 647293
rect 514468 647209 514502 647225
rect 514468 647137 514502 647157
rect 514468 647065 514502 647089
rect 514468 646993 514502 647021
rect 514468 646921 514502 646953
rect 514468 646851 514502 646885
rect 514468 646783 514502 646815
rect 514468 646715 514502 646743
rect 514468 646647 514502 646671
rect 514468 646579 514502 646599
rect 514468 646511 514502 646527
rect 514468 646443 514502 646455
rect 514468 646364 514502 646383
rect 514926 647353 514960 647372
rect 514926 647281 514960 647293
rect 514926 647209 514960 647225
rect 514926 647137 514960 647157
rect 514926 647065 514960 647089
rect 514926 646993 514960 647021
rect 514926 646921 514960 646953
rect 514926 646851 514960 646885
rect 514926 646783 514960 646815
rect 514926 646715 514960 646743
rect 514926 646647 514960 646671
rect 514926 646579 514960 646599
rect 514926 646511 514960 646527
rect 514926 646443 514960 646455
rect 514926 646364 514960 646383
rect 515384 647353 515418 647372
rect 515384 647281 515418 647293
rect 515384 647209 515418 647225
rect 515384 647137 515418 647157
rect 515384 647065 515418 647089
rect 515384 646993 515418 647021
rect 515384 646921 515418 646953
rect 515384 646851 515418 646885
rect 515384 646783 515418 646815
rect 515384 646715 515418 646743
rect 515384 646647 515418 646671
rect 515384 646579 515418 646599
rect 515384 646511 515418 646527
rect 515384 646443 515418 646455
rect 515384 646364 515418 646383
rect 515842 647353 515876 647372
rect 515842 647281 515876 647293
rect 515842 647209 515876 647225
rect 515842 647137 515876 647157
rect 515842 647065 515876 647089
rect 515842 646993 515876 647021
rect 515842 646921 515876 646953
rect 515842 646851 515876 646885
rect 515842 646783 515876 646815
rect 515842 646715 515876 646743
rect 515842 646647 515876 646671
rect 515842 646579 515876 646599
rect 515842 646511 515876 646527
rect 515842 646443 515876 646455
rect 515842 646364 515876 646383
rect 516300 647353 516334 647372
rect 516300 647281 516334 647293
rect 516300 647209 516334 647225
rect 516300 647137 516334 647157
rect 516300 647065 516334 647089
rect 516300 646993 516334 647021
rect 516300 646921 516334 646953
rect 516300 646851 516334 646885
rect 516300 646783 516334 646815
rect 516300 646715 516334 646743
rect 516300 646647 516334 646671
rect 516300 646579 516334 646599
rect 516300 646511 516334 646527
rect 516300 646443 516334 646455
rect 516300 646364 516334 646383
rect 516758 647353 516792 647372
rect 516758 647281 516792 647293
rect 516758 647209 516792 647225
rect 516758 647137 516792 647157
rect 516758 647065 516792 647089
rect 516758 646993 516792 647021
rect 516758 646921 516792 646953
rect 516758 646851 516792 646885
rect 516758 646783 516792 646815
rect 516758 646715 516792 646743
rect 516758 646647 516792 646671
rect 516758 646579 516792 646599
rect 516758 646511 516792 646527
rect 516758 646443 516792 646455
rect 516758 646364 516792 646383
rect 517216 647353 517250 647372
rect 517216 647281 517250 647293
rect 517216 647209 517250 647225
rect 517216 647137 517250 647157
rect 517216 647065 517250 647089
rect 517216 646993 517250 647021
rect 517216 646921 517250 646953
rect 517216 646851 517250 646885
rect 517216 646783 517250 646815
rect 517216 646715 517250 646743
rect 517216 646647 517250 646671
rect 517216 646579 517250 646599
rect 517216 646511 517250 646527
rect 517216 646443 517250 646455
rect 517216 646364 517250 646383
rect 517374 646250 517414 647552
rect 514304 646232 517414 646250
rect 514304 646136 514380 646232
rect 513414 646130 514380 646136
rect 517338 646136 517414 646232
rect 518264 646136 518304 647666
rect 517338 646130 518304 646136
rect 513414 646112 518304 646130
<< viali >>
rect 508033 649443 508427 649693
rect 512492 649443 512886 649693
rect 508033 648913 508427 649163
rect 512492 648913 512886 649163
rect 508030 648383 508424 648633
rect 512489 648383 512883 648633
rect 508030 647853 508424 648103
rect 512489 647853 512883 648103
rect 508030 647323 508424 647573
rect 512489 647323 512883 647573
rect 508030 646793 508424 647043
rect 512489 646793 512883 647043
rect 508030 646263 508424 646513
rect 512489 646263 512883 646513
rect 513147 646159 513253 649793
rect 514309 649529 514343 649531
rect 514309 649497 514343 649529
rect 514309 649427 514343 649459
rect 514309 649425 514343 649427
rect 517367 649529 517401 649531
rect 517367 649497 517401 649529
rect 517367 649427 517401 649459
rect 517367 649425 517401 649427
rect 514398 649297 514410 649331
rect 514410 649297 514432 649331
rect 514470 649297 514478 649331
rect 514478 649297 514504 649331
rect 514542 649297 514546 649331
rect 514546 649297 514576 649331
rect 514614 649297 514648 649331
rect 514686 649297 514716 649331
rect 514716 649297 514720 649331
rect 514758 649297 514784 649331
rect 514784 649297 514792 649331
rect 514830 649297 514852 649331
rect 514852 649297 514864 649331
rect 514902 649297 514920 649331
rect 514920 649297 514936 649331
rect 514974 649297 514988 649331
rect 514988 649297 515008 649331
rect 515046 649297 515056 649331
rect 515056 649297 515080 649331
rect 515118 649297 515124 649331
rect 515124 649297 515152 649331
rect 515190 649297 515192 649331
rect 515192 649297 515224 649331
rect 515262 649297 515294 649331
rect 515294 649297 515296 649331
rect 515334 649297 515362 649331
rect 515362 649297 515368 649331
rect 515406 649297 515430 649331
rect 515430 649297 515440 649331
rect 515478 649297 515498 649331
rect 515498 649297 515512 649331
rect 515550 649297 515566 649331
rect 515566 649297 515584 649331
rect 515622 649297 515634 649331
rect 515634 649297 515656 649331
rect 515694 649297 515702 649331
rect 515702 649297 515728 649331
rect 515766 649297 515770 649331
rect 515770 649297 515800 649331
rect 515838 649297 515872 649331
rect 515910 649297 515940 649331
rect 515940 649297 515944 649331
rect 515982 649297 516008 649331
rect 516008 649297 516016 649331
rect 516054 649297 516076 649331
rect 516076 649297 516088 649331
rect 516126 649297 516144 649331
rect 516144 649297 516160 649331
rect 516198 649297 516212 649331
rect 516212 649297 516232 649331
rect 516270 649297 516280 649331
rect 516280 649297 516304 649331
rect 516342 649297 516348 649331
rect 516348 649297 516376 649331
rect 516414 649297 516416 649331
rect 516416 649297 516448 649331
rect 516486 649297 516518 649331
rect 516518 649297 516520 649331
rect 516558 649297 516586 649331
rect 516586 649297 516592 649331
rect 516630 649297 516654 649331
rect 516654 649297 516664 649331
rect 516702 649297 516722 649331
rect 516722 649297 516736 649331
rect 516774 649297 516790 649331
rect 516790 649297 516808 649331
rect 516846 649297 516858 649331
rect 516858 649297 516880 649331
rect 516918 649297 516926 649331
rect 516926 649297 516952 649331
rect 516990 649297 516994 649331
rect 516994 649297 517024 649331
rect 517062 649297 517096 649331
rect 517134 649297 517164 649331
rect 517164 649297 517168 649331
rect 517206 649297 517232 649331
rect 517232 649297 517240 649331
rect 517278 649297 517300 649331
rect 517300 649297 517312 649331
rect 513663 649172 513697 649198
rect 513663 649164 513697 649172
rect 513663 649104 513697 649126
rect 513663 649092 513697 649104
rect 513663 649036 513697 649054
rect 513663 649020 513697 649036
rect 513663 648968 513697 648982
rect 513663 648948 513697 648968
rect 513663 648900 513697 648910
rect 513663 648876 513697 648900
rect 513663 648832 513697 648838
rect 513663 648804 513697 648832
rect 513663 648764 513697 648766
rect 513663 648732 513697 648764
rect 513663 648662 513697 648694
rect 513663 648660 513697 648662
rect 513663 648594 513697 648622
rect 513663 648588 513697 648594
rect 513663 648526 513697 648550
rect 513663 648516 513697 648526
rect 513663 648458 513697 648478
rect 513663 648444 513697 648458
rect 513663 648390 513697 648406
rect 513663 648372 513697 648390
rect 513663 648322 513697 648334
rect 513663 648300 513697 648322
rect 513663 648254 513697 648262
rect 513663 648228 513697 648254
rect 514121 649172 514155 649198
rect 514121 649164 514155 649172
rect 514121 649104 514155 649126
rect 514121 649092 514155 649104
rect 514121 649036 514155 649054
rect 514121 649020 514155 649036
rect 514121 648968 514155 648982
rect 514121 648948 514155 648968
rect 514121 648900 514155 648910
rect 514121 648876 514155 648900
rect 514121 648832 514155 648838
rect 514121 648804 514155 648832
rect 514121 648764 514155 648766
rect 514121 648732 514155 648764
rect 514121 648662 514155 648694
rect 514121 648660 514155 648662
rect 514121 648594 514155 648622
rect 514121 648588 514155 648594
rect 514121 648526 514155 648550
rect 514121 648516 514155 648526
rect 514121 648458 514155 648478
rect 514121 648444 514155 648458
rect 514121 648390 514155 648406
rect 514121 648372 514155 648390
rect 514121 648322 514155 648334
rect 514121 648300 514155 648322
rect 514121 648254 514155 648262
rect 514121 648228 514155 648254
rect 514579 649172 514613 649198
rect 514579 649164 514613 649172
rect 514579 649104 514613 649126
rect 514579 649092 514613 649104
rect 514579 649036 514613 649054
rect 514579 649020 514613 649036
rect 514579 648968 514613 648982
rect 514579 648948 514613 648968
rect 514579 648900 514613 648910
rect 514579 648876 514613 648900
rect 514579 648832 514613 648838
rect 514579 648804 514613 648832
rect 514579 648764 514613 648766
rect 514579 648732 514613 648764
rect 514579 648662 514613 648694
rect 514579 648660 514613 648662
rect 514579 648594 514613 648622
rect 514579 648588 514613 648594
rect 514579 648526 514613 648550
rect 514579 648516 514613 648526
rect 514579 648458 514613 648478
rect 514579 648444 514613 648458
rect 514579 648390 514613 648406
rect 514579 648372 514613 648390
rect 514579 648322 514613 648334
rect 514579 648300 514613 648322
rect 514579 648254 514613 648262
rect 514579 648228 514613 648254
rect 515037 649172 515071 649198
rect 515037 649164 515071 649172
rect 515037 649104 515071 649126
rect 515037 649092 515071 649104
rect 515037 649036 515071 649054
rect 515037 649020 515071 649036
rect 515037 648968 515071 648982
rect 515037 648948 515071 648968
rect 515037 648900 515071 648910
rect 515037 648876 515071 648900
rect 515037 648832 515071 648838
rect 515037 648804 515071 648832
rect 515037 648764 515071 648766
rect 515037 648732 515071 648764
rect 515037 648662 515071 648694
rect 515037 648660 515071 648662
rect 515037 648594 515071 648622
rect 515037 648588 515071 648594
rect 515037 648526 515071 648550
rect 515037 648516 515071 648526
rect 515037 648458 515071 648478
rect 515037 648444 515071 648458
rect 515037 648390 515071 648406
rect 515037 648372 515071 648390
rect 515037 648322 515071 648334
rect 515037 648300 515071 648322
rect 515037 648254 515071 648262
rect 515037 648228 515071 648254
rect 515495 649172 515529 649198
rect 515495 649164 515529 649172
rect 515495 649104 515529 649126
rect 515495 649092 515529 649104
rect 515495 649036 515529 649054
rect 515495 649020 515529 649036
rect 515495 648968 515529 648982
rect 515495 648948 515529 648968
rect 515495 648900 515529 648910
rect 515495 648876 515529 648900
rect 515495 648832 515529 648838
rect 515495 648804 515529 648832
rect 515495 648764 515529 648766
rect 515495 648732 515529 648764
rect 515495 648662 515529 648694
rect 515495 648660 515529 648662
rect 515495 648594 515529 648622
rect 515495 648588 515529 648594
rect 515495 648526 515529 648550
rect 515495 648516 515529 648526
rect 515495 648458 515529 648478
rect 515495 648444 515529 648458
rect 515495 648390 515529 648406
rect 515495 648372 515529 648390
rect 515495 648322 515529 648334
rect 515495 648300 515529 648322
rect 515495 648254 515529 648262
rect 515495 648228 515529 648254
rect 515613 649172 515647 649198
rect 515613 649164 515647 649172
rect 515613 649104 515647 649126
rect 515613 649092 515647 649104
rect 515613 649036 515647 649054
rect 515613 649020 515647 649036
rect 515613 648968 515647 648982
rect 515613 648948 515647 648968
rect 515613 648900 515647 648910
rect 515613 648876 515647 648900
rect 515613 648832 515647 648838
rect 515613 648804 515647 648832
rect 515613 648764 515647 648766
rect 515613 648732 515647 648764
rect 515613 648662 515647 648694
rect 515613 648660 515647 648662
rect 515613 648594 515647 648622
rect 515613 648588 515647 648594
rect 515613 648526 515647 648550
rect 515613 648516 515647 648526
rect 515613 648458 515647 648478
rect 515613 648444 515647 648458
rect 515613 648390 515647 648406
rect 515613 648372 515647 648390
rect 515613 648322 515647 648334
rect 515613 648300 515647 648322
rect 515613 648254 515647 648262
rect 515613 648228 515647 648254
rect 516071 649172 516105 649198
rect 516071 649164 516105 649172
rect 516071 649104 516105 649126
rect 516071 649092 516105 649104
rect 516071 649036 516105 649054
rect 516071 649020 516105 649036
rect 516071 648968 516105 648982
rect 516071 648948 516105 648968
rect 516071 648900 516105 648910
rect 516071 648876 516105 648900
rect 516071 648832 516105 648838
rect 516071 648804 516105 648832
rect 516071 648764 516105 648766
rect 516071 648732 516105 648764
rect 516071 648662 516105 648694
rect 516071 648660 516105 648662
rect 516071 648594 516105 648622
rect 516071 648588 516105 648594
rect 516071 648526 516105 648550
rect 516071 648516 516105 648526
rect 516071 648458 516105 648478
rect 516071 648444 516105 648458
rect 516071 648390 516105 648406
rect 516071 648372 516105 648390
rect 516071 648322 516105 648334
rect 516071 648300 516105 648322
rect 516071 648254 516105 648262
rect 516071 648228 516105 648254
rect 516529 649172 516563 649198
rect 516529 649164 516563 649172
rect 516529 649104 516563 649126
rect 516529 649092 516563 649104
rect 516529 649036 516563 649054
rect 516529 649020 516563 649036
rect 516529 648968 516563 648982
rect 516529 648948 516563 648968
rect 516529 648900 516563 648910
rect 516529 648876 516563 648900
rect 516529 648832 516563 648838
rect 516529 648804 516563 648832
rect 516529 648764 516563 648766
rect 516529 648732 516563 648764
rect 516529 648662 516563 648694
rect 516529 648660 516563 648662
rect 516529 648594 516563 648622
rect 516529 648588 516563 648594
rect 516529 648526 516563 648550
rect 516529 648516 516563 648526
rect 516529 648458 516563 648478
rect 516529 648444 516563 648458
rect 516529 648390 516563 648406
rect 516529 648372 516563 648390
rect 516529 648322 516563 648334
rect 516529 648300 516563 648322
rect 516529 648254 516563 648262
rect 516529 648228 516563 648254
rect 516987 649172 517021 649198
rect 516987 649164 517021 649172
rect 516987 649104 517021 649126
rect 516987 649092 517021 649104
rect 516987 649036 517021 649054
rect 516987 649020 517021 649036
rect 516987 648968 517021 648982
rect 516987 648948 517021 648968
rect 516987 648900 517021 648910
rect 516987 648876 517021 648900
rect 516987 648832 517021 648838
rect 516987 648804 517021 648832
rect 516987 648764 517021 648766
rect 516987 648732 517021 648764
rect 516987 648662 517021 648694
rect 516987 648660 517021 648662
rect 516987 648594 517021 648622
rect 516987 648588 517021 648594
rect 516987 648526 517021 648550
rect 516987 648516 517021 648526
rect 516987 648458 517021 648478
rect 516987 648444 517021 648458
rect 516987 648390 517021 648406
rect 516987 648372 517021 648390
rect 516987 648322 517021 648334
rect 516987 648300 517021 648322
rect 516987 648254 517021 648262
rect 516987 648228 517021 648254
rect 517445 649172 517479 649198
rect 517445 649164 517479 649172
rect 517445 649104 517479 649126
rect 517445 649092 517479 649104
rect 517445 649036 517479 649054
rect 517445 649020 517479 649036
rect 517445 648968 517479 648982
rect 517445 648948 517479 648968
rect 517445 648900 517479 648910
rect 517445 648876 517479 648900
rect 517445 648832 517479 648838
rect 517445 648804 517479 648832
rect 517445 648764 517479 648766
rect 517445 648732 517479 648764
rect 517445 648662 517479 648694
rect 517445 648660 517479 648662
rect 517445 648594 517479 648622
rect 517445 648588 517479 648594
rect 517445 648526 517479 648550
rect 517445 648516 517479 648526
rect 517445 648458 517479 648478
rect 517445 648444 517479 648458
rect 517445 648390 517479 648406
rect 517445 648372 517479 648390
rect 517445 648322 517479 648334
rect 517445 648300 517479 648322
rect 517445 648254 517479 648262
rect 517445 648228 517479 648254
rect 517563 649172 517597 649198
rect 517563 649164 517597 649172
rect 517563 649104 517597 649126
rect 517563 649092 517597 649104
rect 517563 649036 517597 649054
rect 517563 649020 517597 649036
rect 517563 648968 517597 648982
rect 517563 648948 517597 648968
rect 517563 648900 517597 648910
rect 517563 648876 517597 648900
rect 517563 648832 517597 648838
rect 517563 648804 517597 648832
rect 517563 648764 517597 648766
rect 517563 648732 517597 648764
rect 517563 648662 517597 648694
rect 517563 648660 517597 648662
rect 517563 648594 517597 648622
rect 517563 648588 517597 648594
rect 517563 648526 517597 648550
rect 517563 648516 517597 648526
rect 517563 648458 517597 648478
rect 517563 648444 517597 648458
rect 517563 648390 517597 648406
rect 517563 648372 517597 648390
rect 517563 648322 517597 648334
rect 517563 648300 517597 648322
rect 517563 648254 517597 648262
rect 517563 648228 517597 648254
rect 518021 649172 518055 649198
rect 518021 649164 518055 649172
rect 518021 649104 518055 649126
rect 518021 649092 518055 649104
rect 518021 649036 518055 649054
rect 518021 649020 518055 649036
rect 518021 648968 518055 648982
rect 518021 648948 518055 648968
rect 518021 648900 518055 648910
rect 518021 648876 518055 648900
rect 518021 648832 518055 648838
rect 518021 648804 518055 648832
rect 518021 648764 518055 648766
rect 518021 648732 518055 648764
rect 518021 648662 518055 648694
rect 518021 648660 518055 648662
rect 518021 648594 518055 648622
rect 518021 648588 518055 648594
rect 518021 648526 518055 648550
rect 518021 648516 518055 648526
rect 518021 648458 518055 648478
rect 518021 648444 518055 648458
rect 518021 648390 518055 648406
rect 518021 648372 518055 648390
rect 518021 648322 518055 648334
rect 518021 648300 518055 648322
rect 518021 648254 518055 648262
rect 518021 648228 518055 648254
rect 513748 648132 513756 648166
rect 513756 648132 513782 648166
rect 513820 648132 513824 648166
rect 513824 648132 513854 648166
rect 513892 648132 513926 648166
rect 513964 648132 513994 648166
rect 513994 648132 513998 648166
rect 514036 648132 514062 648166
rect 514062 648132 514070 648166
rect 514206 648132 514214 648166
rect 514214 648132 514240 648166
rect 514278 648132 514282 648166
rect 514282 648132 514312 648166
rect 514350 648132 514384 648166
rect 514422 648132 514452 648166
rect 514452 648132 514456 648166
rect 514494 648132 514520 648166
rect 514520 648132 514528 648166
rect 514664 648132 514672 648166
rect 514672 648132 514698 648166
rect 514736 648132 514740 648166
rect 514740 648132 514770 648166
rect 514808 648132 514842 648166
rect 514880 648132 514910 648166
rect 514910 648132 514914 648166
rect 514952 648132 514978 648166
rect 514978 648132 514986 648166
rect 515122 648132 515130 648166
rect 515130 648132 515156 648166
rect 515194 648132 515198 648166
rect 515198 648132 515228 648166
rect 515266 648132 515300 648166
rect 515338 648132 515368 648166
rect 515368 648132 515372 648166
rect 515410 648132 515436 648166
rect 515436 648132 515444 648166
rect 515698 648132 515706 648166
rect 515706 648132 515732 648166
rect 515770 648132 515774 648166
rect 515774 648132 515804 648166
rect 515842 648132 515876 648166
rect 515914 648132 515944 648166
rect 515944 648132 515948 648166
rect 515986 648132 516012 648166
rect 516012 648132 516020 648166
rect 516156 648132 516164 648166
rect 516164 648132 516190 648166
rect 516228 648132 516232 648166
rect 516232 648132 516262 648166
rect 516300 648132 516334 648166
rect 516372 648132 516402 648166
rect 516402 648132 516406 648166
rect 516444 648132 516470 648166
rect 516470 648132 516478 648166
rect 516614 648132 516622 648166
rect 516622 648132 516648 648166
rect 516686 648132 516690 648166
rect 516690 648132 516720 648166
rect 516758 648132 516792 648166
rect 516830 648132 516860 648166
rect 516860 648132 516864 648166
rect 516902 648132 516928 648166
rect 516928 648132 516936 648166
rect 517072 648132 517080 648166
rect 517080 648132 517106 648166
rect 517144 648132 517148 648166
rect 517148 648132 517178 648166
rect 517216 648132 517250 648166
rect 517288 648132 517318 648166
rect 517318 648132 517322 648166
rect 517360 648132 517386 648166
rect 517386 648132 517394 648166
rect 517648 648132 517656 648166
rect 517656 648132 517682 648166
rect 517720 648132 517724 648166
rect 517724 648132 517754 648166
rect 517792 648132 517826 648166
rect 517864 648132 517894 648166
rect 517894 648132 517898 648166
rect 517936 648132 517962 648166
rect 517962 648132 517970 648166
rect 518219 649614 518253 649648
rect 518219 649542 518253 649576
rect 518219 649470 518253 649504
rect 518218 649054 518252 649088
rect 518218 648982 518252 649016
rect 518218 648910 518252 648944
rect 518218 648838 518252 648872
rect 513610 646459 514148 646709
rect 514553 647406 514561 647440
rect 514561 647406 514587 647440
rect 514625 647406 514629 647440
rect 514629 647406 514659 647440
rect 514697 647406 514731 647440
rect 514769 647406 514799 647440
rect 514799 647406 514803 647440
rect 514841 647406 514867 647440
rect 514867 647406 514875 647440
rect 515011 647406 515019 647440
rect 515019 647406 515045 647440
rect 515083 647406 515087 647440
rect 515087 647406 515117 647440
rect 515155 647406 515189 647440
rect 515227 647406 515257 647440
rect 515257 647406 515261 647440
rect 515299 647406 515325 647440
rect 515325 647406 515333 647440
rect 515469 647406 515477 647440
rect 515477 647406 515503 647440
rect 515541 647406 515545 647440
rect 515545 647406 515575 647440
rect 515613 647406 515647 647440
rect 515685 647406 515715 647440
rect 515715 647406 515719 647440
rect 515757 647406 515783 647440
rect 515783 647406 515791 647440
rect 515927 647406 515935 647440
rect 515935 647406 515961 647440
rect 515999 647406 516003 647440
rect 516003 647406 516033 647440
rect 516071 647406 516105 647440
rect 516143 647406 516173 647440
rect 516173 647406 516177 647440
rect 516215 647406 516241 647440
rect 516241 647406 516249 647440
rect 516385 647406 516393 647440
rect 516393 647406 516419 647440
rect 516457 647406 516461 647440
rect 516461 647406 516491 647440
rect 516529 647406 516563 647440
rect 516601 647406 516631 647440
rect 516631 647406 516635 647440
rect 516673 647406 516699 647440
rect 516699 647406 516707 647440
rect 516843 647406 516851 647440
rect 516851 647406 516877 647440
rect 516915 647406 516919 647440
rect 516919 647406 516949 647440
rect 516987 647406 517021 647440
rect 517059 647406 517089 647440
rect 517089 647406 517093 647440
rect 517131 647406 517157 647440
rect 517157 647406 517165 647440
rect 514468 647327 514502 647353
rect 514468 647319 514502 647327
rect 514468 647259 514502 647281
rect 514468 647247 514502 647259
rect 514468 647191 514502 647209
rect 514468 647175 514502 647191
rect 514468 647123 514502 647137
rect 514468 647103 514502 647123
rect 514468 647055 514502 647065
rect 514468 647031 514502 647055
rect 514468 646987 514502 646993
rect 514468 646959 514502 646987
rect 514468 646919 514502 646921
rect 514468 646887 514502 646919
rect 514468 646817 514502 646849
rect 514468 646815 514502 646817
rect 514468 646749 514502 646777
rect 514468 646743 514502 646749
rect 514468 646681 514502 646705
rect 514468 646671 514502 646681
rect 514468 646613 514502 646633
rect 514468 646599 514502 646613
rect 514468 646545 514502 646561
rect 514468 646527 514502 646545
rect 514468 646477 514502 646489
rect 514468 646455 514502 646477
rect 514468 646409 514502 646417
rect 514468 646383 514502 646409
rect 514926 647327 514960 647353
rect 514926 647319 514960 647327
rect 514926 647259 514960 647281
rect 514926 647247 514960 647259
rect 514926 647191 514960 647209
rect 514926 647175 514960 647191
rect 514926 647123 514960 647137
rect 514926 647103 514960 647123
rect 514926 647055 514960 647065
rect 514926 647031 514960 647055
rect 514926 646987 514960 646993
rect 514926 646959 514960 646987
rect 514926 646919 514960 646921
rect 514926 646887 514960 646919
rect 514926 646817 514960 646849
rect 514926 646815 514960 646817
rect 514926 646749 514960 646777
rect 514926 646743 514960 646749
rect 514926 646681 514960 646705
rect 514926 646671 514960 646681
rect 514926 646613 514960 646633
rect 514926 646599 514960 646613
rect 514926 646545 514960 646561
rect 514926 646527 514960 646545
rect 514926 646477 514960 646489
rect 514926 646455 514960 646477
rect 514926 646409 514960 646417
rect 514926 646383 514960 646409
rect 515384 647327 515418 647353
rect 515384 647319 515418 647327
rect 515384 647259 515418 647281
rect 515384 647247 515418 647259
rect 515384 647191 515418 647209
rect 515384 647175 515418 647191
rect 515384 647123 515418 647137
rect 515384 647103 515418 647123
rect 515384 647055 515418 647065
rect 515384 647031 515418 647055
rect 515384 646987 515418 646993
rect 515384 646959 515418 646987
rect 515384 646919 515418 646921
rect 515384 646887 515418 646919
rect 515384 646817 515418 646849
rect 515384 646815 515418 646817
rect 515384 646749 515418 646777
rect 515384 646743 515418 646749
rect 515384 646681 515418 646705
rect 515384 646671 515418 646681
rect 515384 646613 515418 646633
rect 515384 646599 515418 646613
rect 515384 646545 515418 646561
rect 515384 646527 515418 646545
rect 515384 646477 515418 646489
rect 515384 646455 515418 646477
rect 515384 646409 515418 646417
rect 515384 646383 515418 646409
rect 515842 647327 515876 647353
rect 515842 647319 515876 647327
rect 515842 647259 515876 647281
rect 515842 647247 515876 647259
rect 515842 647191 515876 647209
rect 515842 647175 515876 647191
rect 515842 647123 515876 647137
rect 515842 647103 515876 647123
rect 515842 647055 515876 647065
rect 515842 647031 515876 647055
rect 515842 646987 515876 646993
rect 515842 646959 515876 646987
rect 515842 646919 515876 646921
rect 515842 646887 515876 646919
rect 515842 646817 515876 646849
rect 515842 646815 515876 646817
rect 515842 646749 515876 646777
rect 515842 646743 515876 646749
rect 515842 646681 515876 646705
rect 515842 646671 515876 646681
rect 515842 646613 515876 646633
rect 515842 646599 515876 646613
rect 515842 646545 515876 646561
rect 515842 646527 515876 646545
rect 515842 646477 515876 646489
rect 515842 646455 515876 646477
rect 515842 646409 515876 646417
rect 515842 646383 515876 646409
rect 516300 647327 516334 647353
rect 516300 647319 516334 647327
rect 516300 647259 516334 647281
rect 516300 647247 516334 647259
rect 516300 647191 516334 647209
rect 516300 647175 516334 647191
rect 516300 647123 516334 647137
rect 516300 647103 516334 647123
rect 516300 647055 516334 647065
rect 516300 647031 516334 647055
rect 516300 646987 516334 646993
rect 516300 646959 516334 646987
rect 516300 646919 516334 646921
rect 516300 646887 516334 646919
rect 516300 646817 516334 646849
rect 516300 646815 516334 646817
rect 516300 646749 516334 646777
rect 516300 646743 516334 646749
rect 516300 646681 516334 646705
rect 516300 646671 516334 646681
rect 516300 646613 516334 646633
rect 516300 646599 516334 646613
rect 516300 646545 516334 646561
rect 516300 646527 516334 646545
rect 516300 646477 516334 646489
rect 516300 646455 516334 646477
rect 516300 646409 516334 646417
rect 516300 646383 516334 646409
rect 516758 647327 516792 647353
rect 516758 647319 516792 647327
rect 516758 647259 516792 647281
rect 516758 647247 516792 647259
rect 516758 647191 516792 647209
rect 516758 647175 516792 647191
rect 516758 647123 516792 647137
rect 516758 647103 516792 647123
rect 516758 647055 516792 647065
rect 516758 647031 516792 647055
rect 516758 646987 516792 646993
rect 516758 646959 516792 646987
rect 516758 646919 516792 646921
rect 516758 646887 516792 646919
rect 516758 646817 516792 646849
rect 516758 646815 516792 646817
rect 516758 646749 516792 646777
rect 516758 646743 516792 646749
rect 516758 646681 516792 646705
rect 516758 646671 516792 646681
rect 516758 646613 516792 646633
rect 516758 646599 516792 646613
rect 516758 646545 516792 646561
rect 516758 646527 516792 646545
rect 516758 646477 516792 646489
rect 516758 646455 516792 646477
rect 516758 646409 516792 646417
rect 516758 646383 516792 646409
rect 517216 647327 517250 647353
rect 517216 647319 517250 647327
rect 517216 647259 517250 647281
rect 517216 647247 517250 647259
rect 517216 647191 517250 647209
rect 517216 647175 517250 647191
rect 517216 647123 517250 647137
rect 517216 647103 517250 647123
rect 517216 647055 517250 647065
rect 517216 647031 517250 647055
rect 517216 646987 517250 646993
rect 517216 646959 517250 646987
rect 517216 646919 517250 646921
rect 517216 646887 517250 646919
rect 517216 646817 517250 646849
rect 517216 646815 517250 646817
rect 517216 646749 517250 646777
rect 517216 646743 517250 646749
rect 517216 646681 517250 646705
rect 517216 646671 517250 646681
rect 517216 646613 517250 646633
rect 517216 646599 517250 646613
rect 517216 646545 517250 646561
rect 517216 646527 517250 646545
rect 517216 646477 517250 646489
rect 517216 646455 517250 646477
rect 517216 646409 517250 646417
rect 517216 646383 517250 646409
rect 517566 646459 518104 646709
<< metal1 >>
rect 513107 649794 513293 649842
rect 508019 649693 508440 649699
rect 508019 649443 508033 649693
rect 508427 649443 508440 649693
rect 508019 649437 508440 649443
rect 512478 649693 512899 649699
rect 512478 649443 512492 649693
rect 512886 649443 512899 649693
rect 512478 649437 512899 649443
rect 508150 649169 508310 649437
rect 508019 649163 508440 649169
rect 508019 648913 508033 649163
rect 508427 648913 508440 649163
rect 508019 648907 508440 648913
rect 512478 649163 512899 649169
rect 512478 648913 512492 649163
rect 512886 648913 512899 649163
rect 512478 648907 512899 648913
rect 512609 648639 512769 648907
rect 508017 648633 508438 648639
rect 508017 648383 508030 648633
rect 508424 648383 508438 648633
rect 508017 648377 508438 648383
rect 512476 648633 512897 648639
rect 512476 648383 512489 648633
rect 512883 648383 512897 648633
rect 512476 648377 512897 648383
rect 508147 648109 508307 648377
rect 508017 648103 508438 648109
rect 508017 647853 508030 648103
rect 508424 647853 508438 648103
rect 508017 647847 508438 647853
rect 512476 648103 512897 648109
rect 512476 647853 512489 648103
rect 512883 647853 512897 648103
rect 512476 647847 512897 647853
rect 512606 647579 512766 647847
rect 508017 647573 508438 647579
rect 508017 647323 508030 647573
rect 508424 647323 508438 647573
rect 508017 647317 508438 647323
rect 512476 647573 512897 647579
rect 512476 647323 512489 647573
rect 512883 647323 512897 647573
rect 512476 647317 512897 647323
rect 508147 647049 508307 647317
rect 508017 647043 508438 647049
rect 508017 646793 508030 647043
rect 508424 646793 508438 647043
rect 508017 646787 508438 646793
rect 512476 647043 512897 647049
rect 512476 646793 512489 647043
rect 512883 646793 512897 647043
rect 512476 646787 512897 646793
rect 512606 646519 512766 646787
rect 508017 646513 508438 646519
rect 508017 646263 508030 646513
rect 508424 646263 508438 646513
rect 508017 646257 508438 646263
rect 512476 646513 512897 646519
rect 512476 646263 512489 646513
rect 512883 646263 512897 646513
rect 512476 646257 512897 646263
rect 513107 646158 513142 649794
rect 513258 646158 513293 649794
rect 518182 649649 518288 649690
rect 518182 649597 518210 649649
rect 518262 649597 518288 649649
rect 518182 649585 518288 649597
rect 514303 649542 514349 649578
rect 514295 649536 514359 649542
rect 514295 649484 514301 649536
rect 514353 649484 514359 649536
rect 514295 649472 514359 649484
rect 514295 649420 514301 649472
rect 514353 649420 514359 649472
rect 514295 649414 514359 649420
rect 517361 649531 517407 649578
rect 517361 649497 517367 649531
rect 517401 649497 517407 649531
rect 517361 649459 517407 649497
rect 517361 649425 517367 649459
rect 517401 649425 517407 649459
rect 514303 649378 514349 649414
rect 516450 649349 516642 649355
rect 516450 649337 516456 649349
rect 514359 649331 516456 649337
rect 516508 649331 516520 649349
rect 516572 649331 516584 649349
rect 516636 649337 516642 649349
rect 517361 649337 517407 649425
rect 516636 649331 517407 649337
rect 514359 649297 514398 649331
rect 514432 649297 514470 649331
rect 514504 649297 514542 649331
rect 514576 649297 514614 649331
rect 514648 649297 514686 649331
rect 514720 649297 514758 649331
rect 514792 649297 514830 649331
rect 514864 649297 514902 649331
rect 514936 649297 514974 649331
rect 515008 649297 515046 649331
rect 515080 649297 515118 649331
rect 515152 649297 515190 649331
rect 515224 649297 515262 649331
rect 515296 649297 515334 649331
rect 515368 649297 515406 649331
rect 515440 649297 515478 649331
rect 515512 649297 515550 649331
rect 515584 649297 515622 649331
rect 515656 649297 515694 649331
rect 515728 649297 515766 649331
rect 515800 649297 515838 649331
rect 515872 649297 515910 649331
rect 515944 649297 515982 649331
rect 516016 649297 516054 649331
rect 516088 649297 516126 649331
rect 516160 649297 516198 649331
rect 516232 649297 516270 649331
rect 516304 649297 516342 649331
rect 516376 649297 516414 649331
rect 516448 649297 516456 649331
rect 516664 649297 516702 649331
rect 516736 649297 516774 649331
rect 516808 649297 516846 649331
rect 516880 649297 516918 649331
rect 516952 649297 516990 649331
rect 517024 649297 517062 649331
rect 517096 649297 517134 649331
rect 517168 649297 517206 649331
rect 517240 649297 517278 649331
rect 517312 649297 517407 649331
rect 514359 649291 517407 649297
rect 518182 649533 518210 649585
rect 518262 649533 518288 649585
rect 518182 649521 518288 649533
rect 518182 649469 518210 649521
rect 518262 649469 518288 649521
rect 513657 649198 513703 649213
rect 513657 649164 513663 649198
rect 513697 649164 513703 649198
rect 513657 649126 513703 649164
rect 513657 649092 513663 649126
rect 513697 649092 513703 649126
rect 513657 649054 513703 649092
rect 514115 649198 514161 649213
rect 514115 649164 514121 649198
rect 514155 649164 514161 649198
rect 514115 649126 514161 649164
rect 514115 649092 514121 649126
rect 514155 649092 514161 649126
rect 514115 649091 514161 649092
rect 514573 649198 514619 649213
rect 514573 649164 514579 649198
rect 514613 649164 514619 649198
rect 514573 649126 514619 649164
rect 514573 649092 514579 649126
rect 514613 649092 514619 649126
rect 513657 649020 513663 649054
rect 513697 649020 513703 649054
rect 513657 648982 513703 649020
rect 513657 648948 513663 648982
rect 513697 648948 513703 648982
rect 513657 648910 513703 648948
rect 513657 648876 513663 648910
rect 513697 648876 513703 648910
rect 513657 648838 513703 648876
rect 513657 648804 513663 648838
rect 513697 648804 513703 648838
rect 514106 649085 514170 649091
rect 514106 649033 514112 649085
rect 514164 649033 514170 649085
rect 514106 649021 514121 649033
rect 514155 649021 514170 649033
rect 514106 648969 514112 649021
rect 514164 648969 514170 649021
rect 514106 648957 514121 648969
rect 514155 648957 514170 648969
rect 514106 648905 514112 648957
rect 514164 648905 514170 648957
rect 514106 648893 514121 648905
rect 514155 648893 514170 648905
rect 514106 648841 514112 648893
rect 514164 648841 514170 648893
rect 514106 648838 514170 648841
rect 514106 648835 514121 648838
rect 513657 648766 513703 648804
rect 513657 648732 513663 648766
rect 513697 648732 513703 648766
rect 513657 648694 513703 648732
rect 513657 648660 513663 648694
rect 513697 648660 513703 648694
rect 513657 648622 513703 648660
rect 513657 648597 513663 648622
rect 513648 648591 513663 648597
rect 513697 648597 513703 648622
rect 514115 648804 514121 648835
rect 514155 648835 514170 648838
rect 514573 649054 514619 649092
rect 515031 649198 515077 649213
rect 515031 649164 515037 649198
rect 515071 649164 515077 649198
rect 515031 649126 515077 649164
rect 515031 649092 515037 649126
rect 515071 649092 515077 649126
rect 515031 649091 515077 649092
rect 515489 649198 515535 649213
rect 515489 649164 515495 649198
rect 515529 649164 515535 649198
rect 515489 649126 515535 649164
rect 515489 649092 515495 649126
rect 515529 649092 515535 649126
rect 514573 649020 514579 649054
rect 514613 649020 514619 649054
rect 514573 648982 514619 649020
rect 514573 648948 514579 648982
rect 514613 648948 514619 648982
rect 514573 648910 514619 648948
rect 514573 648876 514579 648910
rect 514613 648876 514619 648910
rect 514573 648838 514619 648876
rect 514155 648804 514161 648835
rect 514115 648766 514161 648804
rect 514115 648732 514121 648766
rect 514155 648732 514161 648766
rect 514115 648694 514161 648732
rect 514115 648660 514121 648694
rect 514155 648660 514161 648694
rect 514115 648622 514161 648660
rect 513697 648591 513712 648597
rect 513648 648539 513654 648591
rect 513706 648539 513712 648591
rect 513648 648527 513663 648539
rect 513697 648527 513712 648539
rect 513648 648475 513654 648527
rect 513706 648475 513712 648527
rect 513648 648463 513663 648475
rect 513697 648463 513712 648475
rect 513648 648411 513654 648463
rect 513706 648411 513712 648463
rect 513648 648406 513712 648411
rect 513648 648399 513663 648406
rect 513697 648399 513712 648406
rect 513648 648347 513654 648399
rect 513706 648347 513712 648399
rect 513648 648341 513712 648347
rect 514115 648588 514121 648622
rect 514155 648588 514161 648622
rect 514573 648804 514579 648838
rect 514613 648804 514619 648838
rect 515022 649085 515086 649091
rect 515022 649033 515028 649085
rect 515080 649033 515086 649085
rect 515022 649021 515037 649033
rect 515071 649021 515086 649033
rect 515022 648969 515028 649021
rect 515080 648969 515086 649021
rect 515022 648957 515037 648969
rect 515071 648957 515086 648969
rect 515022 648905 515028 648957
rect 515080 648905 515086 648957
rect 515022 648893 515037 648905
rect 515071 648893 515086 648905
rect 515022 648841 515028 648893
rect 515080 648841 515086 648893
rect 515022 648838 515086 648841
rect 515022 648835 515037 648838
rect 514573 648766 514619 648804
rect 514573 648732 514579 648766
rect 514613 648732 514619 648766
rect 514573 648694 514619 648732
rect 514573 648660 514579 648694
rect 514613 648660 514619 648694
rect 514573 648622 514619 648660
rect 514573 648597 514579 648622
rect 514115 648550 514161 648588
rect 514115 648516 514121 648550
rect 514155 648516 514161 648550
rect 514115 648478 514161 648516
rect 514115 648444 514121 648478
rect 514155 648444 514161 648478
rect 514115 648406 514161 648444
rect 514115 648372 514121 648406
rect 514155 648372 514161 648406
rect 513657 648334 513703 648341
rect 513657 648300 513663 648334
rect 513697 648300 513703 648334
rect 513657 648262 513703 648300
rect 513657 648228 513663 648262
rect 513697 648228 513703 648262
rect 513657 648213 513703 648228
rect 514115 648334 514161 648372
rect 514564 648591 514579 648597
rect 514613 648597 514619 648622
rect 515031 648804 515037 648835
rect 515071 648835 515086 648838
rect 515489 649054 515535 649092
rect 515607 649198 515653 649213
rect 515607 649164 515613 649198
rect 515647 649164 515653 649198
rect 515607 649126 515653 649164
rect 515607 649092 515613 649126
rect 515647 649092 515653 649126
rect 515607 649091 515653 649092
rect 516065 649198 516111 649213
rect 516065 649164 516071 649198
rect 516105 649164 516111 649198
rect 516065 649126 516111 649164
rect 516065 649092 516071 649126
rect 516105 649092 516111 649126
rect 515489 649020 515495 649054
rect 515529 649020 515535 649054
rect 515489 648982 515535 649020
rect 515489 648948 515495 648982
rect 515529 648948 515535 648982
rect 515489 648910 515535 648948
rect 515489 648876 515495 648910
rect 515529 648876 515535 648910
rect 515489 648838 515535 648876
rect 515071 648804 515077 648835
rect 515031 648766 515077 648804
rect 515031 648732 515037 648766
rect 515071 648732 515077 648766
rect 515031 648694 515077 648732
rect 515031 648660 515037 648694
rect 515071 648660 515077 648694
rect 515031 648622 515077 648660
rect 514613 648591 514628 648597
rect 514564 648539 514570 648591
rect 514622 648539 514628 648591
rect 514564 648527 514579 648539
rect 514613 648527 514628 648539
rect 514564 648475 514570 648527
rect 514622 648475 514628 648527
rect 514564 648463 514579 648475
rect 514613 648463 514628 648475
rect 514564 648411 514570 648463
rect 514622 648411 514628 648463
rect 514564 648406 514628 648411
rect 514564 648399 514579 648406
rect 514613 648399 514628 648406
rect 514564 648347 514570 648399
rect 514622 648347 514628 648399
rect 514564 648341 514628 648347
rect 515031 648588 515037 648622
rect 515071 648588 515077 648622
rect 515489 648804 515495 648838
rect 515529 648804 515535 648838
rect 515598 649085 515662 649091
rect 515598 649033 515604 649085
rect 515656 649033 515662 649085
rect 515598 649021 515613 649033
rect 515647 649021 515662 649033
rect 515598 648969 515604 649021
rect 515656 648969 515662 649021
rect 515598 648957 515613 648969
rect 515647 648957 515662 648969
rect 515598 648905 515604 648957
rect 515656 648905 515662 648957
rect 515598 648893 515613 648905
rect 515647 648893 515662 648905
rect 515598 648841 515604 648893
rect 515656 648841 515662 648893
rect 515598 648838 515662 648841
rect 515598 648835 515613 648838
rect 515489 648766 515535 648804
rect 515489 648732 515495 648766
rect 515529 648732 515535 648766
rect 515489 648694 515535 648732
rect 515489 648660 515495 648694
rect 515529 648660 515535 648694
rect 515489 648622 515535 648660
rect 515489 648597 515495 648622
rect 515031 648550 515077 648588
rect 515031 648516 515037 648550
rect 515071 648516 515077 648550
rect 515031 648478 515077 648516
rect 515031 648444 515037 648478
rect 515071 648444 515077 648478
rect 515031 648406 515077 648444
rect 515031 648372 515037 648406
rect 515071 648372 515077 648406
rect 514115 648300 514121 648334
rect 514155 648300 514161 648334
rect 514115 648262 514161 648300
rect 514115 648228 514121 648262
rect 514155 648228 514161 648262
rect 514115 648213 514161 648228
rect 514573 648334 514619 648341
rect 514573 648300 514579 648334
rect 514613 648300 514619 648334
rect 514573 648262 514619 648300
rect 514573 648228 514579 648262
rect 514613 648228 514619 648262
rect 514573 648213 514619 648228
rect 515031 648334 515077 648372
rect 515480 648591 515495 648597
rect 515529 648597 515535 648622
rect 515607 648804 515613 648835
rect 515647 648835 515662 648838
rect 516065 649054 516111 649092
rect 516523 649198 516569 649213
rect 516523 649164 516529 649198
rect 516563 649164 516569 649198
rect 516523 649126 516569 649164
rect 516523 649092 516529 649126
rect 516563 649092 516569 649126
rect 516523 649091 516569 649092
rect 516981 649198 517027 649213
rect 516981 649164 516987 649198
rect 517021 649164 517027 649198
rect 516981 649126 517027 649164
rect 516981 649092 516987 649126
rect 517021 649092 517027 649126
rect 516065 649020 516071 649054
rect 516105 649020 516111 649054
rect 516065 648982 516111 649020
rect 516065 648948 516071 648982
rect 516105 648948 516111 648982
rect 516065 648910 516111 648948
rect 516065 648876 516071 648910
rect 516105 648876 516111 648910
rect 516065 648838 516111 648876
rect 515647 648804 515653 648835
rect 515607 648766 515653 648804
rect 515607 648732 515613 648766
rect 515647 648732 515653 648766
rect 515607 648694 515653 648732
rect 515607 648660 515613 648694
rect 515647 648660 515653 648694
rect 515607 648622 515653 648660
rect 515529 648591 515544 648597
rect 515480 648539 515486 648591
rect 515538 648539 515544 648591
rect 515480 648527 515495 648539
rect 515529 648527 515544 648539
rect 515480 648475 515486 648527
rect 515538 648475 515544 648527
rect 515480 648463 515495 648475
rect 515529 648463 515544 648475
rect 515480 648411 515486 648463
rect 515538 648411 515544 648463
rect 515480 648406 515544 648411
rect 515480 648399 515495 648406
rect 515529 648399 515544 648406
rect 515480 648347 515486 648399
rect 515538 648347 515544 648399
rect 515480 648341 515544 648347
rect 515607 648588 515613 648622
rect 515647 648588 515653 648622
rect 516065 648804 516071 648838
rect 516105 648804 516111 648838
rect 516514 649085 516578 649091
rect 516514 649033 516520 649085
rect 516572 649033 516578 649085
rect 516514 649021 516529 649033
rect 516563 649021 516578 649033
rect 516514 648969 516520 649021
rect 516572 648969 516578 649021
rect 516514 648957 516529 648969
rect 516563 648957 516578 648969
rect 516514 648905 516520 648957
rect 516572 648905 516578 648957
rect 516514 648893 516529 648905
rect 516563 648893 516578 648905
rect 516514 648841 516520 648893
rect 516572 648841 516578 648893
rect 516514 648838 516578 648841
rect 516514 648835 516529 648838
rect 516065 648766 516111 648804
rect 516065 648732 516071 648766
rect 516105 648732 516111 648766
rect 516065 648694 516111 648732
rect 516065 648660 516071 648694
rect 516105 648660 516111 648694
rect 516065 648622 516111 648660
rect 516065 648597 516071 648622
rect 515607 648550 515653 648588
rect 515607 648516 515613 648550
rect 515647 648516 515653 648550
rect 515607 648478 515653 648516
rect 515607 648444 515613 648478
rect 515647 648444 515653 648478
rect 515607 648406 515653 648444
rect 515607 648372 515613 648406
rect 515647 648372 515653 648406
rect 515031 648300 515037 648334
rect 515071 648300 515077 648334
rect 515031 648262 515077 648300
rect 515031 648228 515037 648262
rect 515071 648228 515077 648262
rect 515031 648213 515077 648228
rect 515489 648334 515535 648341
rect 515489 648300 515495 648334
rect 515529 648300 515535 648334
rect 515489 648262 515535 648300
rect 515489 648228 515495 648262
rect 515529 648228 515535 648262
rect 515489 648213 515535 648228
rect 515607 648334 515653 648372
rect 516056 648591 516071 648597
rect 516105 648597 516111 648622
rect 516523 648804 516529 648835
rect 516563 648835 516578 648838
rect 516981 649054 517027 649092
rect 517439 649198 517485 649213
rect 517439 649164 517445 649198
rect 517479 649164 517485 649198
rect 517439 649126 517485 649164
rect 517439 649092 517445 649126
rect 517479 649092 517485 649126
rect 517439 649091 517485 649092
rect 517557 649198 517603 649213
rect 517557 649164 517563 649198
rect 517597 649164 517603 649198
rect 517557 649126 517603 649164
rect 517557 649092 517563 649126
rect 517597 649092 517603 649126
rect 516981 649020 516987 649054
rect 517021 649020 517027 649054
rect 516981 648982 517027 649020
rect 516981 648948 516987 648982
rect 517021 648948 517027 648982
rect 516981 648910 517027 648948
rect 516981 648876 516987 648910
rect 517021 648876 517027 648910
rect 516981 648838 517027 648876
rect 516563 648804 516569 648835
rect 516523 648766 516569 648804
rect 516523 648732 516529 648766
rect 516563 648732 516569 648766
rect 516523 648694 516569 648732
rect 516523 648660 516529 648694
rect 516563 648660 516569 648694
rect 516523 648622 516569 648660
rect 516105 648591 516120 648597
rect 516056 648539 516062 648591
rect 516114 648539 516120 648591
rect 516056 648527 516071 648539
rect 516105 648527 516120 648539
rect 516056 648475 516062 648527
rect 516114 648475 516120 648527
rect 516056 648463 516071 648475
rect 516105 648463 516120 648475
rect 516056 648411 516062 648463
rect 516114 648411 516120 648463
rect 516056 648406 516120 648411
rect 516056 648399 516071 648406
rect 516105 648399 516120 648406
rect 516056 648347 516062 648399
rect 516114 648347 516120 648399
rect 516056 648341 516120 648347
rect 516523 648588 516529 648622
rect 516563 648588 516569 648622
rect 516981 648804 516987 648838
rect 517021 648804 517027 648838
rect 517430 649085 517494 649091
rect 517430 649033 517436 649085
rect 517488 649033 517494 649085
rect 517430 649021 517445 649033
rect 517479 649021 517494 649033
rect 517430 648969 517436 649021
rect 517488 648969 517494 649021
rect 517430 648957 517445 648969
rect 517479 648957 517494 648969
rect 517430 648905 517436 648957
rect 517488 648905 517494 648957
rect 517430 648893 517445 648905
rect 517479 648893 517494 648905
rect 517430 648841 517436 648893
rect 517488 648841 517494 648893
rect 517430 648838 517494 648841
rect 517430 648835 517445 648838
rect 516981 648766 517027 648804
rect 516981 648732 516987 648766
rect 517021 648732 517027 648766
rect 516981 648694 517027 648732
rect 516981 648660 516987 648694
rect 517021 648660 517027 648694
rect 516981 648622 517027 648660
rect 516981 648597 516987 648622
rect 516523 648550 516569 648588
rect 516523 648516 516529 648550
rect 516563 648516 516569 648550
rect 516523 648478 516569 648516
rect 516523 648444 516529 648478
rect 516563 648444 516569 648478
rect 516523 648406 516569 648444
rect 516523 648372 516529 648406
rect 516563 648372 516569 648406
rect 515607 648300 515613 648334
rect 515647 648300 515653 648334
rect 515607 648262 515653 648300
rect 515607 648228 515613 648262
rect 515647 648228 515653 648262
rect 515607 648213 515653 648228
rect 516065 648334 516111 648341
rect 516065 648300 516071 648334
rect 516105 648300 516111 648334
rect 516065 648262 516111 648300
rect 516065 648228 516071 648262
rect 516105 648228 516111 648262
rect 516065 648213 516111 648228
rect 516523 648334 516569 648372
rect 516972 648591 516987 648597
rect 517021 648597 517027 648622
rect 517439 648804 517445 648835
rect 517479 648835 517494 648838
rect 517557 649054 517603 649092
rect 518015 649198 518061 649213
rect 518015 649164 518021 649198
rect 518055 649164 518061 649198
rect 518015 649126 518061 649164
rect 518015 649092 518021 649126
rect 518055 649092 518061 649126
rect 518015 649091 518061 649092
rect 517557 649020 517563 649054
rect 517597 649020 517603 649054
rect 517557 648982 517603 649020
rect 517557 648948 517563 648982
rect 517597 648948 517603 648982
rect 517557 648910 517603 648948
rect 517557 648876 517563 648910
rect 517597 648876 517603 648910
rect 517557 648838 517603 648876
rect 517479 648804 517485 648835
rect 517439 648766 517485 648804
rect 517439 648732 517445 648766
rect 517479 648732 517485 648766
rect 517439 648694 517485 648732
rect 517439 648660 517445 648694
rect 517479 648660 517485 648694
rect 517439 648622 517485 648660
rect 517021 648591 517036 648597
rect 516972 648539 516978 648591
rect 517030 648539 517036 648591
rect 516972 648527 516987 648539
rect 517021 648527 517036 648539
rect 516972 648475 516978 648527
rect 517030 648475 517036 648527
rect 516972 648463 516987 648475
rect 517021 648463 517036 648475
rect 516972 648411 516978 648463
rect 517030 648411 517036 648463
rect 516972 648406 517036 648411
rect 516972 648399 516987 648406
rect 517021 648399 517036 648406
rect 516972 648347 516978 648399
rect 517030 648347 517036 648399
rect 516972 648341 517036 648347
rect 517439 648588 517445 648622
rect 517479 648588 517485 648622
rect 517557 648804 517563 648838
rect 517597 648804 517603 648838
rect 518006 649085 518070 649091
rect 518006 649033 518012 649085
rect 518064 649033 518070 649085
rect 518006 649021 518021 649033
rect 518055 649021 518070 649033
rect 518006 648969 518012 649021
rect 518064 648969 518070 649021
rect 518006 648957 518021 648969
rect 518055 648957 518070 648969
rect 518006 648905 518012 648957
rect 518064 648905 518070 648957
rect 518006 648893 518021 648905
rect 518055 648893 518070 648905
rect 518006 648841 518012 648893
rect 518064 648841 518070 648893
rect 518006 648838 518070 648841
rect 518006 648835 518021 648838
rect 517557 648766 517603 648804
rect 517557 648732 517563 648766
rect 517597 648732 517603 648766
rect 517557 648694 517603 648732
rect 517557 648660 517563 648694
rect 517597 648660 517603 648694
rect 517557 648622 517603 648660
rect 517557 648597 517563 648622
rect 517439 648550 517485 648588
rect 517439 648516 517445 648550
rect 517479 648516 517485 648550
rect 517439 648478 517485 648516
rect 517439 648444 517445 648478
rect 517479 648444 517485 648478
rect 517439 648406 517485 648444
rect 517439 648372 517445 648406
rect 517479 648372 517485 648406
rect 516523 648300 516529 648334
rect 516563 648300 516569 648334
rect 516523 648262 516569 648300
rect 516523 648228 516529 648262
rect 516563 648228 516569 648262
rect 516523 648213 516569 648228
rect 516981 648334 517027 648341
rect 516981 648300 516987 648334
rect 517021 648300 517027 648334
rect 516981 648262 517027 648300
rect 516981 648228 516987 648262
rect 517021 648228 517027 648262
rect 516981 648213 517027 648228
rect 517439 648334 517485 648372
rect 517548 648591 517563 648597
rect 517597 648597 517603 648622
rect 518015 648804 518021 648835
rect 518055 648835 518070 648838
rect 518182 649088 518288 649469
rect 518182 649085 518218 649088
rect 518252 649085 518288 649088
rect 518182 649033 518209 649085
rect 518261 649033 518288 649085
rect 518182 649021 518288 649033
rect 518182 648969 518209 649021
rect 518261 648969 518288 649021
rect 518182 648957 518288 648969
rect 518182 648905 518209 648957
rect 518261 648905 518288 648957
rect 518182 648893 518288 648905
rect 518182 648841 518209 648893
rect 518261 648841 518288 648893
rect 518182 648838 518218 648841
rect 518252 648838 518288 648841
rect 518055 648804 518061 648835
rect 518182 648825 518288 648838
rect 518015 648766 518061 648804
rect 518015 648732 518021 648766
rect 518055 648732 518061 648766
rect 518015 648694 518061 648732
rect 518015 648660 518021 648694
rect 518055 648660 518061 648694
rect 518015 648622 518061 648660
rect 517597 648591 517612 648597
rect 517548 648539 517554 648591
rect 517606 648539 517612 648591
rect 517548 648527 517563 648539
rect 517597 648527 517612 648539
rect 517548 648475 517554 648527
rect 517606 648475 517612 648527
rect 517548 648463 517563 648475
rect 517597 648463 517612 648475
rect 517548 648411 517554 648463
rect 517606 648411 517612 648463
rect 517548 648406 517612 648411
rect 517548 648399 517563 648406
rect 517597 648399 517612 648406
rect 517548 648347 517554 648399
rect 517606 648347 517612 648399
rect 517548 648341 517612 648347
rect 518015 648588 518021 648622
rect 518055 648588 518061 648622
rect 518015 648550 518061 648588
rect 518015 648516 518021 648550
rect 518055 648516 518061 648550
rect 518015 648478 518061 648516
rect 518015 648444 518021 648478
rect 518055 648444 518061 648478
rect 518015 648406 518061 648444
rect 518015 648372 518021 648406
rect 518055 648372 518061 648406
rect 517439 648300 517445 648334
rect 517479 648300 517485 648334
rect 517439 648262 517485 648300
rect 517439 648228 517445 648262
rect 517479 648228 517485 648262
rect 517439 648213 517485 648228
rect 517557 648334 517603 648341
rect 517557 648300 517563 648334
rect 517597 648300 517603 648334
rect 517557 648262 517603 648300
rect 517557 648228 517563 648262
rect 517597 648228 517603 648262
rect 517557 648213 517603 648228
rect 518015 648334 518061 648372
rect 518015 648300 518021 648334
rect 518055 648300 518061 648334
rect 518015 648262 518061 648300
rect 518015 648228 518021 648262
rect 518055 648228 518061 648262
rect 518015 648213 518061 648228
rect 513713 648166 515479 648172
rect 513713 648132 513748 648166
rect 513782 648132 513820 648166
rect 513854 648132 513892 648166
rect 513926 648132 513964 648166
rect 513998 648132 514036 648166
rect 514070 648132 514206 648166
rect 514240 648132 514278 648166
rect 514312 648132 514350 648166
rect 514384 648132 514422 648166
rect 514456 648132 514474 648166
rect 514528 648132 514538 648166
rect 513713 648126 514474 648132
rect 514468 648114 514474 648126
rect 514526 648114 514538 648132
rect 514590 648114 514602 648166
rect 514654 648132 514664 648166
rect 514718 648132 514736 648166
rect 514770 648132 514808 648166
rect 514842 648132 514880 648166
rect 514914 648132 514952 648166
rect 514986 648132 515122 648166
rect 515156 648132 515194 648166
rect 515228 648132 515266 648166
rect 515300 648132 515338 648166
rect 515372 648132 515410 648166
rect 515444 648132 515479 648166
rect 514654 648114 514666 648132
rect 514718 648126 515479 648132
rect 515663 648166 517429 648172
rect 514718 648114 514724 648126
rect 514468 648108 514724 648114
rect 515663 648114 515669 648166
rect 515732 648132 515733 648166
rect 515876 648132 515914 648166
rect 515948 648132 515986 648166
rect 516020 648132 516156 648166
rect 516190 648132 516228 648166
rect 516262 648132 516300 648166
rect 516334 648132 516372 648166
rect 516406 648132 516444 648166
rect 516478 648132 516614 648166
rect 516648 648132 516686 648166
rect 516720 648132 516758 648166
rect 516792 648132 516830 648166
rect 516864 648132 516902 648166
rect 516936 648132 517072 648166
rect 517106 648132 517144 648166
rect 517178 648132 517216 648166
rect 517250 648132 517288 648166
rect 517322 648132 517360 648166
rect 517394 648132 517429 648166
rect 515721 648114 515733 648132
rect 515785 648114 515797 648132
rect 515849 648126 517429 648132
rect 517613 648166 518005 648172
rect 517613 648132 517648 648166
rect 517682 648132 517719 648166
rect 517613 648126 517719 648132
rect 515849 648114 515855 648126
rect 515663 648108 515855 648114
rect 517713 648114 517719 648126
rect 517771 648114 517783 648166
rect 517835 648114 517847 648166
rect 517899 648132 517936 648166
rect 517970 648132 518005 648166
rect 517899 648126 518005 648132
rect 517899 648114 517905 648126
rect 517713 648108 517905 648114
rect 515076 647458 515268 647464
rect 515076 647446 515082 647458
rect 514462 647440 514910 647446
rect 514462 647406 514553 647440
rect 514587 647406 514625 647440
rect 514659 647406 514697 647440
rect 514731 647406 514769 647440
rect 514803 647406 514841 647440
rect 514875 647406 514910 647440
rect 514462 647400 514910 647406
rect 514976 647440 515082 647446
rect 514976 647406 515011 647440
rect 515045 647406 515082 647440
rect 515134 647406 515146 647458
rect 515198 647406 515210 647458
rect 515262 647446 515268 647458
rect 515534 647458 515726 647464
rect 515534 647446 515540 647458
rect 515262 647440 515368 647446
rect 515262 647406 515299 647440
rect 515333 647406 515368 647440
rect 514976 647400 515368 647406
rect 515434 647440 515540 647446
rect 515434 647406 515469 647440
rect 515503 647406 515540 647440
rect 515592 647406 515604 647458
rect 515656 647406 515668 647458
rect 515720 647446 515726 647458
rect 516450 647458 516642 647464
rect 516450 647446 516456 647458
rect 515720 647440 515826 647446
rect 515720 647406 515757 647440
rect 515791 647406 515826 647440
rect 515434 647400 515826 647406
rect 515892 647440 516284 647446
rect 515892 647406 515927 647440
rect 515961 647406 515999 647440
rect 516033 647406 516071 647440
rect 516105 647406 516143 647440
rect 516177 647406 516215 647440
rect 516249 647406 516284 647440
rect 515892 647400 516284 647406
rect 516350 647440 516456 647446
rect 516350 647406 516385 647440
rect 516419 647406 516456 647440
rect 516508 647406 516520 647458
rect 516572 647406 516584 647458
rect 516636 647446 516642 647458
rect 516636 647440 516742 647446
rect 516636 647406 516673 647440
rect 516707 647406 516742 647440
rect 516350 647400 516742 647406
rect 516808 647440 517256 647446
rect 516808 647406 516843 647440
rect 516877 647406 516915 647440
rect 516949 647406 516987 647440
rect 517021 647406 517059 647440
rect 517093 647406 517131 647440
rect 517165 647406 517256 647440
rect 516808 647400 517256 647406
rect 514462 647353 514508 647400
rect 514976 647368 515022 647400
rect 516238 647368 516284 647400
rect 514462 647319 514468 647353
rect 514502 647319 514508 647353
rect 514462 647281 514508 647319
rect 514462 647247 514468 647281
rect 514502 647247 514508 647281
rect 514462 647209 514508 647247
rect 514920 647353 515022 647368
rect 514920 647319 514926 647353
rect 514960 647322 515022 647353
rect 515378 647353 515424 647368
rect 514960 647319 514966 647322
rect 514920 647281 514966 647319
rect 514920 647247 514926 647281
rect 514960 647247 514966 647281
rect 514920 647236 514966 647247
rect 515378 647319 515384 647353
rect 515418 647319 515424 647353
rect 515378 647281 515424 647319
rect 515378 647247 515384 647281
rect 515418 647247 515424 647281
rect 514462 647175 514468 647209
rect 514502 647175 514508 647209
rect 514462 647137 514508 647175
rect 514462 647103 514468 647137
rect 514502 647103 514508 647137
rect 514462 647065 514508 647103
rect 514462 647031 514468 647065
rect 514502 647031 514508 647065
rect 514462 646993 514508 647031
rect 514462 646959 514468 646993
rect 514502 646959 514508 646993
rect 514911 647230 514975 647236
rect 514911 647178 514917 647230
rect 514969 647178 514975 647230
rect 514911 647175 514926 647178
rect 514960 647175 514975 647178
rect 514911 647166 514975 647175
rect 514911 647114 514917 647166
rect 514969 647114 514975 647166
rect 514911 647103 514926 647114
rect 514960 647103 514975 647114
rect 514911 647102 514975 647103
rect 514911 647050 514917 647102
rect 514969 647050 514975 647102
rect 514911 647038 514926 647050
rect 514960 647038 514975 647050
rect 514911 646986 514917 647038
rect 514969 646986 514975 647038
rect 514911 646980 514926 646986
rect 514462 646921 514508 646959
rect 514462 646887 514468 646921
rect 514502 646887 514508 646921
rect 514462 646849 514508 646887
rect 514462 646815 514468 646849
rect 514502 646815 514508 646849
rect 514462 646777 514508 646815
rect 514462 646743 514468 646777
rect 514502 646743 514508 646777
rect 513598 646709 514160 646721
rect 514462 646712 514508 646743
rect 514920 646959 514926 646980
rect 514960 646980 514975 646986
rect 515378 647209 515424 647247
rect 515836 647353 515882 647368
rect 515836 647319 515842 647353
rect 515876 647319 515882 647353
rect 516238 647353 516340 647368
rect 516238 647322 516300 647353
rect 515836 647281 515882 647319
rect 515836 647247 515842 647281
rect 515876 647247 515882 647281
rect 515836 647236 515882 647247
rect 516294 647319 516300 647322
rect 516334 647319 516340 647353
rect 516294 647281 516340 647319
rect 516294 647247 516300 647281
rect 516334 647247 516340 647281
rect 515378 647175 515384 647209
rect 515418 647175 515424 647209
rect 515378 647137 515424 647175
rect 515378 647103 515384 647137
rect 515418 647103 515424 647137
rect 515378 647065 515424 647103
rect 515378 647031 515384 647065
rect 515418 647031 515424 647065
rect 515378 646993 515424 647031
rect 514960 646959 514966 646980
rect 514920 646921 514966 646959
rect 514920 646887 514926 646921
rect 514960 646887 514966 646921
rect 514920 646849 514966 646887
rect 514920 646815 514926 646849
rect 514960 646815 514966 646849
rect 514920 646777 514966 646815
rect 514920 646743 514926 646777
rect 514960 646743 514966 646777
rect 513598 646459 513610 646709
rect 514148 646459 514160 646709
rect 513598 646447 514160 646459
rect 514453 646706 514517 646712
rect 514453 646654 514459 646706
rect 514511 646654 514517 646706
rect 514453 646642 514517 646654
rect 514453 646590 514459 646642
rect 514511 646590 514517 646642
rect 514453 646578 514517 646590
rect 514453 646526 514459 646578
rect 514511 646526 514517 646578
rect 514453 646514 514517 646526
rect 514453 646462 514459 646514
rect 514511 646462 514517 646514
rect 514453 646456 514468 646462
rect 514462 646455 514468 646456
rect 514502 646456 514517 646462
rect 514920 646705 514966 646743
rect 515378 646959 515384 646993
rect 515418 646959 515424 646993
rect 515827 647230 515891 647236
rect 515827 647178 515833 647230
rect 515885 647178 515891 647230
rect 515827 647175 515842 647178
rect 515876 647175 515891 647178
rect 515827 647166 515891 647175
rect 515827 647114 515833 647166
rect 515885 647114 515891 647166
rect 515827 647103 515842 647114
rect 515876 647103 515891 647114
rect 515827 647102 515891 647103
rect 515827 647050 515833 647102
rect 515885 647050 515891 647102
rect 515827 647038 515842 647050
rect 515876 647038 515891 647050
rect 515827 646986 515833 647038
rect 515885 646986 515891 647038
rect 515827 646980 515842 646986
rect 515378 646921 515424 646959
rect 515378 646887 515384 646921
rect 515418 646887 515424 646921
rect 515378 646849 515424 646887
rect 515378 646815 515384 646849
rect 515418 646815 515424 646849
rect 515378 646777 515424 646815
rect 515378 646743 515384 646777
rect 515418 646743 515424 646777
rect 515378 646712 515424 646743
rect 515836 646959 515842 646980
rect 515876 646980 515891 646986
rect 516294 647209 516340 647247
rect 516752 647353 516798 647368
rect 516752 647319 516758 647353
rect 516792 647319 516798 647353
rect 516752 647281 516798 647319
rect 516752 647247 516758 647281
rect 516792 647247 516798 647281
rect 516752 647236 516798 647247
rect 517210 647353 517256 647400
rect 517210 647319 517216 647353
rect 517250 647319 517256 647353
rect 517210 647281 517256 647319
rect 517210 647247 517216 647281
rect 517250 647247 517256 647281
rect 516294 647175 516300 647209
rect 516334 647175 516340 647209
rect 516294 647137 516340 647175
rect 516294 647103 516300 647137
rect 516334 647103 516340 647137
rect 516294 647065 516340 647103
rect 516294 647031 516300 647065
rect 516334 647031 516340 647065
rect 516294 646993 516340 647031
rect 515876 646959 515882 646980
rect 515836 646921 515882 646959
rect 515836 646887 515842 646921
rect 515876 646887 515882 646921
rect 515836 646849 515882 646887
rect 515836 646815 515842 646849
rect 515876 646815 515882 646849
rect 515836 646777 515882 646815
rect 515836 646743 515842 646777
rect 515876 646743 515882 646777
rect 514920 646671 514926 646705
rect 514960 646671 514966 646705
rect 514920 646633 514966 646671
rect 514920 646599 514926 646633
rect 514960 646599 514966 646633
rect 514920 646561 514966 646599
rect 514920 646527 514926 646561
rect 514960 646527 514966 646561
rect 514920 646489 514966 646527
rect 514502 646455 514508 646456
rect 514462 646417 514508 646455
rect 514462 646383 514468 646417
rect 514502 646383 514508 646417
rect 514462 646368 514508 646383
rect 514920 646455 514926 646489
rect 514960 646455 514966 646489
rect 515369 646706 515433 646712
rect 515369 646654 515375 646706
rect 515427 646654 515433 646706
rect 515369 646642 515433 646654
rect 515369 646590 515375 646642
rect 515427 646590 515433 646642
rect 515369 646578 515433 646590
rect 515369 646526 515375 646578
rect 515427 646526 515433 646578
rect 515369 646514 515433 646526
rect 515369 646462 515375 646514
rect 515427 646462 515433 646514
rect 515369 646456 515384 646462
rect 514920 646417 514966 646455
rect 514920 646383 514926 646417
rect 514960 646383 514966 646417
rect 514920 646368 514966 646383
rect 515378 646455 515384 646456
rect 515418 646456 515433 646462
rect 515836 646705 515882 646743
rect 516294 646959 516300 646993
rect 516334 646959 516340 646993
rect 516743 647230 516807 647236
rect 516743 647178 516749 647230
rect 516801 647178 516807 647230
rect 516743 647175 516758 647178
rect 516792 647175 516807 647178
rect 516743 647166 516807 647175
rect 516743 647114 516749 647166
rect 516801 647114 516807 647166
rect 516743 647103 516758 647114
rect 516792 647103 516807 647114
rect 516743 647102 516807 647103
rect 516743 647050 516749 647102
rect 516801 647050 516807 647102
rect 516743 647038 516758 647050
rect 516792 647038 516807 647050
rect 516743 646986 516749 647038
rect 516801 646986 516807 647038
rect 516743 646980 516758 646986
rect 516294 646921 516340 646959
rect 516294 646887 516300 646921
rect 516334 646887 516340 646921
rect 516294 646849 516340 646887
rect 516294 646815 516300 646849
rect 516334 646815 516340 646849
rect 516294 646777 516340 646815
rect 516294 646743 516300 646777
rect 516334 646743 516340 646777
rect 516294 646712 516340 646743
rect 516752 646959 516758 646980
rect 516792 646980 516807 646986
rect 517210 647209 517256 647247
rect 517210 647175 517216 647209
rect 517250 647175 517256 647209
rect 517210 647137 517256 647175
rect 517210 647103 517216 647137
rect 517250 647103 517256 647137
rect 517210 647065 517256 647103
rect 517210 647031 517216 647065
rect 517250 647031 517256 647065
rect 517210 646993 517256 647031
rect 516792 646959 516798 646980
rect 516752 646921 516798 646959
rect 516752 646887 516758 646921
rect 516792 646887 516798 646921
rect 516752 646849 516798 646887
rect 516752 646815 516758 646849
rect 516792 646815 516798 646849
rect 516752 646777 516798 646815
rect 516752 646743 516758 646777
rect 516792 646743 516798 646777
rect 515836 646671 515842 646705
rect 515876 646671 515882 646705
rect 515836 646633 515882 646671
rect 515836 646599 515842 646633
rect 515876 646599 515882 646633
rect 515836 646561 515882 646599
rect 515836 646527 515842 646561
rect 515876 646527 515882 646561
rect 515836 646489 515882 646527
rect 515418 646455 515424 646456
rect 515378 646417 515424 646455
rect 515378 646383 515384 646417
rect 515418 646383 515424 646417
rect 515378 646368 515424 646383
rect 515836 646455 515842 646489
rect 515876 646455 515882 646489
rect 516285 646706 516349 646712
rect 516285 646654 516291 646706
rect 516343 646654 516349 646706
rect 516285 646642 516349 646654
rect 516285 646590 516291 646642
rect 516343 646590 516349 646642
rect 516285 646578 516349 646590
rect 516285 646526 516291 646578
rect 516343 646526 516349 646578
rect 516285 646514 516349 646526
rect 516285 646462 516291 646514
rect 516343 646462 516349 646514
rect 516285 646456 516300 646462
rect 515836 646417 515882 646455
rect 515836 646383 515842 646417
rect 515876 646383 515882 646417
rect 515836 646368 515882 646383
rect 516294 646455 516300 646456
rect 516334 646456 516349 646462
rect 516752 646705 516798 646743
rect 517210 646959 517216 646993
rect 517250 646959 517256 646993
rect 517210 646921 517256 646959
rect 517210 646887 517216 646921
rect 517250 646887 517256 646921
rect 517210 646849 517256 646887
rect 517210 646815 517216 646849
rect 517250 646815 517256 646849
rect 517210 646777 517256 646815
rect 517210 646743 517216 646777
rect 517250 646743 517256 646777
rect 517210 646712 517256 646743
rect 516752 646671 516758 646705
rect 516792 646671 516798 646705
rect 516752 646633 516798 646671
rect 516752 646599 516758 646633
rect 516792 646599 516798 646633
rect 516752 646561 516798 646599
rect 516752 646527 516758 646561
rect 516792 646527 516798 646561
rect 516752 646489 516798 646527
rect 516334 646455 516340 646456
rect 516294 646417 516340 646455
rect 516294 646383 516300 646417
rect 516334 646383 516340 646417
rect 516294 646368 516340 646383
rect 516752 646455 516758 646489
rect 516792 646455 516798 646489
rect 517201 646706 517265 646712
rect 517201 646654 517207 646706
rect 517259 646654 517265 646706
rect 517201 646642 517265 646654
rect 517201 646590 517207 646642
rect 517259 646590 517265 646642
rect 517201 646578 517265 646590
rect 517201 646526 517207 646578
rect 517259 646526 517265 646578
rect 517201 646514 517265 646526
rect 517201 646462 517207 646514
rect 517259 646462 517265 646514
rect 517201 646456 517216 646462
rect 516752 646417 516798 646455
rect 516752 646383 516758 646417
rect 516792 646383 516798 646417
rect 516752 646368 516798 646383
rect 517210 646455 517216 646456
rect 517250 646456 517265 646462
rect 517554 646709 518116 646721
rect 517554 646459 517566 646709
rect 518104 646459 518116 646709
rect 517250 646455 517256 646456
rect 517210 646417 517256 646455
rect 517554 646447 518116 646459
rect 517210 646383 517216 646417
rect 517250 646383 517256 646417
rect 517210 646368 517256 646383
rect 513107 646108 513293 646158
<< via1 >>
rect 512588 649478 512768 649658
rect 508148 646299 508328 646479
rect 513142 649793 513258 649794
rect 513142 646159 513147 649793
rect 513147 646159 513253 649793
rect 513253 646159 513258 649793
rect 513142 646158 513258 646159
rect 518210 649648 518262 649649
rect 518210 649614 518219 649648
rect 518219 649614 518253 649648
rect 518253 649614 518262 649648
rect 518210 649597 518262 649614
rect 514301 649531 514353 649536
rect 514301 649497 514309 649531
rect 514309 649497 514343 649531
rect 514343 649497 514353 649531
rect 514301 649484 514353 649497
rect 514301 649459 514353 649472
rect 514301 649425 514309 649459
rect 514309 649425 514343 649459
rect 514343 649425 514353 649459
rect 514301 649420 514353 649425
rect 516456 649331 516508 649349
rect 516520 649331 516572 649349
rect 516584 649331 516636 649349
rect 516456 649297 516486 649331
rect 516486 649297 516508 649331
rect 516520 649297 516558 649331
rect 516558 649297 516572 649331
rect 516584 649297 516592 649331
rect 516592 649297 516630 649331
rect 516630 649297 516636 649331
rect 518210 649576 518262 649585
rect 518210 649542 518219 649576
rect 518219 649542 518253 649576
rect 518253 649542 518262 649576
rect 518210 649533 518262 649542
rect 518210 649504 518262 649521
rect 518210 649470 518219 649504
rect 518219 649470 518253 649504
rect 518253 649470 518262 649504
rect 518210 649469 518262 649470
rect 514112 649054 514164 649085
rect 514112 649033 514121 649054
rect 514121 649033 514155 649054
rect 514155 649033 514164 649054
rect 514112 649020 514121 649021
rect 514121 649020 514155 649021
rect 514155 649020 514164 649021
rect 514112 648982 514164 649020
rect 514112 648969 514121 648982
rect 514121 648969 514155 648982
rect 514155 648969 514164 648982
rect 514112 648948 514121 648957
rect 514121 648948 514155 648957
rect 514155 648948 514164 648957
rect 514112 648910 514164 648948
rect 514112 648905 514121 648910
rect 514121 648905 514155 648910
rect 514155 648905 514164 648910
rect 514112 648876 514121 648893
rect 514121 648876 514155 648893
rect 514155 648876 514164 648893
rect 514112 648841 514164 648876
rect 513654 648588 513663 648591
rect 513663 648588 513697 648591
rect 513697 648588 513706 648591
rect 513654 648550 513706 648588
rect 513654 648539 513663 648550
rect 513663 648539 513697 648550
rect 513697 648539 513706 648550
rect 513654 648516 513663 648527
rect 513663 648516 513697 648527
rect 513697 648516 513706 648527
rect 513654 648478 513706 648516
rect 513654 648475 513663 648478
rect 513663 648475 513697 648478
rect 513697 648475 513706 648478
rect 513654 648444 513663 648463
rect 513663 648444 513697 648463
rect 513697 648444 513706 648463
rect 513654 648411 513706 648444
rect 513654 648372 513663 648399
rect 513663 648372 513697 648399
rect 513697 648372 513706 648399
rect 513654 648347 513706 648372
rect 515028 649054 515080 649085
rect 515028 649033 515037 649054
rect 515037 649033 515071 649054
rect 515071 649033 515080 649054
rect 515028 649020 515037 649021
rect 515037 649020 515071 649021
rect 515071 649020 515080 649021
rect 515028 648982 515080 649020
rect 515028 648969 515037 648982
rect 515037 648969 515071 648982
rect 515071 648969 515080 648982
rect 515028 648948 515037 648957
rect 515037 648948 515071 648957
rect 515071 648948 515080 648957
rect 515028 648910 515080 648948
rect 515028 648905 515037 648910
rect 515037 648905 515071 648910
rect 515071 648905 515080 648910
rect 515028 648876 515037 648893
rect 515037 648876 515071 648893
rect 515071 648876 515080 648893
rect 515028 648841 515080 648876
rect 514570 648588 514579 648591
rect 514579 648588 514613 648591
rect 514613 648588 514622 648591
rect 514570 648550 514622 648588
rect 514570 648539 514579 648550
rect 514579 648539 514613 648550
rect 514613 648539 514622 648550
rect 514570 648516 514579 648527
rect 514579 648516 514613 648527
rect 514613 648516 514622 648527
rect 514570 648478 514622 648516
rect 514570 648475 514579 648478
rect 514579 648475 514613 648478
rect 514613 648475 514622 648478
rect 514570 648444 514579 648463
rect 514579 648444 514613 648463
rect 514613 648444 514622 648463
rect 514570 648411 514622 648444
rect 514570 648372 514579 648399
rect 514579 648372 514613 648399
rect 514613 648372 514622 648399
rect 514570 648347 514622 648372
rect 515604 649054 515656 649085
rect 515604 649033 515613 649054
rect 515613 649033 515647 649054
rect 515647 649033 515656 649054
rect 515604 649020 515613 649021
rect 515613 649020 515647 649021
rect 515647 649020 515656 649021
rect 515604 648982 515656 649020
rect 515604 648969 515613 648982
rect 515613 648969 515647 648982
rect 515647 648969 515656 648982
rect 515604 648948 515613 648957
rect 515613 648948 515647 648957
rect 515647 648948 515656 648957
rect 515604 648910 515656 648948
rect 515604 648905 515613 648910
rect 515613 648905 515647 648910
rect 515647 648905 515656 648910
rect 515604 648876 515613 648893
rect 515613 648876 515647 648893
rect 515647 648876 515656 648893
rect 515604 648841 515656 648876
rect 515486 648588 515495 648591
rect 515495 648588 515529 648591
rect 515529 648588 515538 648591
rect 515486 648550 515538 648588
rect 515486 648539 515495 648550
rect 515495 648539 515529 648550
rect 515529 648539 515538 648550
rect 515486 648516 515495 648527
rect 515495 648516 515529 648527
rect 515529 648516 515538 648527
rect 515486 648478 515538 648516
rect 515486 648475 515495 648478
rect 515495 648475 515529 648478
rect 515529 648475 515538 648478
rect 515486 648444 515495 648463
rect 515495 648444 515529 648463
rect 515529 648444 515538 648463
rect 515486 648411 515538 648444
rect 515486 648372 515495 648399
rect 515495 648372 515529 648399
rect 515529 648372 515538 648399
rect 515486 648347 515538 648372
rect 516520 649054 516572 649085
rect 516520 649033 516529 649054
rect 516529 649033 516563 649054
rect 516563 649033 516572 649054
rect 516520 649020 516529 649021
rect 516529 649020 516563 649021
rect 516563 649020 516572 649021
rect 516520 648982 516572 649020
rect 516520 648969 516529 648982
rect 516529 648969 516563 648982
rect 516563 648969 516572 648982
rect 516520 648948 516529 648957
rect 516529 648948 516563 648957
rect 516563 648948 516572 648957
rect 516520 648910 516572 648948
rect 516520 648905 516529 648910
rect 516529 648905 516563 648910
rect 516563 648905 516572 648910
rect 516520 648876 516529 648893
rect 516529 648876 516563 648893
rect 516563 648876 516572 648893
rect 516520 648841 516572 648876
rect 516062 648588 516071 648591
rect 516071 648588 516105 648591
rect 516105 648588 516114 648591
rect 516062 648550 516114 648588
rect 516062 648539 516071 648550
rect 516071 648539 516105 648550
rect 516105 648539 516114 648550
rect 516062 648516 516071 648527
rect 516071 648516 516105 648527
rect 516105 648516 516114 648527
rect 516062 648478 516114 648516
rect 516062 648475 516071 648478
rect 516071 648475 516105 648478
rect 516105 648475 516114 648478
rect 516062 648444 516071 648463
rect 516071 648444 516105 648463
rect 516105 648444 516114 648463
rect 516062 648411 516114 648444
rect 516062 648372 516071 648399
rect 516071 648372 516105 648399
rect 516105 648372 516114 648399
rect 516062 648347 516114 648372
rect 517436 649054 517488 649085
rect 517436 649033 517445 649054
rect 517445 649033 517479 649054
rect 517479 649033 517488 649054
rect 517436 649020 517445 649021
rect 517445 649020 517479 649021
rect 517479 649020 517488 649021
rect 517436 648982 517488 649020
rect 517436 648969 517445 648982
rect 517445 648969 517479 648982
rect 517479 648969 517488 648982
rect 517436 648948 517445 648957
rect 517445 648948 517479 648957
rect 517479 648948 517488 648957
rect 517436 648910 517488 648948
rect 517436 648905 517445 648910
rect 517445 648905 517479 648910
rect 517479 648905 517488 648910
rect 517436 648876 517445 648893
rect 517445 648876 517479 648893
rect 517479 648876 517488 648893
rect 517436 648841 517488 648876
rect 516978 648588 516987 648591
rect 516987 648588 517021 648591
rect 517021 648588 517030 648591
rect 516978 648550 517030 648588
rect 516978 648539 516987 648550
rect 516987 648539 517021 648550
rect 517021 648539 517030 648550
rect 516978 648516 516987 648527
rect 516987 648516 517021 648527
rect 517021 648516 517030 648527
rect 516978 648478 517030 648516
rect 516978 648475 516987 648478
rect 516987 648475 517021 648478
rect 517021 648475 517030 648478
rect 516978 648444 516987 648463
rect 516987 648444 517021 648463
rect 517021 648444 517030 648463
rect 516978 648411 517030 648444
rect 516978 648372 516987 648399
rect 516987 648372 517021 648399
rect 517021 648372 517030 648399
rect 516978 648347 517030 648372
rect 518012 649054 518064 649085
rect 518012 649033 518021 649054
rect 518021 649033 518055 649054
rect 518055 649033 518064 649054
rect 518012 649020 518021 649021
rect 518021 649020 518055 649021
rect 518055 649020 518064 649021
rect 518012 648982 518064 649020
rect 518012 648969 518021 648982
rect 518021 648969 518055 648982
rect 518055 648969 518064 648982
rect 518012 648948 518021 648957
rect 518021 648948 518055 648957
rect 518055 648948 518064 648957
rect 518012 648910 518064 648948
rect 518012 648905 518021 648910
rect 518021 648905 518055 648910
rect 518055 648905 518064 648910
rect 518012 648876 518021 648893
rect 518021 648876 518055 648893
rect 518055 648876 518064 648893
rect 518012 648841 518064 648876
rect 518209 649054 518218 649085
rect 518218 649054 518252 649085
rect 518252 649054 518261 649085
rect 518209 649033 518261 649054
rect 518209 649016 518261 649021
rect 518209 648982 518218 649016
rect 518218 648982 518252 649016
rect 518252 648982 518261 649016
rect 518209 648969 518261 648982
rect 518209 648944 518261 648957
rect 518209 648910 518218 648944
rect 518218 648910 518252 648944
rect 518252 648910 518261 648944
rect 518209 648905 518261 648910
rect 518209 648872 518261 648893
rect 518209 648841 518218 648872
rect 518218 648841 518252 648872
rect 518252 648841 518261 648872
rect 517554 648588 517563 648591
rect 517563 648588 517597 648591
rect 517597 648588 517606 648591
rect 517554 648550 517606 648588
rect 517554 648539 517563 648550
rect 517563 648539 517597 648550
rect 517597 648539 517606 648550
rect 517554 648516 517563 648527
rect 517563 648516 517597 648527
rect 517597 648516 517606 648527
rect 517554 648478 517606 648516
rect 517554 648475 517563 648478
rect 517563 648475 517597 648478
rect 517597 648475 517606 648478
rect 517554 648444 517563 648463
rect 517563 648444 517597 648463
rect 517597 648444 517606 648463
rect 517554 648411 517606 648444
rect 517554 648372 517563 648399
rect 517563 648372 517597 648399
rect 517597 648372 517606 648399
rect 517554 648347 517606 648372
rect 514474 648132 514494 648166
rect 514494 648132 514526 648166
rect 514474 648114 514526 648132
rect 514538 648114 514590 648166
rect 514602 648114 514654 648166
rect 514666 648132 514698 648166
rect 514698 648132 514718 648166
rect 514666 648114 514718 648132
rect 515669 648132 515698 648166
rect 515698 648132 515721 648166
rect 515733 648132 515770 648166
rect 515770 648132 515785 648166
rect 515797 648132 515804 648166
rect 515804 648132 515842 648166
rect 515842 648132 515849 648166
rect 515669 648114 515721 648132
rect 515733 648114 515785 648132
rect 515797 648114 515849 648132
rect 517719 648132 517720 648166
rect 517720 648132 517754 648166
rect 517754 648132 517771 648166
rect 517719 648114 517771 648132
rect 517783 648132 517792 648166
rect 517792 648132 517826 648166
rect 517826 648132 517835 648166
rect 517783 648114 517835 648132
rect 517847 648132 517864 648166
rect 517864 648132 517898 648166
rect 517898 648132 517899 648166
rect 517847 648114 517899 648132
rect 515082 647440 515134 647458
rect 515082 647406 515083 647440
rect 515083 647406 515117 647440
rect 515117 647406 515134 647440
rect 515146 647440 515198 647458
rect 515146 647406 515155 647440
rect 515155 647406 515189 647440
rect 515189 647406 515198 647440
rect 515210 647440 515262 647458
rect 515210 647406 515227 647440
rect 515227 647406 515261 647440
rect 515261 647406 515262 647440
rect 515540 647440 515592 647458
rect 515540 647406 515541 647440
rect 515541 647406 515575 647440
rect 515575 647406 515592 647440
rect 515604 647440 515656 647458
rect 515604 647406 515613 647440
rect 515613 647406 515647 647440
rect 515647 647406 515656 647440
rect 515668 647440 515720 647458
rect 515668 647406 515685 647440
rect 515685 647406 515719 647440
rect 515719 647406 515720 647440
rect 516456 647440 516508 647458
rect 516456 647406 516457 647440
rect 516457 647406 516491 647440
rect 516491 647406 516508 647440
rect 516520 647440 516572 647458
rect 516520 647406 516529 647440
rect 516529 647406 516563 647440
rect 516563 647406 516572 647440
rect 516584 647440 516636 647458
rect 516584 647406 516601 647440
rect 516601 647406 516635 647440
rect 516635 647406 516636 647440
rect 514917 647209 514969 647230
rect 514917 647178 514926 647209
rect 514926 647178 514960 647209
rect 514960 647178 514969 647209
rect 514917 647137 514969 647166
rect 514917 647114 514926 647137
rect 514926 647114 514960 647137
rect 514960 647114 514969 647137
rect 514917 647065 514969 647102
rect 514917 647050 514926 647065
rect 514926 647050 514960 647065
rect 514960 647050 514969 647065
rect 514917 647031 514926 647038
rect 514926 647031 514960 647038
rect 514960 647031 514969 647038
rect 514917 646993 514969 647031
rect 514917 646986 514926 646993
rect 514926 646986 514960 646993
rect 514960 646986 514969 646993
rect 513629 646462 514129 646706
rect 514459 646705 514511 646706
rect 514459 646671 514468 646705
rect 514468 646671 514502 646705
rect 514502 646671 514511 646705
rect 514459 646654 514511 646671
rect 514459 646633 514511 646642
rect 514459 646599 514468 646633
rect 514468 646599 514502 646633
rect 514502 646599 514511 646633
rect 514459 646590 514511 646599
rect 514459 646561 514511 646578
rect 514459 646527 514468 646561
rect 514468 646527 514502 646561
rect 514502 646527 514511 646561
rect 514459 646526 514511 646527
rect 514459 646489 514511 646514
rect 514459 646462 514468 646489
rect 514468 646462 514502 646489
rect 514502 646462 514511 646489
rect 515833 647209 515885 647230
rect 515833 647178 515842 647209
rect 515842 647178 515876 647209
rect 515876 647178 515885 647209
rect 515833 647137 515885 647166
rect 515833 647114 515842 647137
rect 515842 647114 515876 647137
rect 515876 647114 515885 647137
rect 515833 647065 515885 647102
rect 515833 647050 515842 647065
rect 515842 647050 515876 647065
rect 515876 647050 515885 647065
rect 515833 647031 515842 647038
rect 515842 647031 515876 647038
rect 515876 647031 515885 647038
rect 515833 646993 515885 647031
rect 515833 646986 515842 646993
rect 515842 646986 515876 646993
rect 515876 646986 515885 646993
rect 515375 646705 515427 646706
rect 515375 646671 515384 646705
rect 515384 646671 515418 646705
rect 515418 646671 515427 646705
rect 515375 646654 515427 646671
rect 515375 646633 515427 646642
rect 515375 646599 515384 646633
rect 515384 646599 515418 646633
rect 515418 646599 515427 646633
rect 515375 646590 515427 646599
rect 515375 646561 515427 646578
rect 515375 646527 515384 646561
rect 515384 646527 515418 646561
rect 515418 646527 515427 646561
rect 515375 646526 515427 646527
rect 515375 646489 515427 646514
rect 515375 646462 515384 646489
rect 515384 646462 515418 646489
rect 515418 646462 515427 646489
rect 516749 647209 516801 647230
rect 516749 647178 516758 647209
rect 516758 647178 516792 647209
rect 516792 647178 516801 647209
rect 516749 647137 516801 647166
rect 516749 647114 516758 647137
rect 516758 647114 516792 647137
rect 516792 647114 516801 647137
rect 516749 647065 516801 647102
rect 516749 647050 516758 647065
rect 516758 647050 516792 647065
rect 516792 647050 516801 647065
rect 516749 647031 516758 647038
rect 516758 647031 516792 647038
rect 516792 647031 516801 647038
rect 516749 646993 516801 647031
rect 516749 646986 516758 646993
rect 516758 646986 516792 646993
rect 516792 646986 516801 646993
rect 516291 646705 516343 646706
rect 516291 646671 516300 646705
rect 516300 646671 516334 646705
rect 516334 646671 516343 646705
rect 516291 646654 516343 646671
rect 516291 646633 516343 646642
rect 516291 646599 516300 646633
rect 516300 646599 516334 646633
rect 516334 646599 516343 646633
rect 516291 646590 516343 646599
rect 516291 646561 516343 646578
rect 516291 646527 516300 646561
rect 516300 646527 516334 646561
rect 516334 646527 516343 646561
rect 516291 646526 516343 646527
rect 516291 646489 516343 646514
rect 516291 646462 516300 646489
rect 516300 646462 516334 646489
rect 516334 646462 516343 646489
rect 517207 646705 517259 646706
rect 517207 646671 517216 646705
rect 517216 646671 517250 646705
rect 517250 646671 517259 646705
rect 517207 646654 517259 646671
rect 517207 646633 517259 646642
rect 517207 646599 517216 646633
rect 517216 646599 517250 646633
rect 517250 646599 517259 646633
rect 517207 646590 517259 646599
rect 517207 646561 517259 646578
rect 517207 646527 517216 646561
rect 517216 646527 517250 646561
rect 517250 646527 517259 646561
rect 517207 646526 517259 646527
rect 517207 646489 517259 646514
rect 517207 646462 517216 646489
rect 517216 646462 517250 646489
rect 517250 646462 517259 646489
rect 517585 646462 518085 646706
<< metal2 >>
rect 513107 649794 513293 649842
rect 512561 649676 512795 649685
rect 512561 649460 512570 649676
rect 512786 649460 512795 649676
rect 512561 649451 512795 649460
rect 508121 646497 508355 646506
rect 508121 646281 508130 646497
rect 508346 646281 508355 646497
rect 508121 646272 508355 646281
rect 513107 646158 513142 649794
rect 513258 646158 513293 649794
rect 518182 649667 518288 649690
rect 518182 649611 518208 649667
rect 518264 649611 518288 649667
rect 518182 649597 518210 649611
rect 518262 649597 518288 649611
rect 518182 649587 518288 649597
rect 514291 649536 514359 649542
rect 514291 649504 514301 649536
rect 513873 649484 514301 649504
rect 514353 649484 514359 649536
rect 513873 649472 514359 649484
rect 513873 649420 514301 649472
rect 514353 649420 514359 649472
rect 513873 649414 514359 649420
rect 518182 649531 518208 649587
rect 518264 649531 518288 649587
rect 518182 649521 518288 649531
rect 518182 649507 518210 649521
rect 518262 649507 518288 649521
rect 518182 649451 518208 649507
rect 518264 649451 518288 649507
rect 513648 648591 513712 648597
rect 513648 648539 513654 648591
rect 513706 648549 513712 648591
rect 513873 648549 513954 649414
rect 516429 649351 516663 649360
rect 516429 649295 516438 649351
rect 516494 649349 516518 649351
rect 516574 649349 516598 649351
rect 516508 649297 516518 649349
rect 516574 649297 516584 649349
rect 516494 649295 516518 649297
rect 516574 649295 516598 649297
rect 516654 649295 516663 649351
rect 516429 649286 516663 649295
rect 514106 649085 514170 649091
rect 514106 649033 514112 649085
rect 514164 649043 514170 649085
rect 515022 649085 515086 649091
rect 515022 649043 515028 649085
rect 514164 649033 515028 649043
rect 515080 649033 515086 649085
rect 514106 649031 515086 649033
rect 514106 649021 514875 649031
rect 514106 648969 514112 649021
rect 514164 648969 514875 649021
rect 514106 648957 514875 648969
rect 514106 648905 514112 648957
rect 514164 648905 514875 648957
rect 514106 648895 514875 648905
rect 515011 649021 515086 649031
rect 515011 648969 515028 649021
rect 515080 648969 515086 649021
rect 515011 648957 515086 648969
rect 515011 648905 515028 648957
rect 515080 648905 515086 648957
rect 515011 648895 515086 648905
rect 514106 648893 515086 648895
rect 514106 648841 514112 648893
rect 514164 648883 515028 648893
rect 514164 648841 514170 648883
rect 514106 648835 514170 648841
rect 515022 648841 515028 648883
rect 515080 648841 515086 648893
rect 515022 648835 515086 648841
rect 515598 649085 515662 649091
rect 515598 649033 515604 649085
rect 515656 649043 515662 649085
rect 516514 649085 516578 649091
rect 516514 649043 516520 649085
rect 515656 649033 516520 649043
rect 516572 649043 516578 649085
rect 517430 649085 517494 649091
rect 517430 649043 517436 649085
rect 516572 649033 517436 649043
rect 517488 649043 517494 649085
rect 518006 649085 518070 649091
rect 518006 649043 518012 649085
rect 517488 649033 518012 649043
rect 518064 649043 518070 649085
rect 518182 649085 518288 649451
rect 518182 649043 518209 649085
rect 518064 649033 518209 649043
rect 518261 649033 518288 649085
rect 515598 649031 518288 649033
rect 515598 649021 516822 649031
rect 517918 649021 518288 649031
rect 515598 648969 515604 649021
rect 515656 648969 516520 649021
rect 516572 648969 516822 649021
rect 517918 648969 518012 649021
rect 518064 648969 518209 649021
rect 518261 648969 518288 649021
rect 515598 648957 516822 648969
rect 517918 648957 518288 648969
rect 515598 648905 515604 648957
rect 515656 648905 516520 648957
rect 516572 648905 516822 648957
rect 517918 648905 518012 648957
rect 518064 648905 518209 648957
rect 518261 648905 518288 648957
rect 515598 648895 516822 648905
rect 517918 648895 518288 648905
rect 515598 648893 518288 648895
rect 515598 648841 515604 648893
rect 515656 648883 516520 648893
rect 515656 648841 515662 648883
rect 515598 648835 515662 648841
rect 516514 648841 516520 648883
rect 516572 648883 517436 648893
rect 516572 648841 516578 648883
rect 516514 648835 516578 648841
rect 517430 648841 517436 648883
rect 517488 648883 518012 648893
rect 517488 648841 517494 648883
rect 517430 648835 517494 648841
rect 518006 648841 518012 648883
rect 518064 648883 518209 648893
rect 518064 648841 518070 648883
rect 518006 648835 518070 648841
rect 518182 648841 518209 648883
rect 518261 648841 518288 648893
rect 518182 648825 518288 648841
rect 516051 648617 516125 648626
rect 514564 648591 514628 648597
rect 514564 648549 514570 648591
rect 513706 648539 514570 648549
rect 514622 648549 514628 648591
rect 515480 648591 515544 648597
rect 515480 648549 515486 648591
rect 514622 648539 515486 648549
rect 515538 648549 515544 648591
rect 516051 648561 516060 648617
rect 516116 648561 516125 648617
rect 517531 648617 517631 648626
rect 515538 648539 515839 648549
rect 513648 648537 515839 648539
rect 513648 648527 514413 648537
rect 514629 648527 515839 648537
rect 513648 648475 513654 648527
rect 513706 648475 514413 648527
rect 514629 648475 515486 648527
rect 515538 648475 515839 648527
rect 513648 648463 514413 648475
rect 514629 648463 515839 648475
rect 513648 648411 513654 648463
rect 513706 648411 514413 648463
rect 514629 648411 515486 648463
rect 515538 648411 515839 648463
rect 513648 648401 514413 648411
rect 514629 648401 515839 648411
rect 513648 648399 515839 648401
rect 513648 648347 513654 648399
rect 513706 648389 514570 648399
rect 513706 648347 513712 648389
rect 513648 648341 513712 648347
rect 514564 648347 514570 648389
rect 514622 648389 515486 648399
rect 514622 648347 514628 648389
rect 514564 648341 514628 648347
rect 515480 648347 515486 648389
rect 515538 648389 515839 648399
rect 515538 648347 515544 648389
rect 515480 648341 515544 648347
rect 515679 648172 515839 648389
rect 516051 648539 516062 648561
rect 516114 648549 516125 648561
rect 516972 648591 517036 648597
rect 516972 648549 516978 648591
rect 516114 648539 516978 648549
rect 517030 648539 517036 648591
rect 516051 648537 517036 648539
rect 516051 648481 516060 648537
rect 516116 648527 517036 648537
rect 516116 648481 516978 648527
rect 516051 648475 516062 648481
rect 516114 648475 516978 648481
rect 517030 648475 517036 648527
rect 516051 648463 517036 648475
rect 516051 648457 516062 648463
rect 516114 648457 516978 648463
rect 516051 648401 516060 648457
rect 516116 648411 516978 648457
rect 517030 648411 517036 648463
rect 516116 648401 517036 648411
rect 516051 648399 517036 648401
rect 516051 648377 516062 648399
rect 516114 648389 516978 648399
rect 516114 648377 516125 648389
rect 516051 648321 516060 648377
rect 516116 648321 516125 648377
rect 516972 648347 516978 648389
rect 517030 648347 517036 648399
rect 516972 648341 517036 648347
rect 517531 648561 517552 648617
rect 517608 648561 517631 648617
rect 517531 648539 517554 648561
rect 517606 648539 517631 648561
rect 517531 648537 517631 648539
rect 517531 648481 517552 648537
rect 517608 648481 517631 648537
rect 517531 648475 517554 648481
rect 517606 648475 517631 648481
rect 517531 648463 517631 648475
rect 517531 648457 517554 648463
rect 517606 648457 517631 648463
rect 517531 648401 517552 648457
rect 517608 648401 517631 648457
rect 517531 648399 517631 648401
rect 517531 648377 517554 648399
rect 517606 648377 517631 648399
rect 516051 648312 516125 648321
rect 517531 648321 517552 648377
rect 517608 648321 517631 648377
rect 517531 648190 517631 648321
rect 518123 648190 518382 648277
rect 517531 648177 518382 648190
rect 514468 648166 514724 648172
rect 514468 648114 514474 648166
rect 514526 648114 514538 648166
rect 514590 648114 514602 648166
rect 514654 648114 514666 648166
rect 514718 648114 514724 648166
rect 514468 648108 514724 648114
rect 515663 648166 515855 648172
rect 515663 648114 515669 648166
rect 515721 648114 515733 648166
rect 515785 648114 515797 648166
rect 515849 648114 515855 648166
rect 515663 648108 515855 648114
rect 517531 648166 518324 648177
rect 517531 648114 517719 648166
rect 517771 648114 517783 648166
rect 517835 648114 517847 648166
rect 517899 648114 518324 648166
rect 514546 647851 514646 648108
rect 517531 648090 518324 648114
rect 516011 647869 516165 647878
rect 516011 647851 516020 647869
rect 514546 647751 516020 647851
rect 516011 647733 516020 647751
rect 516156 647733 516165 647869
rect 516011 647724 516165 647733
rect 515076 647460 518382 647482
rect 515076 647458 516438 647460
rect 516494 647458 516518 647460
rect 516574 647458 516598 647460
rect 515076 647406 515082 647458
rect 515134 647406 515146 647458
rect 515198 647406 515210 647458
rect 515262 647406 515540 647458
rect 515592 647406 515604 647458
rect 515656 647406 515668 647458
rect 515720 647406 516438 647458
rect 516508 647406 516518 647458
rect 516574 647406 516584 647458
rect 515076 647404 516438 647406
rect 516494 647404 516518 647406
rect 516574 647404 516598 647406
rect 516654 647404 518382 647460
rect 515076 647382 518382 647404
rect 514906 647256 514980 647265
rect 514906 647200 514915 647256
rect 514971 647200 514980 647256
rect 516051 647256 516125 647265
rect 514906 647178 514917 647200
rect 514969 647178 514980 647200
rect 514906 647176 514980 647178
rect 514906 647120 514915 647176
rect 514971 647120 514980 647176
rect 514906 647114 514917 647120
rect 514969 647114 514980 647120
rect 514906 647102 514980 647114
rect 514906 647096 514917 647102
rect 514969 647096 514980 647102
rect 514906 647040 514915 647096
rect 514971 647040 514980 647096
rect 514906 647038 514980 647040
rect 514906 647016 514917 647038
rect 514969 647016 514980 647038
rect 514906 646960 514915 647016
rect 514971 646960 514980 647016
rect 515827 647230 515891 647236
rect 515827 647178 515833 647230
rect 515885 647188 515891 647230
rect 516051 647200 516060 647256
rect 516116 647200 516125 647256
rect 517543 647256 517617 647265
rect 516051 647188 516125 647200
rect 515885 647178 516125 647188
rect 515827 647176 516125 647178
rect 515827 647166 516060 647176
rect 515827 647114 515833 647166
rect 515885 647120 516060 647166
rect 516116 647120 516125 647176
rect 515885 647114 516125 647120
rect 515827 647102 516125 647114
rect 515827 647050 515833 647102
rect 515885 647096 516125 647102
rect 515885 647050 516060 647096
rect 515827 647040 516060 647050
rect 516116 647040 516125 647096
rect 515827 647038 516125 647040
rect 515827 646986 515833 647038
rect 515885 647028 516125 647038
rect 515885 646986 515891 647028
rect 515827 646980 515891 646986
rect 516051 647016 516125 647028
rect 514906 646951 514980 646960
rect 516051 646960 516060 647016
rect 516116 646960 516125 647016
rect 516743 647230 516807 647236
rect 516743 647178 516749 647230
rect 516801 647188 516807 647230
rect 517543 647200 517552 647256
rect 517608 647200 517617 647256
rect 517543 647188 517617 647200
rect 516801 647178 517617 647188
rect 516743 647176 517617 647178
rect 516743 647166 517552 647176
rect 516743 647114 516749 647166
rect 516801 647120 517552 647166
rect 517608 647120 517617 647176
rect 516801 647114 517617 647120
rect 516743 647102 517617 647114
rect 516743 647050 516749 647102
rect 516801 647096 517617 647102
rect 516801 647050 517552 647096
rect 516743 647040 517552 647050
rect 517608 647040 517617 647096
rect 516743 647038 517617 647040
rect 516743 646986 516749 647038
rect 516801 647028 517617 647038
rect 516801 646986 516807 647028
rect 516743 646980 516807 646986
rect 517543 647016 517617 647028
rect 516051 646951 516125 646960
rect 517543 646960 517552 647016
rect 517608 646960 517617 647016
rect 517543 646951 517617 646960
rect 513623 646706 514135 646712
rect 513623 646462 513629 646706
rect 514129 646664 514135 646706
rect 514453 646706 514517 646712
rect 514453 646664 514459 646706
rect 514129 646654 514459 646664
rect 514511 646664 514517 646706
rect 515369 646706 515433 646712
rect 515369 646664 515375 646706
rect 514511 646654 515375 646664
rect 515427 646664 515433 646706
rect 516285 646706 516349 646712
rect 516285 646664 516291 646706
rect 515427 646654 516291 646664
rect 516343 646664 516349 646706
rect 517201 646706 517265 646712
rect 517201 646664 517207 646706
rect 516343 646654 517207 646664
rect 517259 646664 517265 646706
rect 517579 646706 518091 646712
rect 517579 646664 517585 646706
rect 517259 646654 517585 646664
rect 514129 646652 517585 646654
rect 514129 646642 514531 646652
rect 515627 646642 517585 646652
rect 514129 646590 514459 646642
rect 514511 646590 514531 646642
rect 515627 646590 516291 646642
rect 516343 646590 517207 646642
rect 517259 646590 517585 646642
rect 514129 646578 514531 646590
rect 515627 646578 517585 646590
rect 514129 646526 514459 646578
rect 514511 646526 514531 646578
rect 515627 646526 516291 646578
rect 516343 646526 517207 646578
rect 517259 646526 517585 646578
rect 514129 646516 514531 646526
rect 515627 646516 517585 646526
rect 514129 646514 517585 646516
rect 514129 646504 514459 646514
rect 514129 646462 514135 646504
rect 513623 646456 514135 646462
rect 514453 646462 514459 646504
rect 514511 646504 515375 646514
rect 514511 646462 514517 646504
rect 514453 646456 514517 646462
rect 515369 646462 515375 646504
rect 515427 646504 516291 646514
rect 515427 646462 515433 646504
rect 515369 646456 515433 646462
rect 516285 646462 516291 646504
rect 516343 646504 517207 646514
rect 516343 646462 516349 646504
rect 516285 646456 516349 646462
rect 517201 646462 517207 646504
rect 517259 646504 517585 646514
rect 517259 646462 517265 646504
rect 517201 646456 517265 646462
rect 517579 646462 517585 646504
rect 518085 646462 518091 646706
rect 517579 646456 518091 646462
rect 513107 646108 513293 646158
<< via2 >>
rect 512570 649658 512786 649676
rect 512570 649478 512588 649658
rect 512588 649478 512768 649658
rect 512768 649478 512786 649658
rect 512570 649460 512786 649478
rect 508130 646479 508346 646497
rect 508130 646299 508148 646479
rect 508148 646299 508328 646479
rect 508328 646299 508346 646479
rect 508130 646281 508346 646299
rect 513172 649580 513228 649636
rect 513172 649500 513228 649556
rect 518208 649649 518264 649667
rect 518208 649611 518210 649649
rect 518210 649611 518262 649649
rect 518262 649611 518264 649649
rect 518208 649585 518264 649587
rect 518208 649533 518210 649585
rect 518210 649533 518262 649585
rect 518262 649533 518264 649585
rect 518208 649531 518264 649533
rect 518208 649469 518210 649507
rect 518210 649469 518262 649507
rect 518262 649469 518264 649507
rect 518208 649451 518264 649469
rect 516438 649349 516494 649351
rect 516518 649349 516574 649351
rect 516598 649349 516654 649351
rect 516438 649297 516456 649349
rect 516456 649297 516494 649349
rect 516518 649297 516520 649349
rect 516520 649297 516572 649349
rect 516572 649297 516574 649349
rect 516598 649297 516636 649349
rect 516636 649297 516654 649349
rect 516438 649295 516494 649297
rect 516518 649295 516574 649297
rect 516598 649295 516654 649297
rect 514875 648895 515011 649031
rect 516822 649021 517918 649031
rect 516822 648969 517436 649021
rect 517436 648969 517488 649021
rect 517488 648969 517918 649021
rect 516822 648957 517918 648969
rect 516822 648905 517436 648957
rect 517436 648905 517488 648957
rect 517488 648905 517918 648957
rect 516822 648895 517918 648905
rect 516060 648591 516116 648617
rect 516060 648561 516062 648591
rect 516062 648561 516114 648591
rect 516114 648561 516116 648591
rect 514413 648527 514629 648537
rect 514413 648475 514570 648527
rect 514570 648475 514622 648527
rect 514622 648475 514629 648527
rect 514413 648463 514629 648475
rect 514413 648411 514570 648463
rect 514570 648411 514622 648463
rect 514622 648411 514629 648463
rect 514413 648401 514629 648411
rect 516060 648527 516116 648537
rect 516060 648481 516062 648527
rect 516062 648481 516114 648527
rect 516114 648481 516116 648527
rect 516060 648411 516062 648457
rect 516062 648411 516114 648457
rect 516114 648411 516116 648457
rect 516060 648401 516116 648411
rect 516060 648347 516062 648377
rect 516062 648347 516114 648377
rect 516114 648347 516116 648377
rect 516060 648321 516116 648347
rect 517552 648591 517608 648617
rect 517552 648561 517554 648591
rect 517554 648561 517606 648591
rect 517606 648561 517608 648591
rect 517552 648527 517608 648537
rect 517552 648481 517554 648527
rect 517554 648481 517606 648527
rect 517606 648481 517608 648527
rect 517552 648411 517554 648457
rect 517554 648411 517606 648457
rect 517606 648411 517608 648457
rect 517552 648401 517608 648411
rect 517552 648347 517554 648377
rect 517554 648347 517606 648377
rect 517606 648347 517608 648377
rect 517552 648321 517608 648347
rect 516020 647733 516156 647869
rect 516438 647458 516494 647460
rect 516518 647458 516574 647460
rect 516598 647458 516654 647460
rect 516438 647406 516456 647458
rect 516456 647406 516494 647458
rect 516518 647406 516520 647458
rect 516520 647406 516572 647458
rect 516572 647406 516574 647458
rect 516598 647406 516636 647458
rect 516636 647406 516654 647458
rect 516438 647404 516494 647406
rect 516518 647404 516574 647406
rect 516598 647404 516654 647406
rect 514915 647230 514971 647256
rect 514915 647200 514917 647230
rect 514917 647200 514969 647230
rect 514969 647200 514971 647230
rect 514915 647166 514971 647176
rect 514915 647120 514917 647166
rect 514917 647120 514969 647166
rect 514969 647120 514971 647166
rect 514915 647050 514917 647096
rect 514917 647050 514969 647096
rect 514969 647050 514971 647096
rect 514915 647040 514971 647050
rect 514915 646986 514917 647016
rect 514917 646986 514969 647016
rect 514969 646986 514971 647016
rect 514915 646960 514971 646986
rect 516060 647200 516116 647256
rect 516060 647120 516116 647176
rect 516060 647040 516116 647096
rect 516060 646960 516116 647016
rect 517552 647200 517608 647256
rect 517552 647120 517608 647176
rect 517552 647040 517608 647096
rect 517552 646960 517608 647016
rect 514531 646642 515627 646652
rect 514531 646590 515375 646642
rect 515375 646590 515427 646642
rect 515427 646590 515627 646642
rect 514531 646578 515627 646590
rect 514531 646526 515375 646578
rect 515375 646526 515427 646578
rect 515427 646526 515627 646578
rect 514531 646516 515627 646526
<< metal3 >>
rect 512561 649676 512795 649685
rect 512561 649460 512570 649676
rect 512786 649648 512795 649676
rect 518182 649667 518288 649690
rect 513133 649648 513267 649656
rect 518182 649648 518208 649667
rect 512786 649636 518208 649648
rect 512786 649580 513172 649636
rect 513228 649611 518208 649636
rect 518264 649611 518288 649667
rect 513228 649599 518288 649611
rect 513228 649580 516817 649599
rect 512786 649556 516817 649580
rect 512786 649500 513172 649556
rect 513228 649535 516817 649556
rect 516881 649535 516897 649599
rect 516961 649535 516977 649599
rect 517041 649535 517057 649599
rect 517121 649535 517137 649599
rect 517201 649535 517217 649599
rect 517281 649535 517297 649599
rect 517361 649535 517377 649599
rect 517441 649535 517457 649599
rect 517521 649535 517537 649599
rect 517601 649535 517617 649599
rect 517681 649535 517697 649599
rect 517761 649535 517777 649599
rect 517841 649535 517857 649599
rect 517921 649587 518288 649599
rect 517921 649535 518208 649587
rect 513228 649531 518208 649535
rect 518264 649531 518288 649587
rect 513228 649507 518288 649531
rect 513228 649500 518208 649507
rect 512786 649488 518208 649500
rect 512786 649460 512795 649488
rect 513133 649480 513267 649488
rect 512561 649451 512795 649460
rect 516429 649351 516663 649360
rect 516429 649295 516438 649351
rect 516494 649295 516518 649351
rect 516574 649295 516598 649351
rect 516654 649295 516663 649351
rect 516429 649286 516663 649295
rect 514866 649031 515020 649040
rect 514866 648895 514875 649031
rect 515011 648895 515020 649031
rect 514866 648886 515020 648895
rect 513336 648537 514644 648549
rect 513336 648401 514413 648537
rect 514629 648401 514644 648537
rect 513336 648389 514644 648401
rect 508121 646497 508355 646506
rect 508121 646281 508130 646497
rect 508346 646470 508355 646497
rect 513336 646470 513496 648389
rect 514893 647256 514993 648886
rect 516038 648617 516138 648626
rect 516038 648561 516060 648617
rect 516116 648561 516138 648617
rect 516038 648537 516138 648561
rect 516038 648481 516060 648537
rect 516116 648481 516138 648537
rect 516038 648457 516138 648481
rect 516038 648401 516060 648457
rect 516116 648401 516138 648457
rect 516038 648377 516138 648401
rect 516038 648321 516060 648377
rect 516116 648321 516138 648377
rect 516038 647878 516138 648321
rect 516011 647869 516165 647878
rect 516011 647733 516020 647869
rect 516156 647733 516165 647869
rect 516011 647724 516165 647733
rect 514893 647200 514915 647256
rect 514971 647200 514993 647256
rect 514893 647176 514993 647200
rect 514893 647120 514915 647176
rect 514971 647120 514993 647176
rect 514893 647096 514993 647120
rect 514893 647040 514915 647096
rect 514971 647040 514993 647096
rect 514893 647016 514993 647040
rect 514893 646960 514915 647016
rect 514971 646960 514993 647016
rect 514893 646951 514993 646960
rect 516038 647256 516138 647724
rect 516496 647469 516596 649286
rect 516958 649056 517118 649488
rect 518182 649451 518208 649488
rect 518264 649451 518288 649507
rect 518182 649432 518288 649451
rect 516782 649050 517958 649056
rect 516782 648986 516788 649050
rect 516852 649031 516898 649050
rect 516962 649031 517008 649050
rect 517072 649031 517118 649050
rect 517182 649031 517228 649050
rect 517292 649031 517338 649050
rect 517402 649031 517448 649050
rect 517512 649031 517558 649050
rect 517622 649031 517668 649050
rect 517732 649031 517778 649050
rect 517842 649031 517888 649050
rect 517952 648986 517958 649050
rect 516782 648940 516822 648986
rect 517918 648940 517958 648986
rect 516782 648876 516788 648940
rect 516852 648876 516898 648895
rect 516962 648876 517008 648895
rect 517072 648876 517118 648895
rect 517182 648876 517228 648895
rect 517292 648876 517338 648895
rect 517402 648876 517448 648895
rect 517512 648876 517558 648895
rect 517622 648876 517668 648895
rect 517732 648876 517778 648895
rect 517842 648876 517888 648895
rect 517952 648876 517958 648940
rect 516782 648870 517958 648876
rect 517531 648617 517631 648626
rect 517531 648561 517552 648617
rect 517608 648561 517631 648617
rect 517531 648537 517631 648561
rect 517531 648481 517552 648537
rect 517608 648481 517631 648537
rect 517531 648457 517631 648481
rect 517531 648401 517552 648457
rect 517608 648401 517631 648457
rect 517531 648377 517631 648401
rect 517531 648321 517552 648377
rect 517608 648321 517631 648377
rect 516429 647460 516663 647469
rect 516429 647404 516438 647460
rect 516494 647404 516518 647460
rect 516574 647404 516598 647460
rect 516654 647404 516663 647460
rect 516429 647395 516663 647404
rect 516038 647200 516060 647256
rect 516116 647200 516138 647256
rect 516038 647176 516138 647200
rect 516038 647120 516060 647176
rect 516116 647120 516138 647176
rect 516038 647096 516138 647120
rect 516038 647040 516060 647096
rect 516116 647040 516138 647096
rect 516038 647016 516138 647040
rect 516038 646960 516060 647016
rect 516116 646960 516138 647016
rect 516038 646951 516138 646960
rect 514491 646671 515667 646677
rect 514491 646607 514497 646671
rect 514561 646652 514607 646671
rect 514671 646652 514717 646671
rect 514781 646652 514827 646671
rect 514891 646652 514937 646671
rect 515001 646652 515047 646671
rect 515111 646652 515157 646671
rect 515221 646652 515267 646671
rect 515331 646652 515377 646671
rect 515441 646652 515487 646671
rect 515551 646652 515597 646671
rect 515661 646607 515667 646671
rect 514491 646561 514531 646607
rect 515627 646561 515667 646607
rect 514491 646497 514497 646561
rect 514561 646497 514607 646516
rect 514671 646497 514717 646516
rect 514781 646497 514827 646516
rect 514891 646497 514937 646516
rect 515001 646497 515047 646516
rect 515111 646497 515157 646516
rect 515221 646497 515267 646516
rect 515331 646497 515377 646516
rect 515441 646497 515487 646516
rect 515551 646497 515597 646516
rect 515661 646497 515667 646561
rect 514491 646491 515667 646497
rect 508346 646310 513496 646470
rect 508346 646281 508355 646310
rect 508121 646272 508355 646281
rect 516496 646263 516596 647395
rect 517531 647256 517631 648321
rect 517531 647200 517552 647256
rect 517608 647200 517631 647256
rect 517531 647176 517631 647200
rect 517531 647120 517552 647176
rect 517608 647120 517631 647176
rect 517531 647096 517631 647120
rect 517531 647040 517552 647096
rect 517608 647040 517631 647096
rect 517531 647016 517631 647040
rect 517531 646960 517552 647016
rect 517608 646960 517631 647016
rect 517531 646263 517631 646960
<< via3 >>
rect 516817 649535 516881 649599
rect 516897 649535 516961 649599
rect 516977 649535 517041 649599
rect 517057 649535 517121 649599
rect 517137 649535 517201 649599
rect 517217 649535 517281 649599
rect 517297 649535 517361 649599
rect 517377 649535 517441 649599
rect 517457 649535 517521 649599
rect 517537 649535 517601 649599
rect 517617 649535 517681 649599
rect 517697 649535 517761 649599
rect 517777 649535 517841 649599
rect 517857 649535 517921 649599
rect 516788 649031 516852 649050
rect 516898 649031 516962 649050
rect 517008 649031 517072 649050
rect 517118 649031 517182 649050
rect 517228 649031 517292 649050
rect 517338 649031 517402 649050
rect 517448 649031 517512 649050
rect 517558 649031 517622 649050
rect 517668 649031 517732 649050
rect 517778 649031 517842 649050
rect 517888 649031 517952 649050
rect 516788 648986 516822 649031
rect 516822 648986 516852 649031
rect 516898 648986 516962 649031
rect 517008 648986 517072 649031
rect 517118 648986 517182 649031
rect 517228 648986 517292 649031
rect 517338 648986 517402 649031
rect 517448 648986 517512 649031
rect 517558 648986 517622 649031
rect 517668 648986 517732 649031
rect 517778 648986 517842 649031
rect 517888 648986 517918 649031
rect 517918 648986 517952 649031
rect 516788 648895 516822 648940
rect 516822 648895 516852 648940
rect 516898 648895 516962 648940
rect 517008 648895 517072 648940
rect 517118 648895 517182 648940
rect 517228 648895 517292 648940
rect 517338 648895 517402 648940
rect 517448 648895 517512 648940
rect 517558 648895 517622 648940
rect 517668 648895 517732 648940
rect 517778 648895 517842 648940
rect 517888 648895 517918 648940
rect 517918 648895 517952 648940
rect 516788 648876 516852 648895
rect 516898 648876 516962 648895
rect 517008 648876 517072 648895
rect 517118 648876 517182 648895
rect 517228 648876 517292 648895
rect 517338 648876 517402 648895
rect 517448 648876 517512 648895
rect 517558 648876 517622 648895
rect 517668 648876 517732 648895
rect 517778 648876 517842 648895
rect 517888 648876 517952 648895
rect 514497 646652 514561 646671
rect 514607 646652 514671 646671
rect 514717 646652 514781 646671
rect 514827 646652 514891 646671
rect 514937 646652 515001 646671
rect 515047 646652 515111 646671
rect 515157 646652 515221 646671
rect 515267 646652 515331 646671
rect 515377 646652 515441 646671
rect 515487 646652 515551 646671
rect 515597 646652 515661 646671
rect 514497 646607 514531 646652
rect 514531 646607 514561 646652
rect 514607 646607 514671 646652
rect 514717 646607 514781 646652
rect 514827 646607 514891 646652
rect 514937 646607 515001 646652
rect 515047 646607 515111 646652
rect 515157 646607 515221 646652
rect 515267 646607 515331 646652
rect 515377 646607 515441 646652
rect 515487 646607 515551 646652
rect 515597 646607 515627 646652
rect 515627 646607 515661 646652
rect 514497 646516 514531 646561
rect 514531 646516 514561 646561
rect 514607 646516 514671 646561
rect 514717 646516 514781 646561
rect 514827 646516 514891 646561
rect 514937 646516 515001 646561
rect 515047 646516 515111 646561
rect 515157 646516 515221 646561
rect 515267 646516 515331 646561
rect 515377 646516 515441 646561
rect 515487 646516 515551 646561
rect 515597 646516 515627 646561
rect 515627 646516 515661 646561
rect 514497 646497 514561 646516
rect 514607 646497 514671 646516
rect 514717 646497 514781 646516
rect 514827 646497 514891 646516
rect 514937 646497 515001 646516
rect 515047 646497 515111 646516
rect 515157 646497 515221 646516
rect 515267 646497 515331 646516
rect 515377 646497 515441 646516
rect 515487 646497 515551 646516
rect 515597 646497 515661 646516
<< metal4 >>
rect 514484 646671 515684 649891
rect 514484 646607 514497 646671
rect 514561 646607 514607 646671
rect 514671 646607 514717 646671
rect 514781 646607 514827 646671
rect 514891 646607 514937 646671
rect 515001 646607 515047 646671
rect 515111 646607 515157 646671
rect 515221 646607 515267 646671
rect 515331 646607 515377 646671
rect 515441 646607 515487 646671
rect 515551 646607 515597 646671
rect 515661 646607 515684 646671
rect 514484 646561 515684 646607
rect 514484 646497 514497 646561
rect 514561 646497 514607 646561
rect 514671 646497 514717 646561
rect 514781 646497 514827 646561
rect 514891 646497 514937 646561
rect 515001 646497 515047 646561
rect 515111 646497 515157 646561
rect 515221 646497 515267 646561
rect 515331 646497 515377 646561
rect 515441 646497 515487 646561
rect 515551 646497 515597 646561
rect 515661 646497 515684 646561
rect 514484 646078 515684 646497
rect 516769 649599 517969 649891
rect 516769 649535 516817 649599
rect 516881 649535 516897 649599
rect 516961 649535 516977 649599
rect 517041 649535 517057 649599
rect 517121 649535 517137 649599
rect 517201 649535 517217 649599
rect 517281 649535 517297 649599
rect 517361 649535 517377 649599
rect 517441 649535 517457 649599
rect 517521 649535 517537 649599
rect 517601 649535 517617 649599
rect 517681 649535 517697 649599
rect 517761 649535 517777 649599
rect 517841 649535 517857 649599
rect 517921 649535 517969 649599
rect 516769 649050 517969 649535
rect 516769 648986 516788 649050
rect 516852 648986 516898 649050
rect 516962 648986 517008 649050
rect 517072 648986 517118 649050
rect 517182 648986 517228 649050
rect 517292 648986 517338 649050
rect 517402 648986 517448 649050
rect 517512 648986 517558 649050
rect 517622 648986 517668 649050
rect 517732 648986 517778 649050
rect 517842 648986 517888 649050
rect 517952 648986 517969 649050
rect 516769 648940 517969 648986
rect 516769 648876 516788 648940
rect 516852 648876 516898 648940
rect 516962 648876 517008 648940
rect 517072 648876 517118 648940
rect 517182 648876 517228 648940
rect 517292 648876 517338 648940
rect 517402 648876 517448 648940
rect 517512 648876 517558 648940
rect 517622 648876 517668 648940
rect 517732 648876 517778 648940
rect 517842 648876 517888 648940
rect 517952 648876 517969 648940
rect 516769 646078 517969 648876
<< labels >>
flabel metal2 s 518300 647431 518300 647431 0 FreeSans 455 0 0 0 VBN
flabel metal2 s 517339 646584 517339 646584 0 FreeSans 455 0 0 0 VSS
flabel metal2 s 518142 648962 518142 648962 0 FreeSans 455 0 0 0 VDD
flabel metal2 s 518302 648140 518302 648140 0 FreeSans 455 0 0 0 VBP
<< end >>
