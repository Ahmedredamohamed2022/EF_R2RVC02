magic
tech sky130A
magscale 1 2
timestamp 1694080139
<< checkpaint >>
rect -3244 -9876 15464 12536
<< metal1 >>
rect 518 -833 3398 -806
rect 518 -949 524 -833
rect 3392 -949 3398 -833
rect 518 -976 3398 -949
rect 7128 -828 10212 -806
rect 7128 -944 7140 -828
rect 10200 -944 10212 -828
rect 7128 -966 10212 -944
rect 2610 -3843 2814 -3778
rect 2610 -4086 2653 -3843
rect 2600 -4620 2653 -4086
rect 2610 -5047 2653 -4620
rect 2769 -5047 2814 -3843
rect 2610 -5114 2814 -5047
rect 5960 -3827 6146 -3764
rect 5960 -5031 5993 -3827
rect 6109 -5031 6146 -3827
rect 5960 -5098 6146 -5031
rect 9230 -3870 9428 -3804
rect 9230 -5074 9267 -3870
rect 9383 -4022 9428 -3870
rect 12582 -3842 12772 -3784
rect 9383 -4516 9438 -4022
rect 9383 -5074 9428 -4516
rect 9230 -5124 9428 -5074
rect 12582 -5046 12616 -3842
rect 12732 -5046 12772 -3842
rect 12582 -5094 12772 -5046
rect 2834 -7003 12762 -6799
rect 1216 -7670 1734 -7558
rect 8114 -7684 8640 -7570
rect 13236 -7834 13452 -7822
rect -26 -7863 13456 -7834
rect -26 -7979 13254 -7863
rect 13434 -7979 13456 -7863
rect -26 -7998 13456 -7979
rect 11192 -8002 13456 -7998
rect 13236 -8010 13452 -8002
<< via1 >>
rect 524 -949 3392 -833
rect 7140 -944 10200 -828
rect 2653 -5047 2769 -3843
rect 5993 -5031 6109 -3827
rect 9267 -5074 9383 -3870
rect 12616 -5046 12732 -3842
rect 13254 -7979 13434 -7863
<< metal2 >>
rect 12182 5605 13904 5678
rect 12182 5229 13739 5605
rect 13875 5229 13904 5605
rect 12182 5168 13904 5229
rect 11862 4416 11988 4494
rect 12092 4484 14042 4500
rect 12092 4428 13637 4484
rect 13693 4428 13717 4484
rect 13773 4428 13797 4484
rect 13853 4428 13877 4484
rect 13933 4428 13957 4484
rect 14013 4428 14042 4484
rect 12092 4414 14042 4428
rect -216 3590 238 3596
rect -216 3572 244 3590
rect -216 3356 -179 3572
rect 197 3362 244 3572
rect 197 3356 238 3362
rect -216 3324 238 3356
rect 178 3107 410 3176
rect 178 2658 212 3107
rect 182 2571 212 2658
rect 348 2658 410 3107
rect 348 2571 404 2658
rect 182 2486 404 2571
rect 12248 675 13438 710
rect 12248 139 13270 675
rect 13406 139 13438 675
rect 12248 70 13438 139
rect 488 -823 3470 -784
rect 488 -833 530 -823
rect 3386 -833 3470 -823
rect 488 -949 524 -833
rect 3392 -949 3470 -833
rect 488 -959 530 -949
rect 3386 -959 3470 -949
rect 488 -996 3470 -959
rect 7026 -818 10310 -780
rect 7026 -828 7162 -818
rect 10178 -828 10310 -818
rect 7026 -944 7140 -828
rect 10200 -944 10310 -828
rect 7026 -954 7162 -944
rect 10178 -954 10310 -944
rect 7026 -976 10310 -954
rect 2580 -3778 2806 -3772
rect 2580 -3817 2814 -3778
rect 2580 -5073 2643 -3817
rect 2779 -5073 2814 -3817
rect 2580 -5114 2814 -5073
rect 5960 -3827 6146 -3764
rect 5960 -3841 5993 -3827
rect 6109 -3841 6146 -3827
rect 5960 -5017 5983 -3841
rect 6119 -5017 6146 -3841
rect 5960 -5031 5993 -5017
rect 6109 -5031 6146 -5017
rect 5960 -5098 6146 -5031
rect 9230 -3844 9428 -3804
rect 9230 -5100 9257 -3844
rect 9393 -5100 9428 -3844
rect 12582 -3842 12772 -3784
rect 12582 -3856 12616 -3842
rect 12732 -3856 12772 -3842
rect 12582 -5032 12606 -3856
rect 12742 -5032 12772 -3856
rect 12582 -5046 12616 -5032
rect 12732 -5046 12772 -5032
rect 12582 -5094 12772 -5046
rect 2580 -5128 2806 -5114
rect 9230 -5124 9428 -5100
rect 360 -7568 540 -7250
rect 350 -7724 540 -7568
rect 344 -8440 540 -7724
rect 2578 -7791 2798 -7680
rect 2578 -8407 2623 -7791
rect 2759 -7850 2798 -7791
rect 2759 -8407 2804 -7850
rect 344 -8442 534 -8440
rect 344 -8598 528 -8442
rect 2578 -8446 2804 -8407
rect 5956 -8089 6140 -7730
rect 5956 -8385 5982 -8089
rect 6118 -8385 6140 -8089
rect 2578 -8600 2798 -8446
rect 5956 -8604 6140 -8385
rect 6990 -7742 7168 -7186
rect 6990 -8422 7178 -7742
rect 6994 -8616 7178 -8422
rect 9226 -7850 9410 -7720
rect 9226 -7893 9430 -7850
rect 9226 -8349 9256 -7893
rect 9392 -8349 9430 -7893
rect 9226 -8394 9430 -8349
rect 12580 -7852 12764 -7726
rect 12580 -7917 12780 -7852
rect 12580 -8373 12608 -7917
rect 12744 -8373 12780 -7917
rect 13236 -7853 13452 -7822
rect 13236 -7863 13276 -7853
rect 13412 -7863 13452 -7853
rect 13236 -7979 13254 -7863
rect 13434 -7979 13452 -7863
rect 13236 -7989 13276 -7979
rect 13412 -7989 13452 -7979
rect 13236 -8010 13452 -7989
rect 9226 -8594 9410 -8394
rect 12580 -8438 12780 -8373
rect 12580 -8600 12764 -8438
<< via2 >>
rect 13739 5229 13875 5605
rect 13637 4428 13693 4484
rect 13717 4428 13773 4484
rect 13797 4428 13853 4484
rect 13877 4428 13933 4484
rect 13957 4428 14013 4484
rect -179 3356 197 3572
rect 212 2571 348 3107
rect 13270 139 13406 675
rect 530 -833 3386 -823
rect 530 -949 3386 -833
rect 530 -959 3386 -949
rect 7162 -828 10178 -818
rect 7162 -944 10178 -828
rect 7162 -954 10178 -944
rect 2643 -3843 2779 -3817
rect 2643 -5047 2653 -3843
rect 2653 -5047 2769 -3843
rect 2769 -5047 2779 -3843
rect 2643 -5073 2779 -5047
rect 5983 -5017 5993 -3841
rect 5993 -5017 6109 -3841
rect 6109 -5017 6119 -3841
rect 9257 -3870 9393 -3844
rect 9257 -5074 9267 -3870
rect 9267 -5074 9383 -3870
rect 9383 -5074 9393 -3870
rect 9257 -5100 9393 -5074
rect 12606 -5032 12616 -3856
rect 12616 -5032 12732 -3856
rect 12732 -5032 12742 -3856
rect 2623 -8407 2759 -7791
rect 5982 -8385 6118 -8089
rect 9256 -8349 9392 -7893
rect 12608 -8373 12744 -7917
rect 13276 -7863 13412 -7853
rect 13276 -7979 13412 -7863
rect 13276 -7989 13412 -7979
<< metal3 >>
rect -1616 11272 -598 11276
rect -1618 11232 -598 11272
rect -1618 11008 -1572 11232
rect -788 11008 -598 11232
rect -1618 10976 -598 11008
rect -1616 10968 -598 10976
rect -1612 10872 -800 10874
rect -1612 10870 -586 10872
rect -346 10870 4754 10876
rect -1612 10804 4754 10870
rect -1612 10462 -772 10804
rect -820 10180 -772 10462
rect -628 10799 4754 10804
rect -628 10575 3677 10799
rect 4701 10575 4754 10799
rect -628 10448 4754 10575
rect -628 10180 -586 10448
rect -820 10112 -586 10180
rect 13592 5666 13908 5684
rect 13592 5609 14204 5666
rect 13592 5225 13735 5609
rect 13879 5225 14204 5609
rect 13592 5202 14204 5225
rect 13592 5174 13908 5202
rect 13182 4484 14200 4560
rect 13182 4428 13637 4484
rect 13693 4428 13717 4484
rect 13773 4428 13797 4484
rect 13853 4428 13877 4484
rect 13933 4428 13957 4484
rect 14013 4428 14200 4484
rect 13182 4364 14200 4428
rect -216 3572 238 3596
rect -216 3356 -179 3572
rect 197 3356 238 3572
rect -216 3324 238 3356
rect -206 -370 6 3324
rect 182 3107 394 3176
rect 182 2571 212 3107
rect 348 2571 394 3107
rect 182 2 394 2571
rect 13462 716 14196 722
rect 12884 710 14196 716
rect 12248 679 14196 710
rect 12248 135 13266 679
rect 13410 135 14196 679
rect 12248 70 14196 135
rect 12884 68 14196 70
rect 13462 62 14196 68
rect 182 -210 8618 2
rect -206 -582 2008 -370
rect 1450 -784 1998 -582
rect 8212 -780 8618 -210
rect 488 -823 3470 -784
rect 488 -959 530 -823
rect 3386 -959 3470 -823
rect 488 -996 3470 -959
rect 7026 -818 10310 -780
rect 7026 -954 7162 -818
rect 10178 -954 10310 -818
rect 7026 -976 10310 -954
rect -1266 -2687 -1042 -2628
rect -1266 -2915 -1235 -2687
rect -1267 -3141 -1235 -2915
rect -1266 -3471 -1235 -3141
rect -1091 -2915 -1042 -2687
rect -1091 -3141 10085 -2915
rect -1091 -3471 -1042 -3141
rect -1266 -3536 -1042 -3471
rect 2580 -3778 2806 -3772
rect 2580 -3817 2814 -3778
rect 2580 -5073 2643 -3817
rect 2779 -5073 2814 -3817
rect 2580 -5114 2814 -5073
rect 5960 -3837 6146 -3764
rect 5960 -3841 6019 -3837
rect 6083 -3841 6146 -3837
rect 5960 -5017 5983 -3841
rect 6119 -5017 6146 -3841
rect 5960 -5021 6019 -5017
rect 6083 -5021 6146 -5017
rect 5960 -5098 6146 -5021
rect 9230 -3844 9428 -3804
rect 9230 -3880 9257 -3844
rect 9393 -3880 9428 -3844
rect 9230 -5064 9253 -3880
rect 9397 -5064 9428 -3880
rect 9230 -5100 9257 -5064
rect 9393 -5100 9428 -5064
rect 12582 -3852 12772 -3784
rect 12582 -5036 12602 -3852
rect 12746 -5036 12772 -3852
rect 12582 -5094 12772 -5036
rect 2580 -5128 2806 -5114
rect 9230 -5124 9428 -5100
rect 13672 -6216 13952 -6138
rect 13672 -6246 13728 -6216
rect 3211 -6404 13728 -6246
rect 9726 -6426 13728 -6404
rect 13672 -6520 13728 -6426
rect 13872 -6520 13952 -6216
rect 13672 -6614 13952 -6520
rect 2586 -7787 2802 -7686
rect 2586 -8411 2619 -7787
rect 2763 -7850 2802 -7787
rect 13236 -7849 13452 -7822
rect 2763 -8411 2804 -7850
rect 9228 -7889 9430 -7850
rect 2586 -8446 2804 -8411
rect 5956 -8085 6136 -8028
rect 5956 -8389 5978 -8085
rect 6122 -8389 6136 -8085
rect 5956 -8434 6136 -8389
rect 9228 -8353 9252 -7889
rect 9396 -8353 9430 -7889
rect 9228 -8394 9430 -8353
rect 12582 -7913 12780 -7852
rect 12582 -8377 12604 -7913
rect 12748 -8377 12780 -7913
rect 13236 -7993 13272 -7849
rect 13416 -7993 13452 -7849
rect 13236 -8010 13452 -7993
rect 12582 -8438 12780 -8377
<< via3 >>
rect -1572 11008 -788 11232
rect -772 10180 -628 10804
rect 3677 10575 4701 10799
rect 13735 5605 13879 5609
rect 13735 5229 13739 5605
rect 13739 5229 13875 5605
rect 13875 5229 13879 5605
rect 13735 5225 13879 5229
rect 13266 675 13410 679
rect 13266 139 13270 675
rect 13270 139 13406 675
rect 13406 139 13410 675
rect 13266 135 13410 139
rect -1235 -3471 -1091 -2687
rect 2679 -3917 2743 -3853
rect 2679 -3997 2743 -3933
rect 2679 -4077 2743 -4013
rect 2679 -4157 2743 -4093
rect 2679 -4237 2743 -4173
rect 2679 -4317 2743 -4253
rect 2679 -4397 2743 -4333
rect 2679 -4477 2743 -4413
rect 2679 -4557 2743 -4493
rect 2679 -4637 2743 -4573
rect 2679 -4717 2743 -4653
rect 2679 -4797 2743 -4733
rect 2679 -4877 2743 -4813
rect 2679 -4957 2743 -4893
rect 2679 -5037 2743 -4973
rect 6019 -3841 6083 -3837
rect 6019 -3901 6083 -3841
rect 6019 -3981 6083 -3917
rect 6019 -4061 6083 -3997
rect 6019 -4141 6083 -4077
rect 6019 -4221 6083 -4157
rect 6019 -4301 6083 -4237
rect 6019 -4381 6083 -4317
rect 6019 -4461 6083 -4397
rect 6019 -4541 6083 -4477
rect 6019 -4621 6083 -4557
rect 6019 -4701 6083 -4637
rect 6019 -4781 6083 -4717
rect 6019 -4861 6083 -4797
rect 6019 -4941 6083 -4877
rect 6019 -5017 6083 -4957
rect 6019 -5021 6083 -5017
rect 9253 -5064 9257 -3880
rect 9257 -5064 9393 -3880
rect 9393 -5064 9397 -3880
rect 12602 -3856 12746 -3852
rect 12602 -5032 12606 -3856
rect 12606 -5032 12742 -3856
rect 12742 -5032 12746 -3856
rect 12602 -5036 12746 -5032
rect 13728 -6520 13872 -6216
rect 2619 -7791 2763 -7787
rect 2619 -8407 2623 -7791
rect 2623 -8407 2759 -7791
rect 2759 -8407 2763 -7791
rect 2619 -8411 2763 -8407
rect 5978 -8089 6122 -8085
rect 5978 -8385 5982 -8089
rect 5982 -8385 6118 -8089
rect 6118 -8385 6122 -8089
rect 5978 -8389 6122 -8385
rect 9252 -7893 9396 -7889
rect 9252 -8349 9256 -7893
rect 9256 -8349 9392 -7893
rect 9392 -8349 9396 -7893
rect 9252 -8353 9396 -8349
rect 12604 -7917 12748 -7913
rect 12604 -8373 12608 -7917
rect 12608 -8373 12744 -7917
rect 12744 -8373 12748 -7917
rect 12604 -8377 12748 -8373
rect 13272 -7853 13416 -7849
rect 13272 -7989 13276 -7853
rect 13276 -7989 13412 -7853
rect 13412 -7989 13416 -7853
rect 13272 -7993 13416 -7989
<< metal4 >>
rect 1216 11260 2504 11274
rect -1612 11232 2508 11260
rect -1612 11008 -1572 11232
rect -788 11008 2508 11232
rect -1612 10968 2508 11008
rect -1262 10944 2504 10968
rect -1262 -2687 -1038 10944
rect -1262 -3471 -1235 -2687
rect -1091 -3471 -1038 -2687
rect -1262 -8030 -1038 -3471
rect -814 10804 -590 10866
rect 1216 10846 2504 10944
rect 1216 10842 2478 10846
rect -814 10180 -772 10804
rect -628 10180 -590 10804
rect -814 -8006 -590 10180
rect 1284 9978 2478 10842
rect 3570 10799 4764 10866
rect 3570 10575 3677 10799
rect 4701 10575 4764 10799
rect 3570 9912 4764 10575
rect 13246 679 13446 10132
rect 13700 5666 13900 10132
rect 13614 5609 14204 5666
rect 13614 5225 13735 5609
rect 13879 5225 14204 5609
rect 13614 5202 14204 5225
rect 13246 135 13266 679
rect 13410 135 13446 679
rect 2580 -3778 2806 -3772
rect 2580 -3853 2814 -3778
rect 2580 -3917 2679 -3853
rect 2743 -3917 2814 -3853
rect 2580 -3933 2814 -3917
rect 2580 -3997 2679 -3933
rect 2743 -3997 2814 -3933
rect 2580 -4013 2814 -3997
rect 2580 -4077 2679 -4013
rect 2743 -4077 2814 -4013
rect 2580 -4093 2814 -4077
rect 2580 -4157 2679 -4093
rect 2743 -4157 2814 -4093
rect 2580 -4173 2814 -4157
rect 2580 -4237 2679 -4173
rect 2743 -4237 2814 -4173
rect 2580 -4253 2814 -4237
rect 2580 -4317 2679 -4253
rect 2743 -4317 2814 -4253
rect 2580 -4333 2814 -4317
rect 2580 -4397 2679 -4333
rect 2743 -4397 2814 -4333
rect 2580 -4413 2814 -4397
rect 2580 -4477 2679 -4413
rect 2743 -4477 2814 -4413
rect 2580 -4493 2814 -4477
rect 2580 -4557 2679 -4493
rect 2743 -4557 2814 -4493
rect 2580 -4573 2814 -4557
rect 2580 -4637 2679 -4573
rect 2743 -4637 2814 -4573
rect 2580 -4653 2814 -4637
rect 2580 -4717 2679 -4653
rect 2743 -4717 2814 -4653
rect 2580 -4733 2814 -4717
rect 2580 -4797 2679 -4733
rect 2743 -4797 2814 -4733
rect 2580 -4813 2814 -4797
rect 2580 -4877 2679 -4813
rect 2743 -4877 2814 -4813
rect 2580 -4893 2814 -4877
rect 2580 -4957 2679 -4893
rect 2743 -4957 2814 -4893
rect 2580 -4973 2814 -4957
rect 2580 -5037 2679 -4973
rect 2743 -5037 2814 -4973
rect 2580 -5114 2814 -5037
rect 5960 -3837 6146 -3764
rect 5960 -3901 6019 -3837
rect 6083 -3901 6146 -3837
rect 5960 -3917 6146 -3901
rect 5960 -3981 6019 -3917
rect 6083 -3981 6146 -3917
rect 5960 -3997 6146 -3981
rect 5960 -4061 6019 -3997
rect 6083 -4061 6146 -3997
rect 5960 -4077 6146 -4061
rect 5960 -4141 6019 -4077
rect 6083 -4141 6146 -4077
rect 5960 -4157 6146 -4141
rect 5960 -4221 6019 -4157
rect 6083 -4221 6146 -4157
rect 5960 -4237 6146 -4221
rect 5960 -4301 6019 -4237
rect 6083 -4301 6146 -4237
rect 5960 -4317 6146 -4301
rect 5960 -4381 6019 -4317
rect 6083 -4381 6146 -4317
rect 5960 -4397 6146 -4381
rect 5960 -4461 6019 -4397
rect 6083 -4461 6146 -4397
rect 5960 -4477 6146 -4461
rect 5960 -4541 6019 -4477
rect 6083 -4541 6146 -4477
rect 5960 -4557 6146 -4541
rect 5960 -4621 6019 -4557
rect 6083 -4621 6146 -4557
rect 5960 -4637 6146 -4621
rect 5960 -4701 6019 -4637
rect 6083 -4701 6146 -4637
rect 5960 -4717 6146 -4701
rect 5960 -4781 6019 -4717
rect 6083 -4781 6146 -4717
rect 5960 -4797 6146 -4781
rect 5960 -4861 6019 -4797
rect 6083 -4861 6146 -4797
rect 5960 -4877 6146 -4861
rect 5960 -4941 6019 -4877
rect 6083 -4941 6146 -4877
rect 5960 -4957 6146 -4941
rect 5960 -5021 6019 -4957
rect 6083 -5021 6146 -4957
rect 5960 -5098 6146 -5021
rect 9230 -3880 9428 -3804
rect 9230 -5064 9253 -3880
rect 9397 -5064 9428 -3880
rect 12582 -3852 12772 -3784
rect 12582 -4912 12602 -3852
rect 2580 -5128 2810 -5114
rect 2588 -7686 2810 -5128
rect 2586 -7787 2810 -7686
rect 2586 -8411 2619 -7787
rect 2763 -8411 2810 -7787
rect 2586 -8440 2810 -8411
rect 5960 -8085 6140 -5098
rect 9230 -5124 9428 -5064
rect 12572 -5036 12602 -4912
rect 12746 -4912 12772 -3852
rect 12746 -5036 12774 -4912
rect 5960 -8389 5978 -8085
rect 6122 -8389 6140 -8085
rect 2586 -8446 2802 -8440
rect 5960 -8442 6140 -8389
rect 9238 -7889 9424 -5124
rect 9238 -8353 9252 -7889
rect 9396 -8353 9424 -7889
rect 9238 -8406 9424 -8353
rect 12572 -7852 12774 -5036
rect 13246 -7822 13446 135
rect 13700 -6138 13900 5202
rect 13672 -6216 13952 -6138
rect 13672 -6520 13728 -6216
rect 13872 -6520 13952 -6216
rect 13672 -6614 13952 -6520
rect 13236 -7849 13452 -7822
rect 12572 -7913 12780 -7852
rect 12572 -8377 12604 -7913
rect 12748 -8377 12780 -7913
rect 13236 -7993 13272 -7849
rect 13416 -7993 13452 -7849
rect 13700 -7974 13900 -6614
rect 13236 -8010 13452 -7993
rect 13246 -8012 13446 -8010
rect 12572 -8434 12780 -8377
rect 12582 -8438 12780 -8434
use comparator_top  comparator_top_0
timestamp 1694079970
transform 1 0 800 0 1 265
box -1081 -265 11765 10234
use EF_AMUX21m  EF_AMUX21m_1
timestamp 1694079970
transform 1 0 -3364 0 1 -7208
box 1380 -890 10345 6424
use EF_AMUX21m  EF_AMUX21m_2
timestamp 1694079970
transform 1 0 3262 0 1 -7212
box 1380 -890 10345 6424
<< labels >>
flabel metal3 s -1612 10462 -800 10874 0 FreeSans 6104 0 0 0 VSS
port 1 nsew
flabel metal3 s -1616 10968 -598 11276 0 FreeSans 6104 0 0 0 VDD
port 2 nsew
flabel metal2 s 344 -8598 528 -7724 0 FreeSans 6104 0 0 0 SELA
port 3 nsew
flabel metal2 s 5956 -8604 6140 -7730 0 FreeSans 6104 0 0 0 A2
port 4 nsew
flabel metal2 s 6994 -8616 7178 -7742 0 FreeSans 6104 0 0 0 SELB
port 5 nsew
flabel metal2 s 9226 -8594 9410 -7720 0 FreeSans 6104 0 0 0 B1
port 6 nsew
flabel metal2 s 12580 -8600 12764 -7726 0 FreeSans 6104 0 0 0 B2
port 7 nsew
flabel metal3 s 13182 4364 14200 4560 0 FreeSans 6104 0 0 0 VO
port 8 nsew
flabel metal2 s 2578 -8600 2798 -7680 0 FreeSans 4883 0 0 0 A1
port 9 nsew
flabel metal3 s 13462 62 14196 722 0 FreeSans 3906 0 0 0 DVSS
port 10 nsew
flabel metal4 s 13614 5202 14204 5666 0 FreeSans 1000 0 0 0 DVDD
port 11 nsew
<< end >>
