magic
tech sky130A
magscale 1 2
timestamp 1699211738
<< checkpaint >>
rect -3868 -15068 15066 14280
<< metal1 >>
rect 1908 -851 2708 -822
rect 1908 -903 1931 -851
rect 1983 -903 1995 -851
rect 2047 -903 2059 -851
rect 2111 -903 2123 -851
rect 2175 -903 2187 -851
rect 2239 -903 2251 -851
rect 2303 -903 2315 -851
rect 2367 -903 2379 -851
rect 2431 -903 2443 -851
rect 2495 -903 2507 -851
rect 2559 -903 2571 -851
rect 2623 -903 2635 -851
rect 2687 -903 2708 -851
rect 1908 -932 2708 -903
rect 8384 -848 9204 -818
rect 8384 -900 8425 -848
rect 8477 -900 8489 -848
rect 8541 -900 8553 -848
rect 8605 -900 8617 -848
rect 8669 -900 8681 -848
rect 8733 -900 8745 -848
rect 8797 -900 8809 -848
rect 8861 -900 8873 -848
rect 8925 -900 8937 -848
rect 8989 -900 9001 -848
rect 9053 -900 9065 -848
rect 9117 -900 9129 -848
rect 9181 -900 9204 -848
rect 8384 -928 9204 -900
rect 1934 -9433 2040 -9390
rect 1934 -9485 1962 -9433
rect 2014 -9485 2040 -9433
rect 1934 -9497 2040 -9485
rect 1934 -9549 1962 -9497
rect 2014 -9549 2040 -9497
rect 1934 -9561 2040 -9549
rect 1934 -9613 1962 -9561
rect 2014 -9613 2040 -9561
rect 1934 -9625 2040 -9613
rect 1934 -9677 1962 -9625
rect 2014 -9677 2040 -9625
rect 1934 -9689 2040 -9677
rect 1934 -9741 1962 -9689
rect 2014 -9741 2040 -9689
rect 1934 -9753 2040 -9741
rect 1934 -9805 1962 -9753
rect 2014 -9805 2040 -9753
rect 1934 -9817 2040 -9805
rect 1934 -9869 1962 -9817
rect 2014 -9869 2040 -9817
rect 1934 -9881 2040 -9869
rect 1934 -9933 1962 -9881
rect 2014 -9933 2040 -9881
rect 1934 -9988 2040 -9933
rect 5332 -9449 5438 -9402
rect 5332 -9501 5358 -9449
rect 5410 -9501 5438 -9449
rect 5332 -9513 5438 -9501
rect 5332 -9565 5358 -9513
rect 5410 -9565 5438 -9513
rect 5332 -9577 5438 -9565
rect 5332 -9629 5358 -9577
rect 5410 -9629 5438 -9577
rect 5332 -9641 5438 -9629
rect 5332 -9693 5358 -9641
rect 5410 -9693 5438 -9641
rect 5332 -9705 5438 -9693
rect 5332 -9757 5358 -9705
rect 5410 -9757 5438 -9705
rect 5332 -9769 5438 -9757
rect 5332 -9821 5358 -9769
rect 5410 -9821 5438 -9769
rect 5332 -9833 5438 -9821
rect 5332 -9885 5358 -9833
rect 5410 -9885 5438 -9833
rect 5332 -9897 5438 -9885
rect 5332 -9949 5358 -9897
rect 5410 -9949 5438 -9897
rect 5332 -10000 5438 -9949
rect 8528 -9443 8634 -9394
rect 8528 -9495 8554 -9443
rect 8606 -9495 8634 -9443
rect 8528 -9507 8634 -9495
rect 8528 -9559 8554 -9507
rect 8606 -9559 8634 -9507
rect 8528 -9571 8634 -9559
rect 8528 -9623 8554 -9571
rect 8606 -9623 8634 -9571
rect 8528 -9635 8634 -9623
rect 8528 -9687 8554 -9635
rect 8606 -9687 8634 -9635
rect 8528 -9699 8634 -9687
rect 8528 -9751 8554 -9699
rect 8606 -9751 8634 -9699
rect 8528 -9763 8634 -9751
rect 8528 -9815 8554 -9763
rect 8606 -9815 8634 -9763
rect 8528 -9827 8634 -9815
rect 8528 -9879 8554 -9827
rect 8606 -9879 8634 -9827
rect 8528 -9891 8634 -9879
rect 8528 -9943 8554 -9891
rect 8606 -9943 8634 -9891
rect 8528 -9992 8634 -9943
rect 11930 -9445 12036 -9396
rect 11930 -9497 11960 -9445
rect 12012 -9497 12036 -9445
rect 11930 -9509 12036 -9497
rect 11930 -9561 11960 -9509
rect 12012 -9561 12036 -9509
rect 11930 -9573 12036 -9561
rect 11930 -9625 11960 -9573
rect 12012 -9625 12036 -9573
rect 11930 -9637 12036 -9625
rect 11930 -9689 11960 -9637
rect 12012 -9689 12036 -9637
rect 11930 -9701 12036 -9689
rect 11930 -9753 11960 -9701
rect 12012 -9753 12036 -9701
rect 11930 -9765 12036 -9753
rect 11930 -9817 11960 -9765
rect 12012 -9817 12036 -9765
rect 11930 -9829 12036 -9817
rect 11930 -9881 11960 -9829
rect 12012 -9881 12036 -9829
rect 11930 -9893 12036 -9881
rect 11930 -9945 11960 -9893
rect 12012 -9945 12036 -9893
rect 11930 -9994 12036 -9945
rect -809 -13000 3389 -12774
rect 4955 -12794 12595 -12770
rect 4955 -12974 12441 -12794
rect 12557 -12974 12595 -12794
rect 4955 -12996 12595 -12974
<< via1 >>
rect 1931 -903 1983 -851
rect 1995 -903 2047 -851
rect 2059 -903 2111 -851
rect 2123 -903 2175 -851
rect 2187 -903 2239 -851
rect 2251 -903 2303 -851
rect 2315 -903 2367 -851
rect 2379 -903 2431 -851
rect 2443 -903 2495 -851
rect 2507 -903 2559 -851
rect 2571 -903 2623 -851
rect 2635 -903 2687 -851
rect 8425 -900 8477 -848
rect 8489 -900 8541 -848
rect 8553 -900 8605 -848
rect 8617 -900 8669 -848
rect 8681 -900 8733 -848
rect 8745 -900 8797 -848
rect 8809 -900 8861 -848
rect 8873 -900 8925 -848
rect 8937 -900 8989 -848
rect 9001 -900 9053 -848
rect 9065 -900 9117 -848
rect 9129 -900 9181 -848
rect 1962 -9485 2014 -9433
rect 1962 -9549 2014 -9497
rect 1962 -9613 2014 -9561
rect 1962 -9677 2014 -9625
rect 1962 -9741 2014 -9689
rect 1962 -9805 2014 -9753
rect 1962 -9869 2014 -9817
rect 1962 -9933 2014 -9881
rect 5358 -9501 5410 -9449
rect 5358 -9565 5410 -9513
rect 5358 -9629 5410 -9577
rect 5358 -9693 5410 -9641
rect 5358 -9757 5410 -9705
rect 5358 -9821 5410 -9769
rect 5358 -9885 5410 -9833
rect 5358 -9949 5410 -9897
rect 8554 -9495 8606 -9443
rect 8554 -9559 8606 -9507
rect 8554 -9623 8606 -9571
rect 8554 -9687 8606 -9635
rect 8554 -9751 8606 -9699
rect 8554 -9815 8606 -9763
rect 8554 -9879 8606 -9827
rect 8554 -9943 8606 -9891
rect 11960 -9497 12012 -9445
rect 11960 -9561 12012 -9509
rect 11960 -9625 12012 -9573
rect 11960 -9689 12012 -9637
rect 11960 -9753 12012 -9701
rect 11960 -9817 12012 -9765
rect 11960 -9881 12012 -9829
rect 11960 -9945 12012 -9893
rect 12441 -12974 12557 -12794
<< metal2 >>
rect -1404 949 -1204 1004
rect -1404 653 -1382 949
rect -1246 899 -1204 949
rect -1246 739 4640 899
rect -1246 653 -1204 739
rect -1404 600 -1204 653
rect 1908 -849 2708 -822
rect 1908 -851 1961 -849
rect 2017 -851 2041 -849
rect 2097 -851 2121 -849
rect 2177 -851 2201 -849
rect 2257 -851 2281 -849
rect 2337 -851 2361 -849
rect 2417 -851 2441 -849
rect 2497 -851 2521 -849
rect 2577 -851 2601 -849
rect 2657 -851 2708 -849
rect 1908 -903 1931 -851
rect 2111 -903 2121 -851
rect 2177 -903 2187 -851
rect 2431 -903 2441 -851
rect 2497 -903 2507 -851
rect 2687 -903 2708 -851
rect 1908 -905 1961 -903
rect 2017 -905 2041 -903
rect 2097 -905 2121 -903
rect 2177 -905 2201 -903
rect 2257 -905 2281 -903
rect 2337 -905 2361 -903
rect 2417 -905 2441 -903
rect 2497 -905 2521 -903
rect 2577 -905 2601 -903
rect 2657 -905 2708 -903
rect 1908 -932 2708 -905
rect 8384 -846 9204 -818
rect 8384 -902 8415 -846
rect 8471 -848 8495 -846
rect 8551 -848 8575 -846
rect 8631 -848 8655 -846
rect 8711 -848 8735 -846
rect 8791 -848 8815 -846
rect 8871 -848 8895 -846
rect 8951 -848 8975 -846
rect 9031 -848 9055 -846
rect 9111 -848 9135 -846
rect 8477 -900 8489 -848
rect 8551 -900 8553 -848
rect 8733 -900 8735 -848
rect 8797 -900 8809 -848
rect 8871 -900 8873 -848
rect 9053 -900 9055 -848
rect 9117 -900 9129 -848
rect 8471 -902 8495 -900
rect 8551 -902 8575 -900
rect 8631 -902 8655 -900
rect 8711 -902 8735 -900
rect 8791 -902 8815 -900
rect 8871 -902 8895 -900
rect 8951 -902 8975 -900
rect 9031 -902 9055 -900
rect 9111 -902 9135 -900
rect 9191 -902 9204 -846
rect 8384 -928 9204 -902
rect 1934 -9415 2040 -9390
rect 1934 -9471 1960 -9415
rect 2016 -9471 2040 -9415
rect 1934 -9485 1962 -9471
rect 2014 -9485 2040 -9471
rect 1934 -9495 2040 -9485
rect 1934 -9551 1960 -9495
rect 2016 -9551 2040 -9495
rect 1934 -9561 2040 -9551
rect 1934 -9575 1962 -9561
rect 2014 -9575 2040 -9561
rect 1934 -9631 1960 -9575
rect 2016 -9631 2040 -9575
rect 1934 -9655 1962 -9631
rect 2014 -9655 2040 -9631
rect 1934 -9711 1960 -9655
rect 2016 -9711 2040 -9655
rect 1934 -9735 1962 -9711
rect 2014 -9735 2040 -9711
rect 1934 -9791 1960 -9735
rect 2016 -9791 2040 -9735
rect 1934 -9805 1962 -9791
rect 2014 -9805 2040 -9791
rect 1934 -9815 2040 -9805
rect 1934 -9871 1960 -9815
rect 2016 -9871 2040 -9815
rect 1934 -9881 2040 -9871
rect 1934 -9895 1962 -9881
rect 2014 -9895 2040 -9881
rect 1934 -9951 1960 -9895
rect 2016 -9951 2040 -9895
rect 1934 -9988 2040 -9951
rect 5332 -9431 5438 -9402
rect 5332 -9487 5356 -9431
rect 5412 -9487 5438 -9431
rect 5332 -9501 5358 -9487
rect 5410 -9501 5438 -9487
rect 5332 -9511 5438 -9501
rect 5332 -9567 5356 -9511
rect 5412 -9567 5438 -9511
rect 5332 -9577 5438 -9567
rect 5332 -9591 5358 -9577
rect 5410 -9591 5438 -9577
rect 5332 -9647 5356 -9591
rect 5412 -9647 5438 -9591
rect 5332 -9671 5358 -9647
rect 5410 -9671 5438 -9647
rect 5332 -9727 5356 -9671
rect 5412 -9727 5438 -9671
rect 5332 -9751 5358 -9727
rect 5410 -9751 5438 -9727
rect 5332 -9807 5356 -9751
rect 5412 -9807 5438 -9751
rect 5332 -9821 5358 -9807
rect 5410 -9821 5438 -9807
rect 5332 -9831 5438 -9821
rect 5332 -9887 5356 -9831
rect 5412 -9887 5438 -9831
rect 5332 -9897 5438 -9887
rect 5332 -9911 5358 -9897
rect 5410 -9911 5438 -9897
rect 5332 -9967 5356 -9911
rect 5412 -9967 5438 -9911
rect 5332 -10000 5438 -9967
rect 8528 -9425 8634 -9394
rect 8528 -9481 8552 -9425
rect 8608 -9481 8634 -9425
rect 8528 -9495 8554 -9481
rect 8606 -9495 8634 -9481
rect 8528 -9505 8634 -9495
rect 8528 -9561 8552 -9505
rect 8608 -9561 8634 -9505
rect 8528 -9571 8634 -9561
rect 8528 -9585 8554 -9571
rect 8606 -9585 8634 -9571
rect 8528 -9641 8552 -9585
rect 8608 -9641 8634 -9585
rect 8528 -9665 8554 -9641
rect 8606 -9665 8634 -9641
rect 8528 -9721 8552 -9665
rect 8608 -9721 8634 -9665
rect 8528 -9745 8554 -9721
rect 8606 -9745 8634 -9721
rect 8528 -9801 8552 -9745
rect 8608 -9801 8634 -9745
rect 8528 -9815 8554 -9801
rect 8606 -9815 8634 -9801
rect 8528 -9825 8634 -9815
rect 8528 -9881 8552 -9825
rect 8608 -9881 8634 -9825
rect 8528 -9891 8634 -9881
rect 8528 -9905 8554 -9891
rect 8606 -9905 8634 -9891
rect 8528 -9961 8552 -9905
rect 8608 -9961 8634 -9905
rect 8528 -9992 8634 -9961
rect 11930 -9427 12036 -9396
rect 11930 -9483 11958 -9427
rect 12014 -9483 12036 -9427
rect 11930 -9497 11960 -9483
rect 12012 -9497 12036 -9483
rect 11930 -9507 12036 -9497
rect 11930 -9563 11958 -9507
rect 12014 -9563 12036 -9507
rect 11930 -9573 12036 -9563
rect 11930 -9587 11960 -9573
rect 12012 -9587 12036 -9573
rect 11930 -9643 11958 -9587
rect 12014 -9643 12036 -9587
rect 11930 -9667 11960 -9643
rect 12012 -9667 12036 -9643
rect 11930 -9723 11958 -9667
rect 12014 -9723 12036 -9667
rect 11930 -9747 11960 -9723
rect 12012 -9747 12036 -9723
rect 11930 -9803 11958 -9747
rect 12014 -9803 12036 -9747
rect 11930 -9817 11960 -9803
rect 12012 -9817 12036 -9803
rect 11930 -9827 12036 -9817
rect 11930 -9883 11958 -9827
rect 12014 -9883 12036 -9827
rect 11930 -9893 12036 -9883
rect 11930 -9907 11960 -9893
rect 12012 -9907 12036 -9893
rect 11930 -9963 11958 -9907
rect 12014 -9963 12036 -9907
rect 11930 -9994 12036 -9963
rect -395 -13184 -265 -12181
rect -400 -13788 -264 -13184
rect 5334 -13198 5446 -13192
rect 1932 -13230 2044 -13198
rect 1932 -13286 1953 -13230
rect 2009 -13286 2044 -13230
rect 1932 -13310 2044 -13286
rect 1932 -13366 1953 -13310
rect 2009 -13366 2044 -13310
rect 1932 -13390 2044 -13366
rect 1932 -13446 1953 -13390
rect 2009 -13446 2044 -13390
rect 1932 -13470 2044 -13446
rect 1932 -13526 1953 -13470
rect 2009 -13526 2044 -13470
rect 1932 -13550 2044 -13526
rect 1932 -13606 1953 -13550
rect 2009 -13606 2044 -13550
rect 1932 -13630 2044 -13606
rect 1932 -13686 1953 -13630
rect 2009 -13686 2044 -13630
rect 1932 -13710 2044 -13686
rect 1932 -13766 1953 -13710
rect 2009 -13766 2044 -13710
rect -395 -13801 -265 -13788
rect 1932 -13804 2044 -13766
rect 5332 -13234 5446 -13198
rect 6203 -13200 6333 -12233
rect 12394 -12794 12600 -12766
rect 12394 -12816 12441 -12794
rect 12557 -12816 12600 -12794
rect 12394 -12952 12431 -12816
rect 12567 -12952 12600 -12816
rect 12394 -12974 12441 -12952
rect 12557 -12974 12600 -12952
rect 12394 -12996 12600 -12974
rect 5332 -13290 5355 -13234
rect 5411 -13290 5446 -13234
rect 5332 -13314 5446 -13290
rect 5332 -13370 5355 -13314
rect 5411 -13370 5446 -13314
rect 5332 -13394 5446 -13370
rect 5332 -13450 5355 -13394
rect 5411 -13450 5446 -13394
rect 5332 -13474 5446 -13450
rect 5332 -13530 5355 -13474
rect 5411 -13530 5446 -13474
rect 5332 -13554 5446 -13530
rect 5332 -13610 5355 -13554
rect 5411 -13610 5446 -13554
rect 5332 -13634 5446 -13610
rect 5332 -13690 5355 -13634
rect 5411 -13690 5446 -13634
rect 5332 -13714 5446 -13690
rect 5332 -13770 5355 -13714
rect 5411 -13770 5446 -13714
rect 5332 -13800 5446 -13770
rect 5334 -13802 5446 -13800
rect 6200 -13808 6338 -13200
rect 8526 -13230 8636 -13190
rect 8526 -13286 8553 -13230
rect 8609 -13286 8636 -13230
rect 8526 -13310 8636 -13286
rect 8526 -13366 8553 -13310
rect 8609 -13366 8636 -13310
rect 8526 -13390 8636 -13366
rect 8526 -13446 8553 -13390
rect 8609 -13446 8636 -13390
rect 8526 -13470 8636 -13446
rect 8526 -13526 8553 -13470
rect 8609 -13526 8636 -13470
rect 8526 -13550 8636 -13526
rect 8526 -13606 8553 -13550
rect 8609 -13606 8636 -13550
rect 8526 -13630 8636 -13606
rect 8526 -13686 8553 -13630
rect 8609 -13686 8636 -13630
rect 8526 -13710 8636 -13686
rect 8526 -13766 8553 -13710
rect 8609 -13766 8636 -13710
rect 8526 -13798 8636 -13766
rect 11932 -13224 12038 -13196
rect 11932 -13280 11962 -13224
rect 12018 -13280 12038 -13224
rect 11932 -13304 12038 -13280
rect 11932 -13360 11962 -13304
rect 12018 -13360 12038 -13304
rect 11932 -13384 12038 -13360
rect 11932 -13440 11962 -13384
rect 12018 -13440 12038 -13384
rect 11932 -13464 12038 -13440
rect 11932 -13520 11962 -13464
rect 12018 -13520 12038 -13464
rect 11932 -13544 12038 -13520
rect 11932 -13600 11962 -13544
rect 12018 -13600 12038 -13544
rect 11932 -13624 12038 -13600
rect 11932 -13680 11962 -13624
rect 12018 -13680 12038 -13624
rect 11932 -13704 12038 -13680
rect 11932 -13760 11962 -13704
rect 12018 -13760 12038 -13704
rect 11932 -13798 12038 -13760
rect 11938 -13800 12032 -13798
<< via2 >>
rect -1382 653 -1246 949
rect 1961 -851 2017 -849
rect 2041 -851 2097 -849
rect 2121 -851 2177 -849
rect 2201 -851 2257 -849
rect 2281 -851 2337 -849
rect 2361 -851 2417 -849
rect 2441 -851 2497 -849
rect 2521 -851 2577 -849
rect 2601 -851 2657 -849
rect 1961 -903 1983 -851
rect 1983 -903 1995 -851
rect 1995 -903 2017 -851
rect 2041 -903 2047 -851
rect 2047 -903 2059 -851
rect 2059 -903 2097 -851
rect 2121 -903 2123 -851
rect 2123 -903 2175 -851
rect 2175 -903 2177 -851
rect 2201 -903 2239 -851
rect 2239 -903 2251 -851
rect 2251 -903 2257 -851
rect 2281 -903 2303 -851
rect 2303 -903 2315 -851
rect 2315 -903 2337 -851
rect 2361 -903 2367 -851
rect 2367 -903 2379 -851
rect 2379 -903 2417 -851
rect 2441 -903 2443 -851
rect 2443 -903 2495 -851
rect 2495 -903 2497 -851
rect 2521 -903 2559 -851
rect 2559 -903 2571 -851
rect 2571 -903 2577 -851
rect 2601 -903 2623 -851
rect 2623 -903 2635 -851
rect 2635 -903 2657 -851
rect 1961 -905 2017 -903
rect 2041 -905 2097 -903
rect 2121 -905 2177 -903
rect 2201 -905 2257 -903
rect 2281 -905 2337 -903
rect 2361 -905 2417 -903
rect 2441 -905 2497 -903
rect 2521 -905 2577 -903
rect 2601 -905 2657 -903
rect 8415 -848 8471 -846
rect 8495 -848 8551 -846
rect 8575 -848 8631 -846
rect 8655 -848 8711 -846
rect 8735 -848 8791 -846
rect 8815 -848 8871 -846
rect 8895 -848 8951 -846
rect 8975 -848 9031 -846
rect 9055 -848 9111 -846
rect 9135 -848 9191 -846
rect 8415 -900 8425 -848
rect 8425 -900 8471 -848
rect 8495 -900 8541 -848
rect 8541 -900 8551 -848
rect 8575 -900 8605 -848
rect 8605 -900 8617 -848
rect 8617 -900 8631 -848
rect 8655 -900 8669 -848
rect 8669 -900 8681 -848
rect 8681 -900 8711 -848
rect 8735 -900 8745 -848
rect 8745 -900 8791 -848
rect 8815 -900 8861 -848
rect 8861 -900 8871 -848
rect 8895 -900 8925 -848
rect 8925 -900 8937 -848
rect 8937 -900 8951 -848
rect 8975 -900 8989 -848
rect 8989 -900 9001 -848
rect 9001 -900 9031 -848
rect 9055 -900 9065 -848
rect 9065 -900 9111 -848
rect 9135 -900 9181 -848
rect 9181 -900 9191 -848
rect 8415 -902 8471 -900
rect 8495 -902 8551 -900
rect 8575 -902 8631 -900
rect 8655 -902 8711 -900
rect 8735 -902 8791 -900
rect 8815 -902 8871 -900
rect 8895 -902 8951 -900
rect 8975 -902 9031 -900
rect 9055 -902 9111 -900
rect 9135 -902 9191 -900
rect 1960 -9433 2016 -9415
rect 1960 -9471 1962 -9433
rect 1962 -9471 2014 -9433
rect 2014 -9471 2016 -9433
rect 1960 -9497 2016 -9495
rect 1960 -9549 1962 -9497
rect 1962 -9549 2014 -9497
rect 2014 -9549 2016 -9497
rect 1960 -9551 2016 -9549
rect 1960 -9613 1962 -9575
rect 1962 -9613 2014 -9575
rect 2014 -9613 2016 -9575
rect 1960 -9625 2016 -9613
rect 1960 -9631 1962 -9625
rect 1962 -9631 2014 -9625
rect 2014 -9631 2016 -9625
rect 1960 -9677 1962 -9655
rect 1962 -9677 2014 -9655
rect 2014 -9677 2016 -9655
rect 1960 -9689 2016 -9677
rect 1960 -9711 1962 -9689
rect 1962 -9711 2014 -9689
rect 2014 -9711 2016 -9689
rect 1960 -9741 1962 -9735
rect 1962 -9741 2014 -9735
rect 2014 -9741 2016 -9735
rect 1960 -9753 2016 -9741
rect 1960 -9791 1962 -9753
rect 1962 -9791 2014 -9753
rect 2014 -9791 2016 -9753
rect 1960 -9817 2016 -9815
rect 1960 -9869 1962 -9817
rect 1962 -9869 2014 -9817
rect 2014 -9869 2016 -9817
rect 1960 -9871 2016 -9869
rect 1960 -9933 1962 -9895
rect 1962 -9933 2014 -9895
rect 2014 -9933 2016 -9895
rect 1960 -9951 2016 -9933
rect 5356 -9449 5412 -9431
rect 5356 -9487 5358 -9449
rect 5358 -9487 5410 -9449
rect 5410 -9487 5412 -9449
rect 5356 -9513 5412 -9511
rect 5356 -9565 5358 -9513
rect 5358 -9565 5410 -9513
rect 5410 -9565 5412 -9513
rect 5356 -9567 5412 -9565
rect 5356 -9629 5358 -9591
rect 5358 -9629 5410 -9591
rect 5410 -9629 5412 -9591
rect 5356 -9641 5412 -9629
rect 5356 -9647 5358 -9641
rect 5358 -9647 5410 -9641
rect 5410 -9647 5412 -9641
rect 5356 -9693 5358 -9671
rect 5358 -9693 5410 -9671
rect 5410 -9693 5412 -9671
rect 5356 -9705 5412 -9693
rect 5356 -9727 5358 -9705
rect 5358 -9727 5410 -9705
rect 5410 -9727 5412 -9705
rect 5356 -9757 5358 -9751
rect 5358 -9757 5410 -9751
rect 5410 -9757 5412 -9751
rect 5356 -9769 5412 -9757
rect 5356 -9807 5358 -9769
rect 5358 -9807 5410 -9769
rect 5410 -9807 5412 -9769
rect 5356 -9833 5412 -9831
rect 5356 -9885 5358 -9833
rect 5358 -9885 5410 -9833
rect 5410 -9885 5412 -9833
rect 5356 -9887 5412 -9885
rect 5356 -9949 5358 -9911
rect 5358 -9949 5410 -9911
rect 5410 -9949 5412 -9911
rect 5356 -9967 5412 -9949
rect 8552 -9443 8608 -9425
rect 8552 -9481 8554 -9443
rect 8554 -9481 8606 -9443
rect 8606 -9481 8608 -9443
rect 8552 -9507 8608 -9505
rect 8552 -9559 8554 -9507
rect 8554 -9559 8606 -9507
rect 8606 -9559 8608 -9507
rect 8552 -9561 8608 -9559
rect 8552 -9623 8554 -9585
rect 8554 -9623 8606 -9585
rect 8606 -9623 8608 -9585
rect 8552 -9635 8608 -9623
rect 8552 -9641 8554 -9635
rect 8554 -9641 8606 -9635
rect 8606 -9641 8608 -9635
rect 8552 -9687 8554 -9665
rect 8554 -9687 8606 -9665
rect 8606 -9687 8608 -9665
rect 8552 -9699 8608 -9687
rect 8552 -9721 8554 -9699
rect 8554 -9721 8606 -9699
rect 8606 -9721 8608 -9699
rect 8552 -9751 8554 -9745
rect 8554 -9751 8606 -9745
rect 8606 -9751 8608 -9745
rect 8552 -9763 8608 -9751
rect 8552 -9801 8554 -9763
rect 8554 -9801 8606 -9763
rect 8606 -9801 8608 -9763
rect 8552 -9827 8608 -9825
rect 8552 -9879 8554 -9827
rect 8554 -9879 8606 -9827
rect 8606 -9879 8608 -9827
rect 8552 -9881 8608 -9879
rect 8552 -9943 8554 -9905
rect 8554 -9943 8606 -9905
rect 8606 -9943 8608 -9905
rect 8552 -9961 8608 -9943
rect 11958 -9445 12014 -9427
rect 11958 -9483 11960 -9445
rect 11960 -9483 12012 -9445
rect 12012 -9483 12014 -9445
rect 11958 -9509 12014 -9507
rect 11958 -9561 11960 -9509
rect 11960 -9561 12012 -9509
rect 12012 -9561 12014 -9509
rect 11958 -9563 12014 -9561
rect 11958 -9625 11960 -9587
rect 11960 -9625 12012 -9587
rect 12012 -9625 12014 -9587
rect 11958 -9637 12014 -9625
rect 11958 -9643 11960 -9637
rect 11960 -9643 12012 -9637
rect 12012 -9643 12014 -9637
rect 11958 -9689 11960 -9667
rect 11960 -9689 12012 -9667
rect 12012 -9689 12014 -9667
rect 11958 -9701 12014 -9689
rect 11958 -9723 11960 -9701
rect 11960 -9723 12012 -9701
rect 12012 -9723 12014 -9701
rect 11958 -9753 11960 -9747
rect 11960 -9753 12012 -9747
rect 12012 -9753 12014 -9747
rect 11958 -9765 12014 -9753
rect 11958 -9803 11960 -9765
rect 11960 -9803 12012 -9765
rect 12012 -9803 12014 -9765
rect 11958 -9829 12014 -9827
rect 11958 -9881 11960 -9829
rect 11960 -9881 12012 -9829
rect 12012 -9881 12014 -9829
rect 11958 -9883 12014 -9881
rect 11958 -9945 11960 -9907
rect 11960 -9945 12012 -9907
rect 12012 -9945 12014 -9907
rect 11958 -9963 12014 -9945
rect 1953 -13286 2009 -13230
rect 1953 -13366 2009 -13310
rect 1953 -13446 2009 -13390
rect 1953 -13526 2009 -13470
rect 1953 -13606 2009 -13550
rect 1953 -13686 2009 -13630
rect 1953 -13766 2009 -13710
rect 12431 -12952 12441 -12816
rect 12441 -12952 12557 -12816
rect 12557 -12952 12567 -12816
rect 5355 -13290 5411 -13234
rect 5355 -13370 5411 -13314
rect 5355 -13450 5411 -13394
rect 5355 -13530 5411 -13474
rect 5355 -13610 5411 -13554
rect 5355 -13690 5411 -13634
rect 5355 -13770 5411 -13714
rect 8553 -13286 8609 -13230
rect 8553 -13366 8609 -13310
rect 8553 -13446 8609 -13390
rect 8553 -13526 8609 -13470
rect 8553 -13606 8609 -13550
rect 8553 -13686 8609 -13630
rect 8553 -13766 8609 -13710
rect 11962 -13280 12018 -13224
rect 11962 -13360 12018 -13304
rect 11962 -13440 12018 -13384
rect 11962 -13520 12018 -13464
rect 11962 -13600 12018 -13544
rect 11962 -13680 12018 -13624
rect 11962 -13760 12018 -13704
<< metal3 >>
rect -1678 11483 -628 11504
rect -1678 11259 -1654 11483
rect -1510 11259 -628 11483
rect -1678 11240 -628 11259
rect 11502 6847 13806 6888
rect 11502 6383 12707 6847
rect 12851 6383 13806 6847
rect 11502 6360 13806 6383
rect 13196 5770 13802 5774
rect 11402 5596 13802 5770
rect -1110 4466 -578 4688
rect -1404 953 -1204 1004
rect -2608 906 -1996 914
rect -1404 906 -1386 953
rect -2608 700 -1386 906
rect -1404 649 -1386 700
rect -1242 649 -1204 953
rect -1404 600 -1204 649
rect -1110 -381 -888 4466
rect -803 4388 -413 4405
rect -803 4188 -204 4388
rect -803 4183 -413 4188
rect -803 -55 -581 4183
rect 13186 3852 13796 3854
rect 11764 3780 13800 3852
rect 11096 312 13806 338
rect 11096 88 12429 312
rect 12573 88 13806 312
rect 11096 58 13806 88
rect -803 -277 8801 -55
rect -1110 -603 2401 -381
rect 2179 -822 2401 -603
rect 8579 -818 8801 -277
rect 1908 -849 2708 -822
rect 1908 -905 1961 -849
rect 2017 -905 2041 -849
rect 2097 -905 2121 -849
rect 2177 -905 2201 -849
rect 2257 -905 2281 -849
rect 2337 -905 2361 -849
rect 2417 -905 2441 -849
rect 2497 -905 2521 -849
rect 2577 -905 2601 -849
rect 2657 -905 2708 -849
rect 1908 -932 2708 -905
rect 8384 -846 9204 -818
rect 8384 -902 8415 -846
rect 8471 -902 8495 -846
rect 8551 -902 8575 -846
rect 8631 -902 8655 -846
rect 8711 -902 8735 -846
rect 8791 -902 8815 -846
rect 8871 -902 8895 -846
rect 8951 -902 8975 -846
rect 9031 -902 9055 -846
rect 9111 -902 9135 -846
rect 9191 -902 9204 -846
rect 8384 -928 9204 -902
rect 8579 -933 8801 -928
rect -2608 -4954 -1786 -4948
rect -2608 -4980 9072 -4954
rect -2608 -5124 -1646 -4980
rect -1502 -5124 9072 -4980
rect -2608 -5148 9072 -5124
rect -2594 -5154 9072 -5148
rect -2594 -5158 2488 -5154
rect 1934 -9411 2040 -9390
rect 1934 -9475 1956 -9411
rect 2020 -9475 2040 -9411
rect 1934 -9491 2040 -9475
rect 1934 -9555 1956 -9491
rect 2020 -9555 2040 -9491
rect 1934 -9571 2040 -9555
rect 1934 -9635 1956 -9571
rect 2020 -9635 2040 -9571
rect 1934 -9651 2040 -9635
rect 1934 -9715 1956 -9651
rect 2020 -9715 2040 -9651
rect 1934 -9731 2040 -9715
rect 1934 -9795 1956 -9731
rect 2020 -9795 2040 -9731
rect 1934 -9811 2040 -9795
rect 1934 -9875 1956 -9811
rect 2020 -9875 2040 -9811
rect 1934 -9891 2040 -9875
rect 1934 -9955 1956 -9891
rect 2020 -9955 2040 -9891
rect 1934 -9988 2040 -9955
rect 5332 -9427 5438 -9402
rect 5332 -9491 5352 -9427
rect 5416 -9491 5438 -9427
rect 5332 -9507 5438 -9491
rect 5332 -9571 5352 -9507
rect 5416 -9571 5438 -9507
rect 5332 -9587 5438 -9571
rect 5332 -9651 5352 -9587
rect 5416 -9651 5438 -9587
rect 5332 -9667 5438 -9651
rect 5332 -9731 5352 -9667
rect 5416 -9731 5438 -9667
rect 5332 -9747 5438 -9731
rect 5332 -9811 5352 -9747
rect 5416 -9811 5438 -9747
rect 5332 -9827 5438 -9811
rect 5332 -9891 5352 -9827
rect 5416 -9891 5438 -9827
rect 5332 -9907 5438 -9891
rect 5332 -9971 5352 -9907
rect 5416 -9971 5438 -9907
rect 5332 -10000 5438 -9971
rect 8528 -9421 8634 -9394
rect 8528 -9485 8548 -9421
rect 8612 -9485 8634 -9421
rect 8528 -9501 8634 -9485
rect 8528 -9565 8548 -9501
rect 8612 -9565 8634 -9501
rect 8528 -9581 8634 -9565
rect 8528 -9645 8548 -9581
rect 8612 -9645 8634 -9581
rect 8528 -9661 8634 -9645
rect 8528 -9725 8548 -9661
rect 8612 -9725 8634 -9661
rect 8528 -9741 8634 -9725
rect 8528 -9805 8548 -9741
rect 8612 -9805 8634 -9741
rect 8528 -9821 8634 -9805
rect 8528 -9885 8548 -9821
rect 8612 -9885 8634 -9821
rect 8528 -9901 8634 -9885
rect 8528 -9965 8548 -9901
rect 8612 -9965 8634 -9901
rect 8528 -9992 8634 -9965
rect 11930 -9423 12036 -9396
rect 11930 -9487 11954 -9423
rect 12018 -9487 12036 -9423
rect 11930 -9503 12036 -9487
rect 11930 -9567 11954 -9503
rect 12018 -9567 12036 -9503
rect 11930 -9583 12036 -9567
rect 11930 -9647 11954 -9583
rect 12018 -9647 12036 -9583
rect 11930 -9663 12036 -9647
rect 11930 -9727 11954 -9663
rect 12018 -9727 12036 -9663
rect 11930 -9743 12036 -9727
rect 11930 -9807 11954 -9743
rect 12018 -9807 12036 -9743
rect 11930 -9823 12036 -9807
rect 11930 -9887 11954 -9823
rect 12018 -9887 12036 -9823
rect 11930 -9903 12036 -9887
rect 11930 -9967 11954 -9903
rect 12018 -9967 12036 -9903
rect 11930 -9994 12036 -9967
rect 2318 -11109 12898 -11074
rect 2318 -11173 12713 -11109
rect 12777 -11173 12793 -11109
rect 12857 -11173 12898 -11109
rect 2318 -11206 12898 -11173
rect 12394 -12812 12600 -12766
rect 12394 -12956 12427 -12812
rect 12571 -12956 12600 -12812
rect 12394 -12996 12600 -12956
rect 1926 -13226 2032 -13198
rect 1926 -13290 1949 -13226
rect 2013 -13290 2032 -13226
rect 1926 -13306 2032 -13290
rect 1926 -13370 1949 -13306
rect 2013 -13370 2032 -13306
rect 1926 -13386 2032 -13370
rect 1926 -13450 1949 -13386
rect 2013 -13450 2032 -13386
rect 1926 -13466 2032 -13450
rect 1926 -13530 1949 -13466
rect 2013 -13530 2032 -13466
rect 1926 -13546 2032 -13530
rect 1926 -13610 1949 -13546
rect 2013 -13610 2032 -13546
rect 1926 -13626 2032 -13610
rect 1926 -13690 1949 -13626
rect 2013 -13690 2032 -13626
rect 1926 -13706 2032 -13690
rect 1926 -13770 1949 -13706
rect 2013 -13770 2032 -13706
rect 1926 -13800 2032 -13770
rect 5332 -13230 5438 -13198
rect 5332 -13294 5351 -13230
rect 5415 -13294 5438 -13230
rect 5332 -13310 5438 -13294
rect 5332 -13374 5351 -13310
rect 5415 -13374 5438 -13310
rect 5332 -13390 5438 -13374
rect 5332 -13454 5351 -13390
rect 5415 -13454 5438 -13390
rect 5332 -13470 5438 -13454
rect 5332 -13534 5351 -13470
rect 5415 -13534 5438 -13470
rect 5332 -13550 5438 -13534
rect 5332 -13614 5351 -13550
rect 5415 -13614 5438 -13550
rect 5332 -13630 5438 -13614
rect 5332 -13694 5351 -13630
rect 5415 -13694 5438 -13630
rect 5332 -13710 5438 -13694
rect 5332 -13774 5351 -13710
rect 5415 -13774 5438 -13710
rect 5332 -13800 5438 -13774
rect 8526 -13226 8632 -13196
rect 8526 -13290 8549 -13226
rect 8613 -13290 8632 -13226
rect 8526 -13306 8632 -13290
rect 8526 -13370 8549 -13306
rect 8613 -13370 8632 -13306
rect 8526 -13386 8632 -13370
rect 8526 -13450 8549 -13386
rect 8613 -13450 8632 -13386
rect 8526 -13466 8632 -13450
rect 8526 -13530 8549 -13466
rect 8613 -13530 8632 -13466
rect 8526 -13546 8632 -13530
rect 8526 -13610 8549 -13546
rect 8613 -13610 8632 -13546
rect 8526 -13626 8632 -13610
rect 8526 -13690 8549 -13626
rect 8613 -13690 8632 -13626
rect 8526 -13706 8632 -13690
rect 8526 -13770 8549 -13706
rect 8613 -13770 8632 -13706
rect 8526 -13798 8632 -13770
rect 11938 -13220 12040 -13196
rect 11938 -13284 11958 -13220
rect 12022 -13284 12040 -13220
rect 11938 -13300 12040 -13284
rect 11938 -13364 11958 -13300
rect 12022 -13364 12040 -13300
rect 11938 -13380 12040 -13364
rect 11938 -13444 11958 -13380
rect 12022 -13444 12040 -13380
rect 11938 -13460 12040 -13444
rect 11938 -13524 11958 -13460
rect 12022 -13524 12040 -13460
rect 11938 -13540 12040 -13524
rect 11938 -13604 11958 -13540
rect 12022 -13604 12040 -13540
rect 11938 -13620 12040 -13604
rect 11938 -13684 11958 -13620
rect 12022 -13684 12040 -13620
rect 11938 -13700 12040 -13684
rect 11938 -13764 11958 -13700
rect 12022 -13764 12040 -13700
rect 11938 -13796 12040 -13764
<< via3 >>
rect -1654 11259 -1510 11483
rect 12707 6383 12851 6847
rect -1386 949 -1242 953
rect -1386 653 -1382 949
rect -1382 653 -1246 949
rect -1246 653 -1242 949
rect -1386 649 -1242 653
rect 12429 88 12573 312
rect -1646 -5124 -1502 -4980
rect 1956 -9415 2020 -9411
rect 1956 -9471 1960 -9415
rect 1960 -9471 2016 -9415
rect 2016 -9471 2020 -9415
rect 1956 -9475 2020 -9471
rect 1956 -9495 2020 -9491
rect 1956 -9551 1960 -9495
rect 1960 -9551 2016 -9495
rect 2016 -9551 2020 -9495
rect 1956 -9555 2020 -9551
rect 1956 -9575 2020 -9571
rect 1956 -9631 1960 -9575
rect 1960 -9631 2016 -9575
rect 2016 -9631 2020 -9575
rect 1956 -9635 2020 -9631
rect 1956 -9655 2020 -9651
rect 1956 -9711 1960 -9655
rect 1960 -9711 2016 -9655
rect 2016 -9711 2020 -9655
rect 1956 -9715 2020 -9711
rect 1956 -9735 2020 -9731
rect 1956 -9791 1960 -9735
rect 1960 -9791 2016 -9735
rect 2016 -9791 2020 -9735
rect 1956 -9795 2020 -9791
rect 1956 -9815 2020 -9811
rect 1956 -9871 1960 -9815
rect 1960 -9871 2016 -9815
rect 2016 -9871 2020 -9815
rect 1956 -9875 2020 -9871
rect 1956 -9895 2020 -9891
rect 1956 -9951 1960 -9895
rect 1960 -9951 2016 -9895
rect 2016 -9951 2020 -9895
rect 1956 -9955 2020 -9951
rect 5352 -9431 5416 -9427
rect 5352 -9487 5356 -9431
rect 5356 -9487 5412 -9431
rect 5412 -9487 5416 -9431
rect 5352 -9491 5416 -9487
rect 5352 -9511 5416 -9507
rect 5352 -9567 5356 -9511
rect 5356 -9567 5412 -9511
rect 5412 -9567 5416 -9511
rect 5352 -9571 5416 -9567
rect 5352 -9591 5416 -9587
rect 5352 -9647 5356 -9591
rect 5356 -9647 5412 -9591
rect 5412 -9647 5416 -9591
rect 5352 -9651 5416 -9647
rect 5352 -9671 5416 -9667
rect 5352 -9727 5356 -9671
rect 5356 -9727 5412 -9671
rect 5412 -9727 5416 -9671
rect 5352 -9731 5416 -9727
rect 5352 -9751 5416 -9747
rect 5352 -9807 5356 -9751
rect 5356 -9807 5412 -9751
rect 5412 -9807 5416 -9751
rect 5352 -9811 5416 -9807
rect 5352 -9831 5416 -9827
rect 5352 -9887 5356 -9831
rect 5356 -9887 5412 -9831
rect 5412 -9887 5416 -9831
rect 5352 -9891 5416 -9887
rect 5352 -9911 5416 -9907
rect 5352 -9967 5356 -9911
rect 5356 -9967 5412 -9911
rect 5412 -9967 5416 -9911
rect 5352 -9971 5416 -9967
rect 8548 -9425 8612 -9421
rect 8548 -9481 8552 -9425
rect 8552 -9481 8608 -9425
rect 8608 -9481 8612 -9425
rect 8548 -9485 8612 -9481
rect 8548 -9505 8612 -9501
rect 8548 -9561 8552 -9505
rect 8552 -9561 8608 -9505
rect 8608 -9561 8612 -9505
rect 8548 -9565 8612 -9561
rect 8548 -9585 8612 -9581
rect 8548 -9641 8552 -9585
rect 8552 -9641 8608 -9585
rect 8608 -9641 8612 -9585
rect 8548 -9645 8612 -9641
rect 8548 -9665 8612 -9661
rect 8548 -9721 8552 -9665
rect 8552 -9721 8608 -9665
rect 8608 -9721 8612 -9665
rect 8548 -9725 8612 -9721
rect 8548 -9745 8612 -9741
rect 8548 -9801 8552 -9745
rect 8552 -9801 8608 -9745
rect 8608 -9801 8612 -9745
rect 8548 -9805 8612 -9801
rect 8548 -9825 8612 -9821
rect 8548 -9881 8552 -9825
rect 8552 -9881 8608 -9825
rect 8608 -9881 8612 -9825
rect 8548 -9885 8612 -9881
rect 8548 -9905 8612 -9901
rect 8548 -9961 8552 -9905
rect 8552 -9961 8608 -9905
rect 8608 -9961 8612 -9905
rect 8548 -9965 8612 -9961
rect 11954 -9427 12018 -9423
rect 11954 -9483 11958 -9427
rect 11958 -9483 12014 -9427
rect 12014 -9483 12018 -9427
rect 11954 -9487 12018 -9483
rect 11954 -9507 12018 -9503
rect 11954 -9563 11958 -9507
rect 11958 -9563 12014 -9507
rect 12014 -9563 12018 -9507
rect 11954 -9567 12018 -9563
rect 11954 -9587 12018 -9583
rect 11954 -9643 11958 -9587
rect 11958 -9643 12014 -9587
rect 12014 -9643 12018 -9587
rect 11954 -9647 12018 -9643
rect 11954 -9667 12018 -9663
rect 11954 -9723 11958 -9667
rect 11958 -9723 12014 -9667
rect 12014 -9723 12018 -9667
rect 11954 -9727 12018 -9723
rect 11954 -9747 12018 -9743
rect 11954 -9803 11958 -9747
rect 11958 -9803 12014 -9747
rect 12014 -9803 12018 -9747
rect 11954 -9807 12018 -9803
rect 11954 -9827 12018 -9823
rect 11954 -9883 11958 -9827
rect 11958 -9883 12014 -9827
rect 12014 -9883 12018 -9827
rect 11954 -9887 12018 -9883
rect 11954 -9907 12018 -9903
rect 11954 -9963 11958 -9907
rect 11958 -9963 12014 -9907
rect 12014 -9963 12018 -9907
rect 11954 -9967 12018 -9963
rect 12713 -11173 12777 -11109
rect 12793 -11173 12857 -11109
rect 12427 -12816 12571 -12812
rect 12427 -12952 12431 -12816
rect 12431 -12952 12567 -12816
rect 12567 -12952 12571 -12816
rect 12427 -12956 12571 -12952
rect 1949 -13230 2013 -13226
rect 1949 -13286 1953 -13230
rect 1953 -13286 2009 -13230
rect 2009 -13286 2013 -13230
rect 1949 -13290 2013 -13286
rect 1949 -13310 2013 -13306
rect 1949 -13366 1953 -13310
rect 1953 -13366 2009 -13310
rect 2009 -13366 2013 -13310
rect 1949 -13370 2013 -13366
rect 1949 -13390 2013 -13386
rect 1949 -13446 1953 -13390
rect 1953 -13446 2009 -13390
rect 2009 -13446 2013 -13390
rect 1949 -13450 2013 -13446
rect 1949 -13470 2013 -13466
rect 1949 -13526 1953 -13470
rect 1953 -13526 2009 -13470
rect 2009 -13526 2013 -13470
rect 1949 -13530 2013 -13526
rect 1949 -13550 2013 -13546
rect 1949 -13606 1953 -13550
rect 1953 -13606 2009 -13550
rect 2009 -13606 2013 -13550
rect 1949 -13610 2013 -13606
rect 1949 -13630 2013 -13626
rect 1949 -13686 1953 -13630
rect 1953 -13686 2009 -13630
rect 2009 -13686 2013 -13630
rect 1949 -13690 2013 -13686
rect 1949 -13710 2013 -13706
rect 1949 -13766 1953 -13710
rect 1953 -13766 2009 -13710
rect 2009 -13766 2013 -13710
rect 1949 -13770 2013 -13766
rect 5351 -13234 5415 -13230
rect 5351 -13290 5355 -13234
rect 5355 -13290 5411 -13234
rect 5411 -13290 5415 -13234
rect 5351 -13294 5415 -13290
rect 5351 -13314 5415 -13310
rect 5351 -13370 5355 -13314
rect 5355 -13370 5411 -13314
rect 5411 -13370 5415 -13314
rect 5351 -13374 5415 -13370
rect 5351 -13394 5415 -13390
rect 5351 -13450 5355 -13394
rect 5355 -13450 5411 -13394
rect 5411 -13450 5415 -13394
rect 5351 -13454 5415 -13450
rect 5351 -13474 5415 -13470
rect 5351 -13530 5355 -13474
rect 5355 -13530 5411 -13474
rect 5411 -13530 5415 -13474
rect 5351 -13534 5415 -13530
rect 5351 -13554 5415 -13550
rect 5351 -13610 5355 -13554
rect 5355 -13610 5411 -13554
rect 5411 -13610 5415 -13554
rect 5351 -13614 5415 -13610
rect 5351 -13634 5415 -13630
rect 5351 -13690 5355 -13634
rect 5355 -13690 5411 -13634
rect 5411 -13690 5415 -13634
rect 5351 -13694 5415 -13690
rect 5351 -13714 5415 -13710
rect 5351 -13770 5355 -13714
rect 5355 -13770 5411 -13714
rect 5411 -13770 5415 -13714
rect 5351 -13774 5415 -13770
rect 8549 -13230 8613 -13226
rect 8549 -13286 8553 -13230
rect 8553 -13286 8609 -13230
rect 8609 -13286 8613 -13230
rect 8549 -13290 8613 -13286
rect 8549 -13310 8613 -13306
rect 8549 -13366 8553 -13310
rect 8553 -13366 8609 -13310
rect 8609 -13366 8613 -13310
rect 8549 -13370 8613 -13366
rect 8549 -13390 8613 -13386
rect 8549 -13446 8553 -13390
rect 8553 -13446 8609 -13390
rect 8609 -13446 8613 -13390
rect 8549 -13450 8613 -13446
rect 8549 -13470 8613 -13466
rect 8549 -13526 8553 -13470
rect 8553 -13526 8609 -13470
rect 8609 -13526 8613 -13470
rect 8549 -13530 8613 -13526
rect 8549 -13550 8613 -13546
rect 8549 -13606 8553 -13550
rect 8553 -13606 8609 -13550
rect 8609 -13606 8613 -13550
rect 8549 -13610 8613 -13606
rect 8549 -13630 8613 -13626
rect 8549 -13686 8553 -13630
rect 8553 -13686 8609 -13630
rect 8609 -13686 8613 -13630
rect 8549 -13690 8613 -13686
rect 8549 -13710 8613 -13706
rect 8549 -13766 8553 -13710
rect 8553 -13766 8609 -13710
rect 8609 -13766 8613 -13710
rect 8549 -13770 8613 -13766
rect 11958 -13224 12022 -13220
rect 11958 -13280 11962 -13224
rect 11962 -13280 12018 -13224
rect 12018 -13280 12022 -13224
rect 11958 -13284 12022 -13280
rect 11958 -13304 12022 -13300
rect 11958 -13360 11962 -13304
rect 11962 -13360 12018 -13304
rect 12018 -13360 12022 -13304
rect 11958 -13364 12022 -13360
rect 11958 -13384 12022 -13380
rect 11958 -13440 11962 -13384
rect 11962 -13440 12018 -13384
rect 12018 -13440 12022 -13384
rect 11958 -13444 12022 -13440
rect 11958 -13464 12022 -13460
rect 11958 -13520 11962 -13464
rect 11962 -13520 12018 -13464
rect 12018 -13520 12022 -13464
rect 11958 -13524 12022 -13520
rect 11958 -13544 12022 -13540
rect 11958 -13600 11962 -13544
rect 11962 -13600 12018 -13544
rect 12018 -13600 12022 -13544
rect 11958 -13604 12022 -13600
rect 11958 -13624 12022 -13620
rect 11958 -13680 11962 -13624
rect 11962 -13680 12018 -13624
rect 12018 -13680 12022 -13624
rect 11958 -13684 12022 -13680
rect 11958 -13704 12022 -13700
rect 11958 -13760 11962 -13704
rect 11962 -13760 12018 -13704
rect 12018 -13760 12022 -13704
rect 11958 -13764 12022 -13760
<< metal4 >>
rect -1676 11483 -1476 13018
rect -1676 11259 -1654 11483
rect -1510 11259 -1476 11483
rect -1676 -4980 -1476 11259
rect -1676 -5124 -1646 -4980
rect -1502 -5124 -1476 -4980
rect -1676 -12798 -1476 -5124
rect -1402 953 -1202 13020
rect -1402 649 -1386 953
rect -1242 649 -1202 953
rect -1402 -12796 -1202 649
rect 12398 312 12598 12816
rect 12398 88 12429 312
rect 12573 88 12598 312
rect 1934 -9411 2040 -9390
rect 1934 -9475 1956 -9411
rect 2020 -9475 2040 -9411
rect 1934 -9491 2040 -9475
rect 1934 -9555 1956 -9491
rect 2020 -9555 2040 -9491
rect 1934 -9571 2040 -9555
rect 1934 -9635 1956 -9571
rect 2020 -9635 2040 -9571
rect 1934 -9651 2040 -9635
rect 1934 -9715 1956 -9651
rect 2020 -9715 2040 -9651
rect 1934 -9731 2040 -9715
rect 1934 -9795 1956 -9731
rect 2020 -9795 2040 -9731
rect 1934 -9811 2040 -9795
rect 1934 -9875 1956 -9811
rect 2020 -9875 2040 -9811
rect 1934 -9891 2040 -9875
rect 1934 -9955 1956 -9891
rect 2020 -9955 2040 -9891
rect 1934 -9988 2040 -9955
rect 5332 -9427 5438 -9402
rect 5332 -9491 5352 -9427
rect 5416 -9491 5438 -9427
rect 5332 -9507 5438 -9491
rect 5332 -9571 5352 -9507
rect 5416 -9571 5438 -9507
rect 5332 -9587 5438 -9571
rect 5332 -9651 5352 -9587
rect 5416 -9651 5438 -9587
rect 5332 -9667 5438 -9651
rect 5332 -9731 5352 -9667
rect 5416 -9731 5438 -9667
rect 5332 -9747 5438 -9731
rect 5332 -9811 5352 -9747
rect 5416 -9811 5438 -9747
rect 5332 -9827 5438 -9811
rect 5332 -9891 5352 -9827
rect 5416 -9891 5438 -9827
rect 5332 -9907 5438 -9891
rect 5332 -9971 5352 -9907
rect 5416 -9950 5438 -9907
rect 8528 -9421 8634 -9394
rect 8528 -9485 8548 -9421
rect 8612 -9485 8634 -9421
rect 8528 -9501 8634 -9485
rect 8528 -9565 8548 -9501
rect 8612 -9565 8634 -9501
rect 8528 -9581 8634 -9565
rect 8528 -9645 8548 -9581
rect 8612 -9645 8634 -9581
rect 8528 -9661 8634 -9645
rect 8528 -9725 8548 -9661
rect 8612 -9725 8634 -9661
rect 8528 -9741 8634 -9725
rect 8528 -9805 8548 -9741
rect 8612 -9805 8634 -9741
rect 8528 -9821 8634 -9805
rect 8528 -9885 8548 -9821
rect 8612 -9885 8634 -9821
rect 8528 -9901 8634 -9885
rect 5416 -9971 5440 -9950
rect 1934 -13198 2036 -9988
rect 5332 -10026 5440 -9971
rect 8528 -9965 8548 -9901
rect 8612 -9965 8634 -9901
rect 8528 -10008 8634 -9965
rect 11930 -9423 12036 -9396
rect 11930 -9487 11954 -9423
rect 12018 -9487 12036 -9423
rect 11930 -9503 12036 -9487
rect 11930 -9567 11954 -9503
rect 12018 -9567 12036 -9503
rect 11930 -9583 12036 -9567
rect 11930 -9647 11954 -9583
rect 12018 -9647 12036 -9583
rect 11930 -9663 12036 -9647
rect 11930 -9727 11954 -9663
rect 12018 -9727 12036 -9663
rect 11930 -9743 12036 -9727
rect 11930 -9807 11954 -9743
rect 12018 -9807 12036 -9743
rect 11930 -9823 12036 -9807
rect 11930 -9887 11954 -9823
rect 12018 -9887 12036 -9823
rect 11930 -9903 12036 -9887
rect 11930 -9967 11954 -9903
rect 12018 -9967 12036 -9903
rect 11930 -9994 12036 -9967
rect 5340 -13198 5440 -10026
rect 8530 -13196 8630 -10008
rect 1926 -13226 2036 -13198
rect 1926 -13290 1949 -13226
rect 2013 -13290 2036 -13226
rect 1926 -13306 2036 -13290
rect 1926 -13370 1949 -13306
rect 2013 -13370 2036 -13306
rect 1926 -13386 2036 -13370
rect 1926 -13450 1949 -13386
rect 2013 -13450 2036 -13386
rect 1926 -13466 2036 -13450
rect 1926 -13530 1949 -13466
rect 2013 -13530 2036 -13466
rect 1926 -13546 2036 -13530
rect 1926 -13610 1949 -13546
rect 2013 -13610 2036 -13546
rect 1926 -13626 2036 -13610
rect 1926 -13690 1949 -13626
rect 2013 -13690 2036 -13626
rect 1926 -13706 2036 -13690
rect 1926 -13770 1949 -13706
rect 2013 -13770 2036 -13706
rect 1926 -13799 2036 -13770
rect 5332 -13230 5440 -13198
rect 5332 -13294 5351 -13230
rect 5415 -13294 5440 -13230
rect 5332 -13310 5440 -13294
rect 5332 -13374 5351 -13310
rect 5415 -13374 5440 -13310
rect 5332 -13390 5440 -13374
rect 5332 -13454 5351 -13390
rect 5415 -13454 5440 -13390
rect 5332 -13470 5440 -13454
rect 5332 -13534 5351 -13470
rect 5415 -13534 5440 -13470
rect 5332 -13550 5440 -13534
rect 5332 -13614 5351 -13550
rect 5415 -13614 5440 -13550
rect 5332 -13630 5440 -13614
rect 5332 -13694 5351 -13630
rect 5415 -13694 5440 -13630
rect 5332 -13710 5440 -13694
rect 5332 -13774 5351 -13710
rect 5415 -13774 5440 -13710
rect 5332 -13796 5440 -13774
rect 8526 -13226 8632 -13196
rect 8526 -13290 8549 -13226
rect 8613 -13290 8632 -13226
rect 8526 -13306 8632 -13290
rect 8526 -13370 8549 -13306
rect 8613 -13370 8632 -13306
rect 8526 -13386 8632 -13370
rect 8526 -13450 8549 -13386
rect 8613 -13450 8632 -13386
rect 8526 -13466 8632 -13450
rect 8526 -13530 8549 -13466
rect 8613 -13530 8632 -13466
rect 8526 -13546 8632 -13530
rect 8526 -13610 8549 -13546
rect 8613 -13610 8632 -13546
rect 8526 -13626 8632 -13610
rect 8526 -13690 8549 -13626
rect 8613 -13690 8632 -13626
rect 8526 -13706 8632 -13690
rect 8526 -13770 8549 -13706
rect 8613 -13770 8632 -13706
rect 1926 -13800 2032 -13799
rect 5332 -13800 5438 -13796
rect 8526 -13798 8632 -13770
rect 11936 -13220 12036 -9994
rect 12398 -12812 12598 88
rect 12398 -12956 12427 -12812
rect 12571 -12956 12598 -12812
rect 12398 -13000 12598 -12956
rect 12690 6847 12890 12818
rect 12690 6383 12707 6847
rect 12851 6383 12890 6847
rect 12690 -11109 12890 6383
rect 12690 -11173 12713 -11109
rect 12777 -11173 12793 -11109
rect 12857 -11173 12890 -11109
rect 12690 -12998 12890 -11173
rect 11936 -13284 11958 -13220
rect 12022 -13284 12036 -13220
rect 11936 -13300 12036 -13284
rect 11936 -13364 11958 -13300
rect 12022 -13364 12036 -13300
rect 11936 -13380 12036 -13364
rect 11936 -13444 11958 -13380
rect 12022 -13444 12036 -13380
rect 11936 -13460 12036 -13444
rect 11936 -13524 11958 -13460
rect 12022 -13524 12036 -13460
rect 11936 -13540 12036 -13524
rect 11936 -13604 11958 -13540
rect 12022 -13604 12036 -13540
rect 11936 -13620 12036 -13604
rect 11936 -13684 11958 -13620
rect 12022 -13684 12036 -13620
rect 11936 -13700 12036 -13684
rect 11936 -13764 11958 -13700
rect 12022 -13764 12036 -13700
rect 11936 -13802 12036 -13764
use EF_AMUX2to1ISO  EF_AMUX2to1ISO_0
timestamp 1699022965
transform 1 0 -797 0 1 -11804
box -3 -1196 6373 10978
use EF_AMUX2to1ISO  EF_AMUX2to1ISO_1
timestamp 1699022965
transform 1 0 5801 0 1 -11800
box -3 -1196 6373 10978
use EF_R2RVCE  EF_R2RVCE_0
timestamp 1699022965
transform 1 0 4 0 1 1465
box -804 -1465 11921 11144
<< labels >>
flabel metal2 s -400 -13788 -264 -13184 0 FreeSans 1250 0 0 0 SELA
port 1 nsew
flabel metal2 s 6200 -13808 6338 -13200 0 FreeSans 1250 0 0 0 SELB
port 2 nsew
flabel metal2 s 1932 -13804 2044 -13198 0 FreeSans 1250 0 0 0 A1
port 3 nsew
flabel metal2 s 5334 -13802 5446 -13192 0 FreeSans 1250 0 0 0 A2
port 4 nsew
flabel metal2 s 8526 -13798 8636 -13190 0 FreeSans 1250 0 0 0 B1
port 5 nsew
flabel metal2 s 11932 -13798 12038 -13196 0 FreeSans 1250 0 0 0 B2
port 6 nsew
flabel metal3 s -2608 -5148 -1786 -4948 0 FreeSans 1250 0 0 0 VDD
port 7 nsew
flabel metal3 s -2608 700 -1996 914 0 FreeSans 1250 0 0 0 VSS
port 8 nsew
flabel metal3 s 13046 66 13800 336 0 FreeSans 1250 0 0 0 DVSS
port 9 nsew
flabel metal3 s 13184 6370 13800 6886 0 FreeSans 1250 0 0 0 DVDD
port 10 nsew
flabel metal3 s 13196 5598 13802 5774 0 FreeSans 1250 0 0 0 VO
port 11 nsew
flabel metal3 s 13186 3782 13796 3854 0 FreeSans 1250 0 0 0 EN
port 12 nsew
<< end >>
