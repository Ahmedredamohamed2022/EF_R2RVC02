VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_R2RVC02m
  CLASS BLOCK ;
  FOREIGN EF_R2RVC02m ;
  ORIGIN 6.335 40.160 ;
  SIZE 76.095 BY 96.000 ;
  PIN a1
    PORT
      LAYER met1 ;
        RECT 13.000 -23.100 14.040 -20.430 ;
    END
  END a1
  PIN a2
    PORT
      LAYER met1 ;
        RECT 29.810 -25.510 30.770 -18.830 ;
    END
  END a2
  PIN b1
    PORT
      LAYER met1 ;
        RECT 46.210 -22.580 47.190 -20.110 ;
    END
  END b1
  PIN b2
    PORT
      LAYER met1 ;
        RECT 62.920 -22.220 63.900 -18.850 ;
    END
  END b2
  PIN dvss
    PORT
      LAYER met4 ;
        RECT 66.230 -39.245 67.230 0.660 ;
    END
  END dvss
  PIN vdd3p3
    PORT
      LAYER met4 ;
        RECT -6.310 -13.435 -5.190 55.810 ;
    END
  END vdd3p3
  PIN vss
    PORT
      LAYER met3 ;
        RECT -1.730 52.240 18.385 54.380 ;
    END
  END vss
  PIN vo
    PORT
      LAYER met2 ;
        RECT 59.310 22.065 59.940 22.470 ;
    END
  END vo
  PIN sela
    PORT
      LAYER met1 ;
        RECT 6.080 -38.420 8.670 -37.790 ;
    END
  END sela
  PIN selb
    PORT
      LAYER met1 ;
        RECT 40.570 -38.440 43.200 -37.850 ;
    END
  END selb
  PIN vdd1p8
    PORT
      LAYER met4 ;
        RECT 68.500 -39.870 69.500 -32.600 ;
    END
  END vdd1p8
  OBS
      LAYER li1 ;
        RECT 0.330 -39.890 64.300 52.065 ;
      LAYER met1 ;
        RECT -0.130 -18.550 67.280 51.750 ;
        RECT -0.130 -20.150 29.530 -18.550 ;
        RECT -0.130 -23.380 12.720 -20.150 ;
        RECT 14.320 -23.380 29.530 -20.150 ;
        RECT -0.130 -25.790 29.530 -23.380 ;
        RECT 31.050 -18.570 67.280 -18.550 ;
        RECT 31.050 -19.830 62.640 -18.570 ;
        RECT 31.050 -22.860 45.930 -19.830 ;
        RECT 47.470 -22.500 62.640 -19.830 ;
        RECT 64.180 -22.500 67.280 -18.570 ;
        RECT 47.470 -22.860 67.280 -22.500 ;
        RECT 31.050 -25.790 67.280 -22.860 ;
        RECT -0.130 -37.510 67.280 -25.790 ;
        RECT -0.130 -38.700 5.800 -37.510 ;
        RECT 8.950 -37.570 67.280 -37.510 ;
        RECT 8.950 -38.700 40.290 -37.570 ;
        RECT -0.130 -38.720 40.290 -38.700 ;
        RECT 43.480 -38.720 67.280 -37.570 ;
        RECT -0.130 -40.050 67.280 -38.720 ;
      LAYER met2 ;
        RECT -1.080 22.750 69.520 51.750 ;
        RECT -1.080 21.785 59.030 22.750 ;
        RECT 60.220 21.785 69.520 22.750 ;
        RECT -1.080 -40.050 69.520 21.785 ;
      LAYER met3 ;
        RECT -6.335 51.840 -2.130 54.380 ;
        RECT 18.785 51.840 69.760 54.380 ;
        RECT -6.335 -40.050 69.760 51.840 ;
      LAYER met4 ;
        RECT -4.790 1.060 69.760 55.840 ;
        RECT -4.790 -13.835 65.830 1.060 ;
        RECT -6.310 -39.645 65.830 -13.835 ;
        RECT 67.630 -32.200 69.760 1.060 ;
        RECT 67.630 -39.645 68.100 -32.200 ;
        RECT -6.310 -40.150 68.100 -39.645 ;
  END
END EF_R2RVC02m
END LIBRARY

