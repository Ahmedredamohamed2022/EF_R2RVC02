VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_R2RVC02
  CLASS BLOCK ;
  FOREIGN EF_R2RVC02 ;
  ORIGIN 13.040 69.040 ;
  SIZE 82.070 BY 134.140 ;
  PIN SELA
    ANTENNAGATEAREA 4.752000 ;
    PORT
      LAYER met2 ;
        RECT -2.000 -68.940 -1.320 -65.920 ;
    END
  END SELA
  PIN SELB
    ANTENNAGATEAREA 4.752000 ;
    PORT
      LAYER met2 ;
        RECT 31.000 -69.040 31.690 -66.000 ;
    END
  END SELB
  PIN A1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 9.660 -69.020 10.220 -65.990 ;
    END
  END A1
  PIN A2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 26.670 -69.010 27.230 -65.960 ;
    END
  END A2
  PIN B1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 42.630 -68.990 43.180 -65.950 ;
    END
  END B1
  PIN B2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 59.660 -68.990 60.190 -65.980 ;
    END
  END B2
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 598.042908 ;
    PORT
      LAYER met3 ;
        RECT -13.040 -25.740 -8.930 -24.740 ;
    END
  END VDD
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 271.063080 ;
    PORT
      LAYER met3 ;
        RECT -13.040 3.500 -9.980 4.570 ;
    END
  END VSS
  PIN DVSS
    ANTENNADIFFAREA 215.901642 ;
    PORT
      LAYER met3 ;
        RECT 65.230 0.330 69.000 1.680 ;
    END
  END DVSS
  PIN DVDD
    ANTENNADIFFAREA 9.946099 ;
    PORT
      LAYER met3 ;
        RECT 65.920 31.850 69.000 34.430 ;
    END
  END DVDD
  PIN VO
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 65.980 27.990 69.010 28.870 ;
    END
  END VO
  PIN EN
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met3 ;
        RECT 65.930 18.910 68.980 19.270 ;
    END
  END EN
  OBS
      LAYER li1 ;
        RECT -3.655 -64.590 60.445 62.655 ;
      LAYER met1 ;
        RECT -4.045 -65.000 62.975 62.545 ;
      LAYER met2 ;
        RECT -7.020 -65.640 63.000 62.345 ;
        RECT -7.020 -69.005 -2.280 -65.640 ;
        RECT -1.040 -65.670 63.000 -65.640 ;
        RECT -1.040 -65.680 42.350 -65.670 ;
        RECT -1.040 -65.710 26.390 -65.680 ;
        RECT -1.040 -69.005 9.380 -65.710 ;
        RECT 10.500 -69.005 26.390 -65.710 ;
        RECT 27.510 -65.720 42.350 -65.680 ;
        RECT 27.510 -69.005 30.720 -65.720 ;
        RECT 31.970 -69.005 42.350 -65.720 ;
        RECT 43.460 -65.700 63.000 -65.670 ;
        RECT 43.460 -69.005 59.380 -65.700 ;
        RECT 60.470 -69.005 63.000 -65.700 ;
      LAYER met3 ;
        RECT -12.970 34.830 69.030 62.365 ;
        RECT -12.970 31.450 65.520 34.830 ;
        RECT -12.970 29.270 69.030 31.450 ;
        RECT -12.970 27.590 65.580 29.270 ;
        RECT -12.970 19.670 69.030 27.590 ;
        RECT -12.970 18.510 65.530 19.670 ;
        RECT -12.970 4.970 69.030 18.510 ;
        RECT -9.580 3.100 69.030 4.970 ;
        RECT -12.970 2.080 69.030 3.100 ;
        RECT -12.970 -0.070 64.830 2.080 ;
        RECT -12.970 -24.340 69.030 -0.070 ;
        RECT -8.530 -26.140 69.030 -24.340 ;
        RECT -12.970 -69.000 69.030 -26.140 ;
      LAYER met4 ;
        RECT -8.380 -69.010 64.450 65.100 ;
      LAYER met5 ;
        RECT 47.380 2.235 50.380 61.155 ;
  END
END EF_R2RVC02
END LIBRARY

