** NOTE: ngspice DOES NOT handle environment variables used in the test benches. the Makefile handles that for you, if you wish to use your own command make sure you manually update the spice files


V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
C1 VO VSS 1p m=1
V5 DVDD VSS 1.8
.save i(v5)
V3 B1 VSS pulse(0 3.3 0 4.95us 4.95us 0.1us 10us)
.save i(v3)
V4 A1 VSS 1
.save i(v4)
*x1 VO VDD B1 A1 VSS B2 A2 DVDD VSS SELA SELB EF_R2RVC02X
*x1 A1 A2 B1 B2 VO SELA SELB DVDD VSS VSS VDD EF_R2RVC02mf

x2 VSS VO SELB A2 B2 B1 SELA DVSS A1 DVDD VDD EF_R2RVC02

V16 DVSS GND 0
.save i(v16)

V6 B2 VSS pulse(0 2.5 0 4.95us 4.95us 0.1us 10us)
.save i(v6)
V7 A2 VSS 2
.save i(v7)
V8 SELB VSS 0
.save i(v8)
V9 SELA VSS 0
.save i(v9)
**** begin user architecture code


.option wnflag=1
.option TEMP=27
.option TNOM=27
.option wnflag=1
.control
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
save all
run
tran 10n 20e-6 0.1u

plot A1 B1 VO
plot A2 B2 VO

.endc


.lib $PDK_ROOT/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include ../../spice/$SIM/EF_R2RVC02.spice


**.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
**.include /ciic/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /home/ahmedreda/PDK/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /home/ahmedreda/PDK/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl__lsbuflv2hv_1.spice



.GLOBAL GND
.end
