magic
tech sky130A
magscale 1 2
timestamp 1699954036
<< metal1 >>
rect 338 10650 404 10866
rect 42 6609 2578 6670
rect 42 6493 79 6609
rect 195 6556 2578 6609
rect 195 6493 228 6556
rect 42 6424 228 6493
rect 42 6401 734 6424
rect 42 6349 75 6401
rect 127 6349 139 6401
rect 191 6349 734 6401
rect 42 6322 734 6349
rect 52 6318 734 6322
rect 2376 6316 2542 6422
rect 2232 6258 2342 6274
rect 784 6237 2352 6258
rect 784 6185 2257 6237
rect 2309 6185 2352 6237
rect 784 6184 2352 6185
rect 2232 6140 2342 6184
rect 2434 6052 2538 6316
rect 2734 6052 2838 6916
rect 2434 6038 2838 6052
rect 322 5948 2838 6038
rect 322 5934 2542 5948
rect 322 5840 428 5934
rect 2867 4367 2973 7023
rect 2734 1802 2838 1906
rect 2208 1299 2392 1330
rect 2208 1183 2241 1299
rect 2357 1183 2392 1299
rect 2208 1150 2392 1183
rect 1000 589 1200 618
rect 2701 598 2787 658
rect 2867 598 2973 2003
rect 2701 597 2973 598
rect 2701 596 2883 597
rect 1000 537 1043 589
rect 1095 537 1107 589
rect 1159 537 1200 589
rect 1000 500 1200 537
rect 344 246 610 426
<< via1 >>
rect 79 6493 195 6609
rect 75 6349 127 6401
rect 139 6349 191 6401
rect 2257 6185 2309 6237
rect 2241 1183 2357 1299
rect 1043 537 1095 589
rect 1107 537 1159 589
<< metal2 >>
rect 708 8991 880 9010
rect 708 8855 726 8991
rect 862 8855 880 8991
rect 708 8836 880 8855
rect 56 7020 774 7192
rect 56 6609 228 7020
rect 56 6493 79 6609
rect 195 6493 228 6609
rect 56 6401 228 6493
rect 56 6349 75 6401
rect 127 6349 139 6401
rect 191 6349 228 6401
rect 56 2203 228 6349
rect 2230 6239 2344 6282
rect 2230 6183 2255 6239
rect 2311 6183 2344 6239
rect 2230 6150 2344 6183
rect 2232 6140 2342 6150
rect 704 3940 878 3972
rect 704 3884 723 3940
rect 779 3884 803 3940
rect 859 3884 878 3940
rect 704 3852 878 3884
rect 56 2037 787 2203
rect 926 2078 1100 2198
rect 56 1200 228 2037
rect 2208 1309 2392 1330
rect 2208 1173 2231 1309
rect 2367 1173 2392 1309
rect 2208 1150 2392 1173
rect 708 1062 882 1094
rect 708 1006 727 1062
rect 783 1006 807 1062
rect 863 1006 882 1062
rect 708 974 882 1006
rect 1000 591 1200 618
rect 1000 535 1033 591
rect 1089 589 1113 591
rect 1095 537 1107 589
rect 1089 535 1113 537
rect 1169 535 1200 591
rect 1000 500 1200 535
<< via2 >>
rect 726 8855 862 8991
rect 2255 6237 2311 6239
rect 2255 6185 2257 6237
rect 2257 6185 2309 6237
rect 2309 6185 2311 6237
rect 2255 6183 2311 6185
rect 723 3884 779 3940
rect 803 3884 859 3940
rect 2231 1299 2367 1309
rect 2231 1183 2241 1299
rect 2241 1183 2357 1299
rect 2357 1183 2367 1299
rect 2231 1173 2367 1183
rect 727 1006 783 1062
rect 807 1006 863 1062
rect 1033 589 1089 591
rect 1113 589 1169 591
rect 1033 537 1043 589
rect 1043 537 1089 589
rect 1113 537 1159 589
rect 1159 537 1169 589
rect 1033 535 1089 537
rect 1113 535 1169 537
<< metal3 >>
rect 690 8991 890 9024
rect 690 8855 726 8991
rect 862 8855 890 8991
rect 690 3940 890 8855
rect 690 3884 723 3940
rect 779 3884 803 3940
rect 859 3884 890 3940
rect 302 968 618 1092
rect 690 1062 890 3884
rect 2230 6239 2342 6274
rect 2230 6183 2255 6239
rect 2311 6183 2342 6239
rect 2230 1330 2342 6183
rect 2208 1309 2392 1330
rect 2208 1173 2231 1309
rect 2367 1173 2392 1309
rect 2208 1150 2392 1173
rect 690 1006 727 1062
rect 783 1006 807 1062
rect 863 1006 890 1062
rect 690 966 890 1006
rect 1000 591 1200 618
rect 1000 535 1033 591
rect 1089 535 1113 591
rect 1169 535 1200 591
rect 1000 500 1200 535
use single_ls  single_ls_0
timestamp 1699954036
transform 1 0 -2700 0 1 -302
box 2700 202 5594 1958
use single_tg  single_tg_0
timestamp 1699954036
transform -1 0 5076 0 1 6804
box 2103 0 4754 4142
use single_tg  single_tg_1
timestamp 1699954036
transform -1 0 5076 0 1 1802
box 2103 0 4754 4142
use sky130_fd_pr__nfet_g5v0d10v5_RDJSSL  sky130_fd_pr__nfet_g5v0d10v5_RDJSSL_0
timestamp 1699954036
transform 1 0 1552 0 1 6364
box -1018 -298 1018 298
<< labels >>
flabel metal3 s 704 3852 878 3972 0 FreeSans 146 0 0 0 VDD
port 1 nsew
flabel metal2 s 926 2078 1100 2198 0 FreeSans 146 0 0 0 DVSS
port 2 nsew
flabel metal1 s 344 246 610 426 0 FreeSans 146 0 0 0 DINL
port 3 nsew
flabel metal1 s 2734 1802 2838 1906 0 FreeSans 146 0 0 0 VIN
port 4 nsew
flabel metal3 s 1000 502 1200 618 0 FreeSans 146 0 0 0 DVDD
port 5 nsew
flabel metal1 s 338 10650 404 10866 0 FreeSans 374 0 0 0 VOUT
port 6 nsew
<< end >>
