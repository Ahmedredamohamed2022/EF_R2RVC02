VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_R2RVC02
  CLASS BLOCK ;
  FOREIGN EF_R2RVC02 ;
  ORIGIN 9.920 43.080 ;
  SIZE 80.940 BY 99.460 ;
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 263.488281 ;
    PORT
      LAYER met3 ;
        RECT -8.060 52.310 -4.000 54.370 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 433.882782 ;
    PORT
      LAYER met3 ;
        RECT -8.080 54.840 -2.990 56.380 ;
    END
  END VDD
  PIN SELA
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met2 ;
        RECT 1.720 -42.990 2.640 -38.620 ;
    END
  END SELA
  PIN A2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 29.780 -43.020 30.700 -38.650 ;
    END
  END A2
  PIN SELB
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met2 ;
        RECT 34.970 -43.080 35.890 -38.710 ;
    END
  END SELB
  PIN B1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 46.130 -42.970 47.050 -38.600 ;
    END
  END B1
  PIN B2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 62.900 -43.000 63.820 -38.630 ;
    END
  END B2
  PIN VO
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 65.910 21.820 71.000 22.800 ;
    END
  END VO
  PIN A1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 12.890 -43.000 13.990 -38.400 ;
    END
  END A1
  PIN DVSS
    ANTENNADIFFAREA 107.239799 ;
    PORT
      LAYER met3 ;
        RECT 67.310 0.310 70.980 3.610 ;
    END
  END DVSS
  PIN DVDD
    ANTENNADIFFAREA 7.633700 ;
    PORT
      LAYER met4 ;
        RECT 68.070 26.010 71.020 28.330 ;
    END
  END DVDD
  OBS
      LAYER li1 ;
        RECT 0.330 -39.890 64.300 52.065 ;
      LAYER met1 ;
        RECT -0.130 -40.050 67.280 51.750 ;
      LAYER met2 ;
        RECT -1.080 -38.120 70.210 51.750 ;
        RECT -1.080 -38.340 12.610 -38.120 ;
        RECT -1.080 -42.230 1.440 -38.340 ;
        RECT 2.920 -42.230 12.610 -38.340 ;
        RECT 14.270 -38.320 70.210 -38.120 ;
        RECT 14.270 -38.370 45.850 -38.320 ;
        RECT 14.270 -42.230 29.500 -38.370 ;
        RECT 30.980 -38.430 45.850 -38.370 ;
        RECT 30.980 -42.230 34.690 -38.430 ;
        RECT 36.170 -42.230 45.850 -38.430 ;
        RECT 47.330 -38.350 70.210 -38.320 ;
        RECT 47.330 -42.230 62.620 -38.350 ;
        RECT 64.100 -42.230 70.210 -38.350 ;
      LAYER met3 ;
        RECT -2.590 54.440 71.020 56.360 ;
        RECT -3.600 51.910 71.020 54.440 ;
        RECT -8.090 23.200 71.020 51.910 ;
        RECT -8.090 21.420 65.510 23.200 ;
        RECT -8.090 4.010 71.020 21.420 ;
        RECT -8.090 -0.090 66.910 4.010 ;
        RECT -8.090 -42.230 71.020 -0.090 ;
      LAYER met4 ;
        RECT -8.060 28.730 69.760 56.370 ;
        RECT -8.060 25.610 67.670 28.730 ;
        RECT -8.060 -42.230 69.760 25.610 ;
  END
END EF_R2RVC02
END LIBRARY

