magic
tech sky130A
magscale 1 2
timestamp 1699954036
<< dnwell >>
rect -91 5652 10727 10125
rect -91 -1356 9527 5652
<< nwell >>
rect -200 10017 10836 10234
rect -200 -1150 115 10017
rect 10521 6187 10836 10017
rect 5341 5929 10836 6187
rect 9361 5858 10836 5929
rect 9321 5543 10836 5858
rect 9321 -1150 9636 5543
rect -200 -1465 9636 -1150
<< mvnsubdiff >>
rect -134 10148 10770 10168
rect -134 10114 -37 10148
rect -3 10114 31 10148
rect 65 10114 99 10148
rect 133 10114 167 10148
rect 201 10114 235 10148
rect 269 10114 303 10148
rect 337 10114 371 10148
rect 405 10114 439 10148
rect 473 10114 507 10148
rect 541 10114 575 10148
rect 609 10114 643 10148
rect 677 10114 711 10148
rect 745 10114 779 10148
rect 813 10114 847 10148
rect 881 10114 915 10148
rect 949 10114 983 10148
rect 1017 10114 1051 10148
rect 1085 10114 1119 10148
rect 1153 10114 1187 10148
rect 1221 10114 1255 10148
rect 1289 10114 1323 10148
rect 1357 10114 1391 10148
rect 1425 10114 1459 10148
rect 1493 10114 1527 10148
rect 1561 10114 1595 10148
rect 1629 10114 1663 10148
rect 1697 10114 1731 10148
rect 1765 10114 1799 10148
rect 1833 10114 1867 10148
rect 1901 10114 1935 10148
rect 1969 10114 2003 10148
rect 2037 10114 2071 10148
rect 2105 10114 2139 10148
rect 2173 10114 2207 10148
rect 2241 10114 2275 10148
rect 2309 10114 2343 10148
rect 2377 10114 2411 10148
rect 2445 10114 2479 10148
rect 2513 10114 2547 10148
rect 2581 10114 2615 10148
rect 2649 10114 2683 10148
rect 2717 10114 2751 10148
rect 2785 10114 2819 10148
rect 2853 10114 2887 10148
rect 2921 10114 2955 10148
rect 2989 10114 3023 10148
rect 3057 10114 3091 10148
rect 3125 10114 3159 10148
rect 3193 10114 3227 10148
rect 3261 10114 3295 10148
rect 3329 10114 3363 10148
rect 3397 10114 3431 10148
rect 3465 10114 3499 10148
rect 3533 10114 3567 10148
rect 3601 10114 3635 10148
rect 3669 10114 3703 10148
rect 3737 10114 3771 10148
rect 3805 10114 3839 10148
rect 3873 10114 3907 10148
rect 3941 10114 3975 10148
rect 4009 10114 4043 10148
rect 4077 10114 4111 10148
rect 4145 10114 4179 10148
rect 4213 10114 4247 10148
rect 4281 10114 4315 10148
rect 4349 10114 4383 10148
rect 4417 10114 4451 10148
rect 4485 10114 4519 10148
rect 4553 10114 4587 10148
rect 4621 10114 4655 10148
rect 4689 10114 4723 10148
rect 4757 10114 4791 10148
rect 4825 10114 4859 10148
rect 4893 10114 4927 10148
rect 4961 10114 4995 10148
rect 5029 10114 5063 10148
rect 5097 10114 5131 10148
rect 5165 10114 5199 10148
rect 5233 10114 5267 10148
rect 5301 10114 5335 10148
rect 5369 10114 5403 10148
rect 5437 10114 5471 10148
rect 5505 10114 5539 10148
rect 5573 10114 5607 10148
rect 5641 10114 5675 10148
rect 5709 10114 5743 10148
rect 5777 10114 5811 10148
rect 5845 10114 5879 10148
rect 5913 10114 5947 10148
rect 5981 10114 6015 10148
rect 6049 10114 6083 10148
rect 6117 10114 6151 10148
rect 6185 10114 6219 10148
rect 6253 10114 6287 10148
rect 6321 10114 6355 10148
rect 6389 10114 6423 10148
rect 6457 10114 6491 10148
rect 6525 10114 6559 10148
rect 6593 10114 6627 10148
rect 6661 10114 6695 10148
rect 6729 10114 6763 10148
rect 6797 10114 6831 10148
rect 6865 10114 6899 10148
rect 6933 10114 6967 10148
rect 7001 10114 7035 10148
rect 7069 10114 7103 10148
rect 7137 10114 7171 10148
rect 7205 10114 7239 10148
rect 7273 10114 7307 10148
rect 7341 10114 7375 10148
rect 7409 10114 7443 10148
rect 7477 10114 7511 10148
rect 7545 10114 7579 10148
rect 7613 10114 7647 10148
rect 7681 10114 7715 10148
rect 7749 10114 7783 10148
rect 7817 10114 7851 10148
rect 7885 10114 7919 10148
rect 7953 10114 7987 10148
rect 8021 10114 8055 10148
rect 8089 10114 8123 10148
rect 8157 10114 8191 10148
rect 8225 10114 8259 10148
rect 8293 10114 8327 10148
rect 8361 10114 8395 10148
rect 8429 10114 8463 10148
rect 8497 10114 8531 10148
rect 8565 10114 8599 10148
rect 8633 10114 8667 10148
rect 8701 10114 8735 10148
rect 8769 10114 8803 10148
rect 8837 10114 8871 10148
rect 8905 10114 8939 10148
rect 8973 10114 9007 10148
rect 9041 10114 9075 10148
rect 9109 10114 9143 10148
rect 9177 10114 9211 10148
rect 9245 10114 9279 10148
rect 9313 10114 9347 10148
rect 9381 10114 9415 10148
rect 9449 10114 9483 10148
rect 9517 10114 9551 10148
rect 9585 10114 9619 10148
rect 9653 10114 9687 10148
rect 9721 10114 9755 10148
rect 9789 10114 9823 10148
rect 9857 10114 9891 10148
rect 9925 10114 9959 10148
rect 9993 10114 10027 10148
rect 10061 10114 10095 10148
rect 10129 10114 10163 10148
rect 10197 10114 10231 10148
rect 10265 10114 10299 10148
rect 10333 10114 10367 10148
rect 10401 10114 10435 10148
rect 10469 10114 10503 10148
rect 10537 10114 10571 10148
rect 10605 10114 10639 10148
rect 10673 10114 10770 10148
rect -134 10094 10770 10114
rect -134 10067 -60 10094
rect -134 10033 -114 10067
rect -80 10033 -60 10067
rect -134 9999 -60 10033
rect -134 9965 -114 9999
rect -80 9965 -60 9999
rect -134 9931 -60 9965
rect -134 9897 -114 9931
rect -80 9897 -60 9931
rect -134 9863 -60 9897
rect -134 9829 -114 9863
rect -80 9829 -60 9863
rect -134 9795 -60 9829
rect -134 9761 -114 9795
rect -80 9761 -60 9795
rect -134 9727 -60 9761
rect -134 9693 -114 9727
rect -80 9693 -60 9727
rect -134 9659 -60 9693
rect -134 9625 -114 9659
rect -80 9625 -60 9659
rect -134 9591 -60 9625
rect -134 9557 -114 9591
rect -80 9557 -60 9591
rect -134 9523 -60 9557
rect -134 9489 -114 9523
rect -80 9489 -60 9523
rect -134 9455 -60 9489
rect -134 9421 -114 9455
rect -80 9421 -60 9455
rect -134 9387 -60 9421
rect -134 9353 -114 9387
rect -80 9353 -60 9387
rect -134 9319 -60 9353
rect -134 9285 -114 9319
rect -80 9285 -60 9319
rect -134 9251 -60 9285
rect -134 9217 -114 9251
rect -80 9217 -60 9251
rect -134 9183 -60 9217
rect -134 9149 -114 9183
rect -80 9149 -60 9183
rect -134 9115 -60 9149
rect -134 9081 -114 9115
rect -80 9081 -60 9115
rect -134 9047 -60 9081
rect -134 9013 -114 9047
rect -80 9013 -60 9047
rect -134 8979 -60 9013
rect -134 8945 -114 8979
rect -80 8945 -60 8979
rect -134 8911 -60 8945
rect -134 8877 -114 8911
rect -80 8877 -60 8911
rect -134 8843 -60 8877
rect -134 8809 -114 8843
rect -80 8809 -60 8843
rect -134 8775 -60 8809
rect -134 8741 -114 8775
rect -80 8741 -60 8775
rect -134 8707 -60 8741
rect -134 8673 -114 8707
rect -80 8673 -60 8707
rect -134 8639 -60 8673
rect -134 8605 -114 8639
rect -80 8605 -60 8639
rect -134 8571 -60 8605
rect -134 8537 -114 8571
rect -80 8537 -60 8571
rect -134 8503 -60 8537
rect -134 8469 -114 8503
rect -80 8469 -60 8503
rect -134 8435 -60 8469
rect -134 8401 -114 8435
rect -80 8401 -60 8435
rect -134 8367 -60 8401
rect -134 8333 -114 8367
rect -80 8333 -60 8367
rect -134 8299 -60 8333
rect -134 8265 -114 8299
rect -80 8265 -60 8299
rect -134 8231 -60 8265
rect -134 8197 -114 8231
rect -80 8197 -60 8231
rect -134 8163 -60 8197
rect -134 8129 -114 8163
rect -80 8129 -60 8163
rect -134 8095 -60 8129
rect -134 8061 -114 8095
rect -80 8061 -60 8095
rect -134 8027 -60 8061
rect -134 7993 -114 8027
rect -80 7993 -60 8027
rect -134 7959 -60 7993
rect -134 7925 -114 7959
rect -80 7925 -60 7959
rect -134 7891 -60 7925
rect -134 7857 -114 7891
rect -80 7857 -60 7891
rect -134 7823 -60 7857
rect -134 7789 -114 7823
rect -80 7789 -60 7823
rect -134 7755 -60 7789
rect -134 7721 -114 7755
rect -80 7721 -60 7755
rect -134 7687 -60 7721
rect -134 7653 -114 7687
rect -80 7653 -60 7687
rect -134 7619 -60 7653
rect -134 7585 -114 7619
rect -80 7585 -60 7619
rect -134 7551 -60 7585
rect -134 7517 -114 7551
rect -80 7517 -60 7551
rect -134 7483 -60 7517
rect -134 7449 -114 7483
rect -80 7449 -60 7483
rect -134 7415 -60 7449
rect -134 7381 -114 7415
rect -80 7381 -60 7415
rect -134 7347 -60 7381
rect -134 7313 -114 7347
rect -80 7313 -60 7347
rect -134 7279 -60 7313
rect -134 7245 -114 7279
rect -80 7245 -60 7279
rect -134 7211 -60 7245
rect -134 7177 -114 7211
rect -80 7177 -60 7211
rect -134 7143 -60 7177
rect -134 7109 -114 7143
rect -80 7109 -60 7143
rect -134 7075 -60 7109
rect -134 7041 -114 7075
rect -80 7041 -60 7075
rect -134 7007 -60 7041
rect -134 6973 -114 7007
rect -80 6973 -60 7007
rect -134 6939 -60 6973
rect -134 6905 -114 6939
rect -80 6905 -60 6939
rect -134 6871 -60 6905
rect -134 6837 -114 6871
rect -80 6837 -60 6871
rect -134 6803 -60 6837
rect -134 6769 -114 6803
rect -80 6769 -60 6803
rect -134 6735 -60 6769
rect -134 6701 -114 6735
rect -80 6701 -60 6735
rect -134 6667 -60 6701
rect -134 6633 -114 6667
rect -80 6633 -60 6667
rect -134 6599 -60 6633
rect -134 6565 -114 6599
rect -80 6565 -60 6599
rect -134 6531 -60 6565
rect -134 6497 -114 6531
rect -80 6497 -60 6531
rect -134 6463 -60 6497
rect -134 6429 -114 6463
rect -80 6429 -60 6463
rect -134 6395 -60 6429
rect -134 6361 -114 6395
rect -80 6361 -60 6395
rect -134 6327 -60 6361
rect -134 6293 -114 6327
rect -80 6293 -60 6327
rect -134 6259 -60 6293
rect -134 6225 -114 6259
rect -80 6225 -60 6259
rect -134 6191 -60 6225
rect -134 6157 -114 6191
rect -80 6157 -60 6191
rect -134 6123 -60 6157
rect -134 6089 -114 6123
rect -80 6089 -60 6123
rect -134 6055 -60 6089
rect -134 6021 -114 6055
rect -80 6021 -60 6055
rect -134 5987 -60 6021
rect -134 5953 -114 5987
rect -80 5953 -60 5987
rect -134 5919 -60 5953
rect -134 5885 -114 5919
rect -80 5885 -60 5919
rect -134 5851 -60 5885
rect -134 5817 -114 5851
rect -80 5817 -60 5851
rect -134 5783 -60 5817
rect -134 5749 -114 5783
rect -80 5749 -60 5783
rect -134 5715 -60 5749
rect -134 5681 -114 5715
rect -80 5681 -60 5715
rect 10696 10079 10770 10094
rect 10696 10045 10716 10079
rect 10750 10045 10770 10079
rect 10696 10011 10770 10045
rect 10696 9977 10716 10011
rect 10750 9977 10770 10011
rect 10696 9943 10770 9977
rect 10696 9909 10716 9943
rect 10750 9909 10770 9943
rect 10696 9875 10770 9909
rect 10696 9841 10716 9875
rect 10750 9841 10770 9875
rect 10696 9807 10770 9841
rect 10696 9773 10716 9807
rect 10750 9773 10770 9807
rect 10696 9739 10770 9773
rect 10696 9705 10716 9739
rect 10750 9705 10770 9739
rect 10696 9671 10770 9705
rect 10696 9637 10716 9671
rect 10750 9637 10770 9671
rect 10696 9603 10770 9637
rect 10696 9569 10716 9603
rect 10750 9569 10770 9603
rect 10696 9535 10770 9569
rect 10696 9501 10716 9535
rect 10750 9501 10770 9535
rect 10696 9467 10770 9501
rect 10696 9433 10716 9467
rect 10750 9433 10770 9467
rect 10696 9399 10770 9433
rect 10696 9365 10716 9399
rect 10750 9365 10770 9399
rect 10696 9331 10770 9365
rect 10696 9297 10716 9331
rect 10750 9297 10770 9331
rect 10696 9263 10770 9297
rect 10696 9229 10716 9263
rect 10750 9229 10770 9263
rect 10696 9195 10770 9229
rect 10696 9161 10716 9195
rect 10750 9161 10770 9195
rect 10696 9127 10770 9161
rect 10696 9093 10716 9127
rect 10750 9093 10770 9127
rect 10696 9059 10770 9093
rect 10696 9025 10716 9059
rect 10750 9025 10770 9059
rect 10696 8991 10770 9025
rect 10696 8957 10716 8991
rect 10750 8957 10770 8991
rect 10696 8923 10770 8957
rect 10696 8889 10716 8923
rect 10750 8889 10770 8923
rect 10696 8855 10770 8889
rect 10696 8821 10716 8855
rect 10750 8821 10770 8855
rect 10696 8787 10770 8821
rect 10696 8753 10716 8787
rect 10750 8753 10770 8787
rect 10696 8719 10770 8753
rect 10696 8685 10716 8719
rect 10750 8685 10770 8719
rect 10696 8651 10770 8685
rect 10696 8617 10716 8651
rect 10750 8617 10770 8651
rect 10696 8583 10770 8617
rect 10696 8549 10716 8583
rect 10750 8549 10770 8583
rect 10696 8515 10770 8549
rect 10696 8481 10716 8515
rect 10750 8481 10770 8515
rect 10696 8447 10770 8481
rect 10696 8413 10716 8447
rect 10750 8413 10770 8447
rect 10696 8379 10770 8413
rect 10696 8345 10716 8379
rect 10750 8345 10770 8379
rect 10696 8311 10770 8345
rect 10696 8277 10716 8311
rect 10750 8277 10770 8311
rect 10696 8243 10770 8277
rect 10696 8209 10716 8243
rect 10750 8209 10770 8243
rect 10696 8175 10770 8209
rect 10696 8141 10716 8175
rect 10750 8141 10770 8175
rect 10696 8107 10770 8141
rect 10696 8073 10716 8107
rect 10750 8073 10770 8107
rect 10696 8039 10770 8073
rect 10696 8005 10716 8039
rect 10750 8005 10770 8039
rect 10696 7971 10770 8005
rect 10696 7937 10716 7971
rect 10750 7937 10770 7971
rect 10696 7903 10770 7937
rect 10696 7869 10716 7903
rect 10750 7869 10770 7903
rect 10696 7835 10770 7869
rect 10696 7801 10716 7835
rect 10750 7801 10770 7835
rect 10696 7767 10770 7801
rect 10696 7733 10716 7767
rect 10750 7733 10770 7767
rect 10696 7699 10770 7733
rect 10696 7665 10716 7699
rect 10750 7665 10770 7699
rect 10696 7631 10770 7665
rect 10696 7597 10716 7631
rect 10750 7597 10770 7631
rect 10696 7563 10770 7597
rect 10696 7529 10716 7563
rect 10750 7529 10770 7563
rect 10696 7495 10770 7529
rect 10696 7461 10716 7495
rect 10750 7461 10770 7495
rect 10696 7427 10770 7461
rect 10696 7393 10716 7427
rect 10750 7393 10770 7427
rect 10696 7359 10770 7393
rect 10696 7325 10716 7359
rect 10750 7325 10770 7359
rect 10696 7291 10770 7325
rect 10696 7257 10716 7291
rect 10750 7257 10770 7291
rect 10696 7223 10770 7257
rect 10696 7189 10716 7223
rect 10750 7189 10770 7223
rect 10696 7155 10770 7189
rect 10696 7121 10716 7155
rect 10750 7121 10770 7155
rect 10696 7087 10770 7121
rect 10696 7053 10716 7087
rect 10750 7053 10770 7087
rect 10696 7019 10770 7053
rect 10696 6985 10716 7019
rect 10750 6985 10770 7019
rect 10696 6951 10770 6985
rect 10696 6917 10716 6951
rect 10750 6917 10770 6951
rect 10696 6883 10770 6917
rect 10696 6849 10716 6883
rect 10750 6849 10770 6883
rect 10696 6815 10770 6849
rect 10696 6781 10716 6815
rect 10750 6781 10770 6815
rect 10696 6747 10770 6781
rect 10696 6713 10716 6747
rect 10750 6713 10770 6747
rect 10696 6679 10770 6713
rect 10696 6645 10716 6679
rect 10750 6645 10770 6679
rect 10696 6611 10770 6645
rect 10696 6577 10716 6611
rect 10750 6577 10770 6611
rect 10696 6543 10770 6577
rect 10696 6509 10716 6543
rect 10750 6509 10770 6543
rect 10696 6475 10770 6509
rect 10696 6441 10716 6475
rect 10750 6441 10770 6475
rect 10696 6407 10770 6441
rect 10696 6373 10716 6407
rect 10750 6373 10770 6407
rect 10696 6339 10770 6373
rect 10696 6305 10716 6339
rect 10750 6305 10770 6339
rect 10696 6271 10770 6305
rect 10696 6237 10716 6271
rect 10750 6237 10770 6271
rect 10696 6203 10770 6237
rect 10696 6169 10716 6203
rect 10750 6169 10770 6203
rect 10696 6135 10770 6169
rect 10696 6101 10716 6135
rect 10750 6101 10770 6135
rect 10696 6067 10770 6101
rect 10696 6033 10716 6067
rect 10750 6033 10770 6067
rect 10696 5999 10770 6033
rect 10696 5965 10716 5999
rect 10750 5965 10770 5999
rect 10696 5931 10770 5965
rect 10696 5897 10716 5931
rect 10750 5897 10770 5931
rect 10696 5863 10770 5897
rect 10696 5829 10716 5863
rect 10750 5829 10770 5863
rect 10696 5795 10770 5829
rect 10696 5761 10716 5795
rect 10750 5761 10770 5795
rect 10696 5727 10770 5761
rect 10696 5693 10716 5727
rect 10750 5693 10770 5727
rect 10696 5683 10770 5693
rect -134 5647 -60 5681
rect -134 5613 -114 5647
rect -80 5613 -60 5647
rect -134 5579 -60 5613
rect -134 5545 -114 5579
rect -80 5545 -60 5579
rect -134 5511 -60 5545
rect -134 5477 -114 5511
rect -80 5477 -60 5511
rect -134 5443 -60 5477
rect -134 5409 -114 5443
rect -80 5409 -60 5443
rect -134 5375 -60 5409
rect -134 5341 -114 5375
rect -80 5341 -60 5375
rect -134 5307 -60 5341
rect -134 5273 -114 5307
rect -80 5273 -60 5307
rect -134 5239 -60 5273
rect -134 5205 -114 5239
rect -80 5205 -60 5239
rect -134 5171 -60 5205
rect -134 5137 -114 5171
rect -80 5137 -60 5171
rect -134 5103 -60 5137
rect -134 5069 -114 5103
rect -80 5069 -60 5103
rect -134 5035 -60 5069
rect -134 5001 -114 5035
rect -80 5001 -60 5035
rect -134 4967 -60 5001
rect -134 4933 -114 4967
rect -80 4933 -60 4967
rect -134 4899 -60 4933
rect -134 4865 -114 4899
rect -80 4865 -60 4899
rect -134 4831 -60 4865
rect -134 4797 -114 4831
rect -80 4797 -60 4831
rect -134 4763 -60 4797
rect -134 4729 -114 4763
rect -80 4729 -60 4763
rect -134 4695 -60 4729
rect -134 4661 -114 4695
rect -80 4661 -60 4695
rect -134 4627 -60 4661
rect -134 4593 -114 4627
rect -80 4593 -60 4627
rect -134 4559 -60 4593
rect -134 4525 -114 4559
rect -80 4525 -60 4559
rect -134 4491 -60 4525
rect -134 4457 -114 4491
rect -80 4457 -60 4491
rect -134 4423 -60 4457
rect -134 4389 -114 4423
rect -80 4389 -60 4423
rect -134 4355 -60 4389
rect -134 4321 -114 4355
rect -80 4321 -60 4355
rect -134 4287 -60 4321
rect -134 4253 -114 4287
rect -80 4253 -60 4287
rect -134 4219 -60 4253
rect -134 4185 -114 4219
rect -80 4185 -60 4219
rect -134 4151 -60 4185
rect -134 4117 -114 4151
rect -80 4117 -60 4151
rect -134 4083 -60 4117
rect -134 4049 -114 4083
rect -80 4049 -60 4083
rect -134 4015 -60 4049
rect -134 3981 -114 4015
rect -80 3981 -60 4015
rect -134 3947 -60 3981
rect -134 3913 -114 3947
rect -80 3913 -60 3947
rect -134 3879 -60 3913
rect -134 3845 -114 3879
rect -80 3845 -60 3879
rect -134 3811 -60 3845
rect -134 3777 -114 3811
rect -80 3777 -60 3811
rect -134 3743 -60 3777
rect -134 3709 -114 3743
rect -80 3709 -60 3743
rect -134 3675 -60 3709
rect -134 3641 -114 3675
rect -80 3641 -60 3675
rect -134 3607 -60 3641
rect -134 3573 -114 3607
rect -80 3573 -60 3607
rect -134 3539 -60 3573
rect -134 3505 -114 3539
rect -80 3505 -60 3539
rect -134 3471 -60 3505
rect -134 3437 -114 3471
rect -80 3437 -60 3471
rect -134 3403 -60 3437
rect -134 3369 -114 3403
rect -80 3369 -60 3403
rect -134 3335 -60 3369
rect -134 3301 -114 3335
rect -80 3301 -60 3335
rect -134 3267 -60 3301
rect -134 3233 -114 3267
rect -80 3233 -60 3267
rect -134 3199 -60 3233
rect -134 3165 -114 3199
rect -80 3165 -60 3199
rect -134 3131 -60 3165
rect -134 3097 -114 3131
rect -80 3097 -60 3131
rect -134 3063 -60 3097
rect -134 3029 -114 3063
rect -80 3029 -60 3063
rect -134 2995 -60 3029
rect -134 2961 -114 2995
rect -80 2961 -60 2995
rect -134 2927 -60 2961
rect -134 2893 -114 2927
rect -80 2893 -60 2927
rect -134 2859 -60 2893
rect -134 2825 -114 2859
rect -80 2825 -60 2859
rect -134 2791 -60 2825
rect -134 2757 -114 2791
rect -80 2757 -60 2791
rect -134 2723 -60 2757
rect -134 2689 -114 2723
rect -80 2689 -60 2723
rect -134 2655 -60 2689
rect -134 2621 -114 2655
rect -80 2621 -60 2655
rect -134 2587 -60 2621
rect -134 2553 -114 2587
rect -80 2553 -60 2587
rect -134 2519 -60 2553
rect -134 2485 -114 2519
rect -80 2485 -60 2519
rect -134 2451 -60 2485
rect -134 2417 -114 2451
rect -80 2417 -60 2451
rect -134 2383 -60 2417
rect -134 2349 -114 2383
rect -80 2349 -60 2383
rect -134 2315 -60 2349
rect -134 2281 -114 2315
rect -80 2281 -60 2315
rect -134 2247 -60 2281
rect -134 2213 -114 2247
rect -80 2213 -60 2247
rect -134 2179 -60 2213
rect -134 2145 -114 2179
rect -80 2145 -60 2179
rect -134 2111 -60 2145
rect -134 2077 -114 2111
rect -80 2077 -60 2111
rect -134 2043 -60 2077
rect -134 2009 -114 2043
rect -80 2009 -60 2043
rect -134 1975 -60 2009
rect -134 1941 -114 1975
rect -80 1941 -60 1975
rect -134 1907 -60 1941
rect -134 1873 -114 1907
rect -80 1873 -60 1907
rect -134 1839 -60 1873
rect -134 1805 -114 1839
rect -80 1805 -60 1839
rect -134 1771 -60 1805
rect -134 1737 -114 1771
rect -80 1737 -60 1771
rect -134 1703 -60 1737
rect -134 1669 -114 1703
rect -80 1669 -60 1703
rect -134 1635 -60 1669
rect -134 1601 -114 1635
rect -80 1601 -60 1635
rect -134 1567 -60 1601
rect -134 1533 -114 1567
rect -80 1533 -60 1567
rect -134 1499 -60 1533
rect -134 1465 -114 1499
rect -80 1465 -60 1499
rect -134 1431 -60 1465
rect -134 1397 -114 1431
rect -80 1397 -60 1431
rect -134 1363 -60 1397
rect -134 1329 -114 1363
rect -80 1329 -60 1363
rect -134 1295 -60 1329
rect -134 1261 -114 1295
rect -80 1261 -60 1295
rect -134 1227 -60 1261
rect -134 1193 -114 1227
rect -80 1193 -60 1227
rect -134 1159 -60 1193
rect -134 1125 -114 1159
rect -80 1125 -60 1159
rect -134 1091 -60 1125
rect -134 1057 -114 1091
rect -80 1057 -60 1091
rect -134 1023 -60 1057
rect -134 989 -114 1023
rect -80 989 -60 1023
rect -134 955 -60 989
rect -134 921 -114 955
rect -80 921 -60 955
rect -134 887 -60 921
rect -134 853 -114 887
rect -80 853 -60 887
rect -134 819 -60 853
rect -134 785 -114 819
rect -80 785 -60 819
rect -134 751 -60 785
rect -134 717 -114 751
rect -80 717 -60 751
rect -134 683 -60 717
rect -134 649 -114 683
rect -80 649 -60 683
rect -134 615 -60 649
rect -134 581 -114 615
rect -80 581 -60 615
rect -134 547 -60 581
rect -134 513 -114 547
rect -80 513 -60 547
rect -134 479 -60 513
rect -134 445 -114 479
rect -80 445 -60 479
rect -134 411 -60 445
rect -134 377 -114 411
rect -80 377 -60 411
rect -134 343 -60 377
rect -134 309 -114 343
rect -80 309 -60 343
rect -134 275 -60 309
rect -134 241 -114 275
rect -80 241 -60 275
rect -134 207 -60 241
rect -134 173 -114 207
rect -80 173 -60 207
rect -134 139 -60 173
rect -134 105 -114 139
rect -80 105 -60 139
rect -134 49 -60 105
rect -134 15 -114 49
rect -80 15 -60 49
rect -134 -19 -60 15
rect -134 -53 -114 -19
rect -80 -53 -60 -19
rect -134 -87 -60 -53
rect -134 -121 -114 -87
rect -80 -121 -60 -87
rect -134 -155 -60 -121
rect -134 -189 -114 -155
rect -80 -189 -60 -155
rect -134 -223 -60 -189
rect -134 -257 -114 -223
rect -80 -257 -60 -223
rect -134 -291 -60 -257
rect -134 -325 -114 -291
rect -80 -325 -60 -291
rect -134 -359 -60 -325
rect -134 -393 -114 -359
rect -80 -393 -60 -359
rect -134 -427 -60 -393
rect -134 -461 -114 -427
rect -80 -461 -60 -427
rect -134 -495 -60 -461
rect -134 -529 -114 -495
rect -80 -529 -60 -495
rect -134 -563 -60 -529
rect -134 -597 -114 -563
rect -80 -597 -60 -563
rect -134 -631 -60 -597
rect -134 -665 -114 -631
rect -80 -665 -60 -631
rect -134 -699 -60 -665
rect -134 -733 -114 -699
rect -80 -733 -60 -699
rect -134 -767 -60 -733
rect -134 -801 -114 -767
rect -80 -801 -60 -767
rect -134 -835 -60 -801
rect -134 -869 -114 -835
rect -80 -869 -60 -835
rect -134 -903 -60 -869
rect -134 -937 -114 -903
rect -80 -937 -60 -903
rect -134 -971 -60 -937
rect -134 -1005 -114 -971
rect -80 -1005 -60 -971
rect -134 -1039 -60 -1005
rect -134 -1073 -114 -1039
rect -80 -1073 -60 -1039
rect -134 -1107 -60 -1073
rect -134 -1141 -114 -1107
rect -80 -1141 -60 -1107
rect -134 -1197 -60 -1141
rect -134 -1231 -114 -1197
rect -80 -1231 -60 -1197
rect -134 -1265 -60 -1231
rect -134 -1299 -114 -1265
rect -80 -1299 -60 -1265
rect -134 -1325 -60 -1299
rect 9496 5663 10770 5683
rect 9496 5629 9612 5663
rect 9646 5629 9680 5663
rect 9714 5629 9748 5663
rect 9782 5629 9816 5663
rect 9850 5629 9884 5663
rect 9918 5629 9952 5663
rect 9986 5629 10020 5663
rect 10054 5629 10088 5663
rect 10122 5629 10156 5663
rect 10190 5629 10224 5663
rect 10258 5629 10292 5663
rect 10326 5629 10360 5663
rect 10394 5629 10428 5663
rect 10462 5629 10496 5663
rect 10530 5629 10564 5663
rect 10598 5629 10632 5663
rect 10666 5629 10770 5663
rect 9496 5609 10770 5629
rect 9496 5571 9570 5609
rect 9496 5537 9516 5571
rect 9550 5537 9570 5571
rect 9496 5503 9570 5537
rect 9496 5469 9516 5503
rect 9550 5469 9570 5503
rect 9496 5435 9570 5469
rect 9496 5401 9516 5435
rect 9550 5401 9570 5435
rect 9496 5367 9570 5401
rect 9496 5333 9516 5367
rect 9550 5333 9570 5367
rect 9496 5299 9570 5333
rect 9496 5265 9516 5299
rect 9550 5265 9570 5299
rect 9496 5231 9570 5265
rect 9496 5197 9516 5231
rect 9550 5197 9570 5231
rect 9496 5163 9570 5197
rect 9496 5129 9516 5163
rect 9550 5129 9570 5163
rect 9496 5095 9570 5129
rect 9496 5061 9516 5095
rect 9550 5061 9570 5095
rect 9496 5027 9570 5061
rect 9496 4993 9516 5027
rect 9550 4993 9570 5027
rect 9496 4959 9570 4993
rect 9496 4925 9516 4959
rect 9550 4925 9570 4959
rect 9496 4891 9570 4925
rect 9496 4857 9516 4891
rect 9550 4857 9570 4891
rect 9496 4823 9570 4857
rect 9496 4789 9516 4823
rect 9550 4789 9570 4823
rect 9496 4755 9570 4789
rect 9496 4721 9516 4755
rect 9550 4721 9570 4755
rect 9496 4687 9570 4721
rect 9496 4653 9516 4687
rect 9550 4653 9570 4687
rect 9496 4619 9570 4653
rect 9496 4585 9516 4619
rect 9550 4585 9570 4619
rect 9496 4551 9570 4585
rect 9496 4517 9516 4551
rect 9550 4517 9570 4551
rect 9496 4483 9570 4517
rect 9496 4449 9516 4483
rect 9550 4449 9570 4483
rect 9496 4415 9570 4449
rect 9496 4381 9516 4415
rect 9550 4381 9570 4415
rect 9496 4347 9570 4381
rect 9496 4313 9516 4347
rect 9550 4313 9570 4347
rect 9496 4279 9570 4313
rect 9496 4245 9516 4279
rect 9550 4245 9570 4279
rect 9496 4211 9570 4245
rect 9496 4177 9516 4211
rect 9550 4177 9570 4211
rect 9496 4143 9570 4177
rect 9496 4109 9516 4143
rect 9550 4109 9570 4143
rect 9496 4075 9570 4109
rect 9496 4041 9516 4075
rect 9550 4041 9570 4075
rect 9496 4007 9570 4041
rect 9496 3973 9516 4007
rect 9550 3973 9570 4007
rect 9496 3939 9570 3973
rect 9496 3905 9516 3939
rect 9550 3905 9570 3939
rect 9496 3871 9570 3905
rect 9496 3837 9516 3871
rect 9550 3837 9570 3871
rect 9496 3803 9570 3837
rect 9496 3769 9516 3803
rect 9550 3769 9570 3803
rect 9496 3735 9570 3769
rect 9496 3701 9516 3735
rect 9550 3701 9570 3735
rect 9496 3667 9570 3701
rect 9496 3633 9516 3667
rect 9550 3633 9570 3667
rect 9496 3599 9570 3633
rect 9496 3565 9516 3599
rect 9550 3565 9570 3599
rect 9496 3531 9570 3565
rect 9496 3497 9516 3531
rect 9550 3497 9570 3531
rect 9496 3463 9570 3497
rect 9496 3429 9516 3463
rect 9550 3429 9570 3463
rect 9496 3395 9570 3429
rect 9496 3361 9516 3395
rect 9550 3361 9570 3395
rect 9496 3327 9570 3361
rect 9496 3293 9516 3327
rect 9550 3293 9570 3327
rect 9496 3259 9570 3293
rect 9496 3225 9516 3259
rect 9550 3225 9570 3259
rect 9496 3191 9570 3225
rect 9496 3157 9516 3191
rect 9550 3157 9570 3191
rect 9496 3123 9570 3157
rect 9496 3089 9516 3123
rect 9550 3089 9570 3123
rect 9496 3055 9570 3089
rect 9496 3021 9516 3055
rect 9550 3021 9570 3055
rect 9496 2987 9570 3021
rect 9496 2953 9516 2987
rect 9550 2953 9570 2987
rect 9496 2919 9570 2953
rect 9496 2885 9516 2919
rect 9550 2885 9570 2919
rect 9496 2851 9570 2885
rect 9496 2817 9516 2851
rect 9550 2817 9570 2851
rect 9496 2783 9570 2817
rect 9496 2749 9516 2783
rect 9550 2749 9570 2783
rect 9496 2715 9570 2749
rect 9496 2681 9516 2715
rect 9550 2681 9570 2715
rect 9496 2647 9570 2681
rect 9496 2613 9516 2647
rect 9550 2613 9570 2647
rect 9496 2579 9570 2613
rect 9496 2545 9516 2579
rect 9550 2545 9570 2579
rect 9496 2511 9570 2545
rect 9496 2477 9516 2511
rect 9550 2477 9570 2511
rect 9496 2443 9570 2477
rect 9496 2409 9516 2443
rect 9550 2409 9570 2443
rect 9496 2375 9570 2409
rect 9496 2341 9516 2375
rect 9550 2341 9570 2375
rect 9496 2307 9570 2341
rect 9496 2273 9516 2307
rect 9550 2273 9570 2307
rect 9496 2239 9570 2273
rect 9496 2205 9516 2239
rect 9550 2205 9570 2239
rect 9496 2171 9570 2205
rect 9496 2137 9516 2171
rect 9550 2137 9570 2171
rect 9496 2103 9570 2137
rect 9496 2069 9516 2103
rect 9550 2069 9570 2103
rect 9496 2035 9570 2069
rect 9496 2001 9516 2035
rect 9550 2001 9570 2035
rect 9496 1967 9570 2001
rect 9496 1933 9516 1967
rect 9550 1933 9570 1967
rect 9496 1899 9570 1933
rect 9496 1865 9516 1899
rect 9550 1865 9570 1899
rect 9496 1831 9570 1865
rect 9496 1797 9516 1831
rect 9550 1797 9570 1831
rect 9496 1763 9570 1797
rect 9496 1729 9516 1763
rect 9550 1729 9570 1763
rect 9496 1695 9570 1729
rect 9496 1661 9516 1695
rect 9550 1661 9570 1695
rect 9496 1627 9570 1661
rect 9496 1593 9516 1627
rect 9550 1593 9570 1627
rect 9496 1559 9570 1593
rect 9496 1525 9516 1559
rect 9550 1525 9570 1559
rect 9496 1491 9570 1525
rect 9496 1457 9516 1491
rect 9550 1457 9570 1491
rect 9496 1423 9570 1457
rect 9496 1389 9516 1423
rect 9550 1389 9570 1423
rect 9496 1355 9570 1389
rect 9496 1321 9516 1355
rect 9550 1321 9570 1355
rect 9496 1287 9570 1321
rect 9496 1253 9516 1287
rect 9550 1253 9570 1287
rect 9496 1219 9570 1253
rect 9496 1185 9516 1219
rect 9550 1185 9570 1219
rect 9496 1151 9570 1185
rect 9496 1117 9516 1151
rect 9550 1117 9570 1151
rect 9496 1083 9570 1117
rect 9496 1049 9516 1083
rect 9550 1049 9570 1083
rect 9496 1015 9570 1049
rect 9496 981 9516 1015
rect 9550 981 9570 1015
rect 9496 947 9570 981
rect 9496 913 9516 947
rect 9550 913 9570 947
rect 9496 879 9570 913
rect 9496 845 9516 879
rect 9550 845 9570 879
rect 9496 811 9570 845
rect 9496 777 9516 811
rect 9550 777 9570 811
rect 9496 743 9570 777
rect 9496 709 9516 743
rect 9550 709 9570 743
rect 9496 675 9570 709
rect 9496 641 9516 675
rect 9550 641 9570 675
rect 9496 607 9570 641
rect 9496 573 9516 607
rect 9550 573 9570 607
rect 9496 539 9570 573
rect 9496 505 9516 539
rect 9550 505 9570 539
rect 9496 471 9570 505
rect 9496 437 9516 471
rect 9550 437 9570 471
rect 9496 403 9570 437
rect 9496 369 9516 403
rect 9550 369 9570 403
rect 9496 335 9570 369
rect 9496 301 9516 335
rect 9550 301 9570 335
rect 9496 267 9570 301
rect 9496 233 9516 267
rect 9550 233 9570 267
rect 9496 199 9570 233
rect 9496 165 9516 199
rect 9550 165 9570 199
rect 9496 131 9570 165
rect 9496 97 9516 131
rect 9550 97 9570 131
rect 9496 41 9570 97
rect 9496 7 9516 41
rect 9550 7 9570 41
rect 9496 -27 9570 7
rect 9496 -61 9516 -27
rect 9550 -61 9570 -27
rect 9496 -95 9570 -61
rect 9496 -129 9516 -95
rect 9550 -129 9570 -95
rect 9496 -163 9570 -129
rect 9496 -197 9516 -163
rect 9550 -197 9570 -163
rect 9496 -231 9570 -197
rect 9496 -265 9516 -231
rect 9550 -265 9570 -231
rect 9496 -299 9570 -265
rect 9496 -333 9516 -299
rect 9550 -333 9570 -299
rect 9496 -367 9570 -333
rect 9496 -401 9516 -367
rect 9550 -401 9570 -367
rect 9496 -435 9570 -401
rect 9496 -469 9516 -435
rect 9550 -469 9570 -435
rect 9496 -503 9570 -469
rect 9496 -537 9516 -503
rect 9550 -537 9570 -503
rect 9496 -571 9570 -537
rect 9496 -605 9516 -571
rect 9550 -605 9570 -571
rect 9496 -639 9570 -605
rect 9496 -673 9516 -639
rect 9550 -673 9570 -639
rect 9496 -707 9570 -673
rect 9496 -741 9516 -707
rect 9550 -741 9570 -707
rect 9496 -775 9570 -741
rect 9496 -809 9516 -775
rect 9550 -809 9570 -775
rect 9496 -843 9570 -809
rect 9496 -877 9516 -843
rect 9550 -877 9570 -843
rect 9496 -911 9570 -877
rect 9496 -945 9516 -911
rect 9550 -945 9570 -911
rect 9496 -979 9570 -945
rect 9496 -1013 9516 -979
rect 9550 -1013 9570 -979
rect 9496 -1047 9570 -1013
rect 9496 -1081 9516 -1047
rect 9550 -1081 9570 -1047
rect 9496 -1115 9570 -1081
rect 9496 -1149 9516 -1115
rect 9550 -1149 9570 -1115
rect 9496 -1205 9570 -1149
rect 9496 -1239 9516 -1205
rect 9550 -1239 9570 -1205
rect 9496 -1273 9570 -1239
rect 9496 -1307 9516 -1273
rect 9550 -1307 9570 -1273
rect 9496 -1325 9570 -1307
rect -134 -1345 9570 -1325
rect -134 -1379 -30 -1345
rect 4 -1379 38 -1345
rect 72 -1379 106 -1345
rect 140 -1379 174 -1345
rect 208 -1379 242 -1345
rect 276 -1379 310 -1345
rect 344 -1379 378 -1345
rect 412 -1379 446 -1345
rect 480 -1379 514 -1345
rect 548 -1379 582 -1345
rect 616 -1379 650 -1345
rect 684 -1379 718 -1345
rect 752 -1379 786 -1345
rect 820 -1379 854 -1345
rect 888 -1379 922 -1345
rect 956 -1379 990 -1345
rect 1024 -1379 1058 -1345
rect 1092 -1379 1126 -1345
rect 1160 -1379 1194 -1345
rect 1228 -1379 1262 -1345
rect 1296 -1379 1330 -1345
rect 1364 -1379 1398 -1345
rect 1432 -1379 1466 -1345
rect 1500 -1379 1534 -1345
rect 1568 -1379 1602 -1345
rect 1636 -1379 1670 -1345
rect 1704 -1379 1738 -1345
rect 1772 -1379 1806 -1345
rect 1840 -1379 1874 -1345
rect 1908 -1379 1942 -1345
rect 1976 -1379 2010 -1345
rect 2044 -1379 2078 -1345
rect 2112 -1379 2146 -1345
rect 2180 -1379 2214 -1345
rect 2248 -1379 2282 -1345
rect 2316 -1379 2350 -1345
rect 2384 -1379 2418 -1345
rect 2452 -1379 2486 -1345
rect 2520 -1379 2554 -1345
rect 2588 -1379 2622 -1345
rect 2656 -1379 2690 -1345
rect 2724 -1379 2758 -1345
rect 2792 -1379 2826 -1345
rect 2860 -1379 2894 -1345
rect 2928 -1379 2962 -1345
rect 2996 -1379 3030 -1345
rect 3064 -1379 3098 -1345
rect 3132 -1379 3166 -1345
rect 3200 -1379 3234 -1345
rect 3268 -1379 3302 -1345
rect 3336 -1379 3370 -1345
rect 3404 -1379 3438 -1345
rect 3472 -1379 3506 -1345
rect 3540 -1379 3574 -1345
rect 3608 -1379 3642 -1345
rect 3676 -1379 3710 -1345
rect 3744 -1379 3778 -1345
rect 3812 -1379 3846 -1345
rect 3880 -1379 3914 -1345
rect 3948 -1379 3982 -1345
rect 4016 -1379 4050 -1345
rect 4084 -1379 4118 -1345
rect 4152 -1379 4186 -1345
rect 4220 -1379 4254 -1345
rect 4288 -1379 4322 -1345
rect 4356 -1379 4390 -1345
rect 4424 -1379 4458 -1345
rect 4492 -1379 4526 -1345
rect 4560 -1379 4594 -1345
rect 4628 -1379 4662 -1345
rect 4696 -1379 4730 -1345
rect 4764 -1379 4798 -1345
rect 4832 -1379 4866 -1345
rect 4900 -1379 4934 -1345
rect 4968 -1379 5002 -1345
rect 5036 -1379 5070 -1345
rect 5104 -1379 5138 -1345
rect 5172 -1379 5206 -1345
rect 5240 -1379 5274 -1345
rect 5308 -1379 5342 -1345
rect 5376 -1379 5410 -1345
rect 5444 -1379 5478 -1345
rect 5512 -1379 5546 -1345
rect 5580 -1379 5614 -1345
rect 5648 -1379 5682 -1345
rect 5716 -1379 5750 -1345
rect 5784 -1379 5818 -1345
rect 5852 -1379 5886 -1345
rect 5920 -1379 5954 -1345
rect 5988 -1379 6022 -1345
rect 6056 -1379 6090 -1345
rect 6124 -1379 6158 -1345
rect 6192 -1379 6226 -1345
rect 6260 -1379 6294 -1345
rect 6328 -1379 6362 -1345
rect 6396 -1379 6430 -1345
rect 6464 -1379 6498 -1345
rect 6532 -1379 6566 -1345
rect 6600 -1379 6634 -1345
rect 6668 -1379 6702 -1345
rect 6736 -1379 6770 -1345
rect 6804 -1379 6838 -1345
rect 6872 -1379 6906 -1345
rect 6940 -1379 6974 -1345
rect 7008 -1379 7042 -1345
rect 7076 -1379 7110 -1345
rect 7144 -1379 7178 -1345
rect 7212 -1379 7246 -1345
rect 7280 -1379 7314 -1345
rect 7348 -1379 7382 -1345
rect 7416 -1379 7450 -1345
rect 7484 -1379 7518 -1345
rect 7552 -1379 7586 -1345
rect 7620 -1379 7654 -1345
rect 7688 -1379 7722 -1345
rect 7756 -1379 7790 -1345
rect 7824 -1379 7858 -1345
rect 7892 -1379 7926 -1345
rect 7960 -1379 7994 -1345
rect 8028 -1379 8062 -1345
rect 8096 -1379 8130 -1345
rect 8164 -1379 8198 -1345
rect 8232 -1379 8266 -1345
rect 8300 -1379 8334 -1345
rect 8368 -1379 8402 -1345
rect 8436 -1379 8470 -1345
rect 8504 -1379 8538 -1345
rect 8572 -1379 8606 -1345
rect 8640 -1379 8674 -1345
rect 8708 -1379 8742 -1345
rect 8776 -1379 8810 -1345
rect 8844 -1379 8878 -1345
rect 8912 -1379 8946 -1345
rect 8980 -1379 9014 -1345
rect 9048 -1379 9082 -1345
rect 9116 -1379 9150 -1345
rect 9184 -1379 9218 -1345
rect 9252 -1379 9286 -1345
rect 9320 -1379 9354 -1345
rect 9388 -1379 9422 -1345
rect 9456 -1379 9570 -1345
rect -134 -1399 9570 -1379
<< mvnsubdiffcont >>
rect -37 10114 -3 10148
rect 31 10114 65 10148
rect 99 10114 133 10148
rect 167 10114 201 10148
rect 235 10114 269 10148
rect 303 10114 337 10148
rect 371 10114 405 10148
rect 439 10114 473 10148
rect 507 10114 541 10148
rect 575 10114 609 10148
rect 643 10114 677 10148
rect 711 10114 745 10148
rect 779 10114 813 10148
rect 847 10114 881 10148
rect 915 10114 949 10148
rect 983 10114 1017 10148
rect 1051 10114 1085 10148
rect 1119 10114 1153 10148
rect 1187 10114 1221 10148
rect 1255 10114 1289 10148
rect 1323 10114 1357 10148
rect 1391 10114 1425 10148
rect 1459 10114 1493 10148
rect 1527 10114 1561 10148
rect 1595 10114 1629 10148
rect 1663 10114 1697 10148
rect 1731 10114 1765 10148
rect 1799 10114 1833 10148
rect 1867 10114 1901 10148
rect 1935 10114 1969 10148
rect 2003 10114 2037 10148
rect 2071 10114 2105 10148
rect 2139 10114 2173 10148
rect 2207 10114 2241 10148
rect 2275 10114 2309 10148
rect 2343 10114 2377 10148
rect 2411 10114 2445 10148
rect 2479 10114 2513 10148
rect 2547 10114 2581 10148
rect 2615 10114 2649 10148
rect 2683 10114 2717 10148
rect 2751 10114 2785 10148
rect 2819 10114 2853 10148
rect 2887 10114 2921 10148
rect 2955 10114 2989 10148
rect 3023 10114 3057 10148
rect 3091 10114 3125 10148
rect 3159 10114 3193 10148
rect 3227 10114 3261 10148
rect 3295 10114 3329 10148
rect 3363 10114 3397 10148
rect 3431 10114 3465 10148
rect 3499 10114 3533 10148
rect 3567 10114 3601 10148
rect 3635 10114 3669 10148
rect 3703 10114 3737 10148
rect 3771 10114 3805 10148
rect 3839 10114 3873 10148
rect 3907 10114 3941 10148
rect 3975 10114 4009 10148
rect 4043 10114 4077 10148
rect 4111 10114 4145 10148
rect 4179 10114 4213 10148
rect 4247 10114 4281 10148
rect 4315 10114 4349 10148
rect 4383 10114 4417 10148
rect 4451 10114 4485 10148
rect 4519 10114 4553 10148
rect 4587 10114 4621 10148
rect 4655 10114 4689 10148
rect 4723 10114 4757 10148
rect 4791 10114 4825 10148
rect 4859 10114 4893 10148
rect 4927 10114 4961 10148
rect 4995 10114 5029 10148
rect 5063 10114 5097 10148
rect 5131 10114 5165 10148
rect 5199 10114 5233 10148
rect 5267 10114 5301 10148
rect 5335 10114 5369 10148
rect 5403 10114 5437 10148
rect 5471 10114 5505 10148
rect 5539 10114 5573 10148
rect 5607 10114 5641 10148
rect 5675 10114 5709 10148
rect 5743 10114 5777 10148
rect 5811 10114 5845 10148
rect 5879 10114 5913 10148
rect 5947 10114 5981 10148
rect 6015 10114 6049 10148
rect 6083 10114 6117 10148
rect 6151 10114 6185 10148
rect 6219 10114 6253 10148
rect 6287 10114 6321 10148
rect 6355 10114 6389 10148
rect 6423 10114 6457 10148
rect 6491 10114 6525 10148
rect 6559 10114 6593 10148
rect 6627 10114 6661 10148
rect 6695 10114 6729 10148
rect 6763 10114 6797 10148
rect 6831 10114 6865 10148
rect 6899 10114 6933 10148
rect 6967 10114 7001 10148
rect 7035 10114 7069 10148
rect 7103 10114 7137 10148
rect 7171 10114 7205 10148
rect 7239 10114 7273 10148
rect 7307 10114 7341 10148
rect 7375 10114 7409 10148
rect 7443 10114 7477 10148
rect 7511 10114 7545 10148
rect 7579 10114 7613 10148
rect 7647 10114 7681 10148
rect 7715 10114 7749 10148
rect 7783 10114 7817 10148
rect 7851 10114 7885 10148
rect 7919 10114 7953 10148
rect 7987 10114 8021 10148
rect 8055 10114 8089 10148
rect 8123 10114 8157 10148
rect 8191 10114 8225 10148
rect 8259 10114 8293 10148
rect 8327 10114 8361 10148
rect 8395 10114 8429 10148
rect 8463 10114 8497 10148
rect 8531 10114 8565 10148
rect 8599 10114 8633 10148
rect 8667 10114 8701 10148
rect 8735 10114 8769 10148
rect 8803 10114 8837 10148
rect 8871 10114 8905 10148
rect 8939 10114 8973 10148
rect 9007 10114 9041 10148
rect 9075 10114 9109 10148
rect 9143 10114 9177 10148
rect 9211 10114 9245 10148
rect 9279 10114 9313 10148
rect 9347 10114 9381 10148
rect 9415 10114 9449 10148
rect 9483 10114 9517 10148
rect 9551 10114 9585 10148
rect 9619 10114 9653 10148
rect 9687 10114 9721 10148
rect 9755 10114 9789 10148
rect 9823 10114 9857 10148
rect 9891 10114 9925 10148
rect 9959 10114 9993 10148
rect 10027 10114 10061 10148
rect 10095 10114 10129 10148
rect 10163 10114 10197 10148
rect 10231 10114 10265 10148
rect 10299 10114 10333 10148
rect 10367 10114 10401 10148
rect 10435 10114 10469 10148
rect 10503 10114 10537 10148
rect 10571 10114 10605 10148
rect 10639 10114 10673 10148
rect -114 10033 -80 10067
rect -114 9965 -80 9999
rect -114 9897 -80 9931
rect -114 9829 -80 9863
rect -114 9761 -80 9795
rect -114 9693 -80 9727
rect -114 9625 -80 9659
rect -114 9557 -80 9591
rect -114 9489 -80 9523
rect -114 9421 -80 9455
rect -114 9353 -80 9387
rect -114 9285 -80 9319
rect -114 9217 -80 9251
rect -114 9149 -80 9183
rect -114 9081 -80 9115
rect -114 9013 -80 9047
rect -114 8945 -80 8979
rect -114 8877 -80 8911
rect -114 8809 -80 8843
rect -114 8741 -80 8775
rect -114 8673 -80 8707
rect -114 8605 -80 8639
rect -114 8537 -80 8571
rect -114 8469 -80 8503
rect -114 8401 -80 8435
rect -114 8333 -80 8367
rect -114 8265 -80 8299
rect -114 8197 -80 8231
rect -114 8129 -80 8163
rect -114 8061 -80 8095
rect -114 7993 -80 8027
rect -114 7925 -80 7959
rect -114 7857 -80 7891
rect -114 7789 -80 7823
rect -114 7721 -80 7755
rect -114 7653 -80 7687
rect -114 7585 -80 7619
rect -114 7517 -80 7551
rect -114 7449 -80 7483
rect -114 7381 -80 7415
rect -114 7313 -80 7347
rect -114 7245 -80 7279
rect -114 7177 -80 7211
rect -114 7109 -80 7143
rect -114 7041 -80 7075
rect -114 6973 -80 7007
rect -114 6905 -80 6939
rect -114 6837 -80 6871
rect -114 6769 -80 6803
rect -114 6701 -80 6735
rect -114 6633 -80 6667
rect -114 6565 -80 6599
rect -114 6497 -80 6531
rect -114 6429 -80 6463
rect -114 6361 -80 6395
rect -114 6293 -80 6327
rect -114 6225 -80 6259
rect -114 6157 -80 6191
rect -114 6089 -80 6123
rect -114 6021 -80 6055
rect -114 5953 -80 5987
rect -114 5885 -80 5919
rect -114 5817 -80 5851
rect -114 5749 -80 5783
rect -114 5681 -80 5715
rect 10716 10045 10750 10079
rect 10716 9977 10750 10011
rect 10716 9909 10750 9943
rect 10716 9841 10750 9875
rect 10716 9773 10750 9807
rect 10716 9705 10750 9739
rect 10716 9637 10750 9671
rect 10716 9569 10750 9603
rect 10716 9501 10750 9535
rect 10716 9433 10750 9467
rect 10716 9365 10750 9399
rect 10716 9297 10750 9331
rect 10716 9229 10750 9263
rect 10716 9161 10750 9195
rect 10716 9093 10750 9127
rect 10716 9025 10750 9059
rect 10716 8957 10750 8991
rect 10716 8889 10750 8923
rect 10716 8821 10750 8855
rect 10716 8753 10750 8787
rect 10716 8685 10750 8719
rect 10716 8617 10750 8651
rect 10716 8549 10750 8583
rect 10716 8481 10750 8515
rect 10716 8413 10750 8447
rect 10716 8345 10750 8379
rect 10716 8277 10750 8311
rect 10716 8209 10750 8243
rect 10716 8141 10750 8175
rect 10716 8073 10750 8107
rect 10716 8005 10750 8039
rect 10716 7937 10750 7971
rect 10716 7869 10750 7903
rect 10716 7801 10750 7835
rect 10716 7733 10750 7767
rect 10716 7665 10750 7699
rect 10716 7597 10750 7631
rect 10716 7529 10750 7563
rect 10716 7461 10750 7495
rect 10716 7393 10750 7427
rect 10716 7325 10750 7359
rect 10716 7257 10750 7291
rect 10716 7189 10750 7223
rect 10716 7121 10750 7155
rect 10716 7053 10750 7087
rect 10716 6985 10750 7019
rect 10716 6917 10750 6951
rect 10716 6849 10750 6883
rect 10716 6781 10750 6815
rect 10716 6713 10750 6747
rect 10716 6645 10750 6679
rect 10716 6577 10750 6611
rect 10716 6509 10750 6543
rect 10716 6441 10750 6475
rect 10716 6373 10750 6407
rect 10716 6305 10750 6339
rect 10716 6237 10750 6271
rect 10716 6169 10750 6203
rect 10716 6101 10750 6135
rect 10716 6033 10750 6067
rect 10716 5965 10750 5999
rect 10716 5897 10750 5931
rect 10716 5829 10750 5863
rect 10716 5761 10750 5795
rect 10716 5693 10750 5727
rect -114 5613 -80 5647
rect -114 5545 -80 5579
rect -114 5477 -80 5511
rect -114 5409 -80 5443
rect -114 5341 -80 5375
rect -114 5273 -80 5307
rect -114 5205 -80 5239
rect -114 5137 -80 5171
rect -114 5069 -80 5103
rect -114 5001 -80 5035
rect -114 4933 -80 4967
rect -114 4865 -80 4899
rect -114 4797 -80 4831
rect -114 4729 -80 4763
rect -114 4661 -80 4695
rect -114 4593 -80 4627
rect -114 4525 -80 4559
rect -114 4457 -80 4491
rect -114 4389 -80 4423
rect -114 4321 -80 4355
rect -114 4253 -80 4287
rect -114 4185 -80 4219
rect -114 4117 -80 4151
rect -114 4049 -80 4083
rect -114 3981 -80 4015
rect -114 3913 -80 3947
rect -114 3845 -80 3879
rect -114 3777 -80 3811
rect -114 3709 -80 3743
rect -114 3641 -80 3675
rect -114 3573 -80 3607
rect -114 3505 -80 3539
rect -114 3437 -80 3471
rect -114 3369 -80 3403
rect -114 3301 -80 3335
rect -114 3233 -80 3267
rect -114 3165 -80 3199
rect -114 3097 -80 3131
rect -114 3029 -80 3063
rect -114 2961 -80 2995
rect -114 2893 -80 2927
rect -114 2825 -80 2859
rect -114 2757 -80 2791
rect -114 2689 -80 2723
rect -114 2621 -80 2655
rect -114 2553 -80 2587
rect -114 2485 -80 2519
rect -114 2417 -80 2451
rect -114 2349 -80 2383
rect -114 2281 -80 2315
rect -114 2213 -80 2247
rect -114 2145 -80 2179
rect -114 2077 -80 2111
rect -114 2009 -80 2043
rect -114 1941 -80 1975
rect -114 1873 -80 1907
rect -114 1805 -80 1839
rect -114 1737 -80 1771
rect -114 1669 -80 1703
rect -114 1601 -80 1635
rect -114 1533 -80 1567
rect -114 1465 -80 1499
rect -114 1397 -80 1431
rect -114 1329 -80 1363
rect -114 1261 -80 1295
rect -114 1193 -80 1227
rect -114 1125 -80 1159
rect -114 1057 -80 1091
rect -114 989 -80 1023
rect -114 921 -80 955
rect -114 853 -80 887
rect -114 785 -80 819
rect -114 717 -80 751
rect -114 649 -80 683
rect -114 581 -80 615
rect -114 513 -80 547
rect -114 445 -80 479
rect -114 377 -80 411
rect -114 309 -80 343
rect -114 241 -80 275
rect -114 173 -80 207
rect -114 105 -80 139
rect -114 15 -80 49
rect -114 -53 -80 -19
rect -114 -121 -80 -87
rect -114 -189 -80 -155
rect -114 -257 -80 -223
rect -114 -325 -80 -291
rect -114 -393 -80 -359
rect -114 -461 -80 -427
rect -114 -529 -80 -495
rect -114 -597 -80 -563
rect -114 -665 -80 -631
rect -114 -733 -80 -699
rect -114 -801 -80 -767
rect -114 -869 -80 -835
rect -114 -937 -80 -903
rect -114 -1005 -80 -971
rect -114 -1073 -80 -1039
rect -114 -1141 -80 -1107
rect -114 -1231 -80 -1197
rect -114 -1299 -80 -1265
rect 9612 5629 9646 5663
rect 9680 5629 9714 5663
rect 9748 5629 9782 5663
rect 9816 5629 9850 5663
rect 9884 5629 9918 5663
rect 9952 5629 9986 5663
rect 10020 5629 10054 5663
rect 10088 5629 10122 5663
rect 10156 5629 10190 5663
rect 10224 5629 10258 5663
rect 10292 5629 10326 5663
rect 10360 5629 10394 5663
rect 10428 5629 10462 5663
rect 10496 5629 10530 5663
rect 10564 5629 10598 5663
rect 10632 5629 10666 5663
rect 9516 5537 9550 5571
rect 9516 5469 9550 5503
rect 9516 5401 9550 5435
rect 9516 5333 9550 5367
rect 9516 5265 9550 5299
rect 9516 5197 9550 5231
rect 9516 5129 9550 5163
rect 9516 5061 9550 5095
rect 9516 4993 9550 5027
rect 9516 4925 9550 4959
rect 9516 4857 9550 4891
rect 9516 4789 9550 4823
rect 9516 4721 9550 4755
rect 9516 4653 9550 4687
rect 9516 4585 9550 4619
rect 9516 4517 9550 4551
rect 9516 4449 9550 4483
rect 9516 4381 9550 4415
rect 9516 4313 9550 4347
rect 9516 4245 9550 4279
rect 9516 4177 9550 4211
rect 9516 4109 9550 4143
rect 9516 4041 9550 4075
rect 9516 3973 9550 4007
rect 9516 3905 9550 3939
rect 9516 3837 9550 3871
rect 9516 3769 9550 3803
rect 9516 3701 9550 3735
rect 9516 3633 9550 3667
rect 9516 3565 9550 3599
rect 9516 3497 9550 3531
rect 9516 3429 9550 3463
rect 9516 3361 9550 3395
rect 9516 3293 9550 3327
rect 9516 3225 9550 3259
rect 9516 3157 9550 3191
rect 9516 3089 9550 3123
rect 9516 3021 9550 3055
rect 9516 2953 9550 2987
rect 9516 2885 9550 2919
rect 9516 2817 9550 2851
rect 9516 2749 9550 2783
rect 9516 2681 9550 2715
rect 9516 2613 9550 2647
rect 9516 2545 9550 2579
rect 9516 2477 9550 2511
rect 9516 2409 9550 2443
rect 9516 2341 9550 2375
rect 9516 2273 9550 2307
rect 9516 2205 9550 2239
rect 9516 2137 9550 2171
rect 9516 2069 9550 2103
rect 9516 2001 9550 2035
rect 9516 1933 9550 1967
rect 9516 1865 9550 1899
rect 9516 1797 9550 1831
rect 9516 1729 9550 1763
rect 9516 1661 9550 1695
rect 9516 1593 9550 1627
rect 9516 1525 9550 1559
rect 9516 1457 9550 1491
rect 9516 1389 9550 1423
rect 9516 1321 9550 1355
rect 9516 1253 9550 1287
rect 9516 1185 9550 1219
rect 9516 1117 9550 1151
rect 9516 1049 9550 1083
rect 9516 981 9550 1015
rect 9516 913 9550 947
rect 9516 845 9550 879
rect 9516 777 9550 811
rect 9516 709 9550 743
rect 9516 641 9550 675
rect 9516 573 9550 607
rect 9516 505 9550 539
rect 9516 437 9550 471
rect 9516 369 9550 403
rect 9516 301 9550 335
rect 9516 233 9550 267
rect 9516 165 9550 199
rect 9516 97 9550 131
rect 9516 7 9550 41
rect 9516 -61 9550 -27
rect 9516 -129 9550 -95
rect 9516 -197 9550 -163
rect 9516 -265 9550 -231
rect 9516 -333 9550 -299
rect 9516 -401 9550 -367
rect 9516 -469 9550 -435
rect 9516 -537 9550 -503
rect 9516 -605 9550 -571
rect 9516 -673 9550 -639
rect 9516 -741 9550 -707
rect 9516 -809 9550 -775
rect 9516 -877 9550 -843
rect 9516 -945 9550 -911
rect 9516 -1013 9550 -979
rect 9516 -1081 9550 -1047
rect 9516 -1149 9550 -1115
rect 9516 -1239 9550 -1205
rect 9516 -1307 9550 -1273
rect -30 -1379 4 -1345
rect 38 -1379 72 -1345
rect 106 -1379 140 -1345
rect 174 -1379 208 -1345
rect 242 -1379 276 -1345
rect 310 -1379 344 -1345
rect 378 -1379 412 -1345
rect 446 -1379 480 -1345
rect 514 -1379 548 -1345
rect 582 -1379 616 -1345
rect 650 -1379 684 -1345
rect 718 -1379 752 -1345
rect 786 -1379 820 -1345
rect 854 -1379 888 -1345
rect 922 -1379 956 -1345
rect 990 -1379 1024 -1345
rect 1058 -1379 1092 -1345
rect 1126 -1379 1160 -1345
rect 1194 -1379 1228 -1345
rect 1262 -1379 1296 -1345
rect 1330 -1379 1364 -1345
rect 1398 -1379 1432 -1345
rect 1466 -1379 1500 -1345
rect 1534 -1379 1568 -1345
rect 1602 -1379 1636 -1345
rect 1670 -1379 1704 -1345
rect 1738 -1379 1772 -1345
rect 1806 -1379 1840 -1345
rect 1874 -1379 1908 -1345
rect 1942 -1379 1976 -1345
rect 2010 -1379 2044 -1345
rect 2078 -1379 2112 -1345
rect 2146 -1379 2180 -1345
rect 2214 -1379 2248 -1345
rect 2282 -1379 2316 -1345
rect 2350 -1379 2384 -1345
rect 2418 -1379 2452 -1345
rect 2486 -1379 2520 -1345
rect 2554 -1379 2588 -1345
rect 2622 -1379 2656 -1345
rect 2690 -1379 2724 -1345
rect 2758 -1379 2792 -1345
rect 2826 -1379 2860 -1345
rect 2894 -1379 2928 -1345
rect 2962 -1379 2996 -1345
rect 3030 -1379 3064 -1345
rect 3098 -1379 3132 -1345
rect 3166 -1379 3200 -1345
rect 3234 -1379 3268 -1345
rect 3302 -1379 3336 -1345
rect 3370 -1379 3404 -1345
rect 3438 -1379 3472 -1345
rect 3506 -1379 3540 -1345
rect 3574 -1379 3608 -1345
rect 3642 -1379 3676 -1345
rect 3710 -1379 3744 -1345
rect 3778 -1379 3812 -1345
rect 3846 -1379 3880 -1345
rect 3914 -1379 3948 -1345
rect 3982 -1379 4016 -1345
rect 4050 -1379 4084 -1345
rect 4118 -1379 4152 -1345
rect 4186 -1379 4220 -1345
rect 4254 -1379 4288 -1345
rect 4322 -1379 4356 -1345
rect 4390 -1379 4424 -1345
rect 4458 -1379 4492 -1345
rect 4526 -1379 4560 -1345
rect 4594 -1379 4628 -1345
rect 4662 -1379 4696 -1345
rect 4730 -1379 4764 -1345
rect 4798 -1379 4832 -1345
rect 4866 -1379 4900 -1345
rect 4934 -1379 4968 -1345
rect 5002 -1379 5036 -1345
rect 5070 -1379 5104 -1345
rect 5138 -1379 5172 -1345
rect 5206 -1379 5240 -1345
rect 5274 -1379 5308 -1345
rect 5342 -1379 5376 -1345
rect 5410 -1379 5444 -1345
rect 5478 -1379 5512 -1345
rect 5546 -1379 5580 -1345
rect 5614 -1379 5648 -1345
rect 5682 -1379 5716 -1345
rect 5750 -1379 5784 -1345
rect 5818 -1379 5852 -1345
rect 5886 -1379 5920 -1345
rect 5954 -1379 5988 -1345
rect 6022 -1379 6056 -1345
rect 6090 -1379 6124 -1345
rect 6158 -1379 6192 -1345
rect 6226 -1379 6260 -1345
rect 6294 -1379 6328 -1345
rect 6362 -1379 6396 -1345
rect 6430 -1379 6464 -1345
rect 6498 -1379 6532 -1345
rect 6566 -1379 6600 -1345
rect 6634 -1379 6668 -1345
rect 6702 -1379 6736 -1345
rect 6770 -1379 6804 -1345
rect 6838 -1379 6872 -1345
rect 6906 -1379 6940 -1345
rect 6974 -1379 7008 -1345
rect 7042 -1379 7076 -1345
rect 7110 -1379 7144 -1345
rect 7178 -1379 7212 -1345
rect 7246 -1379 7280 -1345
rect 7314 -1379 7348 -1345
rect 7382 -1379 7416 -1345
rect 7450 -1379 7484 -1345
rect 7518 -1379 7552 -1345
rect 7586 -1379 7620 -1345
rect 7654 -1379 7688 -1345
rect 7722 -1379 7756 -1345
rect 7790 -1379 7824 -1345
rect 7858 -1379 7892 -1345
rect 7926 -1379 7960 -1345
rect 7994 -1379 8028 -1345
rect 8062 -1379 8096 -1345
rect 8130 -1379 8164 -1345
rect 8198 -1379 8232 -1345
rect 8266 -1379 8300 -1345
rect 8334 -1379 8368 -1345
rect 8402 -1379 8436 -1345
rect 8470 -1379 8504 -1345
rect 8538 -1379 8572 -1345
rect 8606 -1379 8640 -1345
rect 8674 -1379 8708 -1345
rect 8742 -1379 8776 -1345
rect 8810 -1379 8844 -1345
rect 8878 -1379 8912 -1345
rect 8946 -1379 8980 -1345
rect 9014 -1379 9048 -1345
rect 9082 -1379 9116 -1345
rect 9150 -1379 9184 -1345
rect 9218 -1379 9252 -1345
rect 9286 -1379 9320 -1345
rect 9354 -1379 9388 -1345
rect 9422 -1379 9456 -1345
<< locali >>
rect -114 10114 -37 10148
rect -3 10114 31 10148
rect 65 10114 99 10148
rect 133 10114 167 10148
rect 201 10114 235 10148
rect 269 10114 303 10148
rect 337 10114 371 10148
rect 405 10114 439 10148
rect 473 10114 507 10148
rect 541 10114 575 10148
rect 609 10114 643 10148
rect 677 10114 711 10148
rect 745 10114 779 10148
rect 813 10114 847 10148
rect 881 10114 915 10148
rect 949 10114 983 10148
rect 1017 10114 1051 10148
rect 1085 10114 1119 10148
rect 1153 10114 1187 10148
rect 1221 10114 1255 10148
rect 1289 10114 1323 10148
rect 1357 10114 1391 10148
rect 1425 10114 1459 10148
rect 1493 10114 1527 10148
rect 1561 10114 1595 10148
rect 1629 10114 1663 10148
rect 1697 10114 1731 10148
rect 1765 10114 1799 10148
rect 1833 10114 1867 10148
rect 1901 10114 1935 10148
rect 1969 10114 2003 10148
rect 2037 10114 2071 10148
rect 2105 10114 2139 10148
rect 2173 10114 2207 10148
rect 2241 10114 2275 10148
rect 2309 10114 2343 10148
rect 2377 10114 2411 10148
rect 2445 10114 2479 10148
rect 2513 10114 2547 10148
rect 2581 10114 2615 10148
rect 2649 10114 2683 10148
rect 2717 10114 2751 10148
rect 2785 10114 2819 10148
rect 2853 10114 2887 10148
rect 2921 10114 2955 10148
rect 2989 10114 3023 10148
rect 3057 10114 3091 10148
rect 3125 10114 3159 10148
rect 3193 10114 3227 10148
rect 3261 10114 3295 10148
rect 3329 10114 3363 10148
rect 3397 10114 3431 10148
rect 3465 10114 3499 10148
rect 3533 10114 3567 10148
rect 3601 10114 3635 10148
rect 3669 10114 3703 10148
rect 3737 10114 3771 10148
rect 3805 10114 3839 10148
rect 3873 10114 3907 10148
rect 3941 10114 3975 10148
rect 4009 10114 4043 10148
rect 4077 10114 4111 10148
rect 4145 10114 4179 10148
rect 4213 10114 4247 10148
rect 4281 10114 4315 10148
rect 4349 10114 4383 10148
rect 4417 10114 4451 10148
rect 4485 10114 4519 10148
rect 4553 10114 4587 10148
rect 4621 10114 4655 10148
rect 4689 10114 4723 10148
rect 4757 10114 4791 10148
rect 4825 10114 4859 10148
rect 4893 10114 4927 10148
rect 4961 10114 4995 10148
rect 5029 10114 5063 10148
rect 5097 10114 5131 10148
rect 5165 10114 5199 10148
rect 5233 10114 5267 10148
rect 5301 10114 5335 10148
rect 5369 10114 5403 10148
rect 5437 10114 5471 10148
rect 5505 10114 5539 10148
rect 5573 10114 5607 10148
rect 5641 10114 5675 10148
rect 5709 10114 5743 10148
rect 5777 10114 5811 10148
rect 5845 10114 5879 10148
rect 5913 10114 5947 10148
rect 5981 10114 6015 10148
rect 6049 10114 6083 10148
rect 6117 10114 6151 10148
rect 6185 10114 6219 10148
rect 6253 10114 6287 10148
rect 6321 10114 6355 10148
rect 6389 10114 6423 10148
rect 6457 10114 6491 10148
rect 6525 10114 6559 10148
rect 6593 10114 6627 10148
rect 6661 10114 6695 10148
rect 6729 10114 6763 10148
rect 6797 10114 6831 10148
rect 6865 10114 6899 10148
rect 6933 10114 6967 10148
rect 7001 10114 7035 10148
rect 7069 10114 7103 10148
rect 7137 10114 7171 10148
rect 7205 10114 7239 10148
rect 7273 10114 7307 10148
rect 7341 10114 7375 10148
rect 7409 10114 7443 10148
rect 7477 10114 7511 10148
rect 7545 10114 7579 10148
rect 7613 10114 7647 10148
rect 7681 10114 7715 10148
rect 7749 10114 7783 10148
rect 7817 10114 7851 10148
rect 7885 10114 7919 10148
rect 7953 10114 7987 10148
rect 8021 10114 8055 10148
rect 8089 10114 8123 10148
rect 8157 10114 8191 10148
rect 8225 10114 8259 10148
rect 8293 10114 8327 10148
rect 8361 10114 8395 10148
rect 8429 10114 8463 10148
rect 8497 10114 8531 10148
rect 8565 10114 8599 10148
rect 8633 10114 8667 10148
rect 8701 10114 8735 10148
rect 8769 10114 8803 10148
rect 8837 10114 8871 10148
rect 8905 10114 8939 10148
rect 8973 10114 9007 10148
rect 9041 10114 9075 10148
rect 9109 10114 9143 10148
rect 9177 10114 9211 10148
rect 9245 10114 9279 10148
rect 9313 10114 9347 10148
rect 9381 10114 9415 10148
rect 9449 10114 9483 10148
rect 9517 10114 9551 10148
rect 9585 10114 9619 10148
rect 9653 10114 9687 10148
rect 9721 10114 9755 10148
rect 9789 10114 9823 10148
rect 9857 10114 9891 10148
rect 9925 10114 9959 10148
rect 9993 10114 10027 10148
rect 10061 10114 10095 10148
rect 10129 10114 10163 10148
rect 10197 10114 10231 10148
rect 10265 10114 10299 10148
rect 10333 10114 10367 10148
rect 10401 10114 10435 10148
rect 10469 10114 10503 10148
rect 10537 10114 10571 10148
rect 10605 10114 10639 10148
rect 10673 10114 10750 10148
rect -114 10079 10750 10114
rect -114 10067 10716 10079
rect -80 10057 10716 10067
rect -80 10033 108 10057
rect -114 10023 108 10033
rect 142 10023 180 10057
rect 214 10023 252 10057
rect 286 10023 324 10057
rect 358 10023 396 10057
rect 430 10023 468 10057
rect 502 10023 540 10057
rect 574 10023 612 10057
rect 646 10023 684 10057
rect 718 10023 756 10057
rect 790 10023 828 10057
rect 862 10023 900 10057
rect 934 10023 972 10057
rect 1006 10023 1044 10057
rect 1078 10023 1116 10057
rect 1150 10023 1188 10057
rect 1222 10023 1260 10057
rect 1294 10023 1332 10057
rect 1366 10023 1404 10057
rect 1438 10023 1476 10057
rect 1510 10023 1548 10057
rect 1582 10023 1620 10057
rect 1654 10023 1692 10057
rect 1726 10023 1764 10057
rect 1798 10023 1836 10057
rect 1870 10023 1908 10057
rect 1942 10023 1980 10057
rect 2014 10023 2052 10057
rect 2086 10023 2124 10057
rect 2158 10023 2196 10057
rect 2230 10023 2268 10057
rect 2302 10023 2340 10057
rect 2374 10023 2412 10057
rect 2446 10023 2484 10057
rect 2518 10023 2556 10057
rect 2590 10023 2628 10057
rect 2662 10023 2700 10057
rect 2734 10023 2772 10057
rect 2806 10023 2844 10057
rect 2878 10023 2916 10057
rect 2950 10023 2988 10057
rect 3022 10023 3060 10057
rect 3094 10023 3132 10057
rect 3166 10023 3204 10057
rect 3238 10023 3276 10057
rect 3310 10023 3348 10057
rect 3382 10023 3420 10057
rect 3454 10023 3492 10057
rect 3526 10023 3564 10057
rect 3598 10023 3636 10057
rect 3670 10023 3708 10057
rect 3742 10023 3780 10057
rect 3814 10023 3852 10057
rect 3886 10023 3924 10057
rect 3958 10023 3996 10057
rect 4030 10023 4068 10057
rect 4102 10023 4140 10057
rect 4174 10023 4212 10057
rect 4246 10023 4284 10057
rect 4318 10023 4356 10057
rect 4390 10023 4428 10057
rect 4462 10023 4500 10057
rect 4534 10023 4572 10057
rect 4606 10023 4644 10057
rect 4678 10023 4716 10057
rect 4750 10023 4788 10057
rect 4822 10023 4860 10057
rect 4894 10023 4932 10057
rect 4966 10023 5004 10057
rect 5038 10023 5076 10057
rect 5110 10023 5148 10057
rect 5182 10023 5220 10057
rect 5254 10023 5292 10057
rect 5326 10023 5364 10057
rect 5398 10023 5436 10057
rect 5470 10023 5508 10057
rect 5542 10023 5580 10057
rect 5614 10023 5652 10057
rect 5686 10023 5724 10057
rect 5758 10023 5796 10057
rect 5830 10023 5868 10057
rect 5902 10023 5940 10057
rect 5974 10023 6012 10057
rect 6046 10023 6084 10057
rect 6118 10023 6156 10057
rect 6190 10023 6228 10057
rect 6262 10023 6300 10057
rect 6334 10023 6372 10057
rect 6406 10023 6444 10057
rect 6478 10023 6516 10057
rect 6550 10023 6588 10057
rect 6622 10023 6660 10057
rect 6694 10023 6732 10057
rect 6766 10023 6804 10057
rect 6838 10023 6876 10057
rect 6910 10023 6948 10057
rect 6982 10023 7020 10057
rect 7054 10023 7092 10057
rect 7126 10023 7164 10057
rect 7198 10023 7236 10057
rect 7270 10023 7308 10057
rect 7342 10023 7380 10057
rect 7414 10023 7452 10057
rect 7486 10023 7524 10057
rect 7558 10023 7596 10057
rect 7630 10023 7668 10057
rect 7702 10023 7740 10057
rect 7774 10023 7812 10057
rect 7846 10023 7884 10057
rect 7918 10023 7956 10057
rect 7990 10023 8028 10057
rect 8062 10023 8100 10057
rect 8134 10023 8172 10057
rect 8206 10023 8244 10057
rect 8278 10023 8316 10057
rect 8350 10023 8388 10057
rect 8422 10023 8460 10057
rect 8494 10023 8532 10057
rect 8566 10023 8604 10057
rect 8638 10023 8676 10057
rect 8710 10023 8748 10057
rect 8782 10023 8820 10057
rect 8854 10023 8892 10057
rect 8926 10023 8964 10057
rect 8998 10023 9036 10057
rect 9070 10023 9108 10057
rect 9142 10023 9180 10057
rect 9214 10023 9252 10057
rect 9286 10023 9324 10057
rect 9358 10023 9396 10057
rect 9430 10023 9468 10057
rect 9502 10023 9540 10057
rect 9574 10023 9612 10057
rect 9646 10023 9684 10057
rect 9718 10023 9756 10057
rect 9790 10023 9828 10057
rect 9862 10023 9900 10057
rect 9934 10023 9972 10057
rect 10006 10023 10044 10057
rect 10078 10023 10116 10057
rect 10150 10023 10188 10057
rect 10222 10023 10260 10057
rect 10294 10023 10332 10057
rect 10366 10023 10404 10057
rect 10438 10023 10476 10057
rect 10510 10045 10716 10057
rect 10510 10023 10750 10045
rect -114 10011 10750 10023
rect -114 9999 10716 10011
rect -80 9977 10716 9999
rect -80 9970 10750 9977
rect -80 9965 63 9970
rect -114 9931 63 9965
rect -80 9924 63 9931
rect -80 9897 -49 9924
rect -114 9890 -49 9897
rect -15 9890 63 9924
rect -114 9863 63 9890
rect -80 9852 63 9863
rect -80 9829 -49 9852
rect -114 9818 -49 9829
rect -15 9818 63 9852
rect -114 9795 63 9818
rect -80 9780 63 9795
rect -80 9761 -49 9780
rect -114 9746 -49 9761
rect -15 9746 63 9780
rect -114 9727 63 9746
rect -80 9708 63 9727
rect -80 9693 -49 9708
rect -114 9674 -49 9693
rect -15 9674 63 9708
rect -114 9659 63 9674
rect -80 9636 63 9659
rect -80 9625 -49 9636
rect -114 9602 -49 9625
rect -15 9602 63 9636
rect -114 9591 63 9602
rect -80 9564 63 9591
rect -80 9557 -49 9564
rect -114 9530 -49 9557
rect -15 9530 63 9564
rect -114 9523 63 9530
rect -80 9492 63 9523
rect -80 9489 -49 9492
rect -114 9458 -49 9489
rect -15 9458 63 9492
rect -114 9455 63 9458
rect -80 9421 63 9455
rect -114 9420 63 9421
rect -114 9387 -49 9420
rect -80 9386 -49 9387
rect -15 9386 63 9420
rect -80 9353 63 9386
rect -114 9348 63 9353
rect -114 9319 -49 9348
rect -80 9314 -49 9319
rect -15 9314 63 9348
rect -80 9285 63 9314
rect -114 9276 63 9285
rect -114 9251 -49 9276
rect -80 9242 -49 9251
rect -15 9242 63 9276
rect -80 9217 63 9242
rect -114 9204 63 9217
rect -114 9183 -49 9204
rect -80 9170 -49 9183
rect -15 9170 63 9204
rect -80 9149 63 9170
rect -114 9132 63 9149
rect -114 9115 -49 9132
rect -80 9098 -49 9115
rect -15 9098 63 9132
rect -80 9081 63 9098
rect -114 9060 63 9081
rect -114 9047 -49 9060
rect -80 9026 -49 9047
rect -15 9026 63 9060
rect -80 9013 63 9026
rect -114 8988 63 9013
rect -114 8979 -49 8988
rect -80 8954 -49 8979
rect -15 8954 63 8988
rect -80 8945 63 8954
rect -114 8916 63 8945
rect -114 8911 -49 8916
rect -80 8882 -49 8911
rect -15 8882 63 8916
rect -80 8877 63 8882
rect -114 8844 63 8877
rect -114 8843 -49 8844
rect -80 8810 -49 8843
rect -15 8810 63 8844
rect -80 8809 63 8810
rect -114 8775 63 8809
rect -80 8772 63 8775
rect -80 8741 -49 8772
rect -114 8738 -49 8741
rect -15 8738 63 8772
rect -114 8707 63 8738
rect -80 8700 63 8707
rect -80 8673 -49 8700
rect -114 8666 -49 8673
rect -15 8666 63 8700
rect -114 8639 63 8666
rect -80 8628 63 8639
rect -80 8605 -49 8628
rect -114 8594 -49 8605
rect -15 8594 63 8628
rect -114 8571 63 8594
rect -80 8556 63 8571
rect -80 8537 -49 8556
rect -114 8522 -49 8537
rect -15 8522 63 8556
rect -114 8503 63 8522
rect -80 8484 63 8503
rect -80 8469 -49 8484
rect -114 8450 -49 8469
rect -15 8450 63 8484
rect -114 8435 63 8450
rect -80 8412 63 8435
rect -80 8401 -49 8412
rect -114 8378 -49 8401
rect -15 8378 63 8412
rect -114 8367 63 8378
rect -80 8340 63 8367
rect -80 8333 -49 8340
rect -114 8306 -49 8333
rect -15 8306 63 8340
rect -114 8299 63 8306
rect -80 8268 63 8299
rect -80 8265 -49 8268
rect -114 8234 -49 8265
rect -15 8234 63 8268
rect -114 8231 63 8234
rect -80 8197 63 8231
rect -114 8196 63 8197
rect -114 8163 -49 8196
rect -80 8162 -49 8163
rect -15 8162 63 8196
rect -80 8129 63 8162
rect -114 8124 63 8129
rect -114 8095 -49 8124
rect -80 8090 -49 8095
rect -15 8090 63 8124
rect -80 8061 63 8090
rect -114 8052 63 8061
rect -114 8027 -49 8052
rect -80 8018 -49 8027
rect -15 8018 63 8052
rect -80 7993 63 8018
rect -114 7980 63 7993
rect -114 7959 -49 7980
rect -80 7946 -49 7959
rect -15 7946 63 7980
rect -80 7925 63 7946
rect -114 7908 63 7925
rect -114 7891 -49 7908
rect -80 7874 -49 7891
rect -15 7874 63 7908
rect -80 7857 63 7874
rect -114 7836 63 7857
rect -114 7823 -49 7836
rect -80 7802 -49 7823
rect -15 7802 63 7836
rect -80 7789 63 7802
rect -114 7764 63 7789
rect -114 7755 -49 7764
rect -80 7730 -49 7755
rect -15 7730 63 7764
rect -80 7721 63 7730
rect -114 7692 63 7721
rect -114 7687 -49 7692
rect -80 7658 -49 7687
rect -15 7658 63 7692
rect -80 7653 63 7658
rect -114 7620 63 7653
rect -114 7619 -49 7620
rect -80 7586 -49 7619
rect -15 7586 63 7620
rect -80 7585 63 7586
rect -114 7551 63 7585
rect -80 7548 63 7551
rect -80 7517 -49 7548
rect -114 7514 -49 7517
rect -15 7514 63 7548
rect -114 7483 63 7514
rect -80 7476 63 7483
rect -80 7449 -49 7476
rect -114 7442 -49 7449
rect -15 7442 63 7476
rect -114 7415 63 7442
rect -80 7404 63 7415
rect -80 7381 -49 7404
rect -114 7370 -49 7381
rect -15 7370 63 7404
rect -114 7347 63 7370
rect -80 7332 63 7347
rect -80 7313 -49 7332
rect -114 7298 -49 7313
rect -15 7298 63 7332
rect -114 7279 63 7298
rect -80 7260 63 7279
rect -80 7245 -49 7260
rect -114 7226 -49 7245
rect -15 7226 63 7260
rect -114 7211 63 7226
rect -80 7188 63 7211
rect -80 7177 -49 7188
rect -114 7154 -49 7177
rect -15 7154 63 7188
rect -114 7143 63 7154
rect -80 7116 63 7143
rect -80 7109 -49 7116
rect -114 7082 -49 7109
rect -15 7082 63 7116
rect -114 7075 63 7082
rect -80 7044 63 7075
rect -80 7041 -49 7044
rect -114 7010 -49 7041
rect -15 7010 63 7044
rect -114 7007 63 7010
rect -80 6973 63 7007
rect -114 6972 63 6973
rect -114 6939 -49 6972
rect -80 6938 -49 6939
rect -15 6938 63 6972
rect -80 6905 63 6938
rect -114 6900 63 6905
rect -114 6871 -49 6900
rect -80 6866 -49 6871
rect -15 6866 63 6900
rect -80 6837 63 6866
rect -114 6828 63 6837
rect -114 6803 -49 6828
rect -80 6794 -49 6803
rect -15 6794 63 6828
rect -80 6769 63 6794
rect -114 6756 63 6769
rect -114 6735 -49 6756
rect -80 6722 -49 6735
rect -15 6722 63 6756
rect -80 6701 63 6722
rect -114 6684 63 6701
rect -114 6667 -49 6684
rect -80 6650 -49 6667
rect -15 6650 63 6684
rect -80 6633 63 6650
rect -114 6612 63 6633
rect -114 6599 -49 6612
rect -80 6578 -49 6599
rect -15 6578 63 6612
rect -80 6565 63 6578
rect -114 6540 63 6565
rect -114 6531 -49 6540
rect -80 6506 -49 6531
rect -15 6506 63 6540
rect -80 6497 63 6506
rect -114 6468 63 6497
rect -114 6463 -49 6468
rect -80 6434 -49 6463
rect -15 6434 63 6468
rect -80 6429 63 6434
rect -114 6396 63 6429
rect -114 6395 -49 6396
rect -80 6362 -49 6395
rect -15 6362 63 6396
rect -80 6361 63 6362
rect -114 6327 63 6361
rect -80 6324 63 6327
rect -80 6293 -49 6324
rect -114 6290 -49 6293
rect -15 6290 63 6324
rect -114 6259 63 6290
rect -80 6252 63 6259
rect -80 6225 -49 6252
rect -114 6218 -49 6225
rect -15 6218 63 6252
rect -114 6191 63 6218
rect -80 6180 63 6191
rect -80 6157 -49 6180
rect -114 6146 -49 6157
rect -15 6146 63 6180
rect -114 6123 63 6146
rect -80 6108 63 6123
rect -80 6089 -49 6108
rect -114 6074 -49 6089
rect -15 6074 63 6108
rect -114 6055 63 6074
rect -80 6036 63 6055
rect -80 6021 -49 6036
rect -114 6002 -49 6021
rect -15 6002 63 6036
rect -114 5987 63 6002
rect -80 5964 63 5987
rect -80 5953 -49 5964
rect -114 5930 -49 5953
rect -15 5930 63 5964
rect -114 5919 63 5930
rect -80 5892 63 5919
rect -80 5885 -49 5892
rect -114 5858 -49 5885
rect -15 5858 63 5892
rect -114 5851 63 5858
rect -80 5820 63 5851
rect 10565 9943 10750 9970
rect 10565 9909 10716 9943
rect 10565 9880 10750 9909
rect 10565 9846 10619 9880
rect 10653 9875 10750 9880
rect 10653 9846 10716 9875
rect 10565 9841 10716 9846
rect 10565 9808 10750 9841
rect 10565 9774 10619 9808
rect 10653 9807 10750 9808
rect 10653 9774 10716 9807
rect 10565 9773 10716 9774
rect 10565 9739 10750 9773
rect 10565 9736 10716 9739
rect 10565 9702 10619 9736
rect 10653 9705 10716 9736
rect 10653 9702 10750 9705
rect 10565 9671 10750 9702
rect 10565 9664 10716 9671
rect 10565 9630 10619 9664
rect 10653 9637 10716 9664
rect 10653 9630 10750 9637
rect 10565 9603 10750 9630
rect 10565 9592 10716 9603
rect 10565 9558 10619 9592
rect 10653 9569 10716 9592
rect 10653 9558 10750 9569
rect 10565 9535 10750 9558
rect 10565 9520 10716 9535
rect 10565 9486 10619 9520
rect 10653 9501 10716 9520
rect 10653 9486 10750 9501
rect 10565 9467 10750 9486
rect 10565 9448 10716 9467
rect 10565 9414 10619 9448
rect 10653 9433 10716 9448
rect 10653 9414 10750 9433
rect 10565 9399 10750 9414
rect 10565 9376 10716 9399
rect 10565 9342 10619 9376
rect 10653 9365 10716 9376
rect 10653 9342 10750 9365
rect 10565 9331 10750 9342
rect 10565 9304 10716 9331
rect 10565 9270 10619 9304
rect 10653 9297 10716 9304
rect 10653 9270 10750 9297
rect 10565 9263 10750 9270
rect 10565 9232 10716 9263
rect 10565 9198 10619 9232
rect 10653 9229 10716 9232
rect 10653 9198 10750 9229
rect 10565 9195 10750 9198
rect 10565 9161 10716 9195
rect 10565 9160 10750 9161
rect 10565 9126 10619 9160
rect 10653 9127 10750 9160
rect 10653 9126 10716 9127
rect 10565 9093 10716 9126
rect 10565 9088 10750 9093
rect 10565 9054 10619 9088
rect 10653 9059 10750 9088
rect 10653 9054 10716 9059
rect 10565 9025 10716 9054
rect 10565 9016 10750 9025
rect 10565 8982 10619 9016
rect 10653 8991 10750 9016
rect 10653 8982 10716 8991
rect 10565 8957 10716 8982
rect 10565 8944 10750 8957
rect 10565 8910 10619 8944
rect 10653 8923 10750 8944
rect 10653 8910 10716 8923
rect 10565 8889 10716 8910
rect 10565 8872 10750 8889
rect 10565 8838 10619 8872
rect 10653 8855 10750 8872
rect 10653 8838 10716 8855
rect 10565 8821 10716 8838
rect 10565 8800 10750 8821
rect 10565 8766 10619 8800
rect 10653 8787 10750 8800
rect 10653 8766 10716 8787
rect 10565 8753 10716 8766
rect 10565 8728 10750 8753
rect 10565 8694 10619 8728
rect 10653 8719 10750 8728
rect 10653 8694 10716 8719
rect 10565 8685 10716 8694
rect 10565 8656 10750 8685
rect 10565 8622 10619 8656
rect 10653 8651 10750 8656
rect 10653 8622 10716 8651
rect 10565 8617 10716 8622
rect 10565 8584 10750 8617
rect 10565 8550 10619 8584
rect 10653 8583 10750 8584
rect 10653 8550 10716 8583
rect 10565 8549 10716 8550
rect 10565 8515 10750 8549
rect 10565 8512 10716 8515
rect 10565 8478 10619 8512
rect 10653 8481 10716 8512
rect 10653 8478 10750 8481
rect 10565 8447 10750 8478
rect 10565 8440 10716 8447
rect 10565 8406 10619 8440
rect 10653 8413 10716 8440
rect 10653 8406 10750 8413
rect 10565 8379 10750 8406
rect 10565 8368 10716 8379
rect 10565 8334 10619 8368
rect 10653 8345 10716 8368
rect 10653 8334 10750 8345
rect 10565 8311 10750 8334
rect 10565 8296 10716 8311
rect 10565 8262 10619 8296
rect 10653 8277 10716 8296
rect 10653 8262 10750 8277
rect 10565 8243 10750 8262
rect 10565 8224 10716 8243
rect 10565 8190 10619 8224
rect 10653 8209 10716 8224
rect 10653 8190 10750 8209
rect 10565 8175 10750 8190
rect 10565 8152 10716 8175
rect 10565 8118 10619 8152
rect 10653 8141 10716 8152
rect 10653 8118 10750 8141
rect 10565 8107 10750 8118
rect 10565 8080 10716 8107
rect 10565 8046 10619 8080
rect 10653 8073 10716 8080
rect 10653 8046 10750 8073
rect 10565 8039 10750 8046
rect 10565 8008 10716 8039
rect 10565 7974 10619 8008
rect 10653 8005 10716 8008
rect 10653 7974 10750 8005
rect 10565 7971 10750 7974
rect 10565 7937 10716 7971
rect 10565 7936 10750 7937
rect 10565 7902 10619 7936
rect 10653 7903 10750 7936
rect 10653 7902 10716 7903
rect 10565 7869 10716 7902
rect 10565 7864 10750 7869
rect 10565 7830 10619 7864
rect 10653 7835 10750 7864
rect 10653 7830 10716 7835
rect 10565 7801 10716 7830
rect 10565 7792 10750 7801
rect 10565 7758 10619 7792
rect 10653 7767 10750 7792
rect 10653 7758 10716 7767
rect 10565 7733 10716 7758
rect 10565 7720 10750 7733
rect 10565 7686 10619 7720
rect 10653 7699 10750 7720
rect 10653 7686 10716 7699
rect 10565 7665 10716 7686
rect 10565 7648 10750 7665
rect 10565 7614 10619 7648
rect 10653 7631 10750 7648
rect 10653 7614 10716 7631
rect 10565 7597 10716 7614
rect 10565 7576 10750 7597
rect 10565 7542 10619 7576
rect 10653 7563 10750 7576
rect 10653 7542 10716 7563
rect 10565 7529 10716 7542
rect 10565 7504 10750 7529
rect 10565 7470 10619 7504
rect 10653 7495 10750 7504
rect 10653 7470 10716 7495
rect 10565 7461 10716 7470
rect 10565 7432 10750 7461
rect 10565 7398 10619 7432
rect 10653 7427 10750 7432
rect 10653 7398 10716 7427
rect 10565 7393 10716 7398
rect 10565 7360 10750 7393
rect 10565 7326 10619 7360
rect 10653 7359 10750 7360
rect 10653 7326 10716 7359
rect 10565 7325 10716 7326
rect 10565 7291 10750 7325
rect 10565 7288 10716 7291
rect 10565 7254 10619 7288
rect 10653 7257 10716 7288
rect 10653 7254 10750 7257
rect 10565 7223 10750 7254
rect 10565 7216 10716 7223
rect 10565 7182 10619 7216
rect 10653 7189 10716 7216
rect 10653 7182 10750 7189
rect 10565 7155 10750 7182
rect 10565 7144 10716 7155
rect 10565 7110 10619 7144
rect 10653 7121 10716 7144
rect 10653 7110 10750 7121
rect 10565 7087 10750 7110
rect 10565 7072 10716 7087
rect 10565 7038 10619 7072
rect 10653 7053 10716 7072
rect 10653 7038 10750 7053
rect 10565 7019 10750 7038
rect 10565 7000 10716 7019
rect 10565 6966 10619 7000
rect 10653 6985 10716 7000
rect 10653 6966 10750 6985
rect 10565 6951 10750 6966
rect 10565 6928 10716 6951
rect 10565 6894 10619 6928
rect 10653 6917 10716 6928
rect 10653 6894 10750 6917
rect 10565 6883 10750 6894
rect 10565 6856 10716 6883
rect 10565 6822 10619 6856
rect 10653 6849 10716 6856
rect 10653 6822 10750 6849
rect 10565 6815 10750 6822
rect 10565 6784 10716 6815
rect 10565 6750 10619 6784
rect 10653 6781 10716 6784
rect 10653 6750 10750 6781
rect 10565 6747 10750 6750
rect 10565 6713 10716 6747
rect 10565 6712 10750 6713
rect 10565 6678 10619 6712
rect 10653 6679 10750 6712
rect 10653 6678 10716 6679
rect 10565 6645 10716 6678
rect 10565 6640 10750 6645
rect 10565 6606 10619 6640
rect 10653 6611 10750 6640
rect 10653 6606 10716 6611
rect 10565 6577 10716 6606
rect 10565 6568 10750 6577
rect 10565 6534 10619 6568
rect 10653 6543 10750 6568
rect 10653 6534 10716 6543
rect 10565 6509 10716 6534
rect 10565 6496 10750 6509
rect 10565 6462 10619 6496
rect 10653 6475 10750 6496
rect 10653 6462 10716 6475
rect 10565 6441 10716 6462
rect 10565 6424 10750 6441
rect 10565 6390 10619 6424
rect 10653 6407 10750 6424
rect 10653 6390 10716 6407
rect 10565 6373 10716 6390
rect 10565 6352 10750 6373
rect 10565 6318 10619 6352
rect 10653 6339 10750 6352
rect 10653 6318 10716 6339
rect 10565 6305 10716 6318
rect 10565 6280 10750 6305
rect 10565 6246 10619 6280
rect 10653 6271 10750 6280
rect 10653 6246 10716 6271
rect 10565 6237 10716 6246
rect 10565 6208 10750 6237
rect 10565 6174 10619 6208
rect 10653 6203 10750 6208
rect 10653 6174 10716 6203
rect 10565 6169 10716 6174
rect 10565 6136 10750 6169
rect 10565 6102 10619 6136
rect 10653 6135 10750 6136
rect 10653 6102 10716 6135
rect 10565 6101 10716 6102
rect 10565 6067 10750 6101
rect 10565 6064 10716 6067
rect 10565 6030 10619 6064
rect 10653 6033 10716 6064
rect 10653 6030 10750 6033
rect 10565 5999 10750 6030
rect 10565 5992 10716 5999
rect 10565 5958 10619 5992
rect 10653 5965 10716 5992
rect 10653 5958 10750 5965
rect 10565 5931 10750 5958
rect 10565 5920 10716 5931
rect 10565 5886 10619 5920
rect 10653 5897 10716 5920
rect 10653 5886 10750 5897
rect 10565 5863 10750 5886
rect 10565 5833 10716 5863
rect -80 5817 -49 5820
rect -114 5786 -49 5817
rect -15 5786 63 5820
rect -114 5783 63 5786
rect -80 5749 63 5783
rect -114 5748 63 5749
rect -114 5715 -49 5748
rect -80 5714 -49 5715
rect -15 5714 63 5748
rect -80 5681 63 5714
rect -114 5676 63 5681
rect -114 5647 -49 5676
rect -80 5642 -49 5647
rect -15 5642 63 5676
rect -80 5613 63 5642
rect -114 5604 63 5613
rect -114 5579 -49 5604
rect -80 5570 -49 5579
rect -15 5570 63 5604
rect -80 5545 63 5570
rect -114 5532 63 5545
rect -114 5511 -49 5532
rect -80 5498 -49 5511
rect -15 5498 63 5532
rect -80 5477 63 5498
rect -114 5460 63 5477
rect -114 5443 -49 5460
rect -80 5426 -49 5443
rect -15 5426 63 5460
rect -80 5409 63 5426
rect -114 5388 63 5409
rect -114 5375 -49 5388
rect -80 5354 -49 5375
rect -15 5354 63 5388
rect -80 5341 63 5354
rect -114 5316 63 5341
rect -114 5307 -49 5316
rect -80 5282 -49 5307
rect -15 5282 63 5316
rect -80 5273 63 5282
rect -114 5244 63 5273
rect -114 5239 -49 5244
rect -80 5210 -49 5239
rect -15 5210 63 5244
rect -80 5205 63 5210
rect -114 5172 63 5205
rect -114 5171 -49 5172
rect -80 5138 -49 5171
rect -15 5138 63 5172
rect -80 5137 63 5138
rect -114 5103 63 5137
rect -80 5100 63 5103
rect -80 5069 -49 5100
rect -114 5066 -49 5069
rect -15 5066 63 5100
rect -114 5035 63 5066
rect -80 5028 63 5035
rect -80 5001 -49 5028
rect -114 4994 -49 5001
rect -15 4994 63 5028
rect -114 4967 63 4994
rect -80 4956 63 4967
rect -80 4933 -49 4956
rect -114 4922 -49 4933
rect -15 4922 63 4956
rect -114 4899 63 4922
rect -80 4884 63 4899
rect -80 4865 -49 4884
rect -114 4850 -49 4865
rect -15 4850 63 4884
rect -114 4831 63 4850
rect -80 4812 63 4831
rect -80 4797 -49 4812
rect -114 4778 -49 4797
rect -15 4778 63 4812
rect -114 4763 63 4778
rect -80 4740 63 4763
rect -80 4729 -49 4740
rect -114 4706 -49 4729
rect -15 4706 63 4740
rect -114 4695 63 4706
rect -80 4668 63 4695
rect -80 4661 -49 4668
rect -114 4634 -49 4661
rect -15 4634 63 4668
rect -114 4627 63 4634
rect -80 4596 63 4627
rect -80 4593 -49 4596
rect -114 4562 -49 4593
rect -15 4562 63 4596
rect -114 4559 63 4562
rect -80 4525 63 4559
rect -114 4524 63 4525
rect -114 4491 -49 4524
rect -80 4490 -49 4491
rect -15 4490 63 4524
rect -80 4457 63 4490
rect -114 4452 63 4457
rect -114 4423 -49 4452
rect -80 4418 -49 4423
rect -15 4418 63 4452
rect -80 4389 63 4418
rect -114 4380 63 4389
rect -114 4355 -49 4380
rect -80 4346 -49 4355
rect -15 4346 63 4380
rect -80 4321 63 4346
rect -114 4308 63 4321
rect -114 4287 -49 4308
rect -80 4274 -49 4287
rect -15 4274 63 4308
rect -80 4253 63 4274
rect -114 4236 63 4253
rect -114 4219 -49 4236
rect -80 4202 -49 4219
rect -15 4202 63 4236
rect -80 4185 63 4202
rect -114 4164 63 4185
rect -114 4151 -49 4164
rect -80 4130 -49 4151
rect -15 4130 63 4164
rect -80 4117 63 4130
rect -114 4092 63 4117
rect -114 4083 -49 4092
rect -80 4058 -49 4083
rect -15 4058 63 4092
rect -80 4049 63 4058
rect -114 4020 63 4049
rect -114 4015 -49 4020
rect -80 3986 -49 4015
rect -15 3986 63 4020
rect -80 3981 63 3986
rect -114 3948 63 3981
rect -114 3947 -49 3948
rect -80 3914 -49 3947
rect -15 3914 63 3948
rect -80 3913 63 3914
rect -114 3879 63 3913
rect -80 3876 63 3879
rect -80 3845 -49 3876
rect -114 3842 -49 3845
rect -15 3842 63 3876
rect -114 3811 63 3842
rect -80 3804 63 3811
rect -80 3777 -49 3804
rect -114 3770 -49 3777
rect -15 3770 63 3804
rect -114 3743 63 3770
rect -80 3732 63 3743
rect -80 3709 -49 3732
rect -114 3698 -49 3709
rect -15 3698 63 3732
rect -114 3675 63 3698
rect -80 3660 63 3675
rect -80 3641 -49 3660
rect -114 3626 -49 3641
rect -15 3626 63 3660
rect -114 3607 63 3626
rect -80 3588 63 3607
rect -80 3573 -49 3588
rect -114 3554 -49 3573
rect -15 3554 63 3588
rect -114 3539 63 3554
rect -80 3516 63 3539
rect -80 3505 -49 3516
rect -114 3482 -49 3505
rect -15 3482 63 3516
rect -114 3471 63 3482
rect -80 3444 63 3471
rect -80 3437 -49 3444
rect -114 3410 -49 3437
rect -15 3410 63 3444
rect -114 3403 63 3410
rect -80 3372 63 3403
rect -80 3369 -49 3372
rect -114 3338 -49 3369
rect -15 3338 63 3372
rect -114 3335 63 3338
rect -80 3301 63 3335
rect -114 3300 63 3301
rect -114 3267 -49 3300
rect -80 3266 -49 3267
rect -15 3266 63 3300
rect -80 3233 63 3266
rect -114 3228 63 3233
rect -114 3199 -49 3228
rect -80 3194 -49 3199
rect -15 3194 63 3228
rect -80 3165 63 3194
rect -114 3156 63 3165
rect -114 3131 -49 3156
rect -80 3122 -49 3131
rect -15 3122 63 3156
rect -80 3097 63 3122
rect -114 3084 63 3097
rect -114 3063 -49 3084
rect -80 3050 -49 3063
rect -15 3050 63 3084
rect -80 3029 63 3050
rect -114 3012 63 3029
rect -114 2995 -49 3012
rect -80 2978 -49 2995
rect -15 2978 63 3012
rect -80 2961 63 2978
rect -114 2940 63 2961
rect -114 2927 -49 2940
rect -80 2906 -49 2927
rect -15 2906 63 2940
rect -80 2893 63 2906
rect -114 2868 63 2893
rect -114 2859 -49 2868
rect -80 2834 -49 2859
rect -15 2834 63 2868
rect -80 2825 63 2834
rect -114 2796 63 2825
rect -114 2791 -49 2796
rect -80 2762 -49 2791
rect -15 2762 63 2796
rect -80 2757 63 2762
rect -114 2724 63 2757
rect -114 2723 -49 2724
rect -80 2690 -49 2723
rect -15 2690 63 2724
rect -80 2689 63 2690
rect -114 2655 63 2689
rect -80 2652 63 2655
rect -80 2621 -49 2652
rect -114 2618 -49 2621
rect -15 2618 63 2652
rect -114 2587 63 2618
rect -80 2580 63 2587
rect -80 2553 -49 2580
rect -114 2546 -49 2553
rect -15 2546 63 2580
rect -114 2519 63 2546
rect -80 2508 63 2519
rect -80 2485 -49 2508
rect -114 2474 -49 2485
rect -15 2474 63 2508
rect -114 2451 63 2474
rect -80 2436 63 2451
rect -80 2417 -49 2436
rect -114 2402 -49 2417
rect -15 2402 63 2436
rect -114 2383 63 2402
rect -80 2364 63 2383
rect -80 2349 -49 2364
rect -114 2330 -49 2349
rect -15 2330 63 2364
rect -114 2315 63 2330
rect -80 2292 63 2315
rect -80 2281 -49 2292
rect -114 2258 -49 2281
rect -15 2258 63 2292
rect -114 2247 63 2258
rect -80 2220 63 2247
rect -80 2213 -49 2220
rect -114 2186 -49 2213
rect -15 2186 63 2220
rect -114 2179 63 2186
rect -80 2148 63 2179
rect -80 2145 -49 2148
rect -114 2114 -49 2145
rect -15 2114 63 2148
rect -114 2111 63 2114
rect -80 2077 63 2111
rect -114 2076 63 2077
rect -114 2043 -49 2076
rect -80 2042 -49 2043
rect -15 2042 63 2076
rect -80 2009 63 2042
rect -114 2004 63 2009
rect -114 1975 -49 2004
rect -80 1970 -49 1975
rect -15 1970 63 2004
rect -80 1941 63 1970
rect -114 1932 63 1941
rect -114 1907 -49 1932
rect -80 1898 -49 1907
rect -15 1898 63 1932
rect -80 1873 63 1898
rect -114 1860 63 1873
rect -114 1839 -49 1860
rect -80 1826 -49 1839
rect -15 1826 63 1860
rect -80 1805 63 1826
rect -114 1788 63 1805
rect -114 1771 -49 1788
rect -80 1754 -49 1771
rect -15 1754 63 1788
rect -80 1737 63 1754
rect -114 1716 63 1737
rect -114 1703 -49 1716
rect -80 1682 -49 1703
rect -15 1682 63 1716
rect -80 1669 63 1682
rect -114 1644 63 1669
rect -114 1635 -49 1644
rect -80 1610 -49 1635
rect -15 1610 63 1644
rect -80 1601 63 1610
rect -114 1572 63 1601
rect -114 1567 -49 1572
rect -80 1538 -49 1567
rect -15 1538 63 1572
rect -80 1533 63 1538
rect -114 1500 63 1533
rect -114 1499 -49 1500
rect -80 1466 -49 1499
rect -15 1466 63 1500
rect -80 1465 63 1466
rect -114 1431 63 1465
rect -80 1428 63 1431
rect -80 1397 -49 1428
rect -114 1394 -49 1397
rect -15 1394 63 1428
rect -114 1363 63 1394
rect -80 1356 63 1363
rect -80 1329 -49 1356
rect -114 1322 -49 1329
rect -15 1322 63 1356
rect -114 1295 63 1322
rect -80 1284 63 1295
rect -80 1261 -49 1284
rect -114 1250 -49 1261
rect -15 1250 63 1284
rect -114 1227 63 1250
rect -80 1212 63 1227
rect -80 1193 -49 1212
rect -114 1178 -49 1193
rect -15 1178 63 1212
rect -114 1159 63 1178
rect -80 1140 63 1159
rect -80 1125 -49 1140
rect -114 1106 -49 1125
rect -15 1106 63 1140
rect -114 1091 63 1106
rect -80 1068 63 1091
rect -80 1057 -49 1068
rect -114 1034 -49 1057
rect -15 1034 63 1068
rect -114 1023 63 1034
rect -80 996 63 1023
rect -80 989 -49 996
rect -114 962 -49 989
rect -15 962 63 996
rect -114 955 63 962
rect -80 924 63 955
rect -80 921 -49 924
rect -114 890 -49 921
rect -15 890 63 924
rect -114 887 63 890
rect -80 853 63 887
rect -114 852 63 853
rect -114 819 -49 852
rect -80 818 -49 819
rect -15 818 63 852
rect -80 785 63 818
rect -114 780 63 785
rect -114 751 -49 780
rect -80 746 -49 751
rect -15 746 63 780
rect -80 717 63 746
rect -114 708 63 717
rect -114 683 -49 708
rect -80 674 -49 683
rect -15 674 63 708
rect -80 649 63 674
rect -114 636 63 649
rect -114 615 -49 636
rect -80 602 -49 615
rect -15 602 63 636
rect -80 581 63 602
rect -114 564 63 581
rect -114 547 -49 564
rect -80 530 -49 547
rect -15 530 63 564
rect -80 513 63 530
rect -114 492 63 513
rect -114 479 -49 492
rect -80 458 -49 479
rect -15 458 63 492
rect -80 445 63 458
rect -114 420 63 445
rect -114 411 -49 420
rect -80 386 -49 411
rect -15 386 63 420
rect -80 377 63 386
rect -114 348 63 377
rect -114 343 -49 348
rect -80 314 -49 343
rect -15 314 63 348
rect -80 309 63 314
rect -114 276 63 309
rect -114 275 -49 276
rect -80 242 -49 275
rect -15 242 63 276
rect -80 241 63 242
rect -114 207 63 241
rect -80 204 63 207
rect -80 173 -49 204
rect -114 170 -49 173
rect -15 170 63 204
rect -114 139 63 170
rect -80 132 63 139
rect -80 105 -49 132
rect -114 98 -49 105
rect -15 98 63 132
rect -114 49 63 98
rect -80 15 63 49
rect -114 -19 63 15
rect -80 -53 63 -19
rect -114 -87 63 -53
rect -80 -121 63 -87
rect -114 -155 63 -121
rect -80 -189 63 -155
rect -114 -223 63 -189
rect -80 -257 63 -223
rect -114 -291 63 -257
rect -80 -325 63 -291
rect -114 -359 63 -325
rect -80 -393 63 -359
rect -114 -427 63 -393
rect -80 -461 63 -427
rect -114 -495 63 -461
rect -80 -529 63 -495
rect -114 -563 63 -529
rect -80 -597 63 -563
rect -114 -631 63 -597
rect -80 -665 63 -631
rect -114 -699 63 -665
rect -80 -733 63 -699
rect -114 -767 63 -733
rect -80 -801 63 -767
rect -114 -835 63 -801
rect -80 -869 63 -835
rect -114 -903 63 -869
rect -80 -937 63 -903
rect -114 -971 63 -937
rect -80 -1005 63 -971
rect -114 -1039 63 -1005
rect -80 -1073 63 -1039
rect -114 -1107 63 -1073
rect -80 -1140 63 -1107
rect -80 -1141 -49 -1140
rect -114 -1174 -49 -1141
rect -15 -1174 63 -1140
rect -114 -1190 63 -1174
rect 9360 5829 10716 5833
rect 9360 5795 10750 5829
rect 9360 5774 10716 5795
rect 9360 5740 9510 5774
rect 9544 5740 9582 5774
rect 9616 5740 9654 5774
rect 9688 5740 9726 5774
rect 9760 5740 9798 5774
rect 9832 5740 9870 5774
rect 9904 5740 9942 5774
rect 9976 5740 10014 5774
rect 10048 5740 10086 5774
rect 10120 5740 10158 5774
rect 10192 5740 10230 5774
rect 10264 5740 10302 5774
rect 10336 5740 10374 5774
rect 10408 5740 10446 5774
rect 10480 5740 10518 5774
rect 10552 5761 10716 5774
rect 10552 5740 10750 5761
rect 9360 5727 10750 5740
rect 9360 5693 10716 5727
rect 9360 5683 10750 5693
rect 9360 5649 9417 5683
rect 9451 5663 10750 5683
rect 9451 5649 9612 5663
rect 9360 5629 9612 5649
rect 9646 5629 9680 5663
rect 9714 5629 9748 5663
rect 9782 5629 9816 5663
rect 9850 5629 9884 5663
rect 9918 5629 9952 5663
rect 9986 5629 10020 5663
rect 10054 5629 10088 5663
rect 10122 5629 10156 5663
rect 10190 5629 10224 5663
rect 10258 5629 10292 5663
rect 10326 5629 10360 5663
rect 10394 5629 10428 5663
rect 10462 5629 10496 5663
rect 10530 5629 10564 5663
rect 10598 5629 10632 5663
rect 10666 5629 10750 5663
rect 9360 5611 9550 5629
rect 10565 5627 10730 5629
rect 9360 5577 9417 5611
rect 9451 5577 9550 5611
rect 9360 5571 9550 5577
rect 9360 5539 9516 5571
rect 9360 5505 9417 5539
rect 9451 5537 9516 5539
rect 9451 5505 9550 5537
rect 9360 5503 9550 5505
rect 9360 5469 9516 5503
rect 9360 5467 9550 5469
rect 9360 5433 9417 5467
rect 9451 5435 9550 5467
rect 9451 5433 9516 5435
rect 9360 5401 9516 5433
rect 9360 5395 9550 5401
rect 9360 5361 9417 5395
rect 9451 5367 9550 5395
rect 9451 5361 9516 5367
rect 9360 5333 9516 5361
rect 9360 5323 9550 5333
rect 9360 5289 9417 5323
rect 9451 5299 9550 5323
rect 9451 5289 9516 5299
rect 9360 5265 9516 5289
rect 9360 5251 9550 5265
rect 9360 5217 9417 5251
rect 9451 5231 9550 5251
rect 9451 5217 9516 5231
rect 9360 5197 9516 5217
rect 9360 5179 9550 5197
rect 9360 5145 9417 5179
rect 9451 5163 9550 5179
rect 9451 5145 9516 5163
rect 9360 5129 9516 5145
rect 9360 5107 9550 5129
rect 9360 5073 9417 5107
rect 9451 5095 9550 5107
rect 9451 5073 9516 5095
rect 9360 5061 9516 5073
rect 9360 5035 9550 5061
rect 9360 5001 9417 5035
rect 9451 5027 9550 5035
rect 9451 5001 9516 5027
rect 9360 4993 9516 5001
rect 9360 4963 9550 4993
rect 9360 4929 9417 4963
rect 9451 4959 9550 4963
rect 9451 4929 9516 4959
rect 9360 4925 9516 4929
rect 9360 4891 9550 4925
rect 9360 4857 9417 4891
rect 9451 4857 9516 4891
rect 9360 4823 9550 4857
rect 9360 4819 9516 4823
rect 9360 4785 9417 4819
rect 9451 4789 9516 4819
rect 9451 4785 9550 4789
rect 9360 4755 9550 4785
rect 9360 4747 9516 4755
rect 9360 4713 9417 4747
rect 9451 4721 9516 4747
rect 9451 4713 9550 4721
rect 9360 4687 9550 4713
rect 9360 4675 9516 4687
rect 9360 4641 9417 4675
rect 9451 4653 9516 4675
rect 9451 4641 9550 4653
rect 9360 4619 9550 4641
rect 9360 4603 9516 4619
rect 9360 4569 9417 4603
rect 9451 4585 9516 4603
rect 9451 4569 9550 4585
rect 9360 4551 9550 4569
rect 9360 4531 9516 4551
rect 9360 4497 9417 4531
rect 9451 4517 9516 4531
rect 9451 4497 9550 4517
rect 9360 4483 9550 4497
rect 9360 4459 9516 4483
rect 9360 4425 9417 4459
rect 9451 4449 9516 4459
rect 9451 4425 9550 4449
rect 9360 4415 9550 4425
rect 9360 4387 9516 4415
rect 9360 4353 9417 4387
rect 9451 4381 9516 4387
rect 9451 4353 9550 4381
rect 9360 4347 9550 4353
rect 9360 4315 9516 4347
rect 9360 4281 9417 4315
rect 9451 4313 9516 4315
rect 9451 4281 9550 4313
rect 9360 4279 9550 4281
rect 9360 4245 9516 4279
rect 9360 4243 9550 4245
rect 9360 4209 9417 4243
rect 9451 4211 9550 4243
rect 9451 4209 9516 4211
rect 9360 4177 9516 4209
rect 9360 4171 9550 4177
rect 9360 4137 9417 4171
rect 9451 4143 9550 4171
rect 9451 4137 9516 4143
rect 9360 4109 9516 4137
rect 9360 4099 9550 4109
rect 9360 4065 9417 4099
rect 9451 4075 9550 4099
rect 9451 4065 9516 4075
rect 9360 4041 9516 4065
rect 9360 4027 9550 4041
rect 9360 3993 9417 4027
rect 9451 4007 9550 4027
rect 9451 3993 9516 4007
rect 9360 3973 9516 3993
rect 9360 3955 9550 3973
rect 9360 3921 9417 3955
rect 9451 3939 9550 3955
rect 9451 3921 9516 3939
rect 9360 3905 9516 3921
rect 9360 3883 9550 3905
rect 9360 3849 9417 3883
rect 9451 3871 9550 3883
rect 9451 3849 9516 3871
rect 9360 3837 9516 3849
rect 9360 3811 9550 3837
rect 9360 3777 9417 3811
rect 9451 3803 9550 3811
rect 9451 3777 9516 3803
rect 9360 3769 9516 3777
rect 9360 3739 9550 3769
rect 10233 3809 10532 3828
rect 10233 3775 10257 3809
rect 10291 3775 10329 3809
rect 10363 3775 10401 3809
rect 10435 3775 10473 3809
rect 10507 3775 10532 3809
rect 10233 3756 10532 3775
rect 9360 3705 9417 3739
rect 9451 3735 9550 3739
rect 9451 3705 9516 3735
rect 9360 3701 9516 3705
rect 9360 3667 9550 3701
rect 9360 3633 9417 3667
rect 9451 3633 9516 3667
rect 9360 3599 9550 3633
rect 9360 3595 9516 3599
rect 9360 3561 9417 3595
rect 9451 3565 9516 3595
rect 9451 3561 9550 3565
rect 9360 3531 9550 3561
rect 9360 3523 9516 3531
rect 9360 3489 9417 3523
rect 9451 3497 9516 3523
rect 9451 3489 9550 3497
rect 9360 3463 9550 3489
rect 9360 3451 9516 3463
rect 9360 3417 9417 3451
rect 9451 3429 9516 3451
rect 9451 3417 9550 3429
rect 9360 3395 9550 3417
rect 9360 3379 9516 3395
rect 9360 3345 9417 3379
rect 9451 3361 9516 3379
rect 9451 3345 9550 3361
rect 9360 3327 9550 3345
rect 9360 3307 9516 3327
rect 9360 3273 9417 3307
rect 9451 3293 9516 3307
rect 9451 3273 9550 3293
rect 9360 3259 9550 3273
rect 9360 3235 9516 3259
rect 9360 3201 9417 3235
rect 9451 3225 9516 3235
rect 9451 3201 9550 3225
rect 9360 3191 9550 3201
rect 9360 3163 9516 3191
rect 9360 3129 9417 3163
rect 9451 3157 9516 3163
rect 11025 3288 11082 3304
rect 11025 3254 11036 3288
rect 11070 3254 11082 3288
rect 11025 3216 11082 3254
rect 11025 3182 11036 3216
rect 11070 3182 11082 3216
rect 11025 3174 11082 3182
rect 9451 3129 9550 3157
rect 9360 3123 9550 3129
rect 9360 3091 9516 3123
rect 9360 3057 9417 3091
rect 9451 3089 9516 3091
rect 9451 3057 9550 3089
rect 9360 3055 9550 3057
rect 9360 3021 9516 3055
rect 9360 3019 9550 3021
rect 9360 2985 9417 3019
rect 9451 2987 9550 3019
rect 9451 2985 9516 2987
rect 9360 2953 9516 2985
rect 9360 2947 9550 2953
rect 9360 2913 9417 2947
rect 9451 2919 9550 2947
rect 9451 2913 9516 2919
rect 9360 2885 9516 2913
rect 9360 2875 9550 2885
rect 9360 2841 9417 2875
rect 9451 2851 9550 2875
rect 9451 2841 9516 2851
rect 9360 2817 9516 2841
rect 9360 2803 9550 2817
rect 9360 2769 9417 2803
rect 9451 2783 9550 2803
rect 9451 2769 9516 2783
rect 9360 2749 9516 2769
rect 9360 2731 9550 2749
rect 9360 2697 9417 2731
rect 9451 2715 9550 2731
rect 9451 2697 9516 2715
rect 9360 2681 9516 2697
rect 9360 2659 9550 2681
rect 9360 2625 9417 2659
rect 9451 2647 9550 2659
rect 9451 2625 9516 2647
rect 9360 2613 9516 2625
rect 9360 2587 9550 2613
rect 9360 2553 9417 2587
rect 9451 2579 9550 2587
rect 9451 2553 9516 2579
rect 9360 2545 9516 2553
rect 9360 2515 9550 2545
rect 9360 2481 9417 2515
rect 9451 2511 9550 2515
rect 9451 2481 9516 2511
rect 9360 2477 9516 2481
rect 9360 2443 9550 2477
rect 9360 2409 9417 2443
rect 9451 2409 9516 2443
rect 9360 2375 9550 2409
rect 9360 2371 9516 2375
rect 9360 2337 9417 2371
rect 9451 2341 9516 2371
rect 9451 2337 9550 2341
rect 9360 2307 9550 2337
rect 9360 2299 9516 2307
rect 9360 2265 9417 2299
rect 9451 2273 9516 2299
rect 9451 2265 9550 2273
rect 9360 2239 9550 2265
rect 9360 2227 9516 2239
rect 9360 2193 9417 2227
rect 9451 2205 9516 2227
rect 9451 2193 9550 2205
rect 9360 2171 9550 2193
rect 9360 2155 9516 2171
rect 9360 2121 9417 2155
rect 9451 2137 9516 2155
rect 9451 2121 9550 2137
rect 9360 2103 9550 2121
rect 10366 2182 10476 2220
rect 10366 2148 10404 2182
rect 10438 2148 10476 2182
rect 10366 2110 10476 2148
rect 9360 2083 9516 2103
rect 9360 2049 9417 2083
rect 9451 2069 9516 2083
rect 9451 2049 9550 2069
rect 9360 2035 9550 2049
rect 9360 2011 9516 2035
rect 9360 1977 9417 2011
rect 9451 2001 9516 2011
rect 9451 1977 9550 2001
rect 9360 1967 9550 1977
rect 9360 1939 9516 1967
rect 9360 1905 9417 1939
rect 9451 1933 9516 1939
rect 9451 1905 9550 1933
rect 9360 1899 9550 1905
rect 9360 1867 9516 1899
rect 9360 1833 9417 1867
rect 9451 1865 9516 1867
rect 9451 1833 9550 1865
rect 9360 1831 9550 1833
rect 9360 1797 9516 1831
rect 9360 1795 9550 1797
rect 9360 1761 9417 1795
rect 9451 1763 9550 1795
rect 9451 1761 9516 1763
rect 9360 1729 9516 1761
rect 9360 1723 9550 1729
rect 9360 1689 9417 1723
rect 9451 1695 9550 1723
rect 9451 1689 9516 1695
rect 9360 1661 9516 1689
rect 9360 1651 9550 1661
rect 9360 1617 9417 1651
rect 9451 1627 9550 1651
rect 9451 1617 9516 1627
rect 9360 1593 9516 1617
rect 9360 1579 9550 1593
rect 9360 1545 9417 1579
rect 9451 1559 9550 1579
rect 9451 1545 9516 1559
rect 9360 1525 9516 1545
rect 9360 1507 9550 1525
rect 9360 1473 9417 1507
rect 9451 1491 9550 1507
rect 9451 1473 9516 1491
rect 9360 1457 9516 1473
rect 9360 1435 9550 1457
rect 9360 1401 9417 1435
rect 9451 1423 9550 1435
rect 9451 1401 9516 1423
rect 9360 1389 9516 1401
rect 9360 1363 9550 1389
rect 9360 1329 9417 1363
rect 9451 1355 9550 1363
rect 9451 1329 9516 1355
rect 9360 1321 9516 1329
rect 9360 1291 9550 1321
rect 9360 1257 9417 1291
rect 9451 1287 9550 1291
rect 9451 1257 9516 1287
rect 9360 1253 9516 1257
rect 9360 1219 9550 1253
rect 9360 1185 9417 1219
rect 9451 1185 9516 1219
rect 9360 1151 9550 1185
rect 9360 1147 9516 1151
rect 9360 1113 9417 1147
rect 9451 1117 9516 1147
rect 9451 1113 9550 1117
rect 9360 1083 9550 1113
rect 9360 1075 9516 1083
rect 9360 1041 9417 1075
rect 9451 1049 9516 1075
rect 9451 1041 9550 1049
rect 9360 1015 9550 1041
rect 9360 1003 9516 1015
rect 9360 969 9417 1003
rect 9451 981 9516 1003
rect 9451 969 9550 981
rect 9360 947 9550 969
rect 9360 931 9516 947
rect 9360 897 9417 931
rect 9451 913 9516 931
rect 9451 897 9550 913
rect 9360 879 9550 897
rect 9360 859 9516 879
rect 9360 825 9417 859
rect 9451 845 9516 859
rect 9451 825 9550 845
rect 9360 811 9550 825
rect 9360 787 9516 811
rect 9360 753 9417 787
rect 9451 777 9516 787
rect 9451 753 9550 777
rect 9360 743 9550 753
rect 9360 715 9516 743
rect 9360 681 9417 715
rect 9451 709 9516 715
rect 9451 681 9550 709
rect 9360 675 9550 681
rect 9360 643 9516 675
rect 9360 609 9417 643
rect 9451 641 9516 643
rect 9451 609 9550 641
rect 9360 607 9550 609
rect 9360 573 9516 607
rect 9360 571 9550 573
rect 9360 537 9417 571
rect 9451 539 9550 571
rect 9451 537 9516 539
rect 9360 505 9516 537
rect 11270 581 11384 608
rect 11270 547 11310 581
rect 11344 547 11384 581
rect 11270 510 11384 547
rect 9360 499 9550 505
rect 9360 465 9417 499
rect 9451 471 9550 499
rect 9451 465 9516 471
rect 9360 437 9516 465
rect 9360 427 9550 437
rect 9360 393 9417 427
rect 9451 403 9550 427
rect 9451 393 9516 403
rect 9360 369 9516 393
rect 9360 355 9550 369
rect 9360 321 9417 355
rect 9451 335 9550 355
rect 9451 321 9516 335
rect 9360 301 9516 321
rect 9360 283 9550 301
rect 9360 249 9417 283
rect 9451 267 9550 283
rect 9451 249 9516 267
rect 9360 233 9516 249
rect 9360 211 9550 233
rect 9360 177 9417 211
rect 9451 199 9550 211
rect 9451 177 9516 199
rect 9360 165 9516 177
rect 9360 139 9550 165
rect 9360 105 9417 139
rect 9451 131 9550 139
rect 9451 105 9516 131
rect 9360 97 9516 105
rect 9360 43 9550 97
rect 10414 349 10488 390
rect 10414 315 10434 349
rect 10468 318 10488 349
rect 10468 315 10490 318
rect 10414 277 10490 315
rect 10414 243 10434 277
rect 10468 243 10490 277
rect 10414 205 10490 243
rect 10414 171 10434 205
rect 10468 171 10490 205
rect 10414 80 10490 171
rect 9360 9 9417 43
rect 9451 41 9550 43
rect 9451 9 9516 41
rect 9360 7 9516 9
rect 10416 8 10490 80
rect 9360 -27 9550 7
rect 9360 -29 9516 -27
rect 9360 -63 9417 -29
rect 9451 -61 9516 -29
rect 9451 -63 9550 -61
rect 9360 -95 9550 -63
rect 9360 -101 9516 -95
rect 9360 -135 9417 -101
rect 9451 -129 9516 -101
rect 9451 -135 9550 -129
rect 9360 -163 9550 -135
rect 9360 -173 9516 -163
rect 9360 -207 9417 -173
rect 9451 -197 9516 -173
rect 9451 -207 9550 -197
rect 9360 -231 9550 -207
rect 9360 -245 9516 -231
rect 9360 -279 9417 -245
rect 9451 -265 9516 -245
rect 9451 -279 9550 -265
rect 9360 -299 9550 -279
rect 9360 -317 9516 -299
rect 9360 -351 9417 -317
rect 9451 -333 9516 -317
rect 9451 -351 9550 -333
rect 9360 -367 9550 -351
rect 9360 -389 9516 -367
rect 9360 -423 9417 -389
rect 9451 -401 9516 -389
rect 9451 -423 9550 -401
rect 9360 -435 9550 -423
rect 9360 -461 9516 -435
rect 9360 -495 9417 -461
rect 9451 -469 9516 -461
rect 9451 -495 9550 -469
rect 9360 -503 9550 -495
rect 9360 -533 9516 -503
rect 9360 -567 9417 -533
rect 9451 -537 9516 -533
rect 9451 -567 9550 -537
rect 9360 -571 9550 -567
rect 9360 -605 9516 -571
rect 9360 -639 9417 -605
rect 9451 -639 9550 -605
rect 9360 -673 9516 -639
rect 10424 -507 10534 -462
rect 10424 -541 10460 -507
rect 10494 -541 10534 -507
rect 10424 -579 10534 -541
rect 10424 -613 10460 -579
rect 10494 -613 10534 -579
rect 10424 -666 10534 -613
rect 9360 -677 9550 -673
rect 9360 -711 9417 -677
rect 9451 -707 9550 -677
rect 9451 -711 9516 -707
rect 9360 -741 9516 -711
rect 9360 -749 9550 -741
rect 9360 -783 9417 -749
rect 9451 -775 9550 -749
rect 9451 -783 9516 -775
rect 9360 -809 9516 -783
rect 9360 -821 9550 -809
rect 9360 -855 9417 -821
rect 9451 -843 9550 -821
rect 9451 -855 9516 -843
rect 9360 -877 9516 -855
rect 9360 -893 9550 -877
rect 9360 -927 9417 -893
rect 9451 -911 9550 -893
rect 9451 -927 9516 -911
rect 9360 -945 9516 -927
rect 9360 -965 9550 -945
rect 9360 -999 9417 -965
rect 9451 -979 9550 -965
rect 9451 -999 9516 -979
rect 9360 -1013 9516 -999
rect 9360 -1037 9550 -1013
rect 9360 -1071 9417 -1037
rect 9451 -1047 9550 -1037
rect 9451 -1071 9516 -1047
rect 9360 -1081 9516 -1071
rect 9360 -1109 9550 -1081
rect 9360 -1143 9417 -1109
rect 9451 -1115 9550 -1109
rect 9451 -1143 9516 -1115
rect 9360 -1149 9516 -1143
rect 9360 -1190 9550 -1149
rect -114 -1197 9550 -1190
rect -80 -1205 9550 -1197
rect -80 -1231 9516 -1205
rect -114 -1239 9516 -1231
rect -114 -1262 9550 -1239
rect -114 -1265 32 -1262
rect -80 -1296 32 -1265
rect 66 -1296 104 -1262
rect 138 -1296 176 -1262
rect 210 -1296 248 -1262
rect 282 -1296 320 -1262
rect 354 -1296 392 -1262
rect 426 -1296 464 -1262
rect 498 -1296 536 -1262
rect 570 -1296 608 -1262
rect 642 -1296 680 -1262
rect 714 -1296 752 -1262
rect 786 -1296 824 -1262
rect 858 -1296 896 -1262
rect 930 -1296 968 -1262
rect 1002 -1296 1040 -1262
rect 1074 -1296 1112 -1262
rect 1146 -1296 1184 -1262
rect 1218 -1296 1256 -1262
rect 1290 -1296 1328 -1262
rect 1362 -1296 1400 -1262
rect 1434 -1296 1472 -1262
rect 1506 -1296 1544 -1262
rect 1578 -1296 1616 -1262
rect 1650 -1296 1688 -1262
rect 1722 -1296 1760 -1262
rect 1794 -1296 1832 -1262
rect 1866 -1296 1904 -1262
rect 1938 -1296 1976 -1262
rect 2010 -1296 2048 -1262
rect 2082 -1296 2120 -1262
rect 2154 -1296 2192 -1262
rect 2226 -1296 2264 -1262
rect 2298 -1296 2336 -1262
rect 2370 -1296 2408 -1262
rect 2442 -1296 2480 -1262
rect 2514 -1296 2552 -1262
rect 2586 -1296 2624 -1262
rect 2658 -1296 2696 -1262
rect 2730 -1296 2768 -1262
rect 2802 -1296 2840 -1262
rect 2874 -1296 2912 -1262
rect 2946 -1296 2984 -1262
rect 3018 -1296 3056 -1262
rect 3090 -1296 3128 -1262
rect 3162 -1296 3200 -1262
rect 3234 -1296 3272 -1262
rect 3306 -1296 3344 -1262
rect 3378 -1296 3416 -1262
rect 3450 -1296 3488 -1262
rect 3522 -1296 3560 -1262
rect 3594 -1296 3632 -1262
rect 3666 -1296 3704 -1262
rect 3738 -1296 3776 -1262
rect 3810 -1296 3848 -1262
rect 3882 -1296 3920 -1262
rect 3954 -1296 3992 -1262
rect 4026 -1296 4064 -1262
rect 4098 -1296 4136 -1262
rect 4170 -1296 4208 -1262
rect 4242 -1296 4280 -1262
rect 4314 -1296 4352 -1262
rect 4386 -1296 4424 -1262
rect 4458 -1296 4496 -1262
rect 4530 -1296 4568 -1262
rect 4602 -1296 4640 -1262
rect 4674 -1296 4712 -1262
rect 4746 -1296 4784 -1262
rect 4818 -1296 4856 -1262
rect 4890 -1296 4928 -1262
rect 4962 -1296 5000 -1262
rect 5034 -1296 5072 -1262
rect 5106 -1296 5144 -1262
rect 5178 -1296 5216 -1262
rect 5250 -1296 5288 -1262
rect 5322 -1296 5360 -1262
rect 5394 -1296 5432 -1262
rect 5466 -1296 5504 -1262
rect 5538 -1296 5576 -1262
rect 5610 -1296 5648 -1262
rect 5682 -1296 5720 -1262
rect 5754 -1296 5792 -1262
rect 5826 -1296 5864 -1262
rect 5898 -1296 5936 -1262
rect 5970 -1296 6008 -1262
rect 6042 -1296 6080 -1262
rect 6114 -1296 6152 -1262
rect 6186 -1296 6224 -1262
rect 6258 -1296 6296 -1262
rect 6330 -1296 6368 -1262
rect 6402 -1296 6440 -1262
rect 6474 -1296 6512 -1262
rect 6546 -1296 6584 -1262
rect 6618 -1296 6656 -1262
rect 6690 -1296 6728 -1262
rect 6762 -1296 6800 -1262
rect 6834 -1296 6872 -1262
rect 6906 -1296 6944 -1262
rect 6978 -1296 7016 -1262
rect 7050 -1296 7088 -1262
rect 7122 -1296 7160 -1262
rect 7194 -1296 7232 -1262
rect 7266 -1296 7304 -1262
rect 7338 -1296 7376 -1262
rect 7410 -1296 7448 -1262
rect 7482 -1296 7520 -1262
rect 7554 -1296 7592 -1262
rect 7626 -1296 7664 -1262
rect 7698 -1296 7736 -1262
rect 7770 -1296 7808 -1262
rect 7842 -1296 7880 -1262
rect 7914 -1296 7952 -1262
rect 7986 -1296 8024 -1262
rect 8058 -1296 8096 -1262
rect 8130 -1296 8168 -1262
rect 8202 -1296 8240 -1262
rect 8274 -1296 8312 -1262
rect 8346 -1296 8384 -1262
rect 8418 -1296 8456 -1262
rect 8490 -1296 8528 -1262
rect 8562 -1296 8600 -1262
rect 8634 -1296 8672 -1262
rect 8706 -1296 8744 -1262
rect 8778 -1296 8816 -1262
rect 8850 -1296 8888 -1262
rect 8922 -1296 8960 -1262
rect 8994 -1296 9032 -1262
rect 9066 -1296 9104 -1262
rect 9138 -1296 9176 -1262
rect 9210 -1296 9248 -1262
rect 9282 -1296 9320 -1262
rect 9354 -1273 9550 -1262
rect 9354 -1296 9516 -1273
rect -80 -1299 9516 -1296
rect -114 -1307 9516 -1299
rect -114 -1345 9550 -1307
rect -114 -1379 -30 -1345
rect 4 -1379 38 -1345
rect 72 -1379 106 -1345
rect 140 -1379 174 -1345
rect 208 -1379 242 -1345
rect 276 -1379 310 -1345
rect 344 -1379 378 -1345
rect 412 -1379 446 -1345
rect 480 -1379 514 -1345
rect 548 -1379 582 -1345
rect 616 -1379 650 -1345
rect 684 -1379 718 -1345
rect 752 -1379 786 -1345
rect 820 -1379 854 -1345
rect 888 -1379 922 -1345
rect 956 -1379 990 -1345
rect 1024 -1379 1058 -1345
rect 1092 -1379 1126 -1345
rect 1160 -1379 1194 -1345
rect 1228 -1379 1262 -1345
rect 1296 -1379 1330 -1345
rect 1364 -1379 1398 -1345
rect 1432 -1379 1466 -1345
rect 1500 -1379 1534 -1345
rect 1568 -1379 1602 -1345
rect 1636 -1379 1670 -1345
rect 1704 -1379 1738 -1345
rect 1772 -1379 1806 -1345
rect 1840 -1379 1874 -1345
rect 1908 -1379 1942 -1345
rect 1976 -1379 2010 -1345
rect 2044 -1379 2078 -1345
rect 2112 -1379 2146 -1345
rect 2180 -1379 2214 -1345
rect 2248 -1379 2282 -1345
rect 2316 -1379 2350 -1345
rect 2384 -1379 2418 -1345
rect 2452 -1379 2486 -1345
rect 2520 -1379 2554 -1345
rect 2588 -1379 2622 -1345
rect 2656 -1379 2690 -1345
rect 2724 -1379 2758 -1345
rect 2792 -1379 2826 -1345
rect 2860 -1379 2894 -1345
rect 2928 -1379 2962 -1345
rect 2996 -1379 3030 -1345
rect 3064 -1379 3098 -1345
rect 3132 -1379 3166 -1345
rect 3200 -1379 3234 -1345
rect 3268 -1379 3302 -1345
rect 3336 -1379 3370 -1345
rect 3404 -1379 3438 -1345
rect 3472 -1379 3506 -1345
rect 3540 -1379 3574 -1345
rect 3608 -1379 3642 -1345
rect 3676 -1379 3710 -1345
rect 3744 -1379 3778 -1345
rect 3812 -1379 3846 -1345
rect 3880 -1379 3914 -1345
rect 3948 -1379 3982 -1345
rect 4016 -1379 4050 -1345
rect 4084 -1379 4118 -1345
rect 4152 -1379 4186 -1345
rect 4220 -1379 4254 -1345
rect 4288 -1379 4322 -1345
rect 4356 -1379 4390 -1345
rect 4424 -1379 4458 -1345
rect 4492 -1379 4526 -1345
rect 4560 -1379 4594 -1345
rect 4628 -1379 4662 -1345
rect 4696 -1379 4730 -1345
rect 4764 -1379 4798 -1345
rect 4832 -1379 4866 -1345
rect 4900 -1379 4934 -1345
rect 4968 -1379 5002 -1345
rect 5036 -1379 5070 -1345
rect 5104 -1379 5138 -1345
rect 5172 -1379 5206 -1345
rect 5240 -1379 5274 -1345
rect 5308 -1379 5342 -1345
rect 5376 -1379 5410 -1345
rect 5444 -1379 5478 -1345
rect 5512 -1379 5546 -1345
rect 5580 -1379 5614 -1345
rect 5648 -1379 5682 -1345
rect 5716 -1379 5750 -1345
rect 5784 -1379 5818 -1345
rect 5852 -1379 5886 -1345
rect 5920 -1379 5954 -1345
rect 5988 -1379 6022 -1345
rect 6056 -1379 6090 -1345
rect 6124 -1379 6158 -1345
rect 6192 -1379 6226 -1345
rect 6260 -1379 6294 -1345
rect 6328 -1379 6362 -1345
rect 6396 -1379 6430 -1345
rect 6464 -1379 6498 -1345
rect 6532 -1379 6566 -1345
rect 6600 -1379 6634 -1345
rect 6668 -1379 6702 -1345
rect 6736 -1379 6770 -1345
rect 6804 -1379 6838 -1345
rect 6872 -1379 6906 -1345
rect 6940 -1379 6974 -1345
rect 7008 -1379 7042 -1345
rect 7076 -1379 7110 -1345
rect 7144 -1379 7178 -1345
rect 7212 -1379 7246 -1345
rect 7280 -1379 7314 -1345
rect 7348 -1379 7382 -1345
rect 7416 -1379 7450 -1345
rect 7484 -1379 7518 -1345
rect 7552 -1379 7586 -1345
rect 7620 -1379 7654 -1345
rect 7688 -1379 7722 -1345
rect 7756 -1379 7790 -1345
rect 7824 -1379 7858 -1345
rect 7892 -1379 7926 -1345
rect 7960 -1379 7994 -1345
rect 8028 -1379 8062 -1345
rect 8096 -1379 8130 -1345
rect 8164 -1379 8198 -1345
rect 8232 -1379 8266 -1345
rect 8300 -1379 8334 -1345
rect 8368 -1379 8402 -1345
rect 8436 -1379 8470 -1345
rect 8504 -1379 8538 -1345
rect 8572 -1379 8606 -1345
rect 8640 -1379 8674 -1345
rect 8708 -1379 8742 -1345
rect 8776 -1379 8810 -1345
rect 8844 -1379 8878 -1345
rect 8912 -1379 8946 -1345
rect 8980 -1379 9014 -1345
rect 9048 -1379 9082 -1345
rect 9116 -1379 9150 -1345
rect 9184 -1379 9218 -1345
rect 9252 -1379 9286 -1345
rect 9320 -1379 9354 -1345
rect 9388 -1379 9422 -1345
rect 9456 -1379 9550 -1345
<< viali >>
rect 108 10023 142 10057
rect 180 10023 214 10057
rect 252 10023 286 10057
rect 324 10023 358 10057
rect 396 10023 430 10057
rect 468 10023 502 10057
rect 540 10023 574 10057
rect 612 10023 646 10057
rect 684 10023 718 10057
rect 756 10023 790 10057
rect 828 10023 862 10057
rect 900 10023 934 10057
rect 972 10023 1006 10057
rect 1044 10023 1078 10057
rect 1116 10023 1150 10057
rect 1188 10023 1222 10057
rect 1260 10023 1294 10057
rect 1332 10023 1366 10057
rect 1404 10023 1438 10057
rect 1476 10023 1510 10057
rect 1548 10023 1582 10057
rect 1620 10023 1654 10057
rect 1692 10023 1726 10057
rect 1764 10023 1798 10057
rect 1836 10023 1870 10057
rect 1908 10023 1942 10057
rect 1980 10023 2014 10057
rect 2052 10023 2086 10057
rect 2124 10023 2158 10057
rect 2196 10023 2230 10057
rect 2268 10023 2302 10057
rect 2340 10023 2374 10057
rect 2412 10023 2446 10057
rect 2484 10023 2518 10057
rect 2556 10023 2590 10057
rect 2628 10023 2662 10057
rect 2700 10023 2734 10057
rect 2772 10023 2806 10057
rect 2844 10023 2878 10057
rect 2916 10023 2950 10057
rect 2988 10023 3022 10057
rect 3060 10023 3094 10057
rect 3132 10023 3166 10057
rect 3204 10023 3238 10057
rect 3276 10023 3310 10057
rect 3348 10023 3382 10057
rect 3420 10023 3454 10057
rect 3492 10023 3526 10057
rect 3564 10023 3598 10057
rect 3636 10023 3670 10057
rect 3708 10023 3742 10057
rect 3780 10023 3814 10057
rect 3852 10023 3886 10057
rect 3924 10023 3958 10057
rect 3996 10023 4030 10057
rect 4068 10023 4102 10057
rect 4140 10023 4174 10057
rect 4212 10023 4246 10057
rect 4284 10023 4318 10057
rect 4356 10023 4390 10057
rect 4428 10023 4462 10057
rect 4500 10023 4534 10057
rect 4572 10023 4606 10057
rect 4644 10023 4678 10057
rect 4716 10023 4750 10057
rect 4788 10023 4822 10057
rect 4860 10023 4894 10057
rect 4932 10023 4966 10057
rect 5004 10023 5038 10057
rect 5076 10023 5110 10057
rect 5148 10023 5182 10057
rect 5220 10023 5254 10057
rect 5292 10023 5326 10057
rect 5364 10023 5398 10057
rect 5436 10023 5470 10057
rect 5508 10023 5542 10057
rect 5580 10023 5614 10057
rect 5652 10023 5686 10057
rect 5724 10023 5758 10057
rect 5796 10023 5830 10057
rect 5868 10023 5902 10057
rect 5940 10023 5974 10057
rect 6012 10023 6046 10057
rect 6084 10023 6118 10057
rect 6156 10023 6190 10057
rect 6228 10023 6262 10057
rect 6300 10023 6334 10057
rect 6372 10023 6406 10057
rect 6444 10023 6478 10057
rect 6516 10023 6550 10057
rect 6588 10023 6622 10057
rect 6660 10023 6694 10057
rect 6732 10023 6766 10057
rect 6804 10023 6838 10057
rect 6876 10023 6910 10057
rect 6948 10023 6982 10057
rect 7020 10023 7054 10057
rect 7092 10023 7126 10057
rect 7164 10023 7198 10057
rect 7236 10023 7270 10057
rect 7308 10023 7342 10057
rect 7380 10023 7414 10057
rect 7452 10023 7486 10057
rect 7524 10023 7558 10057
rect 7596 10023 7630 10057
rect 7668 10023 7702 10057
rect 7740 10023 7774 10057
rect 7812 10023 7846 10057
rect 7884 10023 7918 10057
rect 7956 10023 7990 10057
rect 8028 10023 8062 10057
rect 8100 10023 8134 10057
rect 8172 10023 8206 10057
rect 8244 10023 8278 10057
rect 8316 10023 8350 10057
rect 8388 10023 8422 10057
rect 8460 10023 8494 10057
rect 8532 10023 8566 10057
rect 8604 10023 8638 10057
rect 8676 10023 8710 10057
rect 8748 10023 8782 10057
rect 8820 10023 8854 10057
rect 8892 10023 8926 10057
rect 8964 10023 8998 10057
rect 9036 10023 9070 10057
rect 9108 10023 9142 10057
rect 9180 10023 9214 10057
rect 9252 10023 9286 10057
rect 9324 10023 9358 10057
rect 9396 10023 9430 10057
rect 9468 10023 9502 10057
rect 9540 10023 9574 10057
rect 9612 10023 9646 10057
rect 9684 10023 9718 10057
rect 9756 10023 9790 10057
rect 9828 10023 9862 10057
rect 9900 10023 9934 10057
rect 9972 10023 10006 10057
rect 10044 10023 10078 10057
rect 10116 10023 10150 10057
rect 10188 10023 10222 10057
rect 10260 10023 10294 10057
rect 10332 10023 10366 10057
rect 10404 10023 10438 10057
rect 10476 10023 10510 10057
rect -49 9890 -15 9924
rect -49 9818 -15 9852
rect -49 9746 -15 9780
rect -49 9674 -15 9708
rect -49 9602 -15 9636
rect -49 9530 -15 9564
rect -49 9458 -15 9492
rect -49 9386 -15 9420
rect -49 9314 -15 9348
rect -49 9242 -15 9276
rect -49 9170 -15 9204
rect -49 9098 -15 9132
rect -49 9026 -15 9060
rect -49 8954 -15 8988
rect -49 8882 -15 8916
rect -49 8810 -15 8844
rect -49 8738 -15 8772
rect -49 8666 -15 8700
rect -49 8594 -15 8628
rect -49 8522 -15 8556
rect -49 8450 -15 8484
rect -49 8378 -15 8412
rect -49 8306 -15 8340
rect -49 8234 -15 8268
rect -49 8162 -15 8196
rect -49 8090 -15 8124
rect -49 8018 -15 8052
rect -49 7946 -15 7980
rect -49 7874 -15 7908
rect -49 7802 -15 7836
rect -49 7730 -15 7764
rect -49 7658 -15 7692
rect -49 7586 -15 7620
rect -49 7514 -15 7548
rect -49 7442 -15 7476
rect -49 7370 -15 7404
rect -49 7298 -15 7332
rect -49 7226 -15 7260
rect -49 7154 -15 7188
rect -49 7082 -15 7116
rect -49 7010 -15 7044
rect -49 6938 -15 6972
rect -49 6866 -15 6900
rect -49 6794 -15 6828
rect -49 6722 -15 6756
rect -49 6650 -15 6684
rect -49 6578 -15 6612
rect -49 6506 -15 6540
rect -49 6434 -15 6468
rect -49 6362 -15 6396
rect -49 6290 -15 6324
rect -49 6218 -15 6252
rect -49 6146 -15 6180
rect -49 6074 -15 6108
rect -49 6002 -15 6036
rect -49 5930 -15 5964
rect -49 5858 -15 5892
rect 10619 9846 10653 9880
rect 10619 9774 10653 9808
rect 10619 9702 10653 9736
rect 10619 9630 10653 9664
rect 10619 9558 10653 9592
rect 10619 9486 10653 9520
rect 10619 9414 10653 9448
rect 10619 9342 10653 9376
rect 10619 9270 10653 9304
rect 10619 9198 10653 9232
rect 10619 9126 10653 9160
rect 10619 9054 10653 9088
rect 10619 8982 10653 9016
rect 10619 8910 10653 8944
rect 10619 8838 10653 8872
rect 10619 8766 10653 8800
rect 10619 8694 10653 8728
rect 10619 8622 10653 8656
rect 10619 8550 10653 8584
rect 10619 8478 10653 8512
rect 10619 8406 10653 8440
rect 10619 8334 10653 8368
rect 10619 8262 10653 8296
rect 10619 8190 10653 8224
rect 10619 8118 10653 8152
rect 10619 8046 10653 8080
rect 10619 7974 10653 8008
rect 10619 7902 10653 7936
rect 10619 7830 10653 7864
rect 10619 7758 10653 7792
rect 10619 7686 10653 7720
rect 10619 7614 10653 7648
rect 10619 7542 10653 7576
rect 10619 7470 10653 7504
rect 10619 7398 10653 7432
rect 10619 7326 10653 7360
rect 10619 7254 10653 7288
rect 10619 7182 10653 7216
rect 10619 7110 10653 7144
rect 10619 7038 10653 7072
rect 10619 6966 10653 7000
rect 10619 6894 10653 6928
rect 10619 6822 10653 6856
rect 10619 6750 10653 6784
rect 10619 6678 10653 6712
rect 10619 6606 10653 6640
rect 10619 6534 10653 6568
rect 10619 6462 10653 6496
rect 10619 6390 10653 6424
rect 10619 6318 10653 6352
rect 10619 6246 10653 6280
rect 10619 6174 10653 6208
rect 10619 6102 10653 6136
rect 10619 6030 10653 6064
rect 10619 5958 10653 5992
rect 10619 5886 10653 5920
rect -49 5786 -15 5820
rect -49 5714 -15 5748
rect -49 5642 -15 5676
rect -49 5570 -15 5604
rect -49 5498 -15 5532
rect -49 5426 -15 5460
rect -49 5354 -15 5388
rect -49 5282 -15 5316
rect -49 5210 -15 5244
rect -49 5138 -15 5172
rect -49 5066 -15 5100
rect -49 4994 -15 5028
rect -49 4922 -15 4956
rect -49 4850 -15 4884
rect -49 4778 -15 4812
rect -49 4706 -15 4740
rect -49 4634 -15 4668
rect -49 4562 -15 4596
rect -49 4490 -15 4524
rect -49 4418 -15 4452
rect -49 4346 -15 4380
rect -49 4274 -15 4308
rect -49 4202 -15 4236
rect -49 4130 -15 4164
rect -49 4058 -15 4092
rect -49 3986 -15 4020
rect -49 3914 -15 3948
rect -49 3842 -15 3876
rect -49 3770 -15 3804
rect -49 3698 -15 3732
rect -49 3626 -15 3660
rect -49 3554 -15 3588
rect -49 3482 -15 3516
rect -49 3410 -15 3444
rect -49 3338 -15 3372
rect -49 3266 -15 3300
rect -49 3194 -15 3228
rect -49 3122 -15 3156
rect -49 3050 -15 3084
rect -49 2978 -15 3012
rect -49 2906 -15 2940
rect -49 2834 -15 2868
rect -49 2762 -15 2796
rect -49 2690 -15 2724
rect -49 2618 -15 2652
rect -49 2546 -15 2580
rect -49 2474 -15 2508
rect -49 2402 -15 2436
rect -49 2330 -15 2364
rect -49 2258 -15 2292
rect -49 2186 -15 2220
rect -49 2114 -15 2148
rect -49 2042 -15 2076
rect -49 1970 -15 2004
rect -49 1898 -15 1932
rect -49 1826 -15 1860
rect -49 1754 -15 1788
rect -49 1682 -15 1716
rect -49 1610 -15 1644
rect -49 1538 -15 1572
rect -49 1466 -15 1500
rect -49 1394 -15 1428
rect -49 1322 -15 1356
rect -49 1250 -15 1284
rect -49 1178 -15 1212
rect -49 1106 -15 1140
rect -49 1034 -15 1068
rect -49 962 -15 996
rect -49 890 -15 924
rect -49 818 -15 852
rect -49 746 -15 780
rect -49 674 -15 708
rect -49 602 -15 636
rect -49 530 -15 564
rect -49 458 -15 492
rect -49 386 -15 420
rect -49 314 -15 348
rect -49 242 -15 276
rect -49 170 -15 204
rect -49 98 -15 132
rect -49 -1174 -15 -1140
rect 9510 5740 9544 5774
rect 9582 5740 9616 5774
rect 9654 5740 9688 5774
rect 9726 5740 9760 5774
rect 9798 5740 9832 5774
rect 9870 5740 9904 5774
rect 9942 5740 9976 5774
rect 10014 5740 10048 5774
rect 10086 5740 10120 5774
rect 10158 5740 10192 5774
rect 10230 5740 10264 5774
rect 10302 5740 10336 5774
rect 10374 5740 10408 5774
rect 10446 5740 10480 5774
rect 10518 5740 10552 5774
rect 9417 5649 9451 5683
rect 9417 5577 9451 5611
rect 9417 5505 9451 5539
rect 9417 5433 9451 5467
rect 9417 5361 9451 5395
rect 9417 5289 9451 5323
rect 9417 5217 9451 5251
rect 9417 5145 9451 5179
rect 9417 5073 9451 5107
rect 9417 5001 9451 5035
rect 9417 4929 9451 4963
rect 9417 4857 9451 4891
rect 9417 4785 9451 4819
rect 9417 4713 9451 4747
rect 9417 4641 9451 4675
rect 9417 4569 9451 4603
rect 9417 4497 9451 4531
rect 9417 4425 9451 4459
rect 9417 4353 9451 4387
rect 9417 4281 9451 4315
rect 9417 4209 9451 4243
rect 9417 4137 9451 4171
rect 9417 4065 9451 4099
rect 9417 3993 9451 4027
rect 9417 3921 9451 3955
rect 9417 3849 9451 3883
rect 9417 3777 9451 3811
rect 10257 3775 10291 3809
rect 10329 3775 10363 3809
rect 10401 3775 10435 3809
rect 10473 3775 10507 3809
rect 9417 3705 9451 3739
rect 9417 3633 9451 3667
rect 9417 3561 9451 3595
rect 9417 3489 9451 3523
rect 9417 3417 9451 3451
rect 9417 3345 9451 3379
rect 9417 3273 9451 3307
rect 9417 3201 9451 3235
rect 9417 3129 9451 3163
rect 11036 3254 11070 3288
rect 11036 3182 11070 3216
rect 9417 3057 9451 3091
rect 9417 2985 9451 3019
rect 9417 2913 9451 2947
rect 9417 2841 9451 2875
rect 9417 2769 9451 2803
rect 9417 2697 9451 2731
rect 9417 2625 9451 2659
rect 9417 2553 9451 2587
rect 9417 2481 9451 2515
rect 9417 2409 9451 2443
rect 9417 2337 9451 2371
rect 9417 2265 9451 2299
rect 9417 2193 9451 2227
rect 9417 2121 9451 2155
rect 10404 2148 10438 2182
rect 9417 2049 9451 2083
rect 9417 1977 9451 2011
rect 9417 1905 9451 1939
rect 9417 1833 9451 1867
rect 9417 1761 9451 1795
rect 9417 1689 9451 1723
rect 9417 1617 9451 1651
rect 9417 1545 9451 1579
rect 9417 1473 9451 1507
rect 9417 1401 9451 1435
rect 9417 1329 9451 1363
rect 9417 1257 9451 1291
rect 9417 1185 9451 1219
rect 9417 1113 9451 1147
rect 9417 1041 9451 1075
rect 9417 969 9451 1003
rect 9417 897 9451 931
rect 9417 825 9451 859
rect 9417 753 9451 787
rect 9417 681 9451 715
rect 9417 609 9451 643
rect 9417 537 9451 571
rect 11310 547 11344 581
rect 9417 465 9451 499
rect 9417 393 9451 427
rect 9417 321 9451 355
rect 9417 249 9451 283
rect 9417 177 9451 211
rect 9417 105 9451 139
rect 10434 315 10468 349
rect 10434 243 10468 277
rect 10434 171 10468 205
rect 9417 9 9451 43
rect 9417 -63 9451 -29
rect 9417 -135 9451 -101
rect 9417 -207 9451 -173
rect 9417 -279 9451 -245
rect 9417 -351 9451 -317
rect 9417 -423 9451 -389
rect 9417 -495 9451 -461
rect 9417 -567 9451 -533
rect 9417 -639 9451 -605
rect 10460 -541 10494 -507
rect 10460 -613 10494 -579
rect 9417 -711 9451 -677
rect 9417 -783 9451 -749
rect 9417 -855 9451 -821
rect 9417 -927 9451 -893
rect 9417 -999 9451 -965
rect 9417 -1071 9451 -1037
rect 9417 -1143 9451 -1109
rect 32 -1296 66 -1262
rect 104 -1296 138 -1262
rect 176 -1296 210 -1262
rect 248 -1296 282 -1262
rect 320 -1296 354 -1262
rect 392 -1296 426 -1262
rect 464 -1296 498 -1262
rect 536 -1296 570 -1262
rect 608 -1296 642 -1262
rect 680 -1296 714 -1262
rect 752 -1296 786 -1262
rect 824 -1296 858 -1262
rect 896 -1296 930 -1262
rect 968 -1296 1002 -1262
rect 1040 -1296 1074 -1262
rect 1112 -1296 1146 -1262
rect 1184 -1296 1218 -1262
rect 1256 -1296 1290 -1262
rect 1328 -1296 1362 -1262
rect 1400 -1296 1434 -1262
rect 1472 -1296 1506 -1262
rect 1544 -1296 1578 -1262
rect 1616 -1296 1650 -1262
rect 1688 -1296 1722 -1262
rect 1760 -1296 1794 -1262
rect 1832 -1296 1866 -1262
rect 1904 -1296 1938 -1262
rect 1976 -1296 2010 -1262
rect 2048 -1296 2082 -1262
rect 2120 -1296 2154 -1262
rect 2192 -1296 2226 -1262
rect 2264 -1296 2298 -1262
rect 2336 -1296 2370 -1262
rect 2408 -1296 2442 -1262
rect 2480 -1296 2514 -1262
rect 2552 -1296 2586 -1262
rect 2624 -1296 2658 -1262
rect 2696 -1296 2730 -1262
rect 2768 -1296 2802 -1262
rect 2840 -1296 2874 -1262
rect 2912 -1296 2946 -1262
rect 2984 -1296 3018 -1262
rect 3056 -1296 3090 -1262
rect 3128 -1296 3162 -1262
rect 3200 -1296 3234 -1262
rect 3272 -1296 3306 -1262
rect 3344 -1296 3378 -1262
rect 3416 -1296 3450 -1262
rect 3488 -1296 3522 -1262
rect 3560 -1296 3594 -1262
rect 3632 -1296 3666 -1262
rect 3704 -1296 3738 -1262
rect 3776 -1296 3810 -1262
rect 3848 -1296 3882 -1262
rect 3920 -1296 3954 -1262
rect 3992 -1296 4026 -1262
rect 4064 -1296 4098 -1262
rect 4136 -1296 4170 -1262
rect 4208 -1296 4242 -1262
rect 4280 -1296 4314 -1262
rect 4352 -1296 4386 -1262
rect 4424 -1296 4458 -1262
rect 4496 -1296 4530 -1262
rect 4568 -1296 4602 -1262
rect 4640 -1296 4674 -1262
rect 4712 -1296 4746 -1262
rect 4784 -1296 4818 -1262
rect 4856 -1296 4890 -1262
rect 4928 -1296 4962 -1262
rect 5000 -1296 5034 -1262
rect 5072 -1296 5106 -1262
rect 5144 -1296 5178 -1262
rect 5216 -1296 5250 -1262
rect 5288 -1296 5322 -1262
rect 5360 -1296 5394 -1262
rect 5432 -1296 5466 -1262
rect 5504 -1296 5538 -1262
rect 5576 -1296 5610 -1262
rect 5648 -1296 5682 -1262
rect 5720 -1296 5754 -1262
rect 5792 -1296 5826 -1262
rect 5864 -1296 5898 -1262
rect 5936 -1296 5970 -1262
rect 6008 -1296 6042 -1262
rect 6080 -1296 6114 -1262
rect 6152 -1296 6186 -1262
rect 6224 -1296 6258 -1262
rect 6296 -1296 6330 -1262
rect 6368 -1296 6402 -1262
rect 6440 -1296 6474 -1262
rect 6512 -1296 6546 -1262
rect 6584 -1296 6618 -1262
rect 6656 -1296 6690 -1262
rect 6728 -1296 6762 -1262
rect 6800 -1296 6834 -1262
rect 6872 -1296 6906 -1262
rect 6944 -1296 6978 -1262
rect 7016 -1296 7050 -1262
rect 7088 -1296 7122 -1262
rect 7160 -1296 7194 -1262
rect 7232 -1296 7266 -1262
rect 7304 -1296 7338 -1262
rect 7376 -1296 7410 -1262
rect 7448 -1296 7482 -1262
rect 7520 -1296 7554 -1262
rect 7592 -1296 7626 -1262
rect 7664 -1296 7698 -1262
rect 7736 -1296 7770 -1262
rect 7808 -1296 7842 -1262
rect 7880 -1296 7914 -1262
rect 7952 -1296 7986 -1262
rect 8024 -1296 8058 -1262
rect 8096 -1296 8130 -1262
rect 8168 -1296 8202 -1262
rect 8240 -1296 8274 -1262
rect 8312 -1296 8346 -1262
rect 8384 -1296 8418 -1262
rect 8456 -1296 8490 -1262
rect 8528 -1296 8562 -1262
rect 8600 -1296 8634 -1262
rect 8672 -1296 8706 -1262
rect 8744 -1296 8778 -1262
rect 8816 -1296 8850 -1262
rect 8888 -1296 8922 -1262
rect 8960 -1296 8994 -1262
rect 9032 -1296 9066 -1262
rect 9104 -1296 9138 -1262
rect 9176 -1296 9210 -1262
rect 9248 -1296 9282 -1262
rect 9320 -1296 9354 -1262
<< metal1 >>
rect 448 10983 4458 10998
rect 448 10931 470 10983
rect 522 10931 534 10983
rect 586 10931 598 10983
rect 650 10931 662 10983
rect 714 10931 726 10983
rect 778 10931 790 10983
rect 842 10931 854 10983
rect 906 10931 918 10983
rect 970 10931 982 10983
rect 1034 10931 1046 10983
rect 1098 10931 1110 10983
rect 1162 10931 1174 10983
rect 1226 10931 1238 10983
rect 1290 10931 1302 10983
rect 1354 10931 1366 10983
rect 1418 10931 1430 10983
rect 1482 10931 1494 10983
rect 1546 10931 1558 10983
rect 1610 10931 1622 10983
rect 1674 10931 1686 10983
rect 1738 10931 1750 10983
rect 1802 10931 1814 10983
rect 1866 10931 1878 10983
rect 1930 10931 1942 10983
rect 1994 10931 2006 10983
rect 2058 10931 2070 10983
rect 2122 10931 2134 10983
rect 2186 10931 2198 10983
rect 2250 10931 2262 10983
rect 2314 10931 2326 10983
rect 2378 10931 2390 10983
rect 2442 10931 2454 10983
rect 2506 10931 2518 10983
rect 2570 10931 2582 10983
rect 2634 10931 2646 10983
rect 2698 10931 2710 10983
rect 2762 10931 2774 10983
rect 2826 10931 2838 10983
rect 2890 10931 2902 10983
rect 2954 10931 2966 10983
rect 3018 10931 3030 10983
rect 3082 10931 3094 10983
rect 3146 10931 3158 10983
rect 3210 10931 3222 10983
rect 3274 10931 3286 10983
rect 3338 10931 3350 10983
rect 3402 10931 3414 10983
rect 3466 10931 3478 10983
rect 3530 10931 3542 10983
rect 3594 10931 3606 10983
rect 3658 10931 3670 10983
rect 3722 10931 3734 10983
rect 3786 10931 3798 10983
rect 3850 10931 3862 10983
rect 3914 10931 3926 10983
rect 3978 10931 3990 10983
rect 4042 10931 4054 10983
rect 4106 10931 4118 10983
rect 4170 10931 4182 10983
rect 4234 10931 4246 10983
rect 4298 10931 4310 10983
rect 4362 10931 4374 10983
rect 4426 10931 4458 10983
rect 448 10910 4458 10931
rect -200 10760 270 10802
rect -200 10644 -172 10760
rect 200 10644 270 10760
rect -200 10602 270 10644
rect 4492 10788 4758 10812
rect 4492 10544 4535 10788
rect 4715 10544 4758 10788
rect 4492 10514 4758 10544
rect 452 10453 4462 10472
rect 452 10401 486 10453
rect 538 10401 550 10453
rect 602 10401 614 10453
rect 666 10401 678 10453
rect 730 10401 742 10453
rect 794 10401 806 10453
rect 858 10401 870 10453
rect 922 10401 934 10453
rect 986 10401 998 10453
rect 1050 10401 1062 10453
rect 1114 10401 1126 10453
rect 1178 10401 1190 10453
rect 1242 10401 1254 10453
rect 1306 10401 1318 10453
rect 1370 10401 1382 10453
rect 1434 10401 1446 10453
rect 1498 10401 1510 10453
rect 1562 10401 1574 10453
rect 1626 10401 1638 10453
rect 1690 10401 1702 10453
rect 1754 10401 1766 10453
rect 1818 10401 1830 10453
rect 1882 10401 1894 10453
rect 1946 10401 1958 10453
rect 2010 10401 2022 10453
rect 2074 10401 2086 10453
rect 2138 10401 2150 10453
rect 2202 10401 2214 10453
rect 2266 10401 2278 10453
rect 2330 10401 2342 10453
rect 2394 10401 2406 10453
rect 2458 10401 2470 10453
rect 2522 10401 2534 10453
rect 2586 10401 2598 10453
rect 2650 10401 2662 10453
rect 2714 10401 2726 10453
rect 2778 10401 2790 10453
rect 2842 10401 2854 10453
rect 2906 10401 2918 10453
rect 2970 10401 2982 10453
rect 3034 10401 3046 10453
rect 3098 10401 3110 10453
rect 3162 10401 3174 10453
rect 3226 10401 3238 10453
rect 3290 10401 3302 10453
rect 3354 10401 3366 10453
rect 3418 10401 3430 10453
rect 3482 10401 3494 10453
rect 3546 10401 3558 10453
rect 3610 10401 3622 10453
rect 3674 10401 3686 10453
rect 3738 10401 3750 10453
rect 3802 10401 3814 10453
rect 3866 10401 3878 10453
rect 3930 10401 3942 10453
rect 3994 10401 4006 10453
rect 4058 10401 4070 10453
rect 4122 10401 4134 10453
rect 4186 10401 4198 10453
rect 4250 10401 4262 10453
rect 4314 10401 4326 10453
rect 4378 10401 4390 10453
rect 4442 10401 4462 10453
rect 452 10384 4462 10401
rect -72 10057 10680 10085
rect -72 10023 108 10057
rect 142 10023 180 10057
rect 214 10023 252 10057
rect 286 10023 324 10057
rect 358 10023 396 10057
rect 430 10023 468 10057
rect 502 10023 540 10057
rect 574 10023 612 10057
rect 646 10023 684 10057
rect 718 10023 756 10057
rect 790 10023 828 10057
rect 862 10023 900 10057
rect 934 10023 972 10057
rect 1006 10023 1044 10057
rect 1078 10023 1116 10057
rect 1150 10023 1188 10057
rect 1222 10023 1260 10057
rect 1294 10023 1332 10057
rect 1366 10023 1404 10057
rect 1438 10023 1476 10057
rect 1510 10023 1548 10057
rect 1582 10023 1620 10057
rect 1654 10023 1692 10057
rect 1726 10023 1764 10057
rect 1798 10023 1836 10057
rect 1870 10023 1908 10057
rect 1942 10023 1980 10057
rect 2014 10023 2052 10057
rect 2086 10023 2124 10057
rect 2158 10023 2196 10057
rect 2230 10023 2268 10057
rect 2302 10023 2340 10057
rect 2374 10023 2412 10057
rect 2446 10023 2484 10057
rect 2518 10023 2556 10057
rect 2590 10023 2628 10057
rect 2662 10023 2700 10057
rect 2734 10023 2772 10057
rect 2806 10023 2844 10057
rect 2878 10023 2916 10057
rect 2950 10023 2988 10057
rect 3022 10023 3060 10057
rect 3094 10023 3132 10057
rect 3166 10023 3204 10057
rect 3238 10023 3276 10057
rect 3310 10023 3348 10057
rect 3382 10023 3420 10057
rect 3454 10023 3492 10057
rect 3526 10023 3564 10057
rect 3598 10023 3636 10057
rect 3670 10023 3708 10057
rect 3742 10023 3780 10057
rect 3814 10023 3852 10057
rect 3886 10023 3924 10057
rect 3958 10023 3996 10057
rect 4030 10023 4068 10057
rect 4102 10023 4140 10057
rect 4174 10023 4212 10057
rect 4246 10023 4284 10057
rect 4318 10023 4356 10057
rect 4390 10023 4428 10057
rect 4462 10023 4500 10057
rect 4534 10023 4572 10057
rect 4606 10023 4644 10057
rect 4678 10023 4716 10057
rect 4750 10023 4788 10057
rect 4822 10023 4860 10057
rect 4894 10023 4932 10057
rect 4966 10023 5004 10057
rect 5038 10023 5076 10057
rect 5110 10023 5148 10057
rect 5182 10023 5220 10057
rect 5254 10023 5292 10057
rect 5326 10023 5364 10057
rect 5398 10023 5436 10057
rect 5470 10023 5508 10057
rect 5542 10023 5580 10057
rect 5614 10023 5652 10057
rect 5686 10023 5724 10057
rect 5758 10023 5796 10057
rect 5830 10023 5868 10057
rect 5902 10023 5940 10057
rect 5974 10023 6012 10057
rect 6046 10023 6084 10057
rect 6118 10023 6156 10057
rect 6190 10023 6228 10057
rect 6262 10023 6300 10057
rect 6334 10023 6372 10057
rect 6406 10023 6444 10057
rect 6478 10023 6516 10057
rect 6550 10023 6588 10057
rect 6622 10023 6660 10057
rect 6694 10023 6732 10057
rect 6766 10023 6804 10057
rect 6838 10023 6876 10057
rect 6910 10023 6948 10057
rect 6982 10023 7020 10057
rect 7054 10023 7092 10057
rect 7126 10023 7164 10057
rect 7198 10023 7236 10057
rect 7270 10023 7308 10057
rect 7342 10023 7380 10057
rect 7414 10023 7452 10057
rect 7486 10023 7524 10057
rect 7558 10023 7596 10057
rect 7630 10023 7668 10057
rect 7702 10023 7740 10057
rect 7774 10023 7812 10057
rect 7846 10023 7884 10057
rect 7918 10023 7956 10057
rect 7990 10023 8028 10057
rect 8062 10023 8100 10057
rect 8134 10023 8172 10057
rect 8206 10023 8244 10057
rect 8278 10023 8316 10057
rect 8350 10023 8388 10057
rect 8422 10023 8460 10057
rect 8494 10023 8532 10057
rect 8566 10023 8604 10057
rect 8638 10023 8676 10057
rect 8710 10023 8748 10057
rect 8782 10023 8820 10057
rect 8854 10023 8892 10057
rect 8926 10023 8964 10057
rect 8998 10023 9036 10057
rect 9070 10023 9108 10057
rect 9142 10023 9180 10057
rect 9214 10023 9252 10057
rect 9286 10023 9324 10057
rect 9358 10023 9396 10057
rect 9430 10023 9468 10057
rect 9502 10023 9540 10057
rect 9574 10023 9612 10057
rect 9646 10023 9684 10057
rect 9718 10023 9756 10057
rect 9790 10023 9828 10057
rect 9862 10023 9900 10057
rect 9934 10023 9972 10057
rect 10006 10023 10044 10057
rect 10078 10023 10116 10057
rect 10150 10023 10188 10057
rect 10222 10023 10260 10057
rect 10294 10023 10332 10057
rect 10366 10023 10404 10057
rect 10438 10023 10476 10057
rect 10510 10023 10680 10057
rect -72 10002 10680 10023
rect -72 9924 11 10002
rect 5161 9987 5347 10002
rect -72 9890 -49 9924
rect -15 9890 11 9924
rect -72 9852 11 9890
rect -72 9818 -49 9852
rect -15 9818 11 9852
rect -72 9780 11 9818
rect -72 9746 -49 9780
rect -15 9746 11 9780
rect -72 9708 11 9746
rect -72 9674 -49 9708
rect -15 9674 11 9708
rect -72 9636 11 9674
rect -72 9602 -49 9636
rect -15 9602 11 9636
rect -72 9564 11 9602
rect -72 9530 -49 9564
rect -15 9530 11 9564
rect -72 9492 11 9530
rect -72 9458 -49 9492
rect -15 9458 11 9492
rect -72 9420 11 9458
rect -72 9386 -49 9420
rect -15 9386 11 9420
rect -72 9348 11 9386
rect -72 9314 -49 9348
rect -15 9314 11 9348
rect -72 9276 11 9314
rect -72 9242 -49 9276
rect -15 9242 11 9276
rect -72 9204 11 9242
rect -72 9170 -49 9204
rect -15 9170 11 9204
rect -72 9132 11 9170
rect -72 9098 -49 9132
rect -15 9098 11 9132
rect -72 9060 11 9098
rect -72 9026 -49 9060
rect -15 9026 11 9060
rect -72 8988 11 9026
rect -72 8954 -49 8988
rect -15 8954 11 8988
rect -72 8916 11 8954
rect -72 8882 -49 8916
rect -15 8882 11 8916
rect -72 8844 11 8882
rect -72 8810 -49 8844
rect -15 8810 11 8844
rect -72 8772 11 8810
rect -72 8738 -49 8772
rect -15 8738 11 8772
rect -72 8700 11 8738
rect -72 8666 -49 8700
rect -15 8666 11 8700
rect -72 8628 11 8666
rect -72 8594 -49 8628
rect -15 8594 11 8628
rect -72 8556 11 8594
rect -72 8522 -49 8556
rect -15 8522 11 8556
rect -72 8484 11 8522
rect -72 8450 -49 8484
rect -15 8450 11 8484
rect -72 8412 11 8450
rect -72 8378 -49 8412
rect -15 8378 11 8412
rect -72 8340 11 8378
rect -72 8306 -49 8340
rect -15 8306 11 8340
rect -72 8268 11 8306
rect -72 8234 -49 8268
rect -15 8234 11 8268
rect -72 8196 11 8234
rect -72 8162 -49 8196
rect -15 8162 11 8196
rect -72 8124 11 8162
rect -72 8090 -49 8124
rect -15 8090 11 8124
rect -72 8052 11 8090
rect -72 8018 -49 8052
rect -15 8018 11 8052
rect -72 7980 11 8018
rect -72 7946 -49 7980
rect -15 7946 11 7980
rect -72 7908 11 7946
rect -72 7874 -49 7908
rect -15 7874 11 7908
rect -72 7836 11 7874
rect -72 7802 -49 7836
rect -15 7802 11 7836
rect -72 7764 11 7802
rect -72 7730 -49 7764
rect -15 7730 11 7764
rect -72 7692 11 7730
rect -72 7658 -49 7692
rect -15 7658 11 7692
rect -72 7620 11 7658
rect -72 7586 -49 7620
rect -15 7586 11 7620
rect -72 7548 11 7586
rect -72 7514 -49 7548
rect -15 7514 11 7548
rect -72 7476 11 7514
rect -72 7442 -49 7476
rect -15 7442 11 7476
rect -72 7404 11 7442
rect -72 7370 -49 7404
rect -15 7370 11 7404
rect -72 7332 11 7370
rect -72 7298 -49 7332
rect -15 7298 11 7332
rect -72 7260 11 7298
rect -72 7226 -49 7260
rect -15 7226 11 7260
rect -72 7188 11 7226
rect -72 7154 -49 7188
rect -15 7154 11 7188
rect -72 7116 11 7154
rect -72 7082 -49 7116
rect -15 7082 11 7116
rect -72 7044 11 7082
rect -72 7010 -49 7044
rect -15 7010 11 7044
rect -72 6972 11 7010
rect -72 6938 -49 6972
rect -15 6938 11 6972
rect -72 6900 11 6938
rect -72 6866 -49 6900
rect -15 6866 11 6900
rect -72 6828 11 6866
rect -72 6794 -49 6828
rect -15 6794 11 6828
rect -72 6756 11 6794
rect -72 6722 -49 6756
rect -15 6722 11 6756
rect -72 6684 11 6722
rect -72 6650 -49 6684
rect -15 6650 11 6684
rect -72 6612 11 6650
rect -72 6578 -49 6612
rect -15 6578 11 6612
rect -72 6540 11 6578
rect -72 6506 -49 6540
rect -15 6506 11 6540
rect -72 6468 11 6506
rect -72 6434 -49 6468
rect -15 6434 11 6468
rect -72 6396 11 6434
rect -72 6362 -49 6396
rect -15 6362 11 6396
rect -72 6324 11 6362
rect -72 6290 -49 6324
rect -15 6290 11 6324
rect -72 6252 11 6290
rect -72 6218 -49 6252
rect -15 6218 11 6252
rect -72 6180 11 6218
rect -72 6146 -49 6180
rect -15 6146 11 6180
rect -72 6108 11 6146
rect -72 6074 -49 6108
rect -15 6074 11 6108
rect -72 6036 11 6074
rect -72 6002 -49 6036
rect -15 6002 11 6036
rect -72 5964 11 6002
rect -72 5930 -49 5964
rect -15 5930 11 5964
rect -72 5892 11 5930
rect -72 5858 -49 5892
rect -15 5858 11 5892
rect -72 5820 11 5858
rect -72 5786 -49 5820
rect -15 5786 11 5820
rect 10597 9880 10680 10002
rect 10597 9846 10619 9880
rect 10653 9846 10680 9880
rect 10597 9808 10680 9846
rect 10597 9774 10619 9808
rect 10653 9774 10680 9808
rect 10597 9736 10680 9774
rect 10597 9702 10619 9736
rect 10653 9702 10680 9736
rect 10597 9664 10680 9702
rect 10597 9630 10619 9664
rect 10653 9630 10680 9664
rect 10597 9592 10680 9630
rect 10597 9558 10619 9592
rect 10653 9558 10680 9592
rect 10597 9520 10680 9558
rect 10597 9486 10619 9520
rect 10653 9486 10680 9520
rect 10597 9448 10680 9486
rect 10597 9414 10619 9448
rect 10653 9414 10680 9448
rect 10597 9376 10680 9414
rect 10597 9342 10619 9376
rect 10653 9342 10680 9376
rect 10597 9304 10680 9342
rect 10597 9270 10619 9304
rect 10653 9270 10680 9304
rect 10597 9232 10680 9270
rect 10597 9198 10619 9232
rect 10653 9198 10680 9232
rect 10597 9160 10680 9198
rect 10597 9126 10619 9160
rect 10653 9126 10680 9160
rect 10597 9088 10680 9126
rect 10597 9054 10619 9088
rect 10653 9054 10680 9088
rect 10597 9016 10680 9054
rect 10597 8982 10619 9016
rect 10653 8982 10680 9016
rect 10597 8944 10680 8982
rect 10597 8910 10619 8944
rect 10653 8910 10680 8944
rect 10597 8872 10680 8910
rect 10597 8838 10619 8872
rect 10653 8838 10680 8872
rect 10597 8800 10680 8838
rect 10597 8766 10619 8800
rect 10653 8766 10680 8800
rect 10597 8728 10680 8766
rect 10597 8694 10619 8728
rect 10653 8694 10680 8728
rect 10597 8656 10680 8694
rect 10597 8622 10619 8656
rect 10653 8622 10680 8656
rect 10597 8584 10680 8622
rect 10597 8550 10619 8584
rect 10653 8550 10680 8584
rect 10597 8512 10680 8550
rect 10597 8478 10619 8512
rect 10653 8478 10680 8512
rect 10597 8440 10680 8478
rect 10597 8406 10619 8440
rect 10653 8406 10680 8440
rect 10597 8368 10680 8406
rect 10597 8334 10619 8368
rect 10653 8334 10680 8368
rect 10597 8296 10680 8334
rect 10597 8262 10619 8296
rect 10653 8262 10680 8296
rect 10597 8224 10680 8262
rect 10597 8190 10619 8224
rect 10653 8190 10680 8224
rect 10597 8152 10680 8190
rect 10597 8118 10619 8152
rect 10653 8118 10680 8152
rect 10597 8080 10680 8118
rect 10597 8046 10619 8080
rect 10653 8046 10680 8080
rect 10597 8008 10680 8046
rect 10597 7974 10619 8008
rect 10653 7974 10680 8008
rect 10597 7936 10680 7974
rect 10597 7902 10619 7936
rect 10653 7902 10680 7936
rect 10597 7864 10680 7902
rect 10597 7830 10619 7864
rect 10653 7830 10680 7864
rect 10597 7792 10680 7830
rect 10597 7758 10619 7792
rect 10653 7758 10680 7792
rect 10597 7720 10680 7758
rect 10597 7686 10619 7720
rect 10653 7686 10680 7720
rect 10597 7648 10680 7686
rect 10597 7614 10619 7648
rect 10653 7614 10680 7648
rect 10597 7576 10680 7614
rect 10597 7542 10619 7576
rect 10653 7542 10680 7576
rect 10597 7504 10680 7542
rect 10597 7470 10619 7504
rect 10653 7470 10680 7504
rect 10597 7432 10680 7470
rect 10597 7398 10619 7432
rect 10653 7398 10680 7432
rect 10597 7360 10680 7398
rect 10597 7326 10619 7360
rect 10653 7326 10680 7360
rect 10597 7288 10680 7326
rect 10597 7254 10619 7288
rect 10653 7254 10680 7288
rect 10597 7216 10680 7254
rect 10597 7182 10619 7216
rect 10653 7182 10680 7216
rect 10597 7144 10680 7182
rect 10597 7110 10619 7144
rect 10653 7110 10680 7144
rect 10597 7072 10680 7110
rect 10597 7038 10619 7072
rect 10653 7038 10680 7072
rect 10597 7000 10680 7038
rect 10597 6966 10619 7000
rect 10653 6966 10680 7000
rect 10597 6928 10680 6966
rect 10597 6894 10619 6928
rect 10653 6894 10680 6928
rect 10597 6856 10680 6894
rect 10597 6822 10619 6856
rect 10653 6822 10680 6856
rect 10597 6784 10680 6822
rect 10597 6750 10619 6784
rect 10653 6750 10680 6784
rect 10597 6712 10680 6750
rect 10597 6678 10619 6712
rect 10653 6678 10680 6712
rect 10597 6640 10680 6678
rect 10597 6606 10619 6640
rect 10653 6606 10680 6640
rect 10597 6568 10680 6606
rect 10597 6534 10619 6568
rect 10653 6534 10680 6568
rect 10597 6496 10680 6534
rect 10597 6462 10619 6496
rect 10653 6462 10680 6496
rect 10597 6424 10680 6462
rect 10597 6390 10619 6424
rect 10653 6390 10680 6424
rect 10597 6352 10680 6390
rect 10597 6318 10619 6352
rect 10653 6318 10680 6352
rect 10597 6280 10680 6318
rect 10597 6246 10619 6280
rect 10653 6246 10680 6280
rect 10597 6208 10680 6246
rect 10597 6174 10619 6208
rect 10653 6174 10680 6208
rect 10597 6136 10680 6174
rect 10597 6102 10619 6136
rect 10653 6102 10680 6136
rect 10597 6064 10680 6102
rect 10597 6030 10619 6064
rect 10653 6030 10680 6064
rect 10597 5992 10680 6030
rect 10597 5958 10619 5992
rect 10653 5958 10680 5992
rect 10597 5920 10680 5958
rect 10597 5886 10619 5920
rect 10653 5886 10680 5920
rect 10597 5798 10680 5886
rect -72 5748 11 5786
rect -72 5714 -49 5748
rect -15 5714 11 5748
rect -72 5676 11 5714
rect -72 5642 -49 5676
rect -15 5642 11 5676
rect -72 5604 11 5642
rect -72 5570 -49 5604
rect -15 5570 11 5604
rect -72 5532 11 5570
rect -72 5498 -49 5532
rect -15 5498 11 5532
rect -72 5460 11 5498
rect -72 5426 -49 5460
rect -15 5426 11 5460
rect -72 5388 11 5426
rect -72 5354 -49 5388
rect -15 5354 11 5388
rect -72 5316 11 5354
rect -72 5282 -49 5316
rect -15 5282 11 5316
rect -72 5244 11 5282
rect -72 5210 -49 5244
rect -15 5210 11 5244
rect -72 5172 11 5210
rect -72 5138 -49 5172
rect -15 5138 11 5172
rect -72 5100 11 5138
rect -72 5066 -49 5100
rect -15 5066 11 5100
rect -72 5028 11 5066
rect -72 4994 -49 5028
rect -15 4994 11 5028
rect -72 4956 11 4994
rect -72 4922 -49 4956
rect -15 4922 11 4956
rect -72 4884 11 4922
rect -72 4850 -49 4884
rect -15 4850 11 4884
rect -72 4812 11 4850
rect -72 4778 -49 4812
rect -15 4778 11 4812
rect -72 4740 11 4778
rect -72 4706 -49 4740
rect -15 4706 11 4740
rect -72 4668 11 4706
rect -72 4634 -49 4668
rect -15 4634 11 4668
rect -72 4596 11 4634
rect -72 4562 -49 4596
rect -15 4562 11 4596
rect -72 4524 11 4562
rect -72 4490 -49 4524
rect -15 4490 11 4524
rect -72 4452 11 4490
rect -72 4418 -49 4452
rect -15 4418 11 4452
rect -72 4380 11 4418
rect -72 4346 -49 4380
rect -15 4346 11 4380
rect -72 4308 11 4346
rect -72 4274 -49 4308
rect -15 4274 11 4308
rect -72 4236 11 4274
rect -72 4202 -49 4236
rect -15 4202 11 4236
rect -72 4164 11 4202
rect -72 4130 -49 4164
rect -15 4130 11 4164
rect -72 4092 11 4130
rect -72 4058 -49 4092
rect -15 4058 11 4092
rect -72 4020 11 4058
rect -72 3986 -49 4020
rect -15 3986 11 4020
rect -72 3948 11 3986
rect -72 3914 -49 3948
rect -15 3914 11 3948
rect -72 3876 11 3914
rect -72 3842 -49 3876
rect -15 3842 11 3876
rect -72 3804 11 3842
rect -72 3770 -49 3804
rect -15 3770 11 3804
rect -72 3732 11 3770
rect -72 3698 -49 3732
rect -15 3698 11 3732
rect -72 3660 11 3698
rect -72 3626 -49 3660
rect -15 3626 11 3660
rect -72 3588 11 3626
rect -72 3554 -49 3588
rect -15 3554 11 3588
rect -72 3516 11 3554
rect -72 3482 -49 3516
rect -15 3482 11 3516
rect -72 3444 11 3482
rect -72 3410 -49 3444
rect -15 3410 11 3444
rect -72 3372 11 3410
rect -72 3338 -49 3372
rect -15 3338 11 3372
rect -72 3300 11 3338
rect -72 3266 -49 3300
rect -15 3266 11 3300
rect -72 3228 11 3266
rect -72 3194 -49 3228
rect -15 3194 11 3228
rect -72 3156 11 3194
rect -72 3122 -49 3156
rect -15 3122 11 3156
rect -72 3084 11 3122
rect -72 3050 -49 3084
rect -15 3050 11 3084
rect -72 3012 11 3050
rect -72 2978 -49 3012
rect -15 2978 11 3012
rect -72 2940 11 2978
rect -72 2906 -49 2940
rect -15 2906 11 2940
rect -72 2868 11 2906
rect -72 2834 -49 2868
rect -15 2834 11 2868
rect -72 2796 11 2834
rect -72 2762 -49 2796
rect -15 2762 11 2796
rect -72 2724 11 2762
rect -72 2690 -49 2724
rect -15 2690 11 2724
rect -72 2652 11 2690
rect -72 2618 -49 2652
rect -15 2618 11 2652
rect -72 2580 11 2618
rect -72 2546 -49 2580
rect -15 2546 11 2580
rect -72 2508 11 2546
rect -72 2474 -49 2508
rect -15 2474 11 2508
rect -72 2436 11 2474
rect -72 2402 -49 2436
rect -15 2402 11 2436
rect -72 2364 11 2402
rect -72 2330 -49 2364
rect -15 2330 11 2364
rect -72 2292 11 2330
rect -72 2258 -49 2292
rect -15 2258 11 2292
rect -72 2220 11 2258
rect -72 2186 -49 2220
rect -15 2186 11 2220
rect -72 2148 11 2186
rect -72 2114 -49 2148
rect -15 2114 11 2148
rect -72 2076 11 2114
rect -72 2042 -49 2076
rect -15 2042 11 2076
rect -72 2004 11 2042
rect -72 1970 -49 2004
rect -15 1970 11 2004
rect -72 1932 11 1970
rect -72 1898 -49 1932
rect -15 1898 11 1932
rect -72 1860 11 1898
rect -72 1826 -49 1860
rect -15 1826 11 1860
rect -72 1788 11 1826
rect -72 1754 -49 1788
rect -15 1754 11 1788
rect -72 1716 11 1754
rect -72 1682 -49 1716
rect -15 1682 11 1716
rect -72 1644 11 1682
rect -72 1610 -49 1644
rect -15 1610 11 1644
rect -72 1572 11 1610
rect -72 1538 -49 1572
rect -15 1538 11 1572
rect -72 1500 11 1538
rect -72 1466 -49 1500
rect -15 1466 11 1500
rect -72 1428 11 1466
rect -72 1394 -49 1428
rect -15 1394 11 1428
rect -72 1356 11 1394
rect -72 1322 -49 1356
rect -15 1322 11 1356
rect -72 1284 11 1322
rect -72 1250 -49 1284
rect -15 1250 11 1284
rect -72 1212 11 1250
rect -72 1178 -49 1212
rect -15 1178 11 1212
rect -72 1140 11 1178
rect -72 1106 -49 1140
rect -15 1106 11 1140
rect -72 1068 11 1106
rect -72 1034 -49 1068
rect -15 1034 11 1068
rect -72 996 11 1034
rect -72 962 -49 996
rect -15 962 11 996
rect -72 924 11 962
rect -72 890 -49 924
rect -15 890 11 924
rect -72 852 11 890
rect -72 818 -49 852
rect -15 818 11 852
rect -72 780 11 818
rect -72 746 -49 780
rect -15 746 11 780
rect -72 708 11 746
rect -72 674 -49 708
rect -15 674 11 708
rect -72 636 11 674
rect -72 602 -49 636
rect -15 602 11 636
rect -72 564 11 602
rect -72 530 -49 564
rect -15 530 11 564
rect -72 492 11 530
rect -72 458 -49 492
rect -15 458 11 492
rect -72 420 11 458
rect -72 386 -49 420
rect -15 386 11 420
rect -72 348 11 386
rect -72 314 -49 348
rect -15 314 11 348
rect -72 276 11 314
rect -72 242 -49 276
rect -15 242 11 276
rect -72 204 11 242
rect -72 170 -49 204
rect -15 170 11 204
rect -72 132 11 170
rect -72 98 -49 132
rect -15 98 11 132
rect -72 -1140 11 98
rect 9393 5774 10680 5798
rect 9393 5740 9510 5774
rect 9544 5740 9582 5774
rect 9616 5740 9654 5774
rect 9688 5740 9726 5774
rect 9760 5740 9798 5774
rect 9832 5740 9870 5774
rect 9904 5740 9942 5774
rect 9976 5740 10014 5774
rect 10048 5740 10086 5774
rect 10120 5740 10158 5774
rect 10192 5740 10230 5774
rect 10264 5740 10302 5774
rect 10336 5740 10374 5774
rect 10408 5740 10446 5774
rect 10480 5740 10518 5774
rect 10552 5740 10680 5774
rect 9393 5715 10680 5740
rect 10739 6144 10990 6176
rect 10739 5964 10774 6144
rect 10954 5964 10990 6144
rect 9393 5683 9476 5715
rect 9393 5649 9417 5683
rect 9451 5649 9476 5683
rect 9393 5611 9476 5649
rect 9393 5577 9417 5611
rect 9451 5577 9476 5611
rect 9393 5539 9476 5577
rect 9393 5505 9417 5539
rect 9451 5505 9476 5539
rect 9393 5467 9476 5505
rect 9393 5433 9417 5467
rect 9451 5433 9476 5467
rect 9393 5395 9476 5433
rect 10739 5506 10990 5964
rect 9393 5361 9417 5395
rect 9451 5361 9476 5395
rect 9393 5323 9476 5361
rect 9393 5289 9417 5323
rect 9451 5289 9476 5323
rect 9393 5251 9476 5289
rect 9393 5217 9417 5251
rect 9451 5217 9476 5251
rect 9393 5179 9476 5217
rect 9393 5145 9417 5179
rect 9451 5145 9476 5179
rect 9393 5107 9476 5145
rect 9393 5073 9417 5107
rect 9451 5073 9476 5107
rect 9393 5035 9476 5073
rect 9393 5001 9417 5035
rect 9451 5001 9476 5035
rect 9393 4963 9476 5001
rect 9393 4929 9417 4963
rect 9451 4929 9476 4963
rect 9393 4891 9476 4929
rect 9393 4857 9417 4891
rect 9451 4857 9476 4891
rect 9393 4819 9476 4857
rect 9393 4785 9417 4819
rect 9451 4785 9476 4819
rect 9393 4747 9476 4785
rect 9393 4713 9417 4747
rect 9451 4713 9476 4747
rect 10654 5407 10711 5421
rect 10654 5355 10656 5407
rect 10708 5355 10711 5407
rect 10654 5343 10711 5355
rect 10654 5291 10656 5343
rect 10708 5291 10711 5343
rect 10654 5279 10711 5291
rect 10654 5227 10656 5279
rect 10708 5227 10711 5279
rect 10654 5215 10711 5227
rect 10654 5163 10656 5215
rect 10708 5163 10711 5215
rect 10654 5151 10711 5163
rect 10654 5099 10656 5151
rect 10708 5099 10711 5151
rect 10654 5087 10711 5099
rect 10654 5035 10656 5087
rect 10708 5035 10711 5087
rect 10654 5023 10711 5035
rect 10654 4971 10656 5023
rect 10708 4971 10711 5023
rect 10654 4959 10711 4971
rect 10654 4907 10656 4959
rect 10708 4907 10711 4959
rect 9393 4675 9476 4713
rect 9393 4641 9417 4675
rect 9451 4641 9476 4675
rect 9393 4603 9476 4641
rect 9393 4569 9417 4603
rect 9451 4569 9476 4603
rect 9393 4531 9476 4569
rect 9393 4497 9417 4531
rect 9451 4497 9476 4531
rect 9393 4459 9476 4497
rect 9393 4425 9417 4459
rect 9451 4425 9476 4459
rect 9393 4387 9476 4425
rect 9393 4353 9417 4387
rect 9451 4353 9476 4387
rect 9393 4315 9476 4353
rect 9393 4281 9417 4315
rect 9451 4281 9476 4315
rect 9393 4243 9476 4281
rect 9393 4209 9417 4243
rect 9451 4209 9476 4243
rect 9393 4171 9476 4209
rect 9393 4137 9417 4171
rect 9451 4137 9476 4171
rect 9393 4099 9476 4137
rect 9393 4065 9417 4099
rect 9451 4065 9476 4099
rect 9393 4027 9476 4065
rect 9393 3993 9417 4027
rect 9451 3993 9476 4027
rect 9393 3955 9476 3993
rect 9393 3921 9417 3955
rect 9451 3921 9476 3955
rect 9393 3883 9476 3921
rect 9393 3849 9417 3883
rect 9451 3849 9476 3883
rect 9393 3811 9476 3849
rect 9393 3777 9417 3811
rect 9451 3777 9476 3811
rect 9393 3739 9476 3777
rect 9393 3705 9417 3739
rect 9451 3705 9476 3739
rect 9393 3667 9476 3705
rect 9393 3633 9417 3667
rect 9451 3633 9476 3667
rect 9393 3595 9476 3633
rect 9393 3561 9417 3595
rect 9451 3561 9476 3595
rect 9393 3523 9476 3561
rect 9393 3489 9417 3523
rect 9451 3489 9476 3523
rect 9393 3451 9476 3489
rect 9393 3417 9417 3451
rect 9451 3417 9476 3451
rect 9393 3379 9476 3417
rect 9393 3345 9417 3379
rect 9451 3345 9476 3379
rect 9393 3307 9476 3345
rect 9393 3273 9417 3307
rect 9451 3273 9476 3307
rect 9393 3235 9476 3273
rect 9393 3201 9417 3235
rect 9451 3201 9476 3235
rect 9393 3163 9476 3201
rect 9393 3129 9417 3163
rect 9451 3129 9476 3163
rect 9393 3091 9476 3129
rect 9393 3057 9417 3091
rect 9451 3057 9476 3091
rect 9393 3019 9476 3057
rect 9393 2985 9417 3019
rect 9451 2985 9476 3019
rect 9393 2947 9476 2985
rect 9393 2913 9417 2947
rect 9451 2913 9476 2947
rect 9393 2875 9476 2913
rect 9393 2841 9417 2875
rect 9451 2841 9476 2875
rect 9393 2803 9476 2841
rect 9393 2769 9417 2803
rect 9451 2769 9476 2803
rect 9393 2731 9476 2769
rect 9393 2697 9417 2731
rect 9451 2697 9476 2731
rect 9393 2659 9476 2697
rect 9393 2625 9417 2659
rect 9451 2625 9476 2659
rect 9393 2587 9476 2625
rect 9393 2553 9417 2587
rect 9451 2553 9476 2587
rect 9393 2515 9476 2553
rect 9393 2481 9417 2515
rect 9451 2481 9476 2515
rect 9393 2443 9476 2481
rect 9393 2409 9417 2443
rect 9451 2409 9476 2443
rect 9393 2371 9476 2409
rect 9393 2337 9417 2371
rect 9451 2337 9476 2371
rect 9393 2299 9476 2337
rect 9393 2265 9417 2299
rect 9451 2265 9476 2299
rect 9393 2227 9476 2265
rect 9393 2193 9417 2227
rect 9451 2193 9476 2227
rect 9393 2155 9476 2193
rect 9393 2121 9417 2155
rect 9451 2121 9476 2155
rect 9393 2083 9476 2121
rect 9393 2049 9417 2083
rect 9451 2049 9476 2083
rect 9393 2011 9476 2049
rect 9393 1977 9417 2011
rect 9451 1977 9476 2011
rect 9393 1939 9476 1977
rect 9393 1905 9417 1939
rect 9451 1905 9476 1939
rect 9393 1867 9476 1905
rect 9393 1833 9417 1867
rect 9451 1833 9476 1867
rect 9393 1795 9476 1833
rect 9393 1761 9417 1795
rect 9451 1761 9476 1795
rect 9393 1723 9476 1761
rect 9393 1689 9417 1723
rect 9451 1689 9476 1723
rect 9393 1651 9476 1689
rect 9393 1617 9417 1651
rect 9451 1617 9476 1651
rect 9393 1579 9476 1617
rect 9393 1545 9417 1579
rect 9451 1545 9476 1579
rect 9393 1507 9476 1545
rect 9393 1473 9417 1507
rect 9451 1473 9476 1507
rect 9393 1435 9476 1473
rect 9393 1401 9417 1435
rect 9451 1401 9476 1435
rect 9393 1363 9476 1401
rect 9393 1329 9417 1363
rect 9451 1329 9476 1363
rect 9393 1291 9476 1329
rect 9393 1257 9417 1291
rect 9451 1257 9476 1291
rect 9393 1219 9476 1257
rect 9393 1185 9417 1219
rect 9451 1185 9476 1219
rect 9393 1147 9476 1185
rect 9393 1113 9417 1147
rect 9451 1113 9476 1147
rect 9393 1075 9476 1113
rect 9393 1041 9417 1075
rect 9451 1041 9476 1075
rect 9393 1003 9476 1041
rect 9393 969 9417 1003
rect 9451 969 9476 1003
rect 9393 931 9476 969
rect 9393 897 9417 931
rect 9451 897 9476 931
rect 9393 859 9476 897
rect 9393 825 9417 859
rect 9451 825 9476 859
rect 9393 787 9476 825
rect 9393 753 9417 787
rect 9451 753 9476 787
rect 9393 715 9476 753
rect 9393 681 9417 715
rect 9451 681 9476 715
rect 9393 643 9476 681
rect 9393 609 9417 643
rect 9451 609 9476 643
rect 9393 571 9476 609
rect 9393 537 9417 571
rect 9451 537 9476 571
rect 9393 499 9476 537
rect 9393 465 9417 499
rect 9451 465 9476 499
rect 9393 427 9476 465
rect 9393 393 9417 427
rect 9451 393 9476 427
rect 9393 355 9476 393
rect 9393 321 9417 355
rect 9451 321 9476 355
rect 9393 283 9476 321
rect 9393 249 9417 283
rect 9451 249 9476 283
rect 9393 211 9476 249
rect 9393 177 9417 211
rect 9451 177 9476 211
rect 9393 139 9476 177
rect 9393 105 9417 139
rect 9451 105 9476 139
rect 9393 43 9476 105
rect 9393 9 9417 43
rect 9451 9 9476 43
rect 9393 -29 9476 9
rect 8020 -57 9022 -42
rect 8020 -109 8041 -57
rect 8093 -109 8105 -57
rect 8157 -109 8169 -57
rect 8221 -109 8233 -57
rect 8285 -109 8297 -57
rect 8349 -109 8361 -57
rect 8413 -109 8425 -57
rect 8477 -109 8489 -57
rect 8541 -109 8553 -57
rect 8605 -109 8617 -57
rect 8669 -109 8681 -57
rect 8733 -109 8745 -57
rect 8797 -109 8809 -57
rect 8861 -109 8873 -57
rect 8925 -109 8937 -57
rect 8989 -109 9022 -57
rect 8020 -128 9022 -109
rect 9393 -63 9417 -29
rect 9451 -63 9476 -29
rect 9393 -101 9476 -63
rect 9393 -135 9417 -101
rect 9451 -135 9476 -101
rect 9058 -179 9248 -162
rect 9058 -232 9092 -179
rect 9054 -551 9092 -232
rect 9208 -551 9248 -179
rect 9054 -564 9248 -551
rect 9058 -566 9248 -564
rect 9393 -173 9476 -135
rect 9393 -207 9417 -173
rect 9451 -207 9476 -173
rect 9393 -245 9476 -207
rect 9393 -279 9417 -245
rect 9451 -279 9476 -245
rect 9393 -317 9476 -279
rect 9393 -351 9417 -317
rect 9451 -351 9476 -317
rect 9393 -389 9476 -351
rect 9393 -423 9417 -389
rect 9451 -423 9476 -389
rect 9393 -461 9476 -423
rect 9393 -495 9417 -461
rect 9451 -495 9476 -461
rect 9393 -533 9476 -495
rect 9393 -567 9417 -533
rect 9451 -567 9476 -533
rect 8024 -600 9026 -578
rect 8024 -716 8052 -600
rect 9000 -716 9026 -600
rect 8024 -740 9026 -716
rect 9393 -605 9476 -567
rect 9393 -639 9417 -605
rect 9451 -639 9476 -605
rect 9393 -677 9476 -639
rect 9393 -711 9417 -677
rect 9451 -711 9476 -677
rect -72 -1174 -49 -1140
rect -15 -1174 11 -1140
rect -72 -1234 11 -1174
rect 9393 -749 9476 -711
rect 9393 -783 9417 -749
rect 9451 -783 9476 -749
rect 9393 -821 9476 -783
rect 9393 -855 9417 -821
rect 9451 -855 9476 -821
rect 9393 -893 9476 -855
rect 9393 -927 9417 -893
rect 9451 -927 9476 -893
rect 9393 -965 9476 -927
rect 9393 -999 9417 -965
rect 9451 -999 9476 -965
rect 9393 -1037 9476 -999
rect 9393 -1071 9417 -1037
rect 9451 -1071 9476 -1037
rect 9393 -1109 9476 -1071
rect 9393 -1143 9417 -1109
rect 9451 -1143 9476 -1109
rect 9911 -1116 10174 4739
rect 10654 4656 10711 4907
rect 10739 4673 10813 5506
rect 10841 4673 10887 5506
rect 10915 4673 10989 5506
rect 10378 4330 10444 4344
rect 10378 4278 10385 4330
rect 10437 4278 10444 4330
rect 10378 4266 10444 4278
rect 10378 4214 10385 4266
rect 10437 4214 10444 4266
rect 10378 4202 10444 4214
rect 10378 4150 10385 4202
rect 10437 4150 10444 4202
rect 10378 3840 10444 4150
rect 10208 3809 10549 3840
rect 10208 3775 10257 3809
rect 10291 3775 10329 3809
rect 10363 3775 10401 3809
rect 10435 3775 10473 3809
rect 10507 3775 10549 3809
rect 10208 3745 10549 3775
rect 11019 3288 11088 3310
rect 11019 3254 11036 3288
rect 11070 3254 11088 3288
rect 11019 3216 11088 3254
rect 11019 3182 11036 3216
rect 11070 3182 11088 3216
rect 10656 2636 10708 3090
rect 10742 2646 10810 3068
rect 10842 2644 10886 3128
rect 10916 2632 10988 3066
rect 11019 3065 11088 3182
rect 11019 3013 11027 3065
rect 11079 3013 11088 3065
rect 11019 3001 11088 3013
rect 11019 2949 11027 3001
rect 11079 2949 11088 3001
rect 11019 2907 11088 2949
rect 10366 2394 10478 2416
rect 10366 2342 10396 2394
rect 10448 2342 10478 2394
rect 10366 2330 10478 2342
rect 10366 2278 10396 2330
rect 10448 2278 10478 2330
rect 10366 2266 10478 2278
rect 10366 2220 10396 2266
rect 10364 2214 10396 2220
rect 10448 2214 10478 2266
rect 10364 2202 10478 2214
rect 10364 2150 10396 2202
rect 10448 2150 10478 2202
rect 10364 2148 10404 2150
rect 10438 2148 10478 2150
rect 10364 2122 10478 2148
rect 10366 2110 10476 2122
rect 10748 581 10998 756
rect 10741 540 10998 581
rect 11270 581 11384 608
rect 11270 547 11310 581
rect 11344 547 11384 581
rect 11270 542 11384 547
rect 10394 450 10488 480
rect 10741 460 10995 540
rect 11268 468 11384 542
rect 10394 398 10413 450
rect 10465 398 10488 450
rect 10394 388 10488 398
rect 10394 386 10490 388
rect 10394 334 10413 386
rect 10465 349 10490 386
rect 10394 322 10434 334
rect 10394 270 10413 322
rect 10468 315 10490 349
rect 10465 277 10490 315
rect 10394 243 10434 270
rect 10468 243 10490 277
rect 10394 236 10490 243
rect 10396 205 10490 236
rect 10396 171 10434 205
rect 10468 171 10490 205
rect 10396 62 10490 171
rect 10416 8 10490 62
rect 10420 -466 10534 -462
rect 10416 -507 10534 -466
rect 10416 -541 10460 -507
rect 10494 -541 10534 -507
rect 10416 -579 10534 -541
rect 10416 -613 10460 -579
rect 10494 -613 10534 -579
rect 10416 -666 10534 -613
rect 10804 -616 10946 460
rect 11268 416 11300 468
rect 11352 416 11384 468
rect 11268 404 11384 416
rect 11268 352 11300 404
rect 11352 352 11384 404
rect 11268 340 11384 352
rect 11268 288 11300 340
rect 11352 288 11384 340
rect 11268 258 11384 288
rect 10416 -714 10532 -666
rect 10416 -766 10443 -714
rect 10495 -766 10532 -714
rect 10416 -778 10532 -766
rect 10416 -830 10443 -778
rect 10495 -830 10532 -778
rect 10416 -842 10532 -830
rect 10416 -894 10443 -842
rect 10495 -894 10532 -842
rect 10416 -946 10532 -894
rect 11435 -1116 11698 4716
rect 9393 -1234 9476 -1143
rect -72 -1262 9476 -1234
rect -72 -1296 32 -1262
rect 66 -1296 104 -1262
rect 138 -1296 176 -1262
rect 210 -1296 248 -1262
rect 282 -1296 320 -1262
rect 354 -1296 392 -1262
rect 426 -1296 464 -1262
rect 498 -1296 536 -1262
rect 570 -1296 608 -1262
rect 642 -1296 680 -1262
rect 714 -1296 752 -1262
rect 786 -1296 824 -1262
rect 858 -1296 896 -1262
rect 930 -1296 968 -1262
rect 1002 -1296 1040 -1262
rect 1074 -1296 1112 -1262
rect 1146 -1296 1184 -1262
rect 1218 -1296 1256 -1262
rect 1290 -1296 1328 -1262
rect 1362 -1296 1400 -1262
rect 1434 -1296 1472 -1262
rect 1506 -1296 1544 -1262
rect 1578 -1296 1616 -1262
rect 1650 -1296 1688 -1262
rect 1722 -1296 1760 -1262
rect 1794 -1296 1832 -1262
rect 1866 -1296 1904 -1262
rect 1938 -1296 1976 -1262
rect 2010 -1296 2048 -1262
rect 2082 -1296 2120 -1262
rect 2154 -1296 2192 -1262
rect 2226 -1296 2264 -1262
rect 2298 -1296 2336 -1262
rect 2370 -1296 2408 -1262
rect 2442 -1296 2480 -1262
rect 2514 -1296 2552 -1262
rect 2586 -1296 2624 -1262
rect 2658 -1296 2696 -1262
rect 2730 -1296 2768 -1262
rect 2802 -1296 2840 -1262
rect 2874 -1296 2912 -1262
rect 2946 -1296 2984 -1262
rect 3018 -1296 3056 -1262
rect 3090 -1296 3128 -1262
rect 3162 -1296 3200 -1262
rect 3234 -1296 3272 -1262
rect 3306 -1296 3344 -1262
rect 3378 -1296 3416 -1262
rect 3450 -1296 3488 -1262
rect 3522 -1296 3560 -1262
rect 3594 -1296 3632 -1262
rect 3666 -1296 3704 -1262
rect 3738 -1296 3776 -1262
rect 3810 -1296 3848 -1262
rect 3882 -1296 3920 -1262
rect 3954 -1296 3992 -1262
rect 4026 -1296 4064 -1262
rect 4098 -1296 4136 -1262
rect 4170 -1296 4208 -1262
rect 4242 -1296 4280 -1262
rect 4314 -1296 4352 -1262
rect 4386 -1296 4424 -1262
rect 4458 -1296 4496 -1262
rect 4530 -1296 4568 -1262
rect 4602 -1296 4640 -1262
rect 4674 -1296 4712 -1262
rect 4746 -1296 4784 -1262
rect 4818 -1296 4856 -1262
rect 4890 -1296 4928 -1262
rect 4962 -1296 5000 -1262
rect 5034 -1296 5072 -1262
rect 5106 -1296 5144 -1262
rect 5178 -1296 5216 -1262
rect 5250 -1296 5288 -1262
rect 5322 -1296 5360 -1262
rect 5394 -1296 5432 -1262
rect 5466 -1296 5504 -1262
rect 5538 -1296 5576 -1262
rect 5610 -1296 5648 -1262
rect 5682 -1296 5720 -1262
rect 5754 -1296 5792 -1262
rect 5826 -1296 5864 -1262
rect 5898 -1296 5936 -1262
rect 5970 -1296 6008 -1262
rect 6042 -1296 6080 -1262
rect 6114 -1296 6152 -1262
rect 6186 -1296 6224 -1262
rect 6258 -1296 6296 -1262
rect 6330 -1296 6368 -1262
rect 6402 -1296 6440 -1262
rect 6474 -1296 6512 -1262
rect 6546 -1296 6584 -1262
rect 6618 -1296 6656 -1262
rect 6690 -1296 6728 -1262
rect 6762 -1296 6800 -1262
rect 6834 -1296 6872 -1262
rect 6906 -1296 6944 -1262
rect 6978 -1296 7016 -1262
rect 7050 -1296 7088 -1262
rect 7122 -1296 7160 -1262
rect 7194 -1296 7232 -1262
rect 7266 -1296 7304 -1262
rect 7338 -1296 7376 -1262
rect 7410 -1296 7448 -1262
rect 7482 -1296 7520 -1262
rect 7554 -1296 7592 -1262
rect 7626 -1296 7664 -1262
rect 7698 -1296 7736 -1262
rect 7770 -1296 7808 -1262
rect 7842 -1296 7880 -1262
rect 7914 -1296 7952 -1262
rect 7986 -1296 8024 -1262
rect 8058 -1296 8096 -1262
rect 8130 -1296 8168 -1262
rect 8202 -1296 8240 -1262
rect 8274 -1296 8312 -1262
rect 8346 -1296 8384 -1262
rect 8418 -1296 8456 -1262
rect 8490 -1296 8528 -1262
rect 8562 -1296 8600 -1262
rect 8634 -1296 8672 -1262
rect 8706 -1296 8744 -1262
rect 8778 -1296 8816 -1262
rect 8850 -1296 8888 -1262
rect 8922 -1296 8960 -1262
rect 8994 -1296 9032 -1262
rect 9066 -1296 9104 -1262
rect 9138 -1296 9176 -1262
rect 9210 -1296 9248 -1262
rect 9282 -1296 9320 -1262
rect 9354 -1296 9476 -1262
rect -72 -1317 9476 -1296
rect 9910 -1120 11698 -1116
rect 9910 -1128 11710 -1120
rect 9910 -1372 10001 -1128
rect 11589 -1372 11710 -1128
rect 9910 -1396 11710 -1372
rect 9911 -1401 10174 -1396
<< via1 >>
rect 470 10931 522 10983
rect 534 10931 586 10983
rect 598 10931 650 10983
rect 662 10931 714 10983
rect 726 10931 778 10983
rect 790 10931 842 10983
rect 854 10931 906 10983
rect 918 10931 970 10983
rect 982 10931 1034 10983
rect 1046 10931 1098 10983
rect 1110 10931 1162 10983
rect 1174 10931 1226 10983
rect 1238 10931 1290 10983
rect 1302 10931 1354 10983
rect 1366 10931 1418 10983
rect 1430 10931 1482 10983
rect 1494 10931 1546 10983
rect 1558 10931 1610 10983
rect 1622 10931 1674 10983
rect 1686 10931 1738 10983
rect 1750 10931 1802 10983
rect 1814 10931 1866 10983
rect 1878 10931 1930 10983
rect 1942 10931 1994 10983
rect 2006 10931 2058 10983
rect 2070 10931 2122 10983
rect 2134 10931 2186 10983
rect 2198 10931 2250 10983
rect 2262 10931 2314 10983
rect 2326 10931 2378 10983
rect 2390 10931 2442 10983
rect 2454 10931 2506 10983
rect 2518 10931 2570 10983
rect 2582 10931 2634 10983
rect 2646 10931 2698 10983
rect 2710 10931 2762 10983
rect 2774 10931 2826 10983
rect 2838 10931 2890 10983
rect 2902 10931 2954 10983
rect 2966 10931 3018 10983
rect 3030 10931 3082 10983
rect 3094 10931 3146 10983
rect 3158 10931 3210 10983
rect 3222 10931 3274 10983
rect 3286 10931 3338 10983
rect 3350 10931 3402 10983
rect 3414 10931 3466 10983
rect 3478 10931 3530 10983
rect 3542 10931 3594 10983
rect 3606 10931 3658 10983
rect 3670 10931 3722 10983
rect 3734 10931 3786 10983
rect 3798 10931 3850 10983
rect 3862 10931 3914 10983
rect 3926 10931 3978 10983
rect 3990 10931 4042 10983
rect 4054 10931 4106 10983
rect 4118 10931 4170 10983
rect 4182 10931 4234 10983
rect 4246 10931 4298 10983
rect 4310 10931 4362 10983
rect 4374 10931 4426 10983
rect -172 10644 200 10760
rect 4535 10544 4715 10788
rect 486 10401 538 10453
rect 550 10401 602 10453
rect 614 10401 666 10453
rect 678 10401 730 10453
rect 742 10401 794 10453
rect 806 10401 858 10453
rect 870 10401 922 10453
rect 934 10401 986 10453
rect 998 10401 1050 10453
rect 1062 10401 1114 10453
rect 1126 10401 1178 10453
rect 1190 10401 1242 10453
rect 1254 10401 1306 10453
rect 1318 10401 1370 10453
rect 1382 10401 1434 10453
rect 1446 10401 1498 10453
rect 1510 10401 1562 10453
rect 1574 10401 1626 10453
rect 1638 10401 1690 10453
rect 1702 10401 1754 10453
rect 1766 10401 1818 10453
rect 1830 10401 1882 10453
rect 1894 10401 1946 10453
rect 1958 10401 2010 10453
rect 2022 10401 2074 10453
rect 2086 10401 2138 10453
rect 2150 10401 2202 10453
rect 2214 10401 2266 10453
rect 2278 10401 2330 10453
rect 2342 10401 2394 10453
rect 2406 10401 2458 10453
rect 2470 10401 2522 10453
rect 2534 10401 2586 10453
rect 2598 10401 2650 10453
rect 2662 10401 2714 10453
rect 2726 10401 2778 10453
rect 2790 10401 2842 10453
rect 2854 10401 2906 10453
rect 2918 10401 2970 10453
rect 2982 10401 3034 10453
rect 3046 10401 3098 10453
rect 3110 10401 3162 10453
rect 3174 10401 3226 10453
rect 3238 10401 3290 10453
rect 3302 10401 3354 10453
rect 3366 10401 3418 10453
rect 3430 10401 3482 10453
rect 3494 10401 3546 10453
rect 3558 10401 3610 10453
rect 3622 10401 3674 10453
rect 3686 10401 3738 10453
rect 3750 10401 3802 10453
rect 3814 10401 3866 10453
rect 3878 10401 3930 10453
rect 3942 10401 3994 10453
rect 4006 10401 4058 10453
rect 4070 10401 4122 10453
rect 4134 10401 4186 10453
rect 4198 10401 4250 10453
rect 4262 10401 4314 10453
rect 4326 10401 4378 10453
rect 4390 10401 4442 10453
rect 10774 5964 10954 6144
rect 10656 5355 10708 5407
rect 10656 5291 10708 5343
rect 10656 5227 10708 5279
rect 10656 5163 10708 5215
rect 10656 5099 10708 5151
rect 10656 5035 10708 5087
rect 10656 4971 10708 5023
rect 10656 4907 10708 4959
rect 8041 -109 8093 -57
rect 8105 -109 8157 -57
rect 8169 -109 8221 -57
rect 8233 -109 8285 -57
rect 8297 -109 8349 -57
rect 8361 -109 8413 -57
rect 8425 -109 8477 -57
rect 8489 -109 8541 -57
rect 8553 -109 8605 -57
rect 8617 -109 8669 -57
rect 8681 -109 8733 -57
rect 8745 -109 8797 -57
rect 8809 -109 8861 -57
rect 8873 -109 8925 -57
rect 8937 -109 8989 -57
rect 9092 -551 9208 -179
rect 8052 -716 9000 -600
rect 10385 4278 10437 4330
rect 10385 4214 10437 4266
rect 10385 4150 10437 4202
rect 11027 3013 11079 3065
rect 11027 2949 11079 3001
rect 10396 2342 10448 2394
rect 10396 2278 10448 2330
rect 10396 2214 10448 2266
rect 10396 2182 10448 2202
rect 10396 2150 10404 2182
rect 10404 2150 10438 2182
rect 10438 2150 10448 2182
rect 10413 398 10465 450
rect 10413 349 10465 386
rect 10413 334 10434 349
rect 10434 334 10465 349
rect 10413 315 10434 322
rect 10434 315 10465 322
rect 10413 277 10465 315
rect 10413 270 10434 277
rect 10434 270 10465 277
rect 11300 416 11352 468
rect 11300 352 11352 404
rect 11300 288 11352 340
rect 10443 -766 10495 -714
rect 10443 -830 10495 -778
rect 10443 -894 10495 -842
rect 10001 -1372 11589 -1128
<< metal2 >>
rect 5988 10998 6414 11004
rect 448 10983 6414 10998
rect 448 10931 470 10983
rect 522 10931 534 10983
rect 586 10931 598 10983
rect 650 10931 662 10983
rect 714 10931 726 10983
rect 778 10931 790 10983
rect 842 10931 854 10983
rect 906 10931 918 10983
rect 970 10931 982 10983
rect 1034 10931 1046 10983
rect 1098 10931 1110 10983
rect 1162 10931 1174 10983
rect 1226 10931 1238 10983
rect 1290 10931 1302 10983
rect 1354 10931 1366 10983
rect 1418 10931 1430 10983
rect 1482 10931 1494 10983
rect 1546 10931 1558 10983
rect 1610 10931 1622 10983
rect 1674 10931 1686 10983
rect 1738 10931 1750 10983
rect 1802 10931 1814 10983
rect 1866 10931 1878 10983
rect 1930 10931 1942 10983
rect 1994 10931 2006 10983
rect 2058 10931 2070 10983
rect 2122 10931 2134 10983
rect 2186 10931 2198 10983
rect 2250 10931 2262 10983
rect 2314 10931 2326 10983
rect 2378 10931 2390 10983
rect 2442 10931 2454 10983
rect 2506 10931 2518 10983
rect 2570 10931 2582 10983
rect 2634 10931 2646 10983
rect 2698 10931 2710 10983
rect 2762 10931 2774 10983
rect 2826 10931 2838 10983
rect 2890 10931 2902 10983
rect 2954 10931 2966 10983
rect 3018 10931 3030 10983
rect 3082 10931 3094 10983
rect 3146 10931 3158 10983
rect 3210 10931 3222 10983
rect 3274 10931 3286 10983
rect 3338 10931 3350 10983
rect 3402 10931 3414 10983
rect 3466 10931 3478 10983
rect 3530 10931 3542 10983
rect 3594 10931 3606 10983
rect 3658 10931 3670 10983
rect 3722 10931 3734 10983
rect 3786 10931 3798 10983
rect 3850 10931 3862 10983
rect 3914 10931 3926 10983
rect 3978 10931 3990 10983
rect 4042 10931 4054 10983
rect 4106 10931 4118 10983
rect 4170 10931 4182 10983
rect 4234 10931 4246 10983
rect 4298 10931 4310 10983
rect 4362 10931 4374 10983
rect 4426 10931 6414 10983
rect 448 10929 6414 10931
rect 448 10910 6043 10929
rect 5988 10873 6043 10910
rect 6099 10873 6123 10929
rect 6179 10873 6203 10929
rect 6259 10873 6283 10929
rect 6339 10873 6414 10929
rect 5988 10814 6414 10873
rect -200 10770 270 10802
rect -200 10634 -174 10770
rect 202 10634 270 10770
rect -200 10602 270 10634
rect 4492 10788 4758 10812
rect 4492 10544 4535 10788
rect 4715 10726 4758 10788
rect 9622 10726 9952 10736
rect 4715 10707 9952 10726
rect 4715 10578 9669 10707
rect 4715 10544 4758 10578
rect 4492 10514 4758 10544
rect 9622 10491 9669 10578
rect 9885 10491 9952 10707
rect 4284 10472 5116 10476
rect 452 10453 5116 10472
rect 452 10401 486 10453
rect 538 10401 550 10453
rect 602 10401 614 10453
rect 666 10401 678 10453
rect 730 10401 742 10453
rect 794 10401 806 10453
rect 858 10401 870 10453
rect 922 10401 934 10453
rect 986 10401 998 10453
rect 1050 10401 1062 10453
rect 1114 10401 1126 10453
rect 1178 10401 1190 10453
rect 1242 10401 1254 10453
rect 1306 10401 1318 10453
rect 1370 10401 1382 10453
rect 1434 10401 1446 10453
rect 1498 10401 1510 10453
rect 1562 10401 1574 10453
rect 1626 10401 1638 10453
rect 1690 10401 1702 10453
rect 1754 10401 1766 10453
rect 1818 10401 1830 10453
rect 1882 10401 1894 10453
rect 1946 10401 1958 10453
rect 2010 10401 2022 10453
rect 2074 10401 2086 10453
rect 2138 10401 2150 10453
rect 2202 10401 2214 10453
rect 2266 10401 2278 10453
rect 2330 10401 2342 10453
rect 2394 10401 2406 10453
rect 2458 10401 2470 10453
rect 2522 10401 2534 10453
rect 2586 10401 2598 10453
rect 2650 10401 2662 10453
rect 2714 10401 2726 10453
rect 2778 10401 2790 10453
rect 2842 10401 2854 10453
rect 2906 10401 2918 10453
rect 2970 10401 2982 10453
rect 3034 10401 3046 10453
rect 3098 10401 3110 10453
rect 3162 10401 3174 10453
rect 3226 10401 3238 10453
rect 3290 10401 3302 10453
rect 3354 10401 3366 10453
rect 3418 10401 3430 10453
rect 3482 10401 3494 10453
rect 3546 10401 3558 10453
rect 3610 10401 3622 10453
rect 3674 10401 3686 10453
rect 3738 10401 3750 10453
rect 3802 10401 3814 10453
rect 3866 10401 3878 10453
rect 3930 10401 3942 10453
rect 3994 10401 4006 10453
rect 4058 10401 4070 10453
rect 4122 10401 4134 10453
rect 4186 10401 4198 10453
rect 4250 10401 4262 10453
rect 4314 10401 4326 10453
rect 4378 10401 4390 10453
rect 4442 10401 5116 10453
rect 9622 10434 9952 10491
rect 452 10384 5116 10401
rect 4284 10380 5116 10384
rect 4948 9746 5116 10380
rect 5161 9987 5347 10085
rect 4948 9488 5118 9746
rect 4958 9219 5118 9488
rect 4958 9163 5010 9219
rect 5066 9163 5118 9219
rect 4958 9139 5118 9163
rect 4958 9083 5010 9139
rect 5066 9083 5118 9139
rect 4958 9059 5118 9083
rect 4958 9003 5010 9059
rect 5066 9003 5118 9059
rect 4958 8979 5118 9003
rect 4958 8923 5010 8979
rect 5066 8923 5118 8979
rect 4958 8899 5118 8923
rect 4958 8843 5010 8899
rect 5066 8843 5118 8899
rect 4958 8790 5118 8843
rect 4946 8032 5122 8696
rect 5161 6163 5347 6257
rect 5161 5947 5186 6163
rect 5322 5947 5347 6163
rect 5161 5914 5347 5947
rect 9712 6144 10990 6175
rect 9712 6124 10774 6144
rect 9712 5988 9751 6124
rect 10447 5988 10774 6124
rect 9712 5964 10774 5988
rect 10954 5964 10990 6144
rect 9712 5935 10990 5964
rect 11178 5410 11806 5412
rect 10636 5407 11806 5410
rect 10636 5355 10656 5407
rect 10708 5382 11806 5407
rect 10708 5355 11212 5382
rect 10636 5343 11212 5355
rect 10636 5291 10656 5343
rect 10708 5291 11212 5343
rect 10636 5279 11212 5291
rect 10636 5227 10656 5279
rect 10708 5227 11212 5279
rect 10636 5215 11212 5227
rect 10636 5163 10656 5215
rect 10708 5163 11212 5215
rect 10636 5151 11212 5163
rect 10636 5099 10656 5151
rect 10708 5099 11212 5151
rect 10636 5087 11212 5099
rect 10636 5035 10656 5087
rect 10708 5035 11212 5087
rect 10636 5023 11212 5035
rect 10636 4971 10656 5023
rect 10708 4971 11212 5023
rect 10636 4959 11212 4971
rect 10636 4907 10656 4959
rect 10708 4926 11212 4959
rect 11748 4926 11806 5382
rect 10708 4907 11806 4926
rect 10636 4905 11806 4907
rect 11178 4898 11806 4905
rect 10371 4330 10452 4332
rect 10371 4278 10385 4330
rect 10437 4278 10452 4330
rect 10371 4266 10452 4278
rect 10371 4214 10385 4266
rect 10437 4227 10452 4266
rect 11142 4230 11804 4264
rect 11142 4227 11806 4230
rect 10437 4224 11806 4227
rect 10437 4214 11215 4224
rect 10371 4202 11215 4214
rect 10371 4150 10385 4202
rect 10437 4168 11215 4202
rect 11271 4168 11295 4224
rect 11351 4168 11375 4224
rect 11431 4168 11455 4224
rect 11511 4168 11535 4224
rect 11591 4168 11615 4224
rect 11671 4168 11695 4224
rect 11751 4168 11806 4224
rect 10437 4150 11806 4168
rect 10371 4148 11806 4150
rect 11142 4146 11806 4148
rect 11142 4130 11804 4146
rect 11196 4128 11804 4130
rect -802 3220 -208 3222
rect -802 3214 -202 3220
rect -802 3183 314 3214
rect -802 3047 -736 3183
rect -280 3047 314 3183
rect -802 3000 314 3047
rect 11012 3065 11097 3096
rect 11012 3019 11027 3065
rect 9331 3013 11027 3019
rect 11079 3013 11097 3065
rect -800 2940 -228 2942
rect -800 2938 -198 2940
rect -800 2903 314 2938
rect 7830 2912 7962 3010
rect 8016 2991 8170 3006
rect 8016 2935 8025 2991
rect 8081 2935 8105 2991
rect 8161 2935 8170 2991
rect 8016 2920 8170 2935
rect 9331 3001 11097 3013
rect 9331 2949 11027 3001
rect 11079 2949 11097 3001
rect 9331 2919 11097 2949
rect -800 2767 -750 2903
rect -294 2767 314 2903
rect -800 2724 314 2767
rect -800 2718 -198 2724
rect 10368 2416 10488 2418
rect 10366 2394 10488 2416
rect 10366 2342 10396 2394
rect 10448 2384 10488 2394
rect 10448 2382 10532 2384
rect 10448 2378 11921 2382
rect 10448 2342 11772 2378
rect 10366 2330 11772 2342
rect 10366 2278 10396 2330
rect 10448 2322 11772 2330
rect 11828 2322 11852 2378
rect 11908 2322 11921 2378
rect 10448 2316 11921 2322
rect 10448 2278 10478 2316
rect 10366 2266 10478 2278
rect 10366 2214 10396 2266
rect 10448 2214 10478 2266
rect 10366 2202 10478 2214
rect 10366 2150 10396 2202
rect 10448 2150 10478 2202
rect 10366 2122 10478 2150
rect 4192 -566 4352 605
rect 10394 450 10488 480
rect 10394 398 10413 450
rect 10465 424 10488 450
rect 11266 468 11380 490
rect 11266 424 11300 468
rect 10465 416 11300 424
rect 11352 416 11380 468
rect 10465 404 11380 416
rect 10465 398 11300 404
rect 10394 386 11300 398
rect 10394 334 10413 386
rect 10465 352 11300 386
rect 11352 352 11380 404
rect 10465 340 11380 352
rect 10465 334 11300 340
rect 10394 322 11300 334
rect 10394 270 10413 322
rect 10465 296 11300 322
rect 10465 270 10488 296
rect 10394 236 10488 270
rect 11266 288 11300 296
rect 11352 288 11380 340
rect 11266 260 11380 288
rect 8020 -55 9022 -42
rect 8020 -57 8047 -55
rect 8103 -57 8127 -55
rect 8183 -57 8207 -55
rect 8263 -57 8287 -55
rect 8343 -57 8367 -55
rect 8423 -57 8447 -55
rect 8503 -57 8527 -55
rect 8583 -57 8607 -55
rect 8663 -57 8687 -55
rect 8743 -57 8767 -55
rect 8823 -57 8847 -55
rect 8903 -57 8927 -55
rect 8983 -57 9022 -55
rect 8020 -109 8041 -57
rect 8103 -109 8105 -57
rect 8285 -109 8287 -57
rect 8349 -109 8361 -57
rect 8423 -109 8425 -57
rect 8605 -109 8607 -57
rect 8669 -109 8681 -57
rect 8743 -109 8745 -57
rect 8925 -109 8927 -57
rect 8989 -109 9022 -57
rect 8020 -111 8047 -109
rect 8103 -111 8127 -109
rect 8183 -111 8207 -109
rect 8263 -111 8287 -109
rect 8343 -111 8367 -109
rect 8423 -111 8447 -109
rect 8503 -111 8527 -109
rect 8583 -111 8607 -109
rect 8663 -111 8687 -109
rect 8743 -111 8767 -109
rect 8823 -111 8847 -109
rect 8903 -111 8927 -109
rect 8983 -111 9022 -109
rect 8020 -128 9022 -111
rect 9106 -162 9306 -158
rect 9058 -179 9306 -162
rect 9058 -551 9092 -179
rect 9208 -551 9306 -179
rect 9058 -566 9306 -551
rect 4192 -578 7998 -566
rect 4192 -600 9026 -578
rect 4192 -716 8052 -600
rect 9000 -628 9026 -600
rect 9000 -716 9020 -628
rect 4192 -726 9020 -716
rect 7726 -736 9020 -726
rect 8024 -740 9020 -736
rect 9106 -644 9306 -566
rect 10416 -644 10532 -466
rect 9106 -673 10532 -644
rect 9106 -806 9504 -673
rect 9096 -969 9504 -806
rect 10040 -714 10532 -673
rect 10040 -766 10443 -714
rect 10495 -766 10532 -714
rect 10040 -778 10532 -766
rect 10040 -830 10443 -778
rect 10495 -804 10532 -778
rect 10495 -830 10534 -804
rect 10040 -842 10534 -830
rect 10040 -894 10443 -842
rect 10495 -894 10534 -842
rect 10040 -969 10534 -894
rect 9096 -1076 10534 -969
rect 9096 -1078 10440 -1076
rect 9910 -1120 11698 -1116
rect 9910 -1128 11710 -1120
rect 9910 -1167 10001 -1128
rect 11589 -1138 11710 -1128
rect 11589 -1167 11808 -1138
rect 9910 -1383 9984 -1167
rect 11720 -1383 11808 -1167
rect 9910 -1396 11808 -1383
rect 10796 -1404 11808 -1396
<< via2 >>
rect 6043 10873 6099 10929
rect 6123 10873 6179 10929
rect 6203 10873 6259 10929
rect 6283 10873 6339 10929
rect -174 10760 202 10770
rect -174 10644 -172 10760
rect -172 10644 200 10760
rect 200 10644 202 10760
rect -174 10634 202 10644
rect 9669 10491 9885 10707
rect 5010 9163 5066 9219
rect 5010 9083 5066 9139
rect 5010 9003 5066 9059
rect 5010 8923 5066 8979
rect 5010 8843 5066 8899
rect 5186 5947 5322 6163
rect 9751 5988 10447 6124
rect 11212 4926 11748 5382
rect 11215 4168 11271 4224
rect 11295 4168 11351 4224
rect 11375 4168 11431 4224
rect 11455 4168 11511 4224
rect 11535 4168 11591 4224
rect 11615 4168 11671 4224
rect 11695 4168 11751 4224
rect -736 3047 -280 3183
rect 8025 2935 8081 2991
rect 8105 2935 8161 2991
rect -750 2767 -294 2903
rect 11772 2322 11828 2378
rect 11852 2322 11908 2378
rect 8047 -57 8103 -55
rect 8127 -57 8183 -55
rect 8207 -57 8263 -55
rect 8287 -57 8343 -55
rect 8367 -57 8423 -55
rect 8447 -57 8503 -55
rect 8527 -57 8583 -55
rect 8607 -57 8663 -55
rect 8687 -57 8743 -55
rect 8767 -57 8823 -55
rect 8847 -57 8903 -55
rect 8927 -57 8983 -55
rect 8047 -109 8093 -57
rect 8093 -109 8103 -57
rect 8127 -109 8157 -57
rect 8157 -109 8169 -57
rect 8169 -109 8183 -57
rect 8207 -109 8221 -57
rect 8221 -109 8233 -57
rect 8233 -109 8263 -57
rect 8287 -109 8297 -57
rect 8297 -109 8343 -57
rect 8367 -109 8413 -57
rect 8413 -109 8423 -57
rect 8447 -109 8477 -57
rect 8477 -109 8489 -57
rect 8489 -109 8503 -57
rect 8527 -109 8541 -57
rect 8541 -109 8553 -57
rect 8553 -109 8583 -57
rect 8607 -109 8617 -57
rect 8617 -109 8663 -57
rect 8687 -109 8733 -57
rect 8733 -109 8743 -57
rect 8767 -109 8797 -57
rect 8797 -109 8809 -57
rect 8809 -109 8823 -57
rect 8847 -109 8861 -57
rect 8861 -109 8873 -57
rect 8873 -109 8903 -57
rect 8927 -109 8937 -57
rect 8937 -109 8983 -57
rect 8047 -111 8103 -109
rect 8127 -111 8183 -109
rect 8207 -111 8263 -109
rect 8287 -111 8343 -109
rect 8367 -111 8423 -109
rect 8447 -111 8503 -109
rect 8527 -111 8583 -109
rect 8607 -111 8663 -109
rect 8687 -111 8743 -109
rect 8767 -111 8823 -109
rect 8847 -111 8903 -109
rect 8927 -111 8983 -109
rect 9504 -969 10040 -673
rect 9984 -1372 10001 -1167
rect 10001 -1372 11589 -1167
rect 11589 -1372 11720 -1167
rect 9984 -1383 11720 -1372
<< metal3 >>
rect 6206 11004 6366 11008
rect 5988 10929 6414 11004
rect 5988 10873 6043 10929
rect 6099 10873 6123 10929
rect 6179 10873 6203 10929
rect 6259 10873 6283 10929
rect 6339 10873 6414 10929
rect 5988 10814 6414 10873
rect -200 10774 270 10802
rect -200 10630 -178 10774
rect 206 10630 270 10774
rect -200 10602 270 10630
rect -804 10030 -206 10038
rect -804 9976 -198 10030
rect -804 9832 -781 9976
rect -237 9832 -198 9976
rect -804 9788 -198 9832
rect -804 9778 -200 9788
rect 4958 9219 5118 9270
rect 4958 9163 5010 9219
rect 5066 9163 5118 9219
rect 4958 9139 5118 9163
rect 4958 9083 5010 9139
rect 5066 9083 5118 9139
rect 4958 9059 5118 9083
rect 4958 9003 5010 9059
rect 5066 9003 5118 9059
rect 4958 8979 5118 9003
rect 4958 8923 5010 8979
rect 5066 8923 5118 8979
rect 4958 8899 5118 8923
rect 4958 8843 5010 8899
rect 5066 8843 5118 8899
rect 4958 8696 5118 8843
rect 4946 8694 5122 8696
rect 4774 8534 5122 8694
rect 4946 8032 5122 8534
rect 840 5782 900 6482
rect 1884 6137 1944 6464
rect 6206 6455 6366 10814
rect 9622 10711 9956 10748
rect 9622 10487 9665 10711
rect 9889 10487 9956 10711
rect 9622 10434 9956 10487
rect 11002 10004 11800 10006
rect 11000 9973 11800 10004
rect 11000 9829 11040 9973
rect 11744 9829 11800 9973
rect 11000 9770 11800 9829
rect 5154 6175 5358 6184
rect 1137 6077 1944 6137
rect 2077 6163 10490 6175
rect 2077 6126 5186 6163
rect 1137 5787 1197 6077
rect 2077 5982 2097 6126
rect 2481 5982 5186 6126
rect 2077 5947 5186 5982
rect 5322 6124 10490 6163
rect 5322 5988 9751 6124
rect 10447 5988 10490 6124
rect 5322 5947 10490 5988
rect 2077 5935 10490 5947
rect 5154 5927 5358 5935
rect 11186 5382 11810 5418
rect 11186 4926 11212 5382
rect 11748 4926 11810 5382
rect 11186 4896 11810 4926
rect 11138 4264 11800 4300
rect 11138 4224 11804 4264
rect 11138 4168 11215 4224
rect 11271 4168 11295 4224
rect 11351 4168 11375 4224
rect 11431 4168 11455 4224
rect 11511 4168 11535 4224
rect 11591 4168 11615 4224
rect 11671 4168 11695 4224
rect 11751 4168 11804 4224
rect 11138 4128 11804 4168
rect 11138 4122 11800 4128
rect -802 3220 -208 3222
rect -804 3214 -202 3220
rect -804 3183 -198 3214
rect -804 3047 -736 3183
rect -280 3047 -198 3183
rect -804 3002 -198 3047
rect -804 3000 -204 3002
rect 7994 2991 8180 3012
rect -804 2903 -198 2940
rect 7994 2935 8025 2991
rect 8081 2935 8105 2991
rect 8161 2935 8180 2991
rect 7994 2912 8180 2935
rect -804 2767 -750 2903
rect -294 2767 -198 2903
rect 8042 2884 8132 2912
rect -804 2720 -198 2767
rect -796 2718 -198 2720
rect 8046 -40 8130 2884
rect 11762 2378 11918 2384
rect 11762 2322 11772 2378
rect 11828 2322 11852 2378
rect 11908 2322 11918 2378
rect 11762 2316 11918 2322
rect 8020 -55 9022 -40
rect 8020 -111 8047 -55
rect 8103 -111 8127 -55
rect 8183 -111 8207 -55
rect 8263 -111 8287 -55
rect 8343 -111 8367 -55
rect 8423 -111 8447 -55
rect 8503 -111 8527 -55
rect 8583 -111 8607 -55
rect 8663 -111 8687 -55
rect 8743 -111 8767 -55
rect 8823 -111 8847 -55
rect 8903 -111 8927 -55
rect 8983 -111 9022 -55
rect 8020 -126 9022 -111
rect 9472 -669 10072 -644
rect 9472 -973 9500 -669
rect 10044 -973 10072 -669
rect 9472 -1018 10072 -973
rect 9920 -1136 11710 -1120
rect 9906 -1167 11818 -1136
rect 9906 -1383 9984 -1167
rect 11720 -1383 11818 -1167
rect 9906 -1404 11818 -1383
rect 9906 -1412 11814 -1404
<< via3 >>
rect -178 10770 206 10774
rect -178 10634 -174 10770
rect -174 10634 202 10770
rect 202 10634 206 10770
rect -178 10630 206 10634
rect -781 9832 -237 9976
rect 9665 10707 9889 10711
rect 9665 10491 9669 10707
rect 9669 10491 9885 10707
rect 9885 10491 9889 10707
rect 9665 10487 9889 10491
rect 11040 9829 11744 9973
rect 2097 5982 2481 6126
rect 9500 -673 10044 -669
rect 9500 -969 9504 -673
rect 9504 -969 10040 -673
rect 10040 -969 10044 -673
rect 9500 -973 10044 -969
<< metal4 >>
rect -276 10774 270 10802
rect -276 10630 -178 10774
rect 206 10630 270 10774
rect -276 10602 270 10630
rect 9622 10717 9956 10748
rect -276 10032 -170 10602
rect 9622 10481 9659 10717
rect 9895 10481 9956 10717
rect 9622 10434 9956 10481
rect 485 10032 1685 10036
rect -804 9976 1685 10032
rect -804 9832 -781 9976
rect -237 9832 1685 9976
rect -804 9784 1685 9832
rect 485 9775 1685 9784
rect 2770 10004 3970 10036
rect 2770 9973 11796 10004
rect 2770 9829 11040 9973
rect 11744 9829 11796 9973
rect 2770 9770 11796 9829
rect 485 6173 1685 6232
rect 485 6126 2501 6173
rect 2769 6136 5221 6856
rect 485 5982 2097 6126
rect 2481 5982 2501 6126
rect 485 5934 2501 5982
rect 485 5604 1685 5934
rect 4501 5601 5221 6136
rect 9472 -669 10072 -644
rect 9472 -973 9500 -669
rect 10044 -973 10072 -669
rect 9472 -1018 10072 -973
<< via4 >>
rect 9659 10711 9895 10717
rect 9659 10487 9665 10711
rect 9665 10487 9889 10711
rect 9889 10487 9895 10711
rect 9659 10481 9895 10487
rect 9652 -942 9888 -706
<< metal5 >>
rect 9622 10717 9960 10766
rect 9622 10481 9659 10717
rect 9895 10481 9960 10717
rect 9622 10434 9960 10481
rect 9626 -644 9948 10434
rect 9472 -706 10072 -644
rect 9472 -942 9652 -706
rect 9888 -942 10072 -706
rect 9472 -1018 10072 -942
use comparator  comparator_0
timestamp 1699953975
transform 1 0 -507679 0 1 -639888
box 507669 639956 517124 645817
use comparator_bias  comparator_bias_0
timestamp 1699953975
transform -1 0 518454 0 1 -639855
box 507806 646042 518382 649916
use sky130_fd_pr__nfet_g5v0d10v5_SM3UA9  sky130_fd_pr__nfet_g5v0d10v5_SM3UA9_0
timestamp 1699953975
transform 0 1 8524 -1 0 -362
box -418 -748 418 748
use sky130_fd_pr__pfet_g5v0d10v5_H5W24A  sky130_fd_pr__pfet_g5v0d10v5_H5W24A_0
timestamp 1699953975
transform 0 1 2449 -1 0 10686
box -458 -2297 458 2297
use sky130_fd_sc_hvl__inv_4  sky130_fd_sc_hvl__inv_4_0
timestamp 1699954036
transform 0 1 10115 -1 0 152
box -66 -43 834 897
use sky130_fd_sc_hvl__lsbufhv2lv_1  sky130_fd_sc_hvl__lsbufhv2lv_1_0
timestamp 1699953975
transform 0 1 10050 1 0 3048
box -66 -43 1698 1671
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0
timestamp 1699954036
transform 0 1 10051 -1 0 2650
box -66 -43 2178 1671
<< labels >>
flabel metal3 s -804 9786 -206 10038 0 FreeSans 1455 0 0 0 VDD
port 1 nsew
flabel metal3 s -804 3000 -204 3220 0 FreeSans 1455 0 0 0 VINP
port 2 nsew
flabel metal3 s -804 2720 -204 2940 0 FreeSans 1455 0 0 0 VINM
port 3 nsew
flabel metal3 s 11002 9778 11800 10006 0 FreeSans 1455 0 0 0 VSS
port 4 nsew
flabel metal3 s 11186 4896 11810 5418 0 FreeSans 1455 0 0 0 DVDD
port 5 nsew
flabel metal3 s 11138 4122 11800 4300 0 FreeSans 1455 0 0 0 VOUT
port 6 nsew
flabel metal3 s 10802 -1404 11818 -1136 0 FreeSans 1455 0 0 0 DVSS
port 7 nsew
flabel metal3 s 11762 2316 11918 2384 0 FreeSans 244 0 0 0 EN
port 8 nsew
<< end >>
