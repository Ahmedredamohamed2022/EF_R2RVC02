VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_R2RVC02
  CLASS BLOCK ;
  FOREIGN EF_R2RVC02 ;
  ORIGIN 0.000 0.000 ;
  SIZE 82.070 BY 134.140 ;
  PIN SELA
    ANTENNAGATEAREA 4.752000 ;
    PORT
      LAYER met2 ;
        RECT 11.040 0.100 11.720 3.120 ;
    END
  END SELA
  PIN SELB
    ANTENNAGATEAREA 4.752000 ;
    PORT
      LAYER met2 ;
        RECT 44.040 0.000 44.730 3.040 ;
    END
  END SELB
  PIN A1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 22.700 0.020 23.260 3.050 ;
    END
  END A1
  PIN A2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 39.710 0.030 40.270 3.080 ;
    END
  END A2
  PIN B1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 55.670 0.050 56.220 3.090 ;
    END
  END B1
  PIN B2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met2 ;
        RECT 72.700 0.050 73.230 3.060 ;
    END
  END B2
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 598.042908 ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.300 4.110 44.300 ;
    END
  END VDD
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 271.063080 ;
    PORT
      LAYER met3 ;
        RECT 0.000 72.540 3.060 73.610 ;
    END
  END VSS
  PIN DVSS
    ANTENNADIFFAREA 215.901642 ;
    PORT
      LAYER met3 ;
        RECT 78.270 69.370 82.040 70.720 ;
    END
  END DVSS
  PIN DVDD
    ANTENNADIFFAREA 9.946099 ;
    PORT
      LAYER met3 ;
        RECT 78.960 100.890 82.040 103.470 ;
    END
  END DVDD
  PIN VO
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met3 ;
        RECT 79.020 97.030 82.050 97.910 ;
    END
  END VO
  PIN EN
    ANTENNAGATEAREA 0.252000 ;
    PORT
      LAYER met3 ;
        RECT 78.970 87.950 82.020 88.310 ;
    END
  END EN
  OBS
      LAYER li1 ;
        RECT 9.385 3.950 73.485 131.695 ;
      LAYER met1 ;
        RECT 8.995 3.540 76.015 131.585 ;
      LAYER met2 ;
        RECT 6.020 3.400 76.040 131.385 ;
        RECT 6.020 0.035 10.760 3.400 ;
        RECT 12.000 3.370 76.040 3.400 ;
        RECT 12.000 3.360 55.390 3.370 ;
        RECT 12.000 3.330 39.430 3.360 ;
        RECT 12.000 0.035 22.420 3.330 ;
        RECT 23.540 0.035 39.430 3.330 ;
        RECT 40.550 3.320 55.390 3.360 ;
        RECT 40.550 0.035 43.760 3.320 ;
        RECT 45.010 0.035 55.390 3.320 ;
        RECT 56.500 3.340 76.040 3.370 ;
        RECT 56.500 0.035 72.420 3.340 ;
        RECT 73.510 0.035 76.040 3.340 ;
      LAYER met3 ;
        RECT 0.070 103.870 82.070 131.405 ;
        RECT 0.070 100.490 78.560 103.870 ;
        RECT 0.070 98.310 82.070 100.490 ;
        RECT 0.070 96.630 78.620 98.310 ;
        RECT 0.070 88.710 82.070 96.630 ;
        RECT 0.070 87.550 78.570 88.710 ;
        RECT 0.070 74.010 82.070 87.550 ;
        RECT 3.460 72.140 82.070 74.010 ;
        RECT 0.070 71.120 82.070 72.140 ;
        RECT 0.070 68.970 77.870 71.120 ;
        RECT 0.070 44.700 82.070 68.970 ;
        RECT 4.510 42.900 82.070 44.700 ;
        RECT 0.070 0.040 82.070 42.900 ;
      LAYER met4 ;
        RECT 4.660 0.030 77.490 134.140 ;
      LAYER met5 ;
        RECT 60.420 71.275 63.420 130.195 ;
  END
END EF_R2RVC02
END LIBRARY

