** sch_path: /home/ahmedreda/Project/AR_SAR_ADC/comparator_top_02ch/tb/r2rvc02/r2r_dcsweepvinp.sch
**.subckt r2r_dcsweepvinp
V1 VSS GND 0
.save i(v1)
V2 VDD VSS 3.3
.save i(v2)
C1 VOUT VSS 1p m=1
V5 DVDD VSS 1.8
.save i(v5)
x1 a1 a2 b1 b2 VOUT sela selb DVDD VSS VSS VDD EF_R2RVC02mf
V8 selb VSS 1.8
.save i(v8)
V9 sela VSS 1.8
.save i(v9)
V3 a1 VSS 1.65
.save i(v3)
V4 b1 VSS 1.65
.save i(v4)
V6 b2 VSS 1.65
.save i(v6)
V7 a2 VSS 1.65
.save i(v7)
**** begin user architecture code


**.include /usr/share/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
**.include /ciic/pdk/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /home/ahmedreda/PDK/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl.spice
.include /home/ahmedreda/PDK/sky130A/libs.ref/sky130_fd_sc_hvl/spice/sky130_fd_sc_hvl__lsbuflv2hv_1.spice


.lib /home/ahmedreda/PDK/sky130A/libs.tech/ngspice/sky130.lib.spice tt
.include EF_R2RVC02mf.spice


.option wnflag=1
.option TEMP=27
.option TNOM=27
.option wnflag=1
.control
**set filetype=binary
set filetype=ascii
set color0=white
set color1=black
set color3=blue
set xbrushwidth=3
save all
run
op
dc V3 0 3.3 0.01
let icom=abs(v2#branch)
let ibuf=abs(v5#branch)
let itot=icom+ibuf
let voutdigital=vout
plot vinp voutdigital vinm
meas dc offset1 WHEN vinp=1.65
meas dc offset2 FIND vout AT=1.65

plot itot
meas dc itot_1.65 FIND itot AT=1.65
meas dc itot_0 FIND itot AT=0.01
meas dc itot_3.3 FIND itot AT=3.29
meas dc offset_actual WHEN voutdigital=0.9

print (offset_actual-1.65)*1000


.endc






.GLOBAL GND
.end
