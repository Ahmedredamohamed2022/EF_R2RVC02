VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO EF_R2RVC02
  CLASS BLOCK ;
  FOREIGN EF_R2RVC02 ;
  ORIGIN 6.335 40.265 ;
  SIZE 76.095 BY 96.105 ;
  PIN vo
    ANTENNADIFFAREA 0.492900 ;
    PORT
      LAYER met2 ;
        RECT 59.480 22.190 59.700 22.320 ;
    END
  END vo
  PIN B2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 63.110 -21.940 63.650 -21.250 ;
    END
  END B2
  PIN B1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 46.320 -21.650 46.950 -21.050 ;
    END
  END B1
  PIN A2
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 30.100 -22.570 30.560 -21.850 ;
    END
  END A2
  PIN A1
    ANTENNADIFFAREA 2.610000 ;
    PORT
      LAYER met1 ;
        RECT 13.310 -22.370 13.660 -21.680 ;
    END
  END A1
  PIN SELB
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 41.490 -38.270 41.920 -37.890 ;
    END
  END SELB
  PIN SELA
    ANTENNAGATEAREA 2.502000 ;
    PORT
      LAYER met1 ;
        RECT 7.160 -38.210 7.710 -37.870 ;
    END
  END SELA
  PIN DVSS
    ANTENNADIFFAREA 107.239799 ;
    PORT
      LAYER met4 ;
        RECT 66.650 -35.270 66.910 -34.880 ;
    END
  END DVSS
  PIN DVDD
    ANTENNADIFFAREA 7.633700 ;
    PORT
      LAYER met4 ;
        RECT 68.730 -37.200 69.180 -36.730 ;
    END
  END DVDD
  PIN VSS
    ANTENNAGATEAREA 130.000000 ;
    ANTENNADIFFAREA 263.488281 ;
    PORT
      LAYER met3 ;
        RECT -1.880 53.010 -1.650 53.500 ;
    END
  END VSS
  PIN VDD
    ANTENNAGATEAREA 100.000000 ;
    ANTENNADIFFAREA 433.882782 ;
    PORT
      LAYER met4 ;
        RECT -5.320 55.040 -4.940 55.380 ;
    END
  END VDD
  OBS
      LAYER li1 ;
        RECT 0.330 -39.890 64.300 52.065 ;
      LAYER met1 ;
        RECT -0.130 -20.770 67.280 51.750 ;
        RECT -0.130 -21.400 46.040 -20.770 ;
        RECT -0.130 -22.650 13.030 -21.400 ;
        RECT 13.940 -21.570 46.040 -21.400 ;
        RECT 13.940 -22.650 29.820 -21.570 ;
        RECT -0.130 -22.850 29.820 -22.650 ;
        RECT 30.840 -21.930 46.040 -21.570 ;
        RECT 47.230 -20.970 67.280 -20.770 ;
        RECT 47.230 -21.930 62.830 -20.970 ;
        RECT 30.840 -22.220 62.830 -21.930 ;
        RECT 63.930 -22.220 67.280 -20.970 ;
        RECT 30.840 -22.850 67.280 -22.220 ;
        RECT -0.130 -37.590 67.280 -22.850 ;
        RECT -0.130 -38.490 6.880 -37.590 ;
        RECT 7.990 -37.610 67.280 -37.590 ;
        RECT 7.990 -38.490 41.210 -37.610 ;
        RECT -0.130 -38.550 41.210 -38.490 ;
        RECT 42.200 -38.550 67.280 -37.610 ;
        RECT -0.130 -40.050 67.280 -38.550 ;
      LAYER met2 ;
        RECT -1.080 22.600 69.520 51.750 ;
        RECT -1.080 21.910 59.200 22.600 ;
        RECT 59.980 21.910 69.520 22.600 ;
        RECT -1.080 -40.050 69.520 21.910 ;
      LAYER met3 ;
        RECT -6.335 53.900 69.760 54.380 ;
        RECT -6.335 52.610 -2.280 53.900 ;
        RECT -1.250 52.610 69.760 53.900 ;
        RECT -6.335 -40.050 69.760 52.610 ;
      LAYER met4 ;
        RECT -6.310 55.780 69.760 55.840 ;
        RECT -6.310 54.640 -5.720 55.780 ;
        RECT -4.540 54.640 69.760 55.780 ;
        RECT -6.310 -34.480 69.760 54.640 ;
        RECT -6.310 -35.670 66.250 -34.480 ;
        RECT 67.310 -35.670 69.760 -34.480 ;
        RECT -6.310 -36.330 69.760 -35.670 ;
        RECT -6.310 -37.600 68.330 -36.330 ;
        RECT 69.580 -37.600 69.760 -36.330 ;
        RECT -6.310 -40.150 69.760 -37.600 ;
  END
END EF_R2RVC02
END LIBRARY

