magic
tech sky130A
magscale 1 2
timestamp 1694943448
<< nwell >>
rect 1790 604 2054 660
<< locali >>
rect 2044 1339 2206 1372
rect 2044 1233 2069 1339
rect 2175 1233 2206 1339
rect 2044 1192 2206 1233
rect 282 418 544 452
rect 282 312 322 418
rect 500 312 544 418
rect 282 286 544 312
<< viali >>
rect 2069 1233 2175 1339
rect 322 312 500 418
<< metal1 >>
rect -14 1660 2118 1698
rect -14 1544 17 1660
rect 133 1544 2118 1660
rect -14 1500 2118 1544
rect 2044 1339 2206 1372
rect 2044 1233 2069 1339
rect 2175 1233 2206 1339
rect 2044 1192 2206 1233
rect -14 714 336 942
rect 884 870 1158 936
rect 886 798 1196 836
rect 892 700 1208 762
rect 218 604 482 660
rect 902 606 1204 660
rect 1790 604 2054 660
rect 282 418 544 452
rect 282 312 322 418
rect 500 312 544 418
rect 282 286 544 312
rect -14 94 2126 138
rect -14 -22 15 94
rect 131 -22 2126 94
rect -14 -58 2126 -22
<< via1 >>
rect 17 1544 133 1660
rect 15 -22 131 94
<< metal2 >>
rect -10 1660 162 1696
rect -10 1544 17 1660
rect 133 1544 162 1660
rect -10 94 162 1544
rect -10 -22 15 94
rect 131 -22 162 94
rect -10 -54 162 -22
use sky130_fd_sc_hvl__lsbuflv2hv_1  sky130_fd_sc_hvl__lsbuflv2hv_1_0
timestamp 1694943448
transform 1 0 0 0 1 0
box -66 -43 2178 1671
<< labels >>
flabel metal1 s 358 76 404 96 0 FreeSans 555 0 0 0 vss1p8
port 1 nsew
flabel metal1 s 400 438 418 444 0 FreeSans 555 0 0 0 A
port 2 nsew
flabel metal1 s 2194 1266 2202 1282 0 FreeSans 555 0 0 0 X
port 3 nsew
flabel metal1 s 1896 620 1922 640 0 FreeSans 333 0 0 0 vdd1p8
port 4 nsew
flabel metal1 s 210 806 254 826 0 FreeSans 333 0 0 0 vdd3p3
port 5 nsew
<< end >>
