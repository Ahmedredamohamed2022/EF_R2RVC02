magic
tech sky130A
magscale 1 2
timestamp 1699954036
<< metal1 >>
rect 2103 2840 2454 2946
rect 2103 1 2209 2840
rect 4120 2183 4442 2190
rect 4120 2003 4127 2183
rect 4435 2003 4442 2183
rect 4120 1996 4442 2003
rect 4418 1702 4604 1732
rect 4650 1702 4754 4142
rect 4418 1598 4754 1702
rect 4418 1540 4604 1598
rect 2238 1202 2598 1306
rect 2238 0 2342 1202
rect 3846 420 4488 422
rect 3846 240 3853 420
rect 4481 240 4488 420
rect 3846 238 4488 240
<< via1 >>
rect 4127 2003 4435 2183
rect 3853 240 4481 420
<< metal2 >>
rect 4108 2212 4466 2214
rect 4108 2183 4496 2212
rect 4108 2003 4127 2183
rect 4435 2003 4496 2183
rect 4108 1984 4496 2003
rect 4108 1980 4466 1984
rect 3790 438 4538 450
rect 3788 420 4538 438
rect 3788 240 3853 420
rect 4481 240 4538 420
rect 3788 214 4538 240
use tg4dm  tg4dm_1
timestamp 1699954036
transform 1 0 2091 0 1 2311
box 301 -2311 2543 1830
<< labels >>
flabel metal1 s 2238 0 2342 104 0 FreeSans 48 0 0 0 VIN
port 1 nsew
flabel metal2 s 4198 2048 4370 2158 0 FreeSans 116 0 0 0 VDD
port 2 nsew
flabel metal2 s 4268 288 4440 398 0 FreeSans 116 0 0 0 VSS
port 3 nsew
flabel metal1 s 4650 4038 4754 4142 0 FreeSans 116 0 0 0 VOUT
port 4 nsew
flabel metal1 s 2103 1 2209 107 0 FreeSans 48 0 0 0 SEL
port 5 nsew
<< end >>
