magic
tech sky130A
magscale 1 2
timestamp 1694943448
<< nwell >>
rect 507754 642939 517040 645817
<< pwell >>
rect 507794 639956 517000 642754
<< mvnmos >>
rect 508114 641405 508514 642405
rect 508572 641405 508972 642405
rect 509030 641405 509430 642405
rect 509488 641405 509888 642405
rect 509946 641405 510346 642405
rect 510404 641405 510804 642405
rect 510862 641405 511262 642405
rect 511320 641405 511720 642405
rect 511778 641405 512178 642405
rect 512236 641405 512636 642405
rect 512694 641405 513094 642405
rect 513152 641405 513552 642405
rect 513610 641405 514010 642405
rect 514068 641405 514468 642405
rect 514526 641405 514926 642405
rect 514984 641405 515384 642405
rect 508114 640243 508514 641243
rect 508572 640243 508972 641243
rect 509030 640243 509430 641243
rect 509488 640243 509888 641243
rect 509946 640243 510346 641243
rect 510404 640243 510804 641243
rect 510862 640243 511262 641243
rect 511320 640243 511720 641243
rect 511778 640243 512178 641243
rect 512236 640243 512636 641243
rect 512694 640243 513094 641243
rect 513152 640243 513552 641243
rect 513610 640243 514010 641243
rect 514068 640243 514468 641243
rect 514526 640243 514926 641243
rect 514984 640243 515384 641243
rect 515818 641405 516218 642405
rect 516276 641405 516676 642405
<< mvpmos >>
rect 508114 644503 508514 645503
rect 508572 644503 508972 645503
rect 509030 644503 509430 645503
rect 509488 644503 509888 645503
rect 509946 644503 510346 645503
rect 510404 644503 510804 645503
rect 510862 644503 511262 645503
rect 511320 644503 511720 645503
rect 511778 644503 512178 645503
rect 512236 644503 512636 645503
rect 512694 644503 513094 645503
rect 513152 644503 513552 645503
rect 513610 644503 514010 645503
rect 514068 644503 514468 645503
rect 514526 644503 514926 645503
rect 514984 644503 515384 645503
rect 508114 643337 508514 644337
rect 508572 643337 508972 644337
rect 509030 643337 509430 644337
rect 509488 643337 509888 644337
rect 509946 643337 510346 644337
rect 510404 643337 510804 644337
rect 510862 643337 511262 644337
rect 511320 643337 511720 644337
rect 511778 643337 512178 644337
rect 512236 643337 512636 644337
rect 512694 643337 513094 644337
rect 513152 643337 513552 644337
rect 513610 643337 514010 644337
rect 514068 643337 514468 644337
rect 514526 643337 514926 644337
rect 514984 643337 515384 644337
rect 515818 643337 516218 645337
rect 516276 643337 516676 645337
<< mvndiff >>
rect 508056 642364 508114 642405
rect 508056 642330 508068 642364
rect 508102 642330 508114 642364
rect 508056 642296 508114 642330
rect 508056 642262 508068 642296
rect 508102 642262 508114 642296
rect 508056 642228 508114 642262
rect 508056 642194 508068 642228
rect 508102 642194 508114 642228
rect 508056 642160 508114 642194
rect 508056 642126 508068 642160
rect 508102 642126 508114 642160
rect 508056 642092 508114 642126
rect 508056 642058 508068 642092
rect 508102 642058 508114 642092
rect 508056 642024 508114 642058
rect 508056 641990 508068 642024
rect 508102 641990 508114 642024
rect 508056 641956 508114 641990
rect 508056 641922 508068 641956
rect 508102 641922 508114 641956
rect 508056 641888 508114 641922
rect 508056 641854 508068 641888
rect 508102 641854 508114 641888
rect 508056 641820 508114 641854
rect 508056 641786 508068 641820
rect 508102 641786 508114 641820
rect 508056 641752 508114 641786
rect 508056 641718 508068 641752
rect 508102 641718 508114 641752
rect 508056 641684 508114 641718
rect 508056 641650 508068 641684
rect 508102 641650 508114 641684
rect 508056 641616 508114 641650
rect 508056 641582 508068 641616
rect 508102 641582 508114 641616
rect 508056 641548 508114 641582
rect 508056 641514 508068 641548
rect 508102 641514 508114 641548
rect 508056 641480 508114 641514
rect 508056 641446 508068 641480
rect 508102 641446 508114 641480
rect 508056 641405 508114 641446
rect 508514 642364 508572 642405
rect 508514 642330 508526 642364
rect 508560 642330 508572 642364
rect 508514 642296 508572 642330
rect 508514 642262 508526 642296
rect 508560 642262 508572 642296
rect 508514 642228 508572 642262
rect 508514 642194 508526 642228
rect 508560 642194 508572 642228
rect 508514 642160 508572 642194
rect 508514 642126 508526 642160
rect 508560 642126 508572 642160
rect 508514 642092 508572 642126
rect 508514 642058 508526 642092
rect 508560 642058 508572 642092
rect 508514 642024 508572 642058
rect 508514 641990 508526 642024
rect 508560 641990 508572 642024
rect 508514 641956 508572 641990
rect 508514 641922 508526 641956
rect 508560 641922 508572 641956
rect 508514 641888 508572 641922
rect 508514 641854 508526 641888
rect 508560 641854 508572 641888
rect 508514 641820 508572 641854
rect 508514 641786 508526 641820
rect 508560 641786 508572 641820
rect 508514 641752 508572 641786
rect 508514 641718 508526 641752
rect 508560 641718 508572 641752
rect 508514 641684 508572 641718
rect 508514 641650 508526 641684
rect 508560 641650 508572 641684
rect 508514 641616 508572 641650
rect 508514 641582 508526 641616
rect 508560 641582 508572 641616
rect 508514 641548 508572 641582
rect 508514 641514 508526 641548
rect 508560 641514 508572 641548
rect 508514 641480 508572 641514
rect 508514 641446 508526 641480
rect 508560 641446 508572 641480
rect 508514 641405 508572 641446
rect 508972 642364 509030 642405
rect 508972 642330 508984 642364
rect 509018 642330 509030 642364
rect 508972 642296 509030 642330
rect 508972 642262 508984 642296
rect 509018 642262 509030 642296
rect 508972 642228 509030 642262
rect 508972 642194 508984 642228
rect 509018 642194 509030 642228
rect 508972 642160 509030 642194
rect 508972 642126 508984 642160
rect 509018 642126 509030 642160
rect 508972 642092 509030 642126
rect 508972 642058 508984 642092
rect 509018 642058 509030 642092
rect 508972 642024 509030 642058
rect 508972 641990 508984 642024
rect 509018 641990 509030 642024
rect 508972 641956 509030 641990
rect 508972 641922 508984 641956
rect 509018 641922 509030 641956
rect 508972 641888 509030 641922
rect 508972 641854 508984 641888
rect 509018 641854 509030 641888
rect 508972 641820 509030 641854
rect 508972 641786 508984 641820
rect 509018 641786 509030 641820
rect 508972 641752 509030 641786
rect 508972 641718 508984 641752
rect 509018 641718 509030 641752
rect 508972 641684 509030 641718
rect 508972 641650 508984 641684
rect 509018 641650 509030 641684
rect 508972 641616 509030 641650
rect 508972 641582 508984 641616
rect 509018 641582 509030 641616
rect 508972 641548 509030 641582
rect 508972 641514 508984 641548
rect 509018 641514 509030 641548
rect 508972 641480 509030 641514
rect 508972 641446 508984 641480
rect 509018 641446 509030 641480
rect 508972 641405 509030 641446
rect 509430 642364 509488 642405
rect 509430 642330 509442 642364
rect 509476 642330 509488 642364
rect 509430 642296 509488 642330
rect 509430 642262 509442 642296
rect 509476 642262 509488 642296
rect 509430 642228 509488 642262
rect 509430 642194 509442 642228
rect 509476 642194 509488 642228
rect 509430 642160 509488 642194
rect 509430 642126 509442 642160
rect 509476 642126 509488 642160
rect 509430 642092 509488 642126
rect 509430 642058 509442 642092
rect 509476 642058 509488 642092
rect 509430 642024 509488 642058
rect 509430 641990 509442 642024
rect 509476 641990 509488 642024
rect 509430 641956 509488 641990
rect 509430 641922 509442 641956
rect 509476 641922 509488 641956
rect 509430 641888 509488 641922
rect 509430 641854 509442 641888
rect 509476 641854 509488 641888
rect 509430 641820 509488 641854
rect 509430 641786 509442 641820
rect 509476 641786 509488 641820
rect 509430 641752 509488 641786
rect 509430 641718 509442 641752
rect 509476 641718 509488 641752
rect 509430 641684 509488 641718
rect 509430 641650 509442 641684
rect 509476 641650 509488 641684
rect 509430 641616 509488 641650
rect 509430 641582 509442 641616
rect 509476 641582 509488 641616
rect 509430 641548 509488 641582
rect 509430 641514 509442 641548
rect 509476 641514 509488 641548
rect 509430 641480 509488 641514
rect 509430 641446 509442 641480
rect 509476 641446 509488 641480
rect 509430 641405 509488 641446
rect 509888 642364 509946 642405
rect 509888 642330 509900 642364
rect 509934 642330 509946 642364
rect 509888 642296 509946 642330
rect 509888 642262 509900 642296
rect 509934 642262 509946 642296
rect 509888 642228 509946 642262
rect 509888 642194 509900 642228
rect 509934 642194 509946 642228
rect 509888 642160 509946 642194
rect 509888 642126 509900 642160
rect 509934 642126 509946 642160
rect 509888 642092 509946 642126
rect 509888 642058 509900 642092
rect 509934 642058 509946 642092
rect 509888 642024 509946 642058
rect 509888 641990 509900 642024
rect 509934 641990 509946 642024
rect 509888 641956 509946 641990
rect 509888 641922 509900 641956
rect 509934 641922 509946 641956
rect 509888 641888 509946 641922
rect 509888 641854 509900 641888
rect 509934 641854 509946 641888
rect 509888 641820 509946 641854
rect 509888 641786 509900 641820
rect 509934 641786 509946 641820
rect 509888 641752 509946 641786
rect 509888 641718 509900 641752
rect 509934 641718 509946 641752
rect 509888 641684 509946 641718
rect 509888 641650 509900 641684
rect 509934 641650 509946 641684
rect 509888 641616 509946 641650
rect 509888 641582 509900 641616
rect 509934 641582 509946 641616
rect 509888 641548 509946 641582
rect 509888 641514 509900 641548
rect 509934 641514 509946 641548
rect 509888 641480 509946 641514
rect 509888 641446 509900 641480
rect 509934 641446 509946 641480
rect 509888 641405 509946 641446
rect 510346 642364 510404 642405
rect 510346 642330 510358 642364
rect 510392 642330 510404 642364
rect 510346 642296 510404 642330
rect 510346 642262 510358 642296
rect 510392 642262 510404 642296
rect 510346 642228 510404 642262
rect 510346 642194 510358 642228
rect 510392 642194 510404 642228
rect 510346 642160 510404 642194
rect 510346 642126 510358 642160
rect 510392 642126 510404 642160
rect 510346 642092 510404 642126
rect 510346 642058 510358 642092
rect 510392 642058 510404 642092
rect 510346 642024 510404 642058
rect 510346 641990 510358 642024
rect 510392 641990 510404 642024
rect 510346 641956 510404 641990
rect 510346 641922 510358 641956
rect 510392 641922 510404 641956
rect 510346 641888 510404 641922
rect 510346 641854 510358 641888
rect 510392 641854 510404 641888
rect 510346 641820 510404 641854
rect 510346 641786 510358 641820
rect 510392 641786 510404 641820
rect 510346 641752 510404 641786
rect 510346 641718 510358 641752
rect 510392 641718 510404 641752
rect 510346 641684 510404 641718
rect 510346 641650 510358 641684
rect 510392 641650 510404 641684
rect 510346 641616 510404 641650
rect 510346 641582 510358 641616
rect 510392 641582 510404 641616
rect 510346 641548 510404 641582
rect 510346 641514 510358 641548
rect 510392 641514 510404 641548
rect 510346 641480 510404 641514
rect 510346 641446 510358 641480
rect 510392 641446 510404 641480
rect 510346 641405 510404 641446
rect 510804 642364 510862 642405
rect 510804 642330 510816 642364
rect 510850 642330 510862 642364
rect 510804 642296 510862 642330
rect 510804 642262 510816 642296
rect 510850 642262 510862 642296
rect 510804 642228 510862 642262
rect 510804 642194 510816 642228
rect 510850 642194 510862 642228
rect 510804 642160 510862 642194
rect 510804 642126 510816 642160
rect 510850 642126 510862 642160
rect 510804 642092 510862 642126
rect 510804 642058 510816 642092
rect 510850 642058 510862 642092
rect 510804 642024 510862 642058
rect 510804 641990 510816 642024
rect 510850 641990 510862 642024
rect 510804 641956 510862 641990
rect 510804 641922 510816 641956
rect 510850 641922 510862 641956
rect 510804 641888 510862 641922
rect 510804 641854 510816 641888
rect 510850 641854 510862 641888
rect 510804 641820 510862 641854
rect 510804 641786 510816 641820
rect 510850 641786 510862 641820
rect 510804 641752 510862 641786
rect 510804 641718 510816 641752
rect 510850 641718 510862 641752
rect 510804 641684 510862 641718
rect 510804 641650 510816 641684
rect 510850 641650 510862 641684
rect 510804 641616 510862 641650
rect 510804 641582 510816 641616
rect 510850 641582 510862 641616
rect 510804 641548 510862 641582
rect 510804 641514 510816 641548
rect 510850 641514 510862 641548
rect 510804 641480 510862 641514
rect 510804 641446 510816 641480
rect 510850 641446 510862 641480
rect 510804 641405 510862 641446
rect 511262 642364 511320 642405
rect 511262 642330 511274 642364
rect 511308 642330 511320 642364
rect 511262 642296 511320 642330
rect 511262 642262 511274 642296
rect 511308 642262 511320 642296
rect 511262 642228 511320 642262
rect 511262 642194 511274 642228
rect 511308 642194 511320 642228
rect 511262 642160 511320 642194
rect 511262 642126 511274 642160
rect 511308 642126 511320 642160
rect 511262 642092 511320 642126
rect 511262 642058 511274 642092
rect 511308 642058 511320 642092
rect 511262 642024 511320 642058
rect 511262 641990 511274 642024
rect 511308 641990 511320 642024
rect 511262 641956 511320 641990
rect 511262 641922 511274 641956
rect 511308 641922 511320 641956
rect 511262 641888 511320 641922
rect 511262 641854 511274 641888
rect 511308 641854 511320 641888
rect 511262 641820 511320 641854
rect 511262 641786 511274 641820
rect 511308 641786 511320 641820
rect 511262 641752 511320 641786
rect 511262 641718 511274 641752
rect 511308 641718 511320 641752
rect 511262 641684 511320 641718
rect 511262 641650 511274 641684
rect 511308 641650 511320 641684
rect 511262 641616 511320 641650
rect 511262 641582 511274 641616
rect 511308 641582 511320 641616
rect 511262 641548 511320 641582
rect 511262 641514 511274 641548
rect 511308 641514 511320 641548
rect 511262 641480 511320 641514
rect 511262 641446 511274 641480
rect 511308 641446 511320 641480
rect 511262 641405 511320 641446
rect 511720 642364 511778 642405
rect 511720 642330 511732 642364
rect 511766 642330 511778 642364
rect 511720 642296 511778 642330
rect 511720 642262 511732 642296
rect 511766 642262 511778 642296
rect 511720 642228 511778 642262
rect 511720 642194 511732 642228
rect 511766 642194 511778 642228
rect 511720 642160 511778 642194
rect 511720 642126 511732 642160
rect 511766 642126 511778 642160
rect 511720 642092 511778 642126
rect 511720 642058 511732 642092
rect 511766 642058 511778 642092
rect 511720 642024 511778 642058
rect 511720 641990 511732 642024
rect 511766 641990 511778 642024
rect 511720 641956 511778 641990
rect 511720 641922 511732 641956
rect 511766 641922 511778 641956
rect 511720 641888 511778 641922
rect 511720 641854 511732 641888
rect 511766 641854 511778 641888
rect 511720 641820 511778 641854
rect 511720 641786 511732 641820
rect 511766 641786 511778 641820
rect 511720 641752 511778 641786
rect 511720 641718 511732 641752
rect 511766 641718 511778 641752
rect 511720 641684 511778 641718
rect 511720 641650 511732 641684
rect 511766 641650 511778 641684
rect 511720 641616 511778 641650
rect 511720 641582 511732 641616
rect 511766 641582 511778 641616
rect 511720 641548 511778 641582
rect 511720 641514 511732 641548
rect 511766 641514 511778 641548
rect 511720 641480 511778 641514
rect 511720 641446 511732 641480
rect 511766 641446 511778 641480
rect 511720 641405 511778 641446
rect 512178 642364 512236 642405
rect 512178 642330 512190 642364
rect 512224 642330 512236 642364
rect 512178 642296 512236 642330
rect 512178 642262 512190 642296
rect 512224 642262 512236 642296
rect 512178 642228 512236 642262
rect 512178 642194 512190 642228
rect 512224 642194 512236 642228
rect 512178 642160 512236 642194
rect 512178 642126 512190 642160
rect 512224 642126 512236 642160
rect 512178 642092 512236 642126
rect 512178 642058 512190 642092
rect 512224 642058 512236 642092
rect 512178 642024 512236 642058
rect 512178 641990 512190 642024
rect 512224 641990 512236 642024
rect 512178 641956 512236 641990
rect 512178 641922 512190 641956
rect 512224 641922 512236 641956
rect 512178 641888 512236 641922
rect 512178 641854 512190 641888
rect 512224 641854 512236 641888
rect 512178 641820 512236 641854
rect 512178 641786 512190 641820
rect 512224 641786 512236 641820
rect 512178 641752 512236 641786
rect 512178 641718 512190 641752
rect 512224 641718 512236 641752
rect 512178 641684 512236 641718
rect 512178 641650 512190 641684
rect 512224 641650 512236 641684
rect 512178 641616 512236 641650
rect 512178 641582 512190 641616
rect 512224 641582 512236 641616
rect 512178 641548 512236 641582
rect 512178 641514 512190 641548
rect 512224 641514 512236 641548
rect 512178 641480 512236 641514
rect 512178 641446 512190 641480
rect 512224 641446 512236 641480
rect 512178 641405 512236 641446
rect 512636 642364 512694 642405
rect 512636 642330 512648 642364
rect 512682 642330 512694 642364
rect 512636 642296 512694 642330
rect 512636 642262 512648 642296
rect 512682 642262 512694 642296
rect 512636 642228 512694 642262
rect 512636 642194 512648 642228
rect 512682 642194 512694 642228
rect 512636 642160 512694 642194
rect 512636 642126 512648 642160
rect 512682 642126 512694 642160
rect 512636 642092 512694 642126
rect 512636 642058 512648 642092
rect 512682 642058 512694 642092
rect 512636 642024 512694 642058
rect 512636 641990 512648 642024
rect 512682 641990 512694 642024
rect 512636 641956 512694 641990
rect 512636 641922 512648 641956
rect 512682 641922 512694 641956
rect 512636 641888 512694 641922
rect 512636 641854 512648 641888
rect 512682 641854 512694 641888
rect 512636 641820 512694 641854
rect 512636 641786 512648 641820
rect 512682 641786 512694 641820
rect 512636 641752 512694 641786
rect 512636 641718 512648 641752
rect 512682 641718 512694 641752
rect 512636 641684 512694 641718
rect 512636 641650 512648 641684
rect 512682 641650 512694 641684
rect 512636 641616 512694 641650
rect 512636 641582 512648 641616
rect 512682 641582 512694 641616
rect 512636 641548 512694 641582
rect 512636 641514 512648 641548
rect 512682 641514 512694 641548
rect 512636 641480 512694 641514
rect 512636 641446 512648 641480
rect 512682 641446 512694 641480
rect 512636 641405 512694 641446
rect 513094 642364 513152 642405
rect 513094 642330 513106 642364
rect 513140 642330 513152 642364
rect 513094 642296 513152 642330
rect 513094 642262 513106 642296
rect 513140 642262 513152 642296
rect 513094 642228 513152 642262
rect 513094 642194 513106 642228
rect 513140 642194 513152 642228
rect 513094 642160 513152 642194
rect 513094 642126 513106 642160
rect 513140 642126 513152 642160
rect 513094 642092 513152 642126
rect 513094 642058 513106 642092
rect 513140 642058 513152 642092
rect 513094 642024 513152 642058
rect 513094 641990 513106 642024
rect 513140 641990 513152 642024
rect 513094 641956 513152 641990
rect 513094 641922 513106 641956
rect 513140 641922 513152 641956
rect 513094 641888 513152 641922
rect 513094 641854 513106 641888
rect 513140 641854 513152 641888
rect 513094 641820 513152 641854
rect 513094 641786 513106 641820
rect 513140 641786 513152 641820
rect 513094 641752 513152 641786
rect 513094 641718 513106 641752
rect 513140 641718 513152 641752
rect 513094 641684 513152 641718
rect 513094 641650 513106 641684
rect 513140 641650 513152 641684
rect 513094 641616 513152 641650
rect 513094 641582 513106 641616
rect 513140 641582 513152 641616
rect 513094 641548 513152 641582
rect 513094 641514 513106 641548
rect 513140 641514 513152 641548
rect 513094 641480 513152 641514
rect 513094 641446 513106 641480
rect 513140 641446 513152 641480
rect 513094 641405 513152 641446
rect 513552 642364 513610 642405
rect 513552 642330 513564 642364
rect 513598 642330 513610 642364
rect 513552 642296 513610 642330
rect 513552 642262 513564 642296
rect 513598 642262 513610 642296
rect 513552 642228 513610 642262
rect 513552 642194 513564 642228
rect 513598 642194 513610 642228
rect 513552 642160 513610 642194
rect 513552 642126 513564 642160
rect 513598 642126 513610 642160
rect 513552 642092 513610 642126
rect 513552 642058 513564 642092
rect 513598 642058 513610 642092
rect 513552 642024 513610 642058
rect 513552 641990 513564 642024
rect 513598 641990 513610 642024
rect 513552 641956 513610 641990
rect 513552 641922 513564 641956
rect 513598 641922 513610 641956
rect 513552 641888 513610 641922
rect 513552 641854 513564 641888
rect 513598 641854 513610 641888
rect 513552 641820 513610 641854
rect 513552 641786 513564 641820
rect 513598 641786 513610 641820
rect 513552 641752 513610 641786
rect 513552 641718 513564 641752
rect 513598 641718 513610 641752
rect 513552 641684 513610 641718
rect 513552 641650 513564 641684
rect 513598 641650 513610 641684
rect 513552 641616 513610 641650
rect 513552 641582 513564 641616
rect 513598 641582 513610 641616
rect 513552 641548 513610 641582
rect 513552 641514 513564 641548
rect 513598 641514 513610 641548
rect 513552 641480 513610 641514
rect 513552 641446 513564 641480
rect 513598 641446 513610 641480
rect 513552 641405 513610 641446
rect 514010 642364 514068 642405
rect 514010 642330 514022 642364
rect 514056 642330 514068 642364
rect 514010 642296 514068 642330
rect 514010 642262 514022 642296
rect 514056 642262 514068 642296
rect 514010 642228 514068 642262
rect 514010 642194 514022 642228
rect 514056 642194 514068 642228
rect 514010 642160 514068 642194
rect 514010 642126 514022 642160
rect 514056 642126 514068 642160
rect 514010 642092 514068 642126
rect 514010 642058 514022 642092
rect 514056 642058 514068 642092
rect 514010 642024 514068 642058
rect 514010 641990 514022 642024
rect 514056 641990 514068 642024
rect 514010 641956 514068 641990
rect 514010 641922 514022 641956
rect 514056 641922 514068 641956
rect 514010 641888 514068 641922
rect 514010 641854 514022 641888
rect 514056 641854 514068 641888
rect 514010 641820 514068 641854
rect 514010 641786 514022 641820
rect 514056 641786 514068 641820
rect 514010 641752 514068 641786
rect 514010 641718 514022 641752
rect 514056 641718 514068 641752
rect 514010 641684 514068 641718
rect 514010 641650 514022 641684
rect 514056 641650 514068 641684
rect 514010 641616 514068 641650
rect 514010 641582 514022 641616
rect 514056 641582 514068 641616
rect 514010 641548 514068 641582
rect 514010 641514 514022 641548
rect 514056 641514 514068 641548
rect 514010 641480 514068 641514
rect 514010 641446 514022 641480
rect 514056 641446 514068 641480
rect 514010 641405 514068 641446
rect 514468 642364 514526 642405
rect 514468 642330 514480 642364
rect 514514 642330 514526 642364
rect 514468 642296 514526 642330
rect 514468 642262 514480 642296
rect 514514 642262 514526 642296
rect 514468 642228 514526 642262
rect 514468 642194 514480 642228
rect 514514 642194 514526 642228
rect 514468 642160 514526 642194
rect 514468 642126 514480 642160
rect 514514 642126 514526 642160
rect 514468 642092 514526 642126
rect 514468 642058 514480 642092
rect 514514 642058 514526 642092
rect 514468 642024 514526 642058
rect 514468 641990 514480 642024
rect 514514 641990 514526 642024
rect 514468 641956 514526 641990
rect 514468 641922 514480 641956
rect 514514 641922 514526 641956
rect 514468 641888 514526 641922
rect 514468 641854 514480 641888
rect 514514 641854 514526 641888
rect 514468 641820 514526 641854
rect 514468 641786 514480 641820
rect 514514 641786 514526 641820
rect 514468 641752 514526 641786
rect 514468 641718 514480 641752
rect 514514 641718 514526 641752
rect 514468 641684 514526 641718
rect 514468 641650 514480 641684
rect 514514 641650 514526 641684
rect 514468 641616 514526 641650
rect 514468 641582 514480 641616
rect 514514 641582 514526 641616
rect 514468 641548 514526 641582
rect 514468 641514 514480 641548
rect 514514 641514 514526 641548
rect 514468 641480 514526 641514
rect 514468 641446 514480 641480
rect 514514 641446 514526 641480
rect 514468 641405 514526 641446
rect 514926 642364 514984 642405
rect 514926 642330 514938 642364
rect 514972 642330 514984 642364
rect 514926 642296 514984 642330
rect 514926 642262 514938 642296
rect 514972 642262 514984 642296
rect 514926 642228 514984 642262
rect 514926 642194 514938 642228
rect 514972 642194 514984 642228
rect 514926 642160 514984 642194
rect 514926 642126 514938 642160
rect 514972 642126 514984 642160
rect 514926 642092 514984 642126
rect 514926 642058 514938 642092
rect 514972 642058 514984 642092
rect 514926 642024 514984 642058
rect 514926 641990 514938 642024
rect 514972 641990 514984 642024
rect 514926 641956 514984 641990
rect 514926 641922 514938 641956
rect 514972 641922 514984 641956
rect 514926 641888 514984 641922
rect 514926 641854 514938 641888
rect 514972 641854 514984 641888
rect 514926 641820 514984 641854
rect 514926 641786 514938 641820
rect 514972 641786 514984 641820
rect 514926 641752 514984 641786
rect 514926 641718 514938 641752
rect 514972 641718 514984 641752
rect 514926 641684 514984 641718
rect 514926 641650 514938 641684
rect 514972 641650 514984 641684
rect 514926 641616 514984 641650
rect 514926 641582 514938 641616
rect 514972 641582 514984 641616
rect 514926 641548 514984 641582
rect 514926 641514 514938 641548
rect 514972 641514 514984 641548
rect 514926 641480 514984 641514
rect 514926 641446 514938 641480
rect 514972 641446 514984 641480
rect 514926 641405 514984 641446
rect 515384 642364 515442 642405
rect 515384 642330 515396 642364
rect 515430 642330 515442 642364
rect 515384 642296 515442 642330
rect 515384 642262 515396 642296
rect 515430 642262 515442 642296
rect 515384 642228 515442 642262
rect 515384 642194 515396 642228
rect 515430 642194 515442 642228
rect 515384 642160 515442 642194
rect 515384 642126 515396 642160
rect 515430 642126 515442 642160
rect 515384 642092 515442 642126
rect 515384 642058 515396 642092
rect 515430 642058 515442 642092
rect 515384 642024 515442 642058
rect 515384 641990 515396 642024
rect 515430 641990 515442 642024
rect 515384 641956 515442 641990
rect 515384 641922 515396 641956
rect 515430 641922 515442 641956
rect 515384 641888 515442 641922
rect 515384 641854 515396 641888
rect 515430 641854 515442 641888
rect 515384 641820 515442 641854
rect 515384 641786 515396 641820
rect 515430 641786 515442 641820
rect 515384 641752 515442 641786
rect 515384 641718 515396 641752
rect 515430 641718 515442 641752
rect 515384 641684 515442 641718
rect 515384 641650 515396 641684
rect 515430 641650 515442 641684
rect 515384 641616 515442 641650
rect 515384 641582 515396 641616
rect 515430 641582 515442 641616
rect 515384 641548 515442 641582
rect 515384 641514 515396 641548
rect 515430 641514 515442 641548
rect 515384 641480 515442 641514
rect 515384 641446 515396 641480
rect 515430 641446 515442 641480
rect 515384 641405 515442 641446
rect 508056 641202 508114 641243
rect 508056 641168 508068 641202
rect 508102 641168 508114 641202
rect 508056 641134 508114 641168
rect 508056 641100 508068 641134
rect 508102 641100 508114 641134
rect 508056 641066 508114 641100
rect 508056 641032 508068 641066
rect 508102 641032 508114 641066
rect 508056 640998 508114 641032
rect 508056 640964 508068 640998
rect 508102 640964 508114 640998
rect 508056 640930 508114 640964
rect 508056 640896 508068 640930
rect 508102 640896 508114 640930
rect 508056 640862 508114 640896
rect 508056 640828 508068 640862
rect 508102 640828 508114 640862
rect 508056 640794 508114 640828
rect 508056 640760 508068 640794
rect 508102 640760 508114 640794
rect 508056 640726 508114 640760
rect 508056 640692 508068 640726
rect 508102 640692 508114 640726
rect 508056 640658 508114 640692
rect 508056 640624 508068 640658
rect 508102 640624 508114 640658
rect 508056 640590 508114 640624
rect 508056 640556 508068 640590
rect 508102 640556 508114 640590
rect 508056 640522 508114 640556
rect 508056 640488 508068 640522
rect 508102 640488 508114 640522
rect 508056 640454 508114 640488
rect 508056 640420 508068 640454
rect 508102 640420 508114 640454
rect 508056 640386 508114 640420
rect 508056 640352 508068 640386
rect 508102 640352 508114 640386
rect 508056 640318 508114 640352
rect 508056 640284 508068 640318
rect 508102 640284 508114 640318
rect 508056 640243 508114 640284
rect 508514 641202 508572 641243
rect 508514 641168 508526 641202
rect 508560 641168 508572 641202
rect 508514 641134 508572 641168
rect 508514 641100 508526 641134
rect 508560 641100 508572 641134
rect 508514 641066 508572 641100
rect 508514 641032 508526 641066
rect 508560 641032 508572 641066
rect 508514 640998 508572 641032
rect 508514 640964 508526 640998
rect 508560 640964 508572 640998
rect 508514 640930 508572 640964
rect 508514 640896 508526 640930
rect 508560 640896 508572 640930
rect 508514 640862 508572 640896
rect 508514 640828 508526 640862
rect 508560 640828 508572 640862
rect 508514 640794 508572 640828
rect 508514 640760 508526 640794
rect 508560 640760 508572 640794
rect 508514 640726 508572 640760
rect 508514 640692 508526 640726
rect 508560 640692 508572 640726
rect 508514 640658 508572 640692
rect 508514 640624 508526 640658
rect 508560 640624 508572 640658
rect 508514 640590 508572 640624
rect 508514 640556 508526 640590
rect 508560 640556 508572 640590
rect 508514 640522 508572 640556
rect 508514 640488 508526 640522
rect 508560 640488 508572 640522
rect 508514 640454 508572 640488
rect 508514 640420 508526 640454
rect 508560 640420 508572 640454
rect 508514 640386 508572 640420
rect 508514 640352 508526 640386
rect 508560 640352 508572 640386
rect 508514 640318 508572 640352
rect 508514 640284 508526 640318
rect 508560 640284 508572 640318
rect 508514 640243 508572 640284
rect 508972 641202 509030 641243
rect 508972 641168 508984 641202
rect 509018 641168 509030 641202
rect 508972 641134 509030 641168
rect 508972 641100 508984 641134
rect 509018 641100 509030 641134
rect 508972 641066 509030 641100
rect 508972 641032 508984 641066
rect 509018 641032 509030 641066
rect 508972 640998 509030 641032
rect 508972 640964 508984 640998
rect 509018 640964 509030 640998
rect 508972 640930 509030 640964
rect 508972 640896 508984 640930
rect 509018 640896 509030 640930
rect 508972 640862 509030 640896
rect 508972 640828 508984 640862
rect 509018 640828 509030 640862
rect 508972 640794 509030 640828
rect 508972 640760 508984 640794
rect 509018 640760 509030 640794
rect 508972 640726 509030 640760
rect 508972 640692 508984 640726
rect 509018 640692 509030 640726
rect 508972 640658 509030 640692
rect 508972 640624 508984 640658
rect 509018 640624 509030 640658
rect 508972 640590 509030 640624
rect 508972 640556 508984 640590
rect 509018 640556 509030 640590
rect 508972 640522 509030 640556
rect 508972 640488 508984 640522
rect 509018 640488 509030 640522
rect 508972 640454 509030 640488
rect 508972 640420 508984 640454
rect 509018 640420 509030 640454
rect 508972 640386 509030 640420
rect 508972 640352 508984 640386
rect 509018 640352 509030 640386
rect 508972 640318 509030 640352
rect 508972 640284 508984 640318
rect 509018 640284 509030 640318
rect 508972 640243 509030 640284
rect 509430 641202 509488 641243
rect 509430 641168 509442 641202
rect 509476 641168 509488 641202
rect 509430 641134 509488 641168
rect 509430 641100 509442 641134
rect 509476 641100 509488 641134
rect 509430 641066 509488 641100
rect 509430 641032 509442 641066
rect 509476 641032 509488 641066
rect 509430 640998 509488 641032
rect 509430 640964 509442 640998
rect 509476 640964 509488 640998
rect 509430 640930 509488 640964
rect 509430 640896 509442 640930
rect 509476 640896 509488 640930
rect 509430 640862 509488 640896
rect 509430 640828 509442 640862
rect 509476 640828 509488 640862
rect 509430 640794 509488 640828
rect 509430 640760 509442 640794
rect 509476 640760 509488 640794
rect 509430 640726 509488 640760
rect 509430 640692 509442 640726
rect 509476 640692 509488 640726
rect 509430 640658 509488 640692
rect 509430 640624 509442 640658
rect 509476 640624 509488 640658
rect 509430 640590 509488 640624
rect 509430 640556 509442 640590
rect 509476 640556 509488 640590
rect 509430 640522 509488 640556
rect 509430 640488 509442 640522
rect 509476 640488 509488 640522
rect 509430 640454 509488 640488
rect 509430 640420 509442 640454
rect 509476 640420 509488 640454
rect 509430 640386 509488 640420
rect 509430 640352 509442 640386
rect 509476 640352 509488 640386
rect 509430 640318 509488 640352
rect 509430 640284 509442 640318
rect 509476 640284 509488 640318
rect 509430 640243 509488 640284
rect 509888 641202 509946 641243
rect 509888 641168 509900 641202
rect 509934 641168 509946 641202
rect 509888 641134 509946 641168
rect 509888 641100 509900 641134
rect 509934 641100 509946 641134
rect 509888 641066 509946 641100
rect 509888 641032 509900 641066
rect 509934 641032 509946 641066
rect 509888 640998 509946 641032
rect 509888 640964 509900 640998
rect 509934 640964 509946 640998
rect 509888 640930 509946 640964
rect 509888 640896 509900 640930
rect 509934 640896 509946 640930
rect 509888 640862 509946 640896
rect 509888 640828 509900 640862
rect 509934 640828 509946 640862
rect 509888 640794 509946 640828
rect 509888 640760 509900 640794
rect 509934 640760 509946 640794
rect 509888 640726 509946 640760
rect 509888 640692 509900 640726
rect 509934 640692 509946 640726
rect 509888 640658 509946 640692
rect 509888 640624 509900 640658
rect 509934 640624 509946 640658
rect 509888 640590 509946 640624
rect 509888 640556 509900 640590
rect 509934 640556 509946 640590
rect 509888 640522 509946 640556
rect 509888 640488 509900 640522
rect 509934 640488 509946 640522
rect 509888 640454 509946 640488
rect 509888 640420 509900 640454
rect 509934 640420 509946 640454
rect 509888 640386 509946 640420
rect 509888 640352 509900 640386
rect 509934 640352 509946 640386
rect 509888 640318 509946 640352
rect 509888 640284 509900 640318
rect 509934 640284 509946 640318
rect 509888 640243 509946 640284
rect 510346 641202 510404 641243
rect 510346 641168 510358 641202
rect 510392 641168 510404 641202
rect 510346 641134 510404 641168
rect 510346 641100 510358 641134
rect 510392 641100 510404 641134
rect 510346 641066 510404 641100
rect 510346 641032 510358 641066
rect 510392 641032 510404 641066
rect 510346 640998 510404 641032
rect 510346 640964 510358 640998
rect 510392 640964 510404 640998
rect 510346 640930 510404 640964
rect 510346 640896 510358 640930
rect 510392 640896 510404 640930
rect 510346 640862 510404 640896
rect 510346 640828 510358 640862
rect 510392 640828 510404 640862
rect 510346 640794 510404 640828
rect 510346 640760 510358 640794
rect 510392 640760 510404 640794
rect 510346 640726 510404 640760
rect 510346 640692 510358 640726
rect 510392 640692 510404 640726
rect 510346 640658 510404 640692
rect 510346 640624 510358 640658
rect 510392 640624 510404 640658
rect 510346 640590 510404 640624
rect 510346 640556 510358 640590
rect 510392 640556 510404 640590
rect 510346 640522 510404 640556
rect 510346 640488 510358 640522
rect 510392 640488 510404 640522
rect 510346 640454 510404 640488
rect 510346 640420 510358 640454
rect 510392 640420 510404 640454
rect 510346 640386 510404 640420
rect 510346 640352 510358 640386
rect 510392 640352 510404 640386
rect 510346 640318 510404 640352
rect 510346 640284 510358 640318
rect 510392 640284 510404 640318
rect 510346 640243 510404 640284
rect 510804 641202 510862 641243
rect 510804 641168 510816 641202
rect 510850 641168 510862 641202
rect 510804 641134 510862 641168
rect 510804 641100 510816 641134
rect 510850 641100 510862 641134
rect 510804 641066 510862 641100
rect 510804 641032 510816 641066
rect 510850 641032 510862 641066
rect 510804 640998 510862 641032
rect 510804 640964 510816 640998
rect 510850 640964 510862 640998
rect 510804 640930 510862 640964
rect 510804 640896 510816 640930
rect 510850 640896 510862 640930
rect 510804 640862 510862 640896
rect 510804 640828 510816 640862
rect 510850 640828 510862 640862
rect 510804 640794 510862 640828
rect 510804 640760 510816 640794
rect 510850 640760 510862 640794
rect 510804 640726 510862 640760
rect 510804 640692 510816 640726
rect 510850 640692 510862 640726
rect 510804 640658 510862 640692
rect 510804 640624 510816 640658
rect 510850 640624 510862 640658
rect 510804 640590 510862 640624
rect 510804 640556 510816 640590
rect 510850 640556 510862 640590
rect 510804 640522 510862 640556
rect 510804 640488 510816 640522
rect 510850 640488 510862 640522
rect 510804 640454 510862 640488
rect 510804 640420 510816 640454
rect 510850 640420 510862 640454
rect 510804 640386 510862 640420
rect 510804 640352 510816 640386
rect 510850 640352 510862 640386
rect 510804 640318 510862 640352
rect 510804 640284 510816 640318
rect 510850 640284 510862 640318
rect 510804 640243 510862 640284
rect 511262 641202 511320 641243
rect 511262 641168 511274 641202
rect 511308 641168 511320 641202
rect 511262 641134 511320 641168
rect 511262 641100 511274 641134
rect 511308 641100 511320 641134
rect 511262 641066 511320 641100
rect 511262 641032 511274 641066
rect 511308 641032 511320 641066
rect 511262 640998 511320 641032
rect 511262 640964 511274 640998
rect 511308 640964 511320 640998
rect 511262 640930 511320 640964
rect 511262 640896 511274 640930
rect 511308 640896 511320 640930
rect 511262 640862 511320 640896
rect 511262 640828 511274 640862
rect 511308 640828 511320 640862
rect 511262 640794 511320 640828
rect 511262 640760 511274 640794
rect 511308 640760 511320 640794
rect 511262 640726 511320 640760
rect 511262 640692 511274 640726
rect 511308 640692 511320 640726
rect 511262 640658 511320 640692
rect 511262 640624 511274 640658
rect 511308 640624 511320 640658
rect 511262 640590 511320 640624
rect 511262 640556 511274 640590
rect 511308 640556 511320 640590
rect 511262 640522 511320 640556
rect 511262 640488 511274 640522
rect 511308 640488 511320 640522
rect 511262 640454 511320 640488
rect 511262 640420 511274 640454
rect 511308 640420 511320 640454
rect 511262 640386 511320 640420
rect 511262 640352 511274 640386
rect 511308 640352 511320 640386
rect 511262 640318 511320 640352
rect 511262 640284 511274 640318
rect 511308 640284 511320 640318
rect 511262 640243 511320 640284
rect 511720 641202 511778 641243
rect 511720 641168 511732 641202
rect 511766 641168 511778 641202
rect 511720 641134 511778 641168
rect 511720 641100 511732 641134
rect 511766 641100 511778 641134
rect 511720 641066 511778 641100
rect 511720 641032 511732 641066
rect 511766 641032 511778 641066
rect 511720 640998 511778 641032
rect 511720 640964 511732 640998
rect 511766 640964 511778 640998
rect 511720 640930 511778 640964
rect 511720 640896 511732 640930
rect 511766 640896 511778 640930
rect 511720 640862 511778 640896
rect 511720 640828 511732 640862
rect 511766 640828 511778 640862
rect 511720 640794 511778 640828
rect 511720 640760 511732 640794
rect 511766 640760 511778 640794
rect 511720 640726 511778 640760
rect 511720 640692 511732 640726
rect 511766 640692 511778 640726
rect 511720 640658 511778 640692
rect 511720 640624 511732 640658
rect 511766 640624 511778 640658
rect 511720 640590 511778 640624
rect 511720 640556 511732 640590
rect 511766 640556 511778 640590
rect 511720 640522 511778 640556
rect 511720 640488 511732 640522
rect 511766 640488 511778 640522
rect 511720 640454 511778 640488
rect 511720 640420 511732 640454
rect 511766 640420 511778 640454
rect 511720 640386 511778 640420
rect 511720 640352 511732 640386
rect 511766 640352 511778 640386
rect 511720 640318 511778 640352
rect 511720 640284 511732 640318
rect 511766 640284 511778 640318
rect 511720 640243 511778 640284
rect 512178 641202 512236 641243
rect 512178 641168 512190 641202
rect 512224 641168 512236 641202
rect 512178 641134 512236 641168
rect 512178 641100 512190 641134
rect 512224 641100 512236 641134
rect 512178 641066 512236 641100
rect 512178 641032 512190 641066
rect 512224 641032 512236 641066
rect 512178 640998 512236 641032
rect 512178 640964 512190 640998
rect 512224 640964 512236 640998
rect 512178 640930 512236 640964
rect 512178 640896 512190 640930
rect 512224 640896 512236 640930
rect 512178 640862 512236 640896
rect 512178 640828 512190 640862
rect 512224 640828 512236 640862
rect 512178 640794 512236 640828
rect 512178 640760 512190 640794
rect 512224 640760 512236 640794
rect 512178 640726 512236 640760
rect 512178 640692 512190 640726
rect 512224 640692 512236 640726
rect 512178 640658 512236 640692
rect 512178 640624 512190 640658
rect 512224 640624 512236 640658
rect 512178 640590 512236 640624
rect 512178 640556 512190 640590
rect 512224 640556 512236 640590
rect 512178 640522 512236 640556
rect 512178 640488 512190 640522
rect 512224 640488 512236 640522
rect 512178 640454 512236 640488
rect 512178 640420 512190 640454
rect 512224 640420 512236 640454
rect 512178 640386 512236 640420
rect 512178 640352 512190 640386
rect 512224 640352 512236 640386
rect 512178 640318 512236 640352
rect 512178 640284 512190 640318
rect 512224 640284 512236 640318
rect 512178 640243 512236 640284
rect 512636 641202 512694 641243
rect 512636 641168 512648 641202
rect 512682 641168 512694 641202
rect 512636 641134 512694 641168
rect 512636 641100 512648 641134
rect 512682 641100 512694 641134
rect 512636 641066 512694 641100
rect 512636 641032 512648 641066
rect 512682 641032 512694 641066
rect 512636 640998 512694 641032
rect 512636 640964 512648 640998
rect 512682 640964 512694 640998
rect 512636 640930 512694 640964
rect 512636 640896 512648 640930
rect 512682 640896 512694 640930
rect 512636 640862 512694 640896
rect 512636 640828 512648 640862
rect 512682 640828 512694 640862
rect 512636 640794 512694 640828
rect 512636 640760 512648 640794
rect 512682 640760 512694 640794
rect 512636 640726 512694 640760
rect 512636 640692 512648 640726
rect 512682 640692 512694 640726
rect 512636 640658 512694 640692
rect 512636 640624 512648 640658
rect 512682 640624 512694 640658
rect 512636 640590 512694 640624
rect 512636 640556 512648 640590
rect 512682 640556 512694 640590
rect 512636 640522 512694 640556
rect 512636 640488 512648 640522
rect 512682 640488 512694 640522
rect 512636 640454 512694 640488
rect 512636 640420 512648 640454
rect 512682 640420 512694 640454
rect 512636 640386 512694 640420
rect 512636 640352 512648 640386
rect 512682 640352 512694 640386
rect 512636 640318 512694 640352
rect 512636 640284 512648 640318
rect 512682 640284 512694 640318
rect 512636 640243 512694 640284
rect 513094 641202 513152 641243
rect 513094 641168 513106 641202
rect 513140 641168 513152 641202
rect 513094 641134 513152 641168
rect 513094 641100 513106 641134
rect 513140 641100 513152 641134
rect 513094 641066 513152 641100
rect 513094 641032 513106 641066
rect 513140 641032 513152 641066
rect 513094 640998 513152 641032
rect 513094 640964 513106 640998
rect 513140 640964 513152 640998
rect 513094 640930 513152 640964
rect 513094 640896 513106 640930
rect 513140 640896 513152 640930
rect 513094 640862 513152 640896
rect 513094 640828 513106 640862
rect 513140 640828 513152 640862
rect 513094 640794 513152 640828
rect 513094 640760 513106 640794
rect 513140 640760 513152 640794
rect 513094 640726 513152 640760
rect 513094 640692 513106 640726
rect 513140 640692 513152 640726
rect 513094 640658 513152 640692
rect 513094 640624 513106 640658
rect 513140 640624 513152 640658
rect 513094 640590 513152 640624
rect 513094 640556 513106 640590
rect 513140 640556 513152 640590
rect 513094 640522 513152 640556
rect 513094 640488 513106 640522
rect 513140 640488 513152 640522
rect 513094 640454 513152 640488
rect 513094 640420 513106 640454
rect 513140 640420 513152 640454
rect 513094 640386 513152 640420
rect 513094 640352 513106 640386
rect 513140 640352 513152 640386
rect 513094 640318 513152 640352
rect 513094 640284 513106 640318
rect 513140 640284 513152 640318
rect 513094 640243 513152 640284
rect 513552 641202 513610 641243
rect 513552 641168 513564 641202
rect 513598 641168 513610 641202
rect 513552 641134 513610 641168
rect 513552 641100 513564 641134
rect 513598 641100 513610 641134
rect 513552 641066 513610 641100
rect 513552 641032 513564 641066
rect 513598 641032 513610 641066
rect 513552 640998 513610 641032
rect 513552 640964 513564 640998
rect 513598 640964 513610 640998
rect 513552 640930 513610 640964
rect 513552 640896 513564 640930
rect 513598 640896 513610 640930
rect 513552 640862 513610 640896
rect 513552 640828 513564 640862
rect 513598 640828 513610 640862
rect 513552 640794 513610 640828
rect 513552 640760 513564 640794
rect 513598 640760 513610 640794
rect 513552 640726 513610 640760
rect 513552 640692 513564 640726
rect 513598 640692 513610 640726
rect 513552 640658 513610 640692
rect 513552 640624 513564 640658
rect 513598 640624 513610 640658
rect 513552 640590 513610 640624
rect 513552 640556 513564 640590
rect 513598 640556 513610 640590
rect 513552 640522 513610 640556
rect 513552 640488 513564 640522
rect 513598 640488 513610 640522
rect 513552 640454 513610 640488
rect 513552 640420 513564 640454
rect 513598 640420 513610 640454
rect 513552 640386 513610 640420
rect 513552 640352 513564 640386
rect 513598 640352 513610 640386
rect 513552 640318 513610 640352
rect 513552 640284 513564 640318
rect 513598 640284 513610 640318
rect 513552 640243 513610 640284
rect 514010 641202 514068 641243
rect 514010 641168 514022 641202
rect 514056 641168 514068 641202
rect 514010 641134 514068 641168
rect 514010 641100 514022 641134
rect 514056 641100 514068 641134
rect 514010 641066 514068 641100
rect 514010 641032 514022 641066
rect 514056 641032 514068 641066
rect 514010 640998 514068 641032
rect 514010 640964 514022 640998
rect 514056 640964 514068 640998
rect 514010 640930 514068 640964
rect 514010 640896 514022 640930
rect 514056 640896 514068 640930
rect 514010 640862 514068 640896
rect 514010 640828 514022 640862
rect 514056 640828 514068 640862
rect 514010 640794 514068 640828
rect 514010 640760 514022 640794
rect 514056 640760 514068 640794
rect 514010 640726 514068 640760
rect 514010 640692 514022 640726
rect 514056 640692 514068 640726
rect 514010 640658 514068 640692
rect 514010 640624 514022 640658
rect 514056 640624 514068 640658
rect 514010 640590 514068 640624
rect 514010 640556 514022 640590
rect 514056 640556 514068 640590
rect 514010 640522 514068 640556
rect 514010 640488 514022 640522
rect 514056 640488 514068 640522
rect 514010 640454 514068 640488
rect 514010 640420 514022 640454
rect 514056 640420 514068 640454
rect 514010 640386 514068 640420
rect 514010 640352 514022 640386
rect 514056 640352 514068 640386
rect 514010 640318 514068 640352
rect 514010 640284 514022 640318
rect 514056 640284 514068 640318
rect 514010 640243 514068 640284
rect 514468 641202 514526 641243
rect 514468 641168 514480 641202
rect 514514 641168 514526 641202
rect 514468 641134 514526 641168
rect 514468 641100 514480 641134
rect 514514 641100 514526 641134
rect 514468 641066 514526 641100
rect 514468 641032 514480 641066
rect 514514 641032 514526 641066
rect 514468 640998 514526 641032
rect 514468 640964 514480 640998
rect 514514 640964 514526 640998
rect 514468 640930 514526 640964
rect 514468 640896 514480 640930
rect 514514 640896 514526 640930
rect 514468 640862 514526 640896
rect 514468 640828 514480 640862
rect 514514 640828 514526 640862
rect 514468 640794 514526 640828
rect 514468 640760 514480 640794
rect 514514 640760 514526 640794
rect 514468 640726 514526 640760
rect 514468 640692 514480 640726
rect 514514 640692 514526 640726
rect 514468 640658 514526 640692
rect 514468 640624 514480 640658
rect 514514 640624 514526 640658
rect 514468 640590 514526 640624
rect 514468 640556 514480 640590
rect 514514 640556 514526 640590
rect 514468 640522 514526 640556
rect 514468 640488 514480 640522
rect 514514 640488 514526 640522
rect 514468 640454 514526 640488
rect 514468 640420 514480 640454
rect 514514 640420 514526 640454
rect 514468 640386 514526 640420
rect 514468 640352 514480 640386
rect 514514 640352 514526 640386
rect 514468 640318 514526 640352
rect 514468 640284 514480 640318
rect 514514 640284 514526 640318
rect 514468 640243 514526 640284
rect 514926 641202 514984 641243
rect 514926 641168 514938 641202
rect 514972 641168 514984 641202
rect 514926 641134 514984 641168
rect 514926 641100 514938 641134
rect 514972 641100 514984 641134
rect 514926 641066 514984 641100
rect 514926 641032 514938 641066
rect 514972 641032 514984 641066
rect 514926 640998 514984 641032
rect 514926 640964 514938 640998
rect 514972 640964 514984 640998
rect 514926 640930 514984 640964
rect 514926 640896 514938 640930
rect 514972 640896 514984 640930
rect 514926 640862 514984 640896
rect 514926 640828 514938 640862
rect 514972 640828 514984 640862
rect 514926 640794 514984 640828
rect 514926 640760 514938 640794
rect 514972 640760 514984 640794
rect 514926 640726 514984 640760
rect 514926 640692 514938 640726
rect 514972 640692 514984 640726
rect 514926 640658 514984 640692
rect 514926 640624 514938 640658
rect 514972 640624 514984 640658
rect 514926 640590 514984 640624
rect 514926 640556 514938 640590
rect 514972 640556 514984 640590
rect 514926 640522 514984 640556
rect 514926 640488 514938 640522
rect 514972 640488 514984 640522
rect 514926 640454 514984 640488
rect 514926 640420 514938 640454
rect 514972 640420 514984 640454
rect 514926 640386 514984 640420
rect 514926 640352 514938 640386
rect 514972 640352 514984 640386
rect 514926 640318 514984 640352
rect 514926 640284 514938 640318
rect 514972 640284 514984 640318
rect 514926 640243 514984 640284
rect 515384 641202 515442 641243
rect 515384 641168 515396 641202
rect 515430 641168 515442 641202
rect 515384 641134 515442 641168
rect 515384 641100 515396 641134
rect 515430 641100 515442 641134
rect 515384 641066 515442 641100
rect 515384 641032 515396 641066
rect 515430 641032 515442 641066
rect 515384 640998 515442 641032
rect 515384 640964 515396 640998
rect 515430 640964 515442 640998
rect 515384 640930 515442 640964
rect 515384 640896 515396 640930
rect 515430 640896 515442 640930
rect 515384 640862 515442 640896
rect 515384 640828 515396 640862
rect 515430 640828 515442 640862
rect 515384 640794 515442 640828
rect 515384 640760 515396 640794
rect 515430 640760 515442 640794
rect 515384 640726 515442 640760
rect 515384 640692 515396 640726
rect 515430 640692 515442 640726
rect 515384 640658 515442 640692
rect 515384 640624 515396 640658
rect 515430 640624 515442 640658
rect 515384 640590 515442 640624
rect 515384 640556 515396 640590
rect 515430 640556 515442 640590
rect 515384 640522 515442 640556
rect 515384 640488 515396 640522
rect 515430 640488 515442 640522
rect 515384 640454 515442 640488
rect 515384 640420 515396 640454
rect 515430 640420 515442 640454
rect 515384 640386 515442 640420
rect 515384 640352 515396 640386
rect 515430 640352 515442 640386
rect 515384 640318 515442 640352
rect 515384 640284 515396 640318
rect 515430 640284 515442 640318
rect 515384 640243 515442 640284
rect 515760 642364 515818 642405
rect 515760 642330 515772 642364
rect 515806 642330 515818 642364
rect 515760 642296 515818 642330
rect 515760 642262 515772 642296
rect 515806 642262 515818 642296
rect 515760 642228 515818 642262
rect 515760 642194 515772 642228
rect 515806 642194 515818 642228
rect 515760 642160 515818 642194
rect 515760 642126 515772 642160
rect 515806 642126 515818 642160
rect 515760 642092 515818 642126
rect 515760 642058 515772 642092
rect 515806 642058 515818 642092
rect 515760 642024 515818 642058
rect 515760 641990 515772 642024
rect 515806 641990 515818 642024
rect 515760 641956 515818 641990
rect 515760 641922 515772 641956
rect 515806 641922 515818 641956
rect 515760 641888 515818 641922
rect 515760 641854 515772 641888
rect 515806 641854 515818 641888
rect 515760 641820 515818 641854
rect 515760 641786 515772 641820
rect 515806 641786 515818 641820
rect 515760 641752 515818 641786
rect 515760 641718 515772 641752
rect 515806 641718 515818 641752
rect 515760 641684 515818 641718
rect 515760 641650 515772 641684
rect 515806 641650 515818 641684
rect 515760 641616 515818 641650
rect 515760 641582 515772 641616
rect 515806 641582 515818 641616
rect 515760 641548 515818 641582
rect 515760 641514 515772 641548
rect 515806 641514 515818 641548
rect 515760 641480 515818 641514
rect 515760 641446 515772 641480
rect 515806 641446 515818 641480
rect 515760 641405 515818 641446
rect 516218 642364 516276 642405
rect 516218 642330 516230 642364
rect 516264 642330 516276 642364
rect 516218 642296 516276 642330
rect 516218 642262 516230 642296
rect 516264 642262 516276 642296
rect 516218 642228 516276 642262
rect 516218 642194 516230 642228
rect 516264 642194 516276 642228
rect 516218 642160 516276 642194
rect 516218 642126 516230 642160
rect 516264 642126 516276 642160
rect 516218 642092 516276 642126
rect 516218 642058 516230 642092
rect 516264 642058 516276 642092
rect 516218 642024 516276 642058
rect 516218 641990 516230 642024
rect 516264 641990 516276 642024
rect 516218 641956 516276 641990
rect 516218 641922 516230 641956
rect 516264 641922 516276 641956
rect 516218 641888 516276 641922
rect 516218 641854 516230 641888
rect 516264 641854 516276 641888
rect 516218 641820 516276 641854
rect 516218 641786 516230 641820
rect 516264 641786 516276 641820
rect 516218 641752 516276 641786
rect 516218 641718 516230 641752
rect 516264 641718 516276 641752
rect 516218 641684 516276 641718
rect 516218 641650 516230 641684
rect 516264 641650 516276 641684
rect 516218 641616 516276 641650
rect 516218 641582 516230 641616
rect 516264 641582 516276 641616
rect 516218 641548 516276 641582
rect 516218 641514 516230 641548
rect 516264 641514 516276 641548
rect 516218 641480 516276 641514
rect 516218 641446 516230 641480
rect 516264 641446 516276 641480
rect 516218 641405 516276 641446
rect 516676 642364 516734 642405
rect 516676 642330 516688 642364
rect 516722 642330 516734 642364
rect 516676 642296 516734 642330
rect 516676 642262 516688 642296
rect 516722 642262 516734 642296
rect 516676 642228 516734 642262
rect 516676 642194 516688 642228
rect 516722 642194 516734 642228
rect 516676 642160 516734 642194
rect 516676 642126 516688 642160
rect 516722 642126 516734 642160
rect 516676 642092 516734 642126
rect 516676 642058 516688 642092
rect 516722 642058 516734 642092
rect 516676 642024 516734 642058
rect 516676 641990 516688 642024
rect 516722 641990 516734 642024
rect 516676 641956 516734 641990
rect 516676 641922 516688 641956
rect 516722 641922 516734 641956
rect 516676 641888 516734 641922
rect 516676 641854 516688 641888
rect 516722 641854 516734 641888
rect 516676 641820 516734 641854
rect 516676 641786 516688 641820
rect 516722 641786 516734 641820
rect 516676 641752 516734 641786
rect 516676 641718 516688 641752
rect 516722 641718 516734 641752
rect 516676 641684 516734 641718
rect 516676 641650 516688 641684
rect 516722 641650 516734 641684
rect 516676 641616 516734 641650
rect 516676 641582 516688 641616
rect 516722 641582 516734 641616
rect 516676 641548 516734 641582
rect 516676 641514 516688 641548
rect 516722 641514 516734 641548
rect 516676 641480 516734 641514
rect 516676 641446 516688 641480
rect 516722 641446 516734 641480
rect 516676 641405 516734 641446
<< mvpdiff >>
rect 508056 645462 508114 645503
rect 508056 645428 508068 645462
rect 508102 645428 508114 645462
rect 508056 645394 508114 645428
rect 508056 645360 508068 645394
rect 508102 645360 508114 645394
rect 508056 645326 508114 645360
rect 508056 645292 508068 645326
rect 508102 645292 508114 645326
rect 508056 645258 508114 645292
rect 508056 645224 508068 645258
rect 508102 645224 508114 645258
rect 508056 645190 508114 645224
rect 508056 645156 508068 645190
rect 508102 645156 508114 645190
rect 508056 645122 508114 645156
rect 508056 645088 508068 645122
rect 508102 645088 508114 645122
rect 508056 645054 508114 645088
rect 508056 645020 508068 645054
rect 508102 645020 508114 645054
rect 508056 644986 508114 645020
rect 508056 644952 508068 644986
rect 508102 644952 508114 644986
rect 508056 644918 508114 644952
rect 508056 644884 508068 644918
rect 508102 644884 508114 644918
rect 508056 644850 508114 644884
rect 508056 644816 508068 644850
rect 508102 644816 508114 644850
rect 508056 644782 508114 644816
rect 508056 644748 508068 644782
rect 508102 644748 508114 644782
rect 508056 644714 508114 644748
rect 508056 644680 508068 644714
rect 508102 644680 508114 644714
rect 508056 644646 508114 644680
rect 508056 644612 508068 644646
rect 508102 644612 508114 644646
rect 508056 644578 508114 644612
rect 508056 644544 508068 644578
rect 508102 644544 508114 644578
rect 508056 644503 508114 644544
rect 508514 645462 508572 645503
rect 508514 645428 508526 645462
rect 508560 645428 508572 645462
rect 508514 645394 508572 645428
rect 508514 645360 508526 645394
rect 508560 645360 508572 645394
rect 508514 645326 508572 645360
rect 508514 645292 508526 645326
rect 508560 645292 508572 645326
rect 508514 645258 508572 645292
rect 508514 645224 508526 645258
rect 508560 645224 508572 645258
rect 508514 645190 508572 645224
rect 508514 645156 508526 645190
rect 508560 645156 508572 645190
rect 508514 645122 508572 645156
rect 508514 645088 508526 645122
rect 508560 645088 508572 645122
rect 508514 645054 508572 645088
rect 508514 645020 508526 645054
rect 508560 645020 508572 645054
rect 508514 644986 508572 645020
rect 508514 644952 508526 644986
rect 508560 644952 508572 644986
rect 508514 644918 508572 644952
rect 508514 644884 508526 644918
rect 508560 644884 508572 644918
rect 508514 644850 508572 644884
rect 508514 644816 508526 644850
rect 508560 644816 508572 644850
rect 508514 644782 508572 644816
rect 508514 644748 508526 644782
rect 508560 644748 508572 644782
rect 508514 644714 508572 644748
rect 508514 644680 508526 644714
rect 508560 644680 508572 644714
rect 508514 644646 508572 644680
rect 508514 644612 508526 644646
rect 508560 644612 508572 644646
rect 508514 644578 508572 644612
rect 508514 644544 508526 644578
rect 508560 644544 508572 644578
rect 508514 644503 508572 644544
rect 508972 645462 509030 645503
rect 508972 645428 508984 645462
rect 509018 645428 509030 645462
rect 508972 645394 509030 645428
rect 508972 645360 508984 645394
rect 509018 645360 509030 645394
rect 508972 645326 509030 645360
rect 508972 645292 508984 645326
rect 509018 645292 509030 645326
rect 508972 645258 509030 645292
rect 508972 645224 508984 645258
rect 509018 645224 509030 645258
rect 508972 645190 509030 645224
rect 508972 645156 508984 645190
rect 509018 645156 509030 645190
rect 508972 645122 509030 645156
rect 508972 645088 508984 645122
rect 509018 645088 509030 645122
rect 508972 645054 509030 645088
rect 508972 645020 508984 645054
rect 509018 645020 509030 645054
rect 508972 644986 509030 645020
rect 508972 644952 508984 644986
rect 509018 644952 509030 644986
rect 508972 644918 509030 644952
rect 508972 644884 508984 644918
rect 509018 644884 509030 644918
rect 508972 644850 509030 644884
rect 508972 644816 508984 644850
rect 509018 644816 509030 644850
rect 508972 644782 509030 644816
rect 508972 644748 508984 644782
rect 509018 644748 509030 644782
rect 508972 644714 509030 644748
rect 508972 644680 508984 644714
rect 509018 644680 509030 644714
rect 508972 644646 509030 644680
rect 508972 644612 508984 644646
rect 509018 644612 509030 644646
rect 508972 644578 509030 644612
rect 508972 644544 508984 644578
rect 509018 644544 509030 644578
rect 508972 644503 509030 644544
rect 509430 645462 509488 645503
rect 509430 645428 509442 645462
rect 509476 645428 509488 645462
rect 509430 645394 509488 645428
rect 509430 645360 509442 645394
rect 509476 645360 509488 645394
rect 509430 645326 509488 645360
rect 509430 645292 509442 645326
rect 509476 645292 509488 645326
rect 509430 645258 509488 645292
rect 509430 645224 509442 645258
rect 509476 645224 509488 645258
rect 509430 645190 509488 645224
rect 509430 645156 509442 645190
rect 509476 645156 509488 645190
rect 509430 645122 509488 645156
rect 509430 645088 509442 645122
rect 509476 645088 509488 645122
rect 509430 645054 509488 645088
rect 509430 645020 509442 645054
rect 509476 645020 509488 645054
rect 509430 644986 509488 645020
rect 509430 644952 509442 644986
rect 509476 644952 509488 644986
rect 509430 644918 509488 644952
rect 509430 644884 509442 644918
rect 509476 644884 509488 644918
rect 509430 644850 509488 644884
rect 509430 644816 509442 644850
rect 509476 644816 509488 644850
rect 509430 644782 509488 644816
rect 509430 644748 509442 644782
rect 509476 644748 509488 644782
rect 509430 644714 509488 644748
rect 509430 644680 509442 644714
rect 509476 644680 509488 644714
rect 509430 644646 509488 644680
rect 509430 644612 509442 644646
rect 509476 644612 509488 644646
rect 509430 644578 509488 644612
rect 509430 644544 509442 644578
rect 509476 644544 509488 644578
rect 509430 644503 509488 644544
rect 509888 645462 509946 645503
rect 509888 645428 509900 645462
rect 509934 645428 509946 645462
rect 509888 645394 509946 645428
rect 509888 645360 509900 645394
rect 509934 645360 509946 645394
rect 509888 645326 509946 645360
rect 509888 645292 509900 645326
rect 509934 645292 509946 645326
rect 509888 645258 509946 645292
rect 509888 645224 509900 645258
rect 509934 645224 509946 645258
rect 509888 645190 509946 645224
rect 509888 645156 509900 645190
rect 509934 645156 509946 645190
rect 509888 645122 509946 645156
rect 509888 645088 509900 645122
rect 509934 645088 509946 645122
rect 509888 645054 509946 645088
rect 509888 645020 509900 645054
rect 509934 645020 509946 645054
rect 509888 644986 509946 645020
rect 509888 644952 509900 644986
rect 509934 644952 509946 644986
rect 509888 644918 509946 644952
rect 509888 644884 509900 644918
rect 509934 644884 509946 644918
rect 509888 644850 509946 644884
rect 509888 644816 509900 644850
rect 509934 644816 509946 644850
rect 509888 644782 509946 644816
rect 509888 644748 509900 644782
rect 509934 644748 509946 644782
rect 509888 644714 509946 644748
rect 509888 644680 509900 644714
rect 509934 644680 509946 644714
rect 509888 644646 509946 644680
rect 509888 644612 509900 644646
rect 509934 644612 509946 644646
rect 509888 644578 509946 644612
rect 509888 644544 509900 644578
rect 509934 644544 509946 644578
rect 509888 644503 509946 644544
rect 510346 645462 510404 645503
rect 510346 645428 510358 645462
rect 510392 645428 510404 645462
rect 510346 645394 510404 645428
rect 510346 645360 510358 645394
rect 510392 645360 510404 645394
rect 510346 645326 510404 645360
rect 510346 645292 510358 645326
rect 510392 645292 510404 645326
rect 510346 645258 510404 645292
rect 510346 645224 510358 645258
rect 510392 645224 510404 645258
rect 510346 645190 510404 645224
rect 510346 645156 510358 645190
rect 510392 645156 510404 645190
rect 510346 645122 510404 645156
rect 510346 645088 510358 645122
rect 510392 645088 510404 645122
rect 510346 645054 510404 645088
rect 510346 645020 510358 645054
rect 510392 645020 510404 645054
rect 510346 644986 510404 645020
rect 510346 644952 510358 644986
rect 510392 644952 510404 644986
rect 510346 644918 510404 644952
rect 510346 644884 510358 644918
rect 510392 644884 510404 644918
rect 510346 644850 510404 644884
rect 510346 644816 510358 644850
rect 510392 644816 510404 644850
rect 510346 644782 510404 644816
rect 510346 644748 510358 644782
rect 510392 644748 510404 644782
rect 510346 644714 510404 644748
rect 510346 644680 510358 644714
rect 510392 644680 510404 644714
rect 510346 644646 510404 644680
rect 510346 644612 510358 644646
rect 510392 644612 510404 644646
rect 510346 644578 510404 644612
rect 510346 644544 510358 644578
rect 510392 644544 510404 644578
rect 510346 644503 510404 644544
rect 510804 645462 510862 645503
rect 510804 645428 510816 645462
rect 510850 645428 510862 645462
rect 510804 645394 510862 645428
rect 510804 645360 510816 645394
rect 510850 645360 510862 645394
rect 510804 645326 510862 645360
rect 510804 645292 510816 645326
rect 510850 645292 510862 645326
rect 510804 645258 510862 645292
rect 510804 645224 510816 645258
rect 510850 645224 510862 645258
rect 510804 645190 510862 645224
rect 510804 645156 510816 645190
rect 510850 645156 510862 645190
rect 510804 645122 510862 645156
rect 510804 645088 510816 645122
rect 510850 645088 510862 645122
rect 510804 645054 510862 645088
rect 510804 645020 510816 645054
rect 510850 645020 510862 645054
rect 510804 644986 510862 645020
rect 510804 644952 510816 644986
rect 510850 644952 510862 644986
rect 510804 644918 510862 644952
rect 510804 644884 510816 644918
rect 510850 644884 510862 644918
rect 510804 644850 510862 644884
rect 510804 644816 510816 644850
rect 510850 644816 510862 644850
rect 510804 644782 510862 644816
rect 510804 644748 510816 644782
rect 510850 644748 510862 644782
rect 510804 644714 510862 644748
rect 510804 644680 510816 644714
rect 510850 644680 510862 644714
rect 510804 644646 510862 644680
rect 510804 644612 510816 644646
rect 510850 644612 510862 644646
rect 510804 644578 510862 644612
rect 510804 644544 510816 644578
rect 510850 644544 510862 644578
rect 510804 644503 510862 644544
rect 511262 645462 511320 645503
rect 511262 645428 511274 645462
rect 511308 645428 511320 645462
rect 511262 645394 511320 645428
rect 511262 645360 511274 645394
rect 511308 645360 511320 645394
rect 511262 645326 511320 645360
rect 511262 645292 511274 645326
rect 511308 645292 511320 645326
rect 511262 645258 511320 645292
rect 511262 645224 511274 645258
rect 511308 645224 511320 645258
rect 511262 645190 511320 645224
rect 511262 645156 511274 645190
rect 511308 645156 511320 645190
rect 511262 645122 511320 645156
rect 511262 645088 511274 645122
rect 511308 645088 511320 645122
rect 511262 645054 511320 645088
rect 511262 645020 511274 645054
rect 511308 645020 511320 645054
rect 511262 644986 511320 645020
rect 511262 644952 511274 644986
rect 511308 644952 511320 644986
rect 511262 644918 511320 644952
rect 511262 644884 511274 644918
rect 511308 644884 511320 644918
rect 511262 644850 511320 644884
rect 511262 644816 511274 644850
rect 511308 644816 511320 644850
rect 511262 644782 511320 644816
rect 511262 644748 511274 644782
rect 511308 644748 511320 644782
rect 511262 644714 511320 644748
rect 511262 644680 511274 644714
rect 511308 644680 511320 644714
rect 511262 644646 511320 644680
rect 511262 644612 511274 644646
rect 511308 644612 511320 644646
rect 511262 644578 511320 644612
rect 511262 644544 511274 644578
rect 511308 644544 511320 644578
rect 511262 644503 511320 644544
rect 511720 645462 511778 645503
rect 511720 645428 511732 645462
rect 511766 645428 511778 645462
rect 511720 645394 511778 645428
rect 511720 645360 511732 645394
rect 511766 645360 511778 645394
rect 511720 645326 511778 645360
rect 511720 645292 511732 645326
rect 511766 645292 511778 645326
rect 511720 645258 511778 645292
rect 511720 645224 511732 645258
rect 511766 645224 511778 645258
rect 511720 645190 511778 645224
rect 511720 645156 511732 645190
rect 511766 645156 511778 645190
rect 511720 645122 511778 645156
rect 511720 645088 511732 645122
rect 511766 645088 511778 645122
rect 511720 645054 511778 645088
rect 511720 645020 511732 645054
rect 511766 645020 511778 645054
rect 511720 644986 511778 645020
rect 511720 644952 511732 644986
rect 511766 644952 511778 644986
rect 511720 644918 511778 644952
rect 511720 644884 511732 644918
rect 511766 644884 511778 644918
rect 511720 644850 511778 644884
rect 511720 644816 511732 644850
rect 511766 644816 511778 644850
rect 511720 644782 511778 644816
rect 511720 644748 511732 644782
rect 511766 644748 511778 644782
rect 511720 644714 511778 644748
rect 511720 644680 511732 644714
rect 511766 644680 511778 644714
rect 511720 644646 511778 644680
rect 511720 644612 511732 644646
rect 511766 644612 511778 644646
rect 511720 644578 511778 644612
rect 511720 644544 511732 644578
rect 511766 644544 511778 644578
rect 511720 644503 511778 644544
rect 512178 645462 512236 645503
rect 512178 645428 512190 645462
rect 512224 645428 512236 645462
rect 512178 645394 512236 645428
rect 512178 645360 512190 645394
rect 512224 645360 512236 645394
rect 512178 645326 512236 645360
rect 512178 645292 512190 645326
rect 512224 645292 512236 645326
rect 512178 645258 512236 645292
rect 512178 645224 512190 645258
rect 512224 645224 512236 645258
rect 512178 645190 512236 645224
rect 512178 645156 512190 645190
rect 512224 645156 512236 645190
rect 512178 645122 512236 645156
rect 512178 645088 512190 645122
rect 512224 645088 512236 645122
rect 512178 645054 512236 645088
rect 512178 645020 512190 645054
rect 512224 645020 512236 645054
rect 512178 644986 512236 645020
rect 512178 644952 512190 644986
rect 512224 644952 512236 644986
rect 512178 644918 512236 644952
rect 512178 644884 512190 644918
rect 512224 644884 512236 644918
rect 512178 644850 512236 644884
rect 512178 644816 512190 644850
rect 512224 644816 512236 644850
rect 512178 644782 512236 644816
rect 512178 644748 512190 644782
rect 512224 644748 512236 644782
rect 512178 644714 512236 644748
rect 512178 644680 512190 644714
rect 512224 644680 512236 644714
rect 512178 644646 512236 644680
rect 512178 644612 512190 644646
rect 512224 644612 512236 644646
rect 512178 644578 512236 644612
rect 512178 644544 512190 644578
rect 512224 644544 512236 644578
rect 512178 644503 512236 644544
rect 512636 645462 512694 645503
rect 512636 645428 512648 645462
rect 512682 645428 512694 645462
rect 512636 645394 512694 645428
rect 512636 645360 512648 645394
rect 512682 645360 512694 645394
rect 512636 645326 512694 645360
rect 512636 645292 512648 645326
rect 512682 645292 512694 645326
rect 512636 645258 512694 645292
rect 512636 645224 512648 645258
rect 512682 645224 512694 645258
rect 512636 645190 512694 645224
rect 512636 645156 512648 645190
rect 512682 645156 512694 645190
rect 512636 645122 512694 645156
rect 512636 645088 512648 645122
rect 512682 645088 512694 645122
rect 512636 645054 512694 645088
rect 512636 645020 512648 645054
rect 512682 645020 512694 645054
rect 512636 644986 512694 645020
rect 512636 644952 512648 644986
rect 512682 644952 512694 644986
rect 512636 644918 512694 644952
rect 512636 644884 512648 644918
rect 512682 644884 512694 644918
rect 512636 644850 512694 644884
rect 512636 644816 512648 644850
rect 512682 644816 512694 644850
rect 512636 644782 512694 644816
rect 512636 644748 512648 644782
rect 512682 644748 512694 644782
rect 512636 644714 512694 644748
rect 512636 644680 512648 644714
rect 512682 644680 512694 644714
rect 512636 644646 512694 644680
rect 512636 644612 512648 644646
rect 512682 644612 512694 644646
rect 512636 644578 512694 644612
rect 512636 644544 512648 644578
rect 512682 644544 512694 644578
rect 512636 644503 512694 644544
rect 513094 645462 513152 645503
rect 513094 645428 513106 645462
rect 513140 645428 513152 645462
rect 513094 645394 513152 645428
rect 513094 645360 513106 645394
rect 513140 645360 513152 645394
rect 513094 645326 513152 645360
rect 513094 645292 513106 645326
rect 513140 645292 513152 645326
rect 513094 645258 513152 645292
rect 513094 645224 513106 645258
rect 513140 645224 513152 645258
rect 513094 645190 513152 645224
rect 513094 645156 513106 645190
rect 513140 645156 513152 645190
rect 513094 645122 513152 645156
rect 513094 645088 513106 645122
rect 513140 645088 513152 645122
rect 513094 645054 513152 645088
rect 513094 645020 513106 645054
rect 513140 645020 513152 645054
rect 513094 644986 513152 645020
rect 513094 644952 513106 644986
rect 513140 644952 513152 644986
rect 513094 644918 513152 644952
rect 513094 644884 513106 644918
rect 513140 644884 513152 644918
rect 513094 644850 513152 644884
rect 513094 644816 513106 644850
rect 513140 644816 513152 644850
rect 513094 644782 513152 644816
rect 513094 644748 513106 644782
rect 513140 644748 513152 644782
rect 513094 644714 513152 644748
rect 513094 644680 513106 644714
rect 513140 644680 513152 644714
rect 513094 644646 513152 644680
rect 513094 644612 513106 644646
rect 513140 644612 513152 644646
rect 513094 644578 513152 644612
rect 513094 644544 513106 644578
rect 513140 644544 513152 644578
rect 513094 644503 513152 644544
rect 513552 645462 513610 645503
rect 513552 645428 513564 645462
rect 513598 645428 513610 645462
rect 513552 645394 513610 645428
rect 513552 645360 513564 645394
rect 513598 645360 513610 645394
rect 513552 645326 513610 645360
rect 513552 645292 513564 645326
rect 513598 645292 513610 645326
rect 513552 645258 513610 645292
rect 513552 645224 513564 645258
rect 513598 645224 513610 645258
rect 513552 645190 513610 645224
rect 513552 645156 513564 645190
rect 513598 645156 513610 645190
rect 513552 645122 513610 645156
rect 513552 645088 513564 645122
rect 513598 645088 513610 645122
rect 513552 645054 513610 645088
rect 513552 645020 513564 645054
rect 513598 645020 513610 645054
rect 513552 644986 513610 645020
rect 513552 644952 513564 644986
rect 513598 644952 513610 644986
rect 513552 644918 513610 644952
rect 513552 644884 513564 644918
rect 513598 644884 513610 644918
rect 513552 644850 513610 644884
rect 513552 644816 513564 644850
rect 513598 644816 513610 644850
rect 513552 644782 513610 644816
rect 513552 644748 513564 644782
rect 513598 644748 513610 644782
rect 513552 644714 513610 644748
rect 513552 644680 513564 644714
rect 513598 644680 513610 644714
rect 513552 644646 513610 644680
rect 513552 644612 513564 644646
rect 513598 644612 513610 644646
rect 513552 644578 513610 644612
rect 513552 644544 513564 644578
rect 513598 644544 513610 644578
rect 513552 644503 513610 644544
rect 514010 645462 514068 645503
rect 514010 645428 514022 645462
rect 514056 645428 514068 645462
rect 514010 645394 514068 645428
rect 514010 645360 514022 645394
rect 514056 645360 514068 645394
rect 514010 645326 514068 645360
rect 514010 645292 514022 645326
rect 514056 645292 514068 645326
rect 514010 645258 514068 645292
rect 514010 645224 514022 645258
rect 514056 645224 514068 645258
rect 514010 645190 514068 645224
rect 514010 645156 514022 645190
rect 514056 645156 514068 645190
rect 514010 645122 514068 645156
rect 514010 645088 514022 645122
rect 514056 645088 514068 645122
rect 514010 645054 514068 645088
rect 514010 645020 514022 645054
rect 514056 645020 514068 645054
rect 514010 644986 514068 645020
rect 514010 644952 514022 644986
rect 514056 644952 514068 644986
rect 514010 644918 514068 644952
rect 514010 644884 514022 644918
rect 514056 644884 514068 644918
rect 514010 644850 514068 644884
rect 514010 644816 514022 644850
rect 514056 644816 514068 644850
rect 514010 644782 514068 644816
rect 514010 644748 514022 644782
rect 514056 644748 514068 644782
rect 514010 644714 514068 644748
rect 514010 644680 514022 644714
rect 514056 644680 514068 644714
rect 514010 644646 514068 644680
rect 514010 644612 514022 644646
rect 514056 644612 514068 644646
rect 514010 644578 514068 644612
rect 514010 644544 514022 644578
rect 514056 644544 514068 644578
rect 514010 644503 514068 644544
rect 514468 645462 514526 645503
rect 514468 645428 514480 645462
rect 514514 645428 514526 645462
rect 514468 645394 514526 645428
rect 514468 645360 514480 645394
rect 514514 645360 514526 645394
rect 514468 645326 514526 645360
rect 514468 645292 514480 645326
rect 514514 645292 514526 645326
rect 514468 645258 514526 645292
rect 514468 645224 514480 645258
rect 514514 645224 514526 645258
rect 514468 645190 514526 645224
rect 514468 645156 514480 645190
rect 514514 645156 514526 645190
rect 514468 645122 514526 645156
rect 514468 645088 514480 645122
rect 514514 645088 514526 645122
rect 514468 645054 514526 645088
rect 514468 645020 514480 645054
rect 514514 645020 514526 645054
rect 514468 644986 514526 645020
rect 514468 644952 514480 644986
rect 514514 644952 514526 644986
rect 514468 644918 514526 644952
rect 514468 644884 514480 644918
rect 514514 644884 514526 644918
rect 514468 644850 514526 644884
rect 514468 644816 514480 644850
rect 514514 644816 514526 644850
rect 514468 644782 514526 644816
rect 514468 644748 514480 644782
rect 514514 644748 514526 644782
rect 514468 644714 514526 644748
rect 514468 644680 514480 644714
rect 514514 644680 514526 644714
rect 514468 644646 514526 644680
rect 514468 644612 514480 644646
rect 514514 644612 514526 644646
rect 514468 644578 514526 644612
rect 514468 644544 514480 644578
rect 514514 644544 514526 644578
rect 514468 644503 514526 644544
rect 514926 645462 514984 645503
rect 514926 645428 514938 645462
rect 514972 645428 514984 645462
rect 514926 645394 514984 645428
rect 514926 645360 514938 645394
rect 514972 645360 514984 645394
rect 514926 645326 514984 645360
rect 514926 645292 514938 645326
rect 514972 645292 514984 645326
rect 514926 645258 514984 645292
rect 514926 645224 514938 645258
rect 514972 645224 514984 645258
rect 514926 645190 514984 645224
rect 514926 645156 514938 645190
rect 514972 645156 514984 645190
rect 514926 645122 514984 645156
rect 514926 645088 514938 645122
rect 514972 645088 514984 645122
rect 514926 645054 514984 645088
rect 514926 645020 514938 645054
rect 514972 645020 514984 645054
rect 514926 644986 514984 645020
rect 514926 644952 514938 644986
rect 514972 644952 514984 644986
rect 514926 644918 514984 644952
rect 514926 644884 514938 644918
rect 514972 644884 514984 644918
rect 514926 644850 514984 644884
rect 514926 644816 514938 644850
rect 514972 644816 514984 644850
rect 514926 644782 514984 644816
rect 514926 644748 514938 644782
rect 514972 644748 514984 644782
rect 514926 644714 514984 644748
rect 514926 644680 514938 644714
rect 514972 644680 514984 644714
rect 514926 644646 514984 644680
rect 514926 644612 514938 644646
rect 514972 644612 514984 644646
rect 514926 644578 514984 644612
rect 514926 644544 514938 644578
rect 514972 644544 514984 644578
rect 514926 644503 514984 644544
rect 515384 645462 515442 645503
rect 515384 645428 515396 645462
rect 515430 645428 515442 645462
rect 515384 645394 515442 645428
rect 515384 645360 515396 645394
rect 515430 645360 515442 645394
rect 515384 645326 515442 645360
rect 515384 645292 515396 645326
rect 515430 645292 515442 645326
rect 515384 645258 515442 645292
rect 515384 645224 515396 645258
rect 515430 645224 515442 645258
rect 515384 645190 515442 645224
rect 515384 645156 515396 645190
rect 515430 645156 515442 645190
rect 515384 645122 515442 645156
rect 515384 645088 515396 645122
rect 515430 645088 515442 645122
rect 515384 645054 515442 645088
rect 515384 645020 515396 645054
rect 515430 645020 515442 645054
rect 515384 644986 515442 645020
rect 515384 644952 515396 644986
rect 515430 644952 515442 644986
rect 515384 644918 515442 644952
rect 515384 644884 515396 644918
rect 515430 644884 515442 644918
rect 515384 644850 515442 644884
rect 515384 644816 515396 644850
rect 515430 644816 515442 644850
rect 515384 644782 515442 644816
rect 515384 644748 515396 644782
rect 515430 644748 515442 644782
rect 515384 644714 515442 644748
rect 515384 644680 515396 644714
rect 515430 644680 515442 644714
rect 515384 644646 515442 644680
rect 515384 644612 515396 644646
rect 515430 644612 515442 644646
rect 515384 644578 515442 644612
rect 515384 644544 515396 644578
rect 515430 644544 515442 644578
rect 515384 644503 515442 644544
rect 508056 644296 508114 644337
rect 508056 644262 508068 644296
rect 508102 644262 508114 644296
rect 508056 644228 508114 644262
rect 508056 644194 508068 644228
rect 508102 644194 508114 644228
rect 508056 644160 508114 644194
rect 508056 644126 508068 644160
rect 508102 644126 508114 644160
rect 508056 644092 508114 644126
rect 508056 644058 508068 644092
rect 508102 644058 508114 644092
rect 508056 644024 508114 644058
rect 508056 643990 508068 644024
rect 508102 643990 508114 644024
rect 508056 643956 508114 643990
rect 508056 643922 508068 643956
rect 508102 643922 508114 643956
rect 508056 643888 508114 643922
rect 508056 643854 508068 643888
rect 508102 643854 508114 643888
rect 508056 643820 508114 643854
rect 508056 643786 508068 643820
rect 508102 643786 508114 643820
rect 508056 643752 508114 643786
rect 508056 643718 508068 643752
rect 508102 643718 508114 643752
rect 508056 643684 508114 643718
rect 508056 643650 508068 643684
rect 508102 643650 508114 643684
rect 508056 643616 508114 643650
rect 508056 643582 508068 643616
rect 508102 643582 508114 643616
rect 508056 643548 508114 643582
rect 508056 643514 508068 643548
rect 508102 643514 508114 643548
rect 508056 643480 508114 643514
rect 508056 643446 508068 643480
rect 508102 643446 508114 643480
rect 508056 643412 508114 643446
rect 508056 643378 508068 643412
rect 508102 643378 508114 643412
rect 508056 643337 508114 643378
rect 508514 644296 508572 644337
rect 508514 644262 508526 644296
rect 508560 644262 508572 644296
rect 508514 644228 508572 644262
rect 508514 644194 508526 644228
rect 508560 644194 508572 644228
rect 508514 644160 508572 644194
rect 508514 644126 508526 644160
rect 508560 644126 508572 644160
rect 508514 644092 508572 644126
rect 508514 644058 508526 644092
rect 508560 644058 508572 644092
rect 508514 644024 508572 644058
rect 508514 643990 508526 644024
rect 508560 643990 508572 644024
rect 508514 643956 508572 643990
rect 508514 643922 508526 643956
rect 508560 643922 508572 643956
rect 508514 643888 508572 643922
rect 508514 643854 508526 643888
rect 508560 643854 508572 643888
rect 508514 643820 508572 643854
rect 508514 643786 508526 643820
rect 508560 643786 508572 643820
rect 508514 643752 508572 643786
rect 508514 643718 508526 643752
rect 508560 643718 508572 643752
rect 508514 643684 508572 643718
rect 508514 643650 508526 643684
rect 508560 643650 508572 643684
rect 508514 643616 508572 643650
rect 508514 643582 508526 643616
rect 508560 643582 508572 643616
rect 508514 643548 508572 643582
rect 508514 643514 508526 643548
rect 508560 643514 508572 643548
rect 508514 643480 508572 643514
rect 508514 643446 508526 643480
rect 508560 643446 508572 643480
rect 508514 643412 508572 643446
rect 508514 643378 508526 643412
rect 508560 643378 508572 643412
rect 508514 643337 508572 643378
rect 508972 644296 509030 644337
rect 508972 644262 508984 644296
rect 509018 644262 509030 644296
rect 508972 644228 509030 644262
rect 508972 644194 508984 644228
rect 509018 644194 509030 644228
rect 508972 644160 509030 644194
rect 508972 644126 508984 644160
rect 509018 644126 509030 644160
rect 508972 644092 509030 644126
rect 508972 644058 508984 644092
rect 509018 644058 509030 644092
rect 508972 644024 509030 644058
rect 508972 643990 508984 644024
rect 509018 643990 509030 644024
rect 508972 643956 509030 643990
rect 508972 643922 508984 643956
rect 509018 643922 509030 643956
rect 508972 643888 509030 643922
rect 508972 643854 508984 643888
rect 509018 643854 509030 643888
rect 508972 643820 509030 643854
rect 508972 643786 508984 643820
rect 509018 643786 509030 643820
rect 508972 643752 509030 643786
rect 508972 643718 508984 643752
rect 509018 643718 509030 643752
rect 508972 643684 509030 643718
rect 508972 643650 508984 643684
rect 509018 643650 509030 643684
rect 508972 643616 509030 643650
rect 508972 643582 508984 643616
rect 509018 643582 509030 643616
rect 508972 643548 509030 643582
rect 508972 643514 508984 643548
rect 509018 643514 509030 643548
rect 508972 643480 509030 643514
rect 508972 643446 508984 643480
rect 509018 643446 509030 643480
rect 508972 643412 509030 643446
rect 508972 643378 508984 643412
rect 509018 643378 509030 643412
rect 508972 643337 509030 643378
rect 509430 644296 509488 644337
rect 509430 644262 509442 644296
rect 509476 644262 509488 644296
rect 509430 644228 509488 644262
rect 509430 644194 509442 644228
rect 509476 644194 509488 644228
rect 509430 644160 509488 644194
rect 509430 644126 509442 644160
rect 509476 644126 509488 644160
rect 509430 644092 509488 644126
rect 509430 644058 509442 644092
rect 509476 644058 509488 644092
rect 509430 644024 509488 644058
rect 509430 643990 509442 644024
rect 509476 643990 509488 644024
rect 509430 643956 509488 643990
rect 509430 643922 509442 643956
rect 509476 643922 509488 643956
rect 509430 643888 509488 643922
rect 509430 643854 509442 643888
rect 509476 643854 509488 643888
rect 509430 643820 509488 643854
rect 509430 643786 509442 643820
rect 509476 643786 509488 643820
rect 509430 643752 509488 643786
rect 509430 643718 509442 643752
rect 509476 643718 509488 643752
rect 509430 643684 509488 643718
rect 509430 643650 509442 643684
rect 509476 643650 509488 643684
rect 509430 643616 509488 643650
rect 509430 643582 509442 643616
rect 509476 643582 509488 643616
rect 509430 643548 509488 643582
rect 509430 643514 509442 643548
rect 509476 643514 509488 643548
rect 509430 643480 509488 643514
rect 509430 643446 509442 643480
rect 509476 643446 509488 643480
rect 509430 643412 509488 643446
rect 509430 643378 509442 643412
rect 509476 643378 509488 643412
rect 509430 643337 509488 643378
rect 509888 644296 509946 644337
rect 509888 644262 509900 644296
rect 509934 644262 509946 644296
rect 509888 644228 509946 644262
rect 509888 644194 509900 644228
rect 509934 644194 509946 644228
rect 509888 644160 509946 644194
rect 509888 644126 509900 644160
rect 509934 644126 509946 644160
rect 509888 644092 509946 644126
rect 509888 644058 509900 644092
rect 509934 644058 509946 644092
rect 509888 644024 509946 644058
rect 509888 643990 509900 644024
rect 509934 643990 509946 644024
rect 509888 643956 509946 643990
rect 509888 643922 509900 643956
rect 509934 643922 509946 643956
rect 509888 643888 509946 643922
rect 509888 643854 509900 643888
rect 509934 643854 509946 643888
rect 509888 643820 509946 643854
rect 509888 643786 509900 643820
rect 509934 643786 509946 643820
rect 509888 643752 509946 643786
rect 509888 643718 509900 643752
rect 509934 643718 509946 643752
rect 509888 643684 509946 643718
rect 509888 643650 509900 643684
rect 509934 643650 509946 643684
rect 509888 643616 509946 643650
rect 509888 643582 509900 643616
rect 509934 643582 509946 643616
rect 509888 643548 509946 643582
rect 509888 643514 509900 643548
rect 509934 643514 509946 643548
rect 509888 643480 509946 643514
rect 509888 643446 509900 643480
rect 509934 643446 509946 643480
rect 509888 643412 509946 643446
rect 509888 643378 509900 643412
rect 509934 643378 509946 643412
rect 509888 643337 509946 643378
rect 510346 644296 510404 644337
rect 510346 644262 510358 644296
rect 510392 644262 510404 644296
rect 510346 644228 510404 644262
rect 510346 644194 510358 644228
rect 510392 644194 510404 644228
rect 510346 644160 510404 644194
rect 510346 644126 510358 644160
rect 510392 644126 510404 644160
rect 510346 644092 510404 644126
rect 510346 644058 510358 644092
rect 510392 644058 510404 644092
rect 510346 644024 510404 644058
rect 510346 643990 510358 644024
rect 510392 643990 510404 644024
rect 510346 643956 510404 643990
rect 510346 643922 510358 643956
rect 510392 643922 510404 643956
rect 510346 643888 510404 643922
rect 510346 643854 510358 643888
rect 510392 643854 510404 643888
rect 510346 643820 510404 643854
rect 510346 643786 510358 643820
rect 510392 643786 510404 643820
rect 510346 643752 510404 643786
rect 510346 643718 510358 643752
rect 510392 643718 510404 643752
rect 510346 643684 510404 643718
rect 510346 643650 510358 643684
rect 510392 643650 510404 643684
rect 510346 643616 510404 643650
rect 510346 643582 510358 643616
rect 510392 643582 510404 643616
rect 510346 643548 510404 643582
rect 510346 643514 510358 643548
rect 510392 643514 510404 643548
rect 510346 643480 510404 643514
rect 510346 643446 510358 643480
rect 510392 643446 510404 643480
rect 510346 643412 510404 643446
rect 510346 643378 510358 643412
rect 510392 643378 510404 643412
rect 510346 643337 510404 643378
rect 510804 644296 510862 644337
rect 510804 644262 510816 644296
rect 510850 644262 510862 644296
rect 510804 644228 510862 644262
rect 510804 644194 510816 644228
rect 510850 644194 510862 644228
rect 510804 644160 510862 644194
rect 510804 644126 510816 644160
rect 510850 644126 510862 644160
rect 510804 644092 510862 644126
rect 510804 644058 510816 644092
rect 510850 644058 510862 644092
rect 510804 644024 510862 644058
rect 510804 643990 510816 644024
rect 510850 643990 510862 644024
rect 510804 643956 510862 643990
rect 510804 643922 510816 643956
rect 510850 643922 510862 643956
rect 510804 643888 510862 643922
rect 510804 643854 510816 643888
rect 510850 643854 510862 643888
rect 510804 643820 510862 643854
rect 510804 643786 510816 643820
rect 510850 643786 510862 643820
rect 510804 643752 510862 643786
rect 510804 643718 510816 643752
rect 510850 643718 510862 643752
rect 510804 643684 510862 643718
rect 510804 643650 510816 643684
rect 510850 643650 510862 643684
rect 510804 643616 510862 643650
rect 510804 643582 510816 643616
rect 510850 643582 510862 643616
rect 510804 643548 510862 643582
rect 510804 643514 510816 643548
rect 510850 643514 510862 643548
rect 510804 643480 510862 643514
rect 510804 643446 510816 643480
rect 510850 643446 510862 643480
rect 510804 643412 510862 643446
rect 510804 643378 510816 643412
rect 510850 643378 510862 643412
rect 510804 643337 510862 643378
rect 511262 644296 511320 644337
rect 511262 644262 511274 644296
rect 511308 644262 511320 644296
rect 511262 644228 511320 644262
rect 511262 644194 511274 644228
rect 511308 644194 511320 644228
rect 511262 644160 511320 644194
rect 511262 644126 511274 644160
rect 511308 644126 511320 644160
rect 511262 644092 511320 644126
rect 511262 644058 511274 644092
rect 511308 644058 511320 644092
rect 511262 644024 511320 644058
rect 511262 643990 511274 644024
rect 511308 643990 511320 644024
rect 511262 643956 511320 643990
rect 511262 643922 511274 643956
rect 511308 643922 511320 643956
rect 511262 643888 511320 643922
rect 511262 643854 511274 643888
rect 511308 643854 511320 643888
rect 511262 643820 511320 643854
rect 511262 643786 511274 643820
rect 511308 643786 511320 643820
rect 511262 643752 511320 643786
rect 511262 643718 511274 643752
rect 511308 643718 511320 643752
rect 511262 643684 511320 643718
rect 511262 643650 511274 643684
rect 511308 643650 511320 643684
rect 511262 643616 511320 643650
rect 511262 643582 511274 643616
rect 511308 643582 511320 643616
rect 511262 643548 511320 643582
rect 511262 643514 511274 643548
rect 511308 643514 511320 643548
rect 511262 643480 511320 643514
rect 511262 643446 511274 643480
rect 511308 643446 511320 643480
rect 511262 643412 511320 643446
rect 511262 643378 511274 643412
rect 511308 643378 511320 643412
rect 511262 643337 511320 643378
rect 511720 644296 511778 644337
rect 511720 644262 511732 644296
rect 511766 644262 511778 644296
rect 511720 644228 511778 644262
rect 511720 644194 511732 644228
rect 511766 644194 511778 644228
rect 511720 644160 511778 644194
rect 511720 644126 511732 644160
rect 511766 644126 511778 644160
rect 511720 644092 511778 644126
rect 511720 644058 511732 644092
rect 511766 644058 511778 644092
rect 511720 644024 511778 644058
rect 511720 643990 511732 644024
rect 511766 643990 511778 644024
rect 511720 643956 511778 643990
rect 511720 643922 511732 643956
rect 511766 643922 511778 643956
rect 511720 643888 511778 643922
rect 511720 643854 511732 643888
rect 511766 643854 511778 643888
rect 511720 643820 511778 643854
rect 511720 643786 511732 643820
rect 511766 643786 511778 643820
rect 511720 643752 511778 643786
rect 511720 643718 511732 643752
rect 511766 643718 511778 643752
rect 511720 643684 511778 643718
rect 511720 643650 511732 643684
rect 511766 643650 511778 643684
rect 511720 643616 511778 643650
rect 511720 643582 511732 643616
rect 511766 643582 511778 643616
rect 511720 643548 511778 643582
rect 511720 643514 511732 643548
rect 511766 643514 511778 643548
rect 511720 643480 511778 643514
rect 511720 643446 511732 643480
rect 511766 643446 511778 643480
rect 511720 643412 511778 643446
rect 511720 643378 511732 643412
rect 511766 643378 511778 643412
rect 511720 643337 511778 643378
rect 512178 644296 512236 644337
rect 512178 644262 512190 644296
rect 512224 644262 512236 644296
rect 512178 644228 512236 644262
rect 512178 644194 512190 644228
rect 512224 644194 512236 644228
rect 512178 644160 512236 644194
rect 512178 644126 512190 644160
rect 512224 644126 512236 644160
rect 512178 644092 512236 644126
rect 512178 644058 512190 644092
rect 512224 644058 512236 644092
rect 512178 644024 512236 644058
rect 512178 643990 512190 644024
rect 512224 643990 512236 644024
rect 512178 643956 512236 643990
rect 512178 643922 512190 643956
rect 512224 643922 512236 643956
rect 512178 643888 512236 643922
rect 512178 643854 512190 643888
rect 512224 643854 512236 643888
rect 512178 643820 512236 643854
rect 512178 643786 512190 643820
rect 512224 643786 512236 643820
rect 512178 643752 512236 643786
rect 512178 643718 512190 643752
rect 512224 643718 512236 643752
rect 512178 643684 512236 643718
rect 512178 643650 512190 643684
rect 512224 643650 512236 643684
rect 512178 643616 512236 643650
rect 512178 643582 512190 643616
rect 512224 643582 512236 643616
rect 512178 643548 512236 643582
rect 512178 643514 512190 643548
rect 512224 643514 512236 643548
rect 512178 643480 512236 643514
rect 512178 643446 512190 643480
rect 512224 643446 512236 643480
rect 512178 643412 512236 643446
rect 512178 643378 512190 643412
rect 512224 643378 512236 643412
rect 512178 643337 512236 643378
rect 512636 644296 512694 644337
rect 512636 644262 512648 644296
rect 512682 644262 512694 644296
rect 512636 644228 512694 644262
rect 512636 644194 512648 644228
rect 512682 644194 512694 644228
rect 512636 644160 512694 644194
rect 512636 644126 512648 644160
rect 512682 644126 512694 644160
rect 512636 644092 512694 644126
rect 512636 644058 512648 644092
rect 512682 644058 512694 644092
rect 512636 644024 512694 644058
rect 512636 643990 512648 644024
rect 512682 643990 512694 644024
rect 512636 643956 512694 643990
rect 512636 643922 512648 643956
rect 512682 643922 512694 643956
rect 512636 643888 512694 643922
rect 512636 643854 512648 643888
rect 512682 643854 512694 643888
rect 512636 643820 512694 643854
rect 512636 643786 512648 643820
rect 512682 643786 512694 643820
rect 512636 643752 512694 643786
rect 512636 643718 512648 643752
rect 512682 643718 512694 643752
rect 512636 643684 512694 643718
rect 512636 643650 512648 643684
rect 512682 643650 512694 643684
rect 512636 643616 512694 643650
rect 512636 643582 512648 643616
rect 512682 643582 512694 643616
rect 512636 643548 512694 643582
rect 512636 643514 512648 643548
rect 512682 643514 512694 643548
rect 512636 643480 512694 643514
rect 512636 643446 512648 643480
rect 512682 643446 512694 643480
rect 512636 643412 512694 643446
rect 512636 643378 512648 643412
rect 512682 643378 512694 643412
rect 512636 643337 512694 643378
rect 513094 644296 513152 644337
rect 513094 644262 513106 644296
rect 513140 644262 513152 644296
rect 513094 644228 513152 644262
rect 513094 644194 513106 644228
rect 513140 644194 513152 644228
rect 513094 644160 513152 644194
rect 513094 644126 513106 644160
rect 513140 644126 513152 644160
rect 513094 644092 513152 644126
rect 513094 644058 513106 644092
rect 513140 644058 513152 644092
rect 513094 644024 513152 644058
rect 513094 643990 513106 644024
rect 513140 643990 513152 644024
rect 513094 643956 513152 643990
rect 513094 643922 513106 643956
rect 513140 643922 513152 643956
rect 513094 643888 513152 643922
rect 513094 643854 513106 643888
rect 513140 643854 513152 643888
rect 513094 643820 513152 643854
rect 513094 643786 513106 643820
rect 513140 643786 513152 643820
rect 513094 643752 513152 643786
rect 513094 643718 513106 643752
rect 513140 643718 513152 643752
rect 513094 643684 513152 643718
rect 513094 643650 513106 643684
rect 513140 643650 513152 643684
rect 513094 643616 513152 643650
rect 513094 643582 513106 643616
rect 513140 643582 513152 643616
rect 513094 643548 513152 643582
rect 513094 643514 513106 643548
rect 513140 643514 513152 643548
rect 513094 643480 513152 643514
rect 513094 643446 513106 643480
rect 513140 643446 513152 643480
rect 513094 643412 513152 643446
rect 513094 643378 513106 643412
rect 513140 643378 513152 643412
rect 513094 643337 513152 643378
rect 513552 644296 513610 644337
rect 513552 644262 513564 644296
rect 513598 644262 513610 644296
rect 513552 644228 513610 644262
rect 513552 644194 513564 644228
rect 513598 644194 513610 644228
rect 513552 644160 513610 644194
rect 513552 644126 513564 644160
rect 513598 644126 513610 644160
rect 513552 644092 513610 644126
rect 513552 644058 513564 644092
rect 513598 644058 513610 644092
rect 513552 644024 513610 644058
rect 513552 643990 513564 644024
rect 513598 643990 513610 644024
rect 513552 643956 513610 643990
rect 513552 643922 513564 643956
rect 513598 643922 513610 643956
rect 513552 643888 513610 643922
rect 513552 643854 513564 643888
rect 513598 643854 513610 643888
rect 513552 643820 513610 643854
rect 513552 643786 513564 643820
rect 513598 643786 513610 643820
rect 513552 643752 513610 643786
rect 513552 643718 513564 643752
rect 513598 643718 513610 643752
rect 513552 643684 513610 643718
rect 513552 643650 513564 643684
rect 513598 643650 513610 643684
rect 513552 643616 513610 643650
rect 513552 643582 513564 643616
rect 513598 643582 513610 643616
rect 513552 643548 513610 643582
rect 513552 643514 513564 643548
rect 513598 643514 513610 643548
rect 513552 643480 513610 643514
rect 513552 643446 513564 643480
rect 513598 643446 513610 643480
rect 513552 643412 513610 643446
rect 513552 643378 513564 643412
rect 513598 643378 513610 643412
rect 513552 643337 513610 643378
rect 514010 644296 514068 644337
rect 514010 644262 514022 644296
rect 514056 644262 514068 644296
rect 514010 644228 514068 644262
rect 514010 644194 514022 644228
rect 514056 644194 514068 644228
rect 514010 644160 514068 644194
rect 514010 644126 514022 644160
rect 514056 644126 514068 644160
rect 514010 644092 514068 644126
rect 514010 644058 514022 644092
rect 514056 644058 514068 644092
rect 514010 644024 514068 644058
rect 514010 643990 514022 644024
rect 514056 643990 514068 644024
rect 514010 643956 514068 643990
rect 514010 643922 514022 643956
rect 514056 643922 514068 643956
rect 514010 643888 514068 643922
rect 514010 643854 514022 643888
rect 514056 643854 514068 643888
rect 514010 643820 514068 643854
rect 514010 643786 514022 643820
rect 514056 643786 514068 643820
rect 514010 643752 514068 643786
rect 514010 643718 514022 643752
rect 514056 643718 514068 643752
rect 514010 643684 514068 643718
rect 514010 643650 514022 643684
rect 514056 643650 514068 643684
rect 514010 643616 514068 643650
rect 514010 643582 514022 643616
rect 514056 643582 514068 643616
rect 514010 643548 514068 643582
rect 514010 643514 514022 643548
rect 514056 643514 514068 643548
rect 514010 643480 514068 643514
rect 514010 643446 514022 643480
rect 514056 643446 514068 643480
rect 514010 643412 514068 643446
rect 514010 643378 514022 643412
rect 514056 643378 514068 643412
rect 514010 643337 514068 643378
rect 514468 644296 514526 644337
rect 514468 644262 514480 644296
rect 514514 644262 514526 644296
rect 514468 644228 514526 644262
rect 514468 644194 514480 644228
rect 514514 644194 514526 644228
rect 514468 644160 514526 644194
rect 514468 644126 514480 644160
rect 514514 644126 514526 644160
rect 514468 644092 514526 644126
rect 514468 644058 514480 644092
rect 514514 644058 514526 644092
rect 514468 644024 514526 644058
rect 514468 643990 514480 644024
rect 514514 643990 514526 644024
rect 514468 643956 514526 643990
rect 514468 643922 514480 643956
rect 514514 643922 514526 643956
rect 514468 643888 514526 643922
rect 514468 643854 514480 643888
rect 514514 643854 514526 643888
rect 514468 643820 514526 643854
rect 514468 643786 514480 643820
rect 514514 643786 514526 643820
rect 514468 643752 514526 643786
rect 514468 643718 514480 643752
rect 514514 643718 514526 643752
rect 514468 643684 514526 643718
rect 514468 643650 514480 643684
rect 514514 643650 514526 643684
rect 514468 643616 514526 643650
rect 514468 643582 514480 643616
rect 514514 643582 514526 643616
rect 514468 643548 514526 643582
rect 514468 643514 514480 643548
rect 514514 643514 514526 643548
rect 514468 643480 514526 643514
rect 514468 643446 514480 643480
rect 514514 643446 514526 643480
rect 514468 643412 514526 643446
rect 514468 643378 514480 643412
rect 514514 643378 514526 643412
rect 514468 643337 514526 643378
rect 514926 644296 514984 644337
rect 514926 644262 514938 644296
rect 514972 644262 514984 644296
rect 514926 644228 514984 644262
rect 514926 644194 514938 644228
rect 514972 644194 514984 644228
rect 514926 644160 514984 644194
rect 514926 644126 514938 644160
rect 514972 644126 514984 644160
rect 514926 644092 514984 644126
rect 514926 644058 514938 644092
rect 514972 644058 514984 644092
rect 514926 644024 514984 644058
rect 514926 643990 514938 644024
rect 514972 643990 514984 644024
rect 514926 643956 514984 643990
rect 514926 643922 514938 643956
rect 514972 643922 514984 643956
rect 514926 643888 514984 643922
rect 514926 643854 514938 643888
rect 514972 643854 514984 643888
rect 514926 643820 514984 643854
rect 514926 643786 514938 643820
rect 514972 643786 514984 643820
rect 514926 643752 514984 643786
rect 514926 643718 514938 643752
rect 514972 643718 514984 643752
rect 514926 643684 514984 643718
rect 514926 643650 514938 643684
rect 514972 643650 514984 643684
rect 514926 643616 514984 643650
rect 514926 643582 514938 643616
rect 514972 643582 514984 643616
rect 514926 643548 514984 643582
rect 514926 643514 514938 643548
rect 514972 643514 514984 643548
rect 514926 643480 514984 643514
rect 514926 643446 514938 643480
rect 514972 643446 514984 643480
rect 514926 643412 514984 643446
rect 514926 643378 514938 643412
rect 514972 643378 514984 643412
rect 514926 643337 514984 643378
rect 515384 644296 515442 644337
rect 515384 644262 515396 644296
rect 515430 644262 515442 644296
rect 515384 644228 515442 644262
rect 515384 644194 515396 644228
rect 515430 644194 515442 644228
rect 515384 644160 515442 644194
rect 515384 644126 515396 644160
rect 515430 644126 515442 644160
rect 515384 644092 515442 644126
rect 515384 644058 515396 644092
rect 515430 644058 515442 644092
rect 515384 644024 515442 644058
rect 515384 643990 515396 644024
rect 515430 643990 515442 644024
rect 515384 643956 515442 643990
rect 515384 643922 515396 643956
rect 515430 643922 515442 643956
rect 515384 643888 515442 643922
rect 515384 643854 515396 643888
rect 515430 643854 515442 643888
rect 515384 643820 515442 643854
rect 515384 643786 515396 643820
rect 515430 643786 515442 643820
rect 515384 643752 515442 643786
rect 515384 643718 515396 643752
rect 515430 643718 515442 643752
rect 515384 643684 515442 643718
rect 515384 643650 515396 643684
rect 515430 643650 515442 643684
rect 515384 643616 515442 643650
rect 515384 643582 515396 643616
rect 515430 643582 515442 643616
rect 515384 643548 515442 643582
rect 515384 643514 515396 643548
rect 515430 643514 515442 643548
rect 515384 643480 515442 643514
rect 515384 643446 515396 643480
rect 515430 643446 515442 643480
rect 515384 643412 515442 643446
rect 515384 643378 515396 643412
rect 515430 643378 515442 643412
rect 515384 643337 515442 643378
rect 515760 645306 515818 645337
rect 515760 645272 515772 645306
rect 515806 645272 515818 645306
rect 515760 645238 515818 645272
rect 515760 645204 515772 645238
rect 515806 645204 515818 645238
rect 515760 645170 515818 645204
rect 515760 645136 515772 645170
rect 515806 645136 515818 645170
rect 515760 645102 515818 645136
rect 515760 645068 515772 645102
rect 515806 645068 515818 645102
rect 515760 645034 515818 645068
rect 515760 645000 515772 645034
rect 515806 645000 515818 645034
rect 515760 644966 515818 645000
rect 515760 644932 515772 644966
rect 515806 644932 515818 644966
rect 515760 644898 515818 644932
rect 515760 644864 515772 644898
rect 515806 644864 515818 644898
rect 515760 644830 515818 644864
rect 515760 644796 515772 644830
rect 515806 644796 515818 644830
rect 515760 644762 515818 644796
rect 515760 644728 515772 644762
rect 515806 644728 515818 644762
rect 515760 644694 515818 644728
rect 515760 644660 515772 644694
rect 515806 644660 515818 644694
rect 515760 644626 515818 644660
rect 515760 644592 515772 644626
rect 515806 644592 515818 644626
rect 515760 644558 515818 644592
rect 515760 644524 515772 644558
rect 515806 644524 515818 644558
rect 515760 644490 515818 644524
rect 515760 644456 515772 644490
rect 515806 644456 515818 644490
rect 515760 644422 515818 644456
rect 515760 644388 515772 644422
rect 515806 644388 515818 644422
rect 515760 644354 515818 644388
rect 515760 644320 515772 644354
rect 515806 644320 515818 644354
rect 515760 644286 515818 644320
rect 515760 644252 515772 644286
rect 515806 644252 515818 644286
rect 515760 644218 515818 644252
rect 515760 644184 515772 644218
rect 515806 644184 515818 644218
rect 515760 644150 515818 644184
rect 515760 644116 515772 644150
rect 515806 644116 515818 644150
rect 515760 644082 515818 644116
rect 515760 644048 515772 644082
rect 515806 644048 515818 644082
rect 515760 644014 515818 644048
rect 515760 643980 515772 644014
rect 515806 643980 515818 644014
rect 515760 643946 515818 643980
rect 515760 643912 515772 643946
rect 515806 643912 515818 643946
rect 515760 643878 515818 643912
rect 515760 643844 515772 643878
rect 515806 643844 515818 643878
rect 515760 643810 515818 643844
rect 515760 643776 515772 643810
rect 515806 643776 515818 643810
rect 515760 643742 515818 643776
rect 515760 643708 515772 643742
rect 515806 643708 515818 643742
rect 515760 643674 515818 643708
rect 515760 643640 515772 643674
rect 515806 643640 515818 643674
rect 515760 643606 515818 643640
rect 515760 643572 515772 643606
rect 515806 643572 515818 643606
rect 515760 643538 515818 643572
rect 515760 643504 515772 643538
rect 515806 643504 515818 643538
rect 515760 643470 515818 643504
rect 515760 643436 515772 643470
rect 515806 643436 515818 643470
rect 515760 643402 515818 643436
rect 515760 643368 515772 643402
rect 515806 643368 515818 643402
rect 515760 643337 515818 643368
rect 516218 645306 516276 645337
rect 516218 645272 516230 645306
rect 516264 645272 516276 645306
rect 516218 645238 516276 645272
rect 516218 645204 516230 645238
rect 516264 645204 516276 645238
rect 516218 645170 516276 645204
rect 516218 645136 516230 645170
rect 516264 645136 516276 645170
rect 516218 645102 516276 645136
rect 516218 645068 516230 645102
rect 516264 645068 516276 645102
rect 516218 645034 516276 645068
rect 516218 645000 516230 645034
rect 516264 645000 516276 645034
rect 516218 644966 516276 645000
rect 516218 644932 516230 644966
rect 516264 644932 516276 644966
rect 516218 644898 516276 644932
rect 516218 644864 516230 644898
rect 516264 644864 516276 644898
rect 516218 644830 516276 644864
rect 516218 644796 516230 644830
rect 516264 644796 516276 644830
rect 516218 644762 516276 644796
rect 516218 644728 516230 644762
rect 516264 644728 516276 644762
rect 516218 644694 516276 644728
rect 516218 644660 516230 644694
rect 516264 644660 516276 644694
rect 516218 644626 516276 644660
rect 516218 644592 516230 644626
rect 516264 644592 516276 644626
rect 516218 644558 516276 644592
rect 516218 644524 516230 644558
rect 516264 644524 516276 644558
rect 516218 644490 516276 644524
rect 516218 644456 516230 644490
rect 516264 644456 516276 644490
rect 516218 644422 516276 644456
rect 516218 644388 516230 644422
rect 516264 644388 516276 644422
rect 516218 644354 516276 644388
rect 516218 644320 516230 644354
rect 516264 644320 516276 644354
rect 516218 644286 516276 644320
rect 516218 644252 516230 644286
rect 516264 644252 516276 644286
rect 516218 644218 516276 644252
rect 516218 644184 516230 644218
rect 516264 644184 516276 644218
rect 516218 644150 516276 644184
rect 516218 644116 516230 644150
rect 516264 644116 516276 644150
rect 516218 644082 516276 644116
rect 516218 644048 516230 644082
rect 516264 644048 516276 644082
rect 516218 644014 516276 644048
rect 516218 643980 516230 644014
rect 516264 643980 516276 644014
rect 516218 643946 516276 643980
rect 516218 643912 516230 643946
rect 516264 643912 516276 643946
rect 516218 643878 516276 643912
rect 516218 643844 516230 643878
rect 516264 643844 516276 643878
rect 516218 643810 516276 643844
rect 516218 643776 516230 643810
rect 516264 643776 516276 643810
rect 516218 643742 516276 643776
rect 516218 643708 516230 643742
rect 516264 643708 516276 643742
rect 516218 643674 516276 643708
rect 516218 643640 516230 643674
rect 516264 643640 516276 643674
rect 516218 643606 516276 643640
rect 516218 643572 516230 643606
rect 516264 643572 516276 643606
rect 516218 643538 516276 643572
rect 516218 643504 516230 643538
rect 516264 643504 516276 643538
rect 516218 643470 516276 643504
rect 516218 643436 516230 643470
rect 516264 643436 516276 643470
rect 516218 643402 516276 643436
rect 516218 643368 516230 643402
rect 516264 643368 516276 643402
rect 516218 643337 516276 643368
rect 516676 645306 516734 645337
rect 516676 645272 516688 645306
rect 516722 645272 516734 645306
rect 516676 645238 516734 645272
rect 516676 645204 516688 645238
rect 516722 645204 516734 645238
rect 516676 645170 516734 645204
rect 516676 645136 516688 645170
rect 516722 645136 516734 645170
rect 516676 645102 516734 645136
rect 516676 645068 516688 645102
rect 516722 645068 516734 645102
rect 516676 645034 516734 645068
rect 516676 645000 516688 645034
rect 516722 645000 516734 645034
rect 516676 644966 516734 645000
rect 516676 644932 516688 644966
rect 516722 644932 516734 644966
rect 516676 644898 516734 644932
rect 516676 644864 516688 644898
rect 516722 644864 516734 644898
rect 516676 644830 516734 644864
rect 516676 644796 516688 644830
rect 516722 644796 516734 644830
rect 516676 644762 516734 644796
rect 516676 644728 516688 644762
rect 516722 644728 516734 644762
rect 516676 644694 516734 644728
rect 516676 644660 516688 644694
rect 516722 644660 516734 644694
rect 516676 644626 516734 644660
rect 516676 644592 516688 644626
rect 516722 644592 516734 644626
rect 516676 644558 516734 644592
rect 516676 644524 516688 644558
rect 516722 644524 516734 644558
rect 516676 644490 516734 644524
rect 516676 644456 516688 644490
rect 516722 644456 516734 644490
rect 516676 644422 516734 644456
rect 516676 644388 516688 644422
rect 516722 644388 516734 644422
rect 516676 644354 516734 644388
rect 516676 644320 516688 644354
rect 516722 644320 516734 644354
rect 516676 644286 516734 644320
rect 516676 644252 516688 644286
rect 516722 644252 516734 644286
rect 516676 644218 516734 644252
rect 516676 644184 516688 644218
rect 516722 644184 516734 644218
rect 516676 644150 516734 644184
rect 516676 644116 516688 644150
rect 516722 644116 516734 644150
rect 516676 644082 516734 644116
rect 516676 644048 516688 644082
rect 516722 644048 516734 644082
rect 516676 644014 516734 644048
rect 516676 643980 516688 644014
rect 516722 643980 516734 644014
rect 516676 643946 516734 643980
rect 516676 643912 516688 643946
rect 516722 643912 516734 643946
rect 516676 643878 516734 643912
rect 516676 643844 516688 643878
rect 516722 643844 516734 643878
rect 516676 643810 516734 643844
rect 516676 643776 516688 643810
rect 516722 643776 516734 643810
rect 516676 643742 516734 643776
rect 516676 643708 516688 643742
rect 516722 643708 516734 643742
rect 516676 643674 516734 643708
rect 516676 643640 516688 643674
rect 516722 643640 516734 643674
rect 516676 643606 516734 643640
rect 516676 643572 516688 643606
rect 516722 643572 516734 643606
rect 516676 643538 516734 643572
rect 516676 643504 516688 643538
rect 516722 643504 516734 643538
rect 516676 643470 516734 643504
rect 516676 643436 516688 643470
rect 516722 643436 516734 643470
rect 516676 643402 516734 643436
rect 516676 643368 516688 643402
rect 516722 643368 516734 643402
rect 516676 643337 516734 643368
<< mvndiffc >>
rect 508068 642330 508102 642364
rect 508068 642262 508102 642296
rect 508068 642194 508102 642228
rect 508068 642126 508102 642160
rect 508068 642058 508102 642092
rect 508068 641990 508102 642024
rect 508068 641922 508102 641956
rect 508068 641854 508102 641888
rect 508068 641786 508102 641820
rect 508068 641718 508102 641752
rect 508068 641650 508102 641684
rect 508068 641582 508102 641616
rect 508068 641514 508102 641548
rect 508068 641446 508102 641480
rect 508526 642330 508560 642364
rect 508526 642262 508560 642296
rect 508526 642194 508560 642228
rect 508526 642126 508560 642160
rect 508526 642058 508560 642092
rect 508526 641990 508560 642024
rect 508526 641922 508560 641956
rect 508526 641854 508560 641888
rect 508526 641786 508560 641820
rect 508526 641718 508560 641752
rect 508526 641650 508560 641684
rect 508526 641582 508560 641616
rect 508526 641514 508560 641548
rect 508526 641446 508560 641480
rect 508984 642330 509018 642364
rect 508984 642262 509018 642296
rect 508984 642194 509018 642228
rect 508984 642126 509018 642160
rect 508984 642058 509018 642092
rect 508984 641990 509018 642024
rect 508984 641922 509018 641956
rect 508984 641854 509018 641888
rect 508984 641786 509018 641820
rect 508984 641718 509018 641752
rect 508984 641650 509018 641684
rect 508984 641582 509018 641616
rect 508984 641514 509018 641548
rect 508984 641446 509018 641480
rect 509442 642330 509476 642364
rect 509442 642262 509476 642296
rect 509442 642194 509476 642228
rect 509442 642126 509476 642160
rect 509442 642058 509476 642092
rect 509442 641990 509476 642024
rect 509442 641922 509476 641956
rect 509442 641854 509476 641888
rect 509442 641786 509476 641820
rect 509442 641718 509476 641752
rect 509442 641650 509476 641684
rect 509442 641582 509476 641616
rect 509442 641514 509476 641548
rect 509442 641446 509476 641480
rect 509900 642330 509934 642364
rect 509900 642262 509934 642296
rect 509900 642194 509934 642228
rect 509900 642126 509934 642160
rect 509900 642058 509934 642092
rect 509900 641990 509934 642024
rect 509900 641922 509934 641956
rect 509900 641854 509934 641888
rect 509900 641786 509934 641820
rect 509900 641718 509934 641752
rect 509900 641650 509934 641684
rect 509900 641582 509934 641616
rect 509900 641514 509934 641548
rect 509900 641446 509934 641480
rect 510358 642330 510392 642364
rect 510358 642262 510392 642296
rect 510358 642194 510392 642228
rect 510358 642126 510392 642160
rect 510358 642058 510392 642092
rect 510358 641990 510392 642024
rect 510358 641922 510392 641956
rect 510358 641854 510392 641888
rect 510358 641786 510392 641820
rect 510358 641718 510392 641752
rect 510358 641650 510392 641684
rect 510358 641582 510392 641616
rect 510358 641514 510392 641548
rect 510358 641446 510392 641480
rect 510816 642330 510850 642364
rect 510816 642262 510850 642296
rect 510816 642194 510850 642228
rect 510816 642126 510850 642160
rect 510816 642058 510850 642092
rect 510816 641990 510850 642024
rect 510816 641922 510850 641956
rect 510816 641854 510850 641888
rect 510816 641786 510850 641820
rect 510816 641718 510850 641752
rect 510816 641650 510850 641684
rect 510816 641582 510850 641616
rect 510816 641514 510850 641548
rect 510816 641446 510850 641480
rect 511274 642330 511308 642364
rect 511274 642262 511308 642296
rect 511274 642194 511308 642228
rect 511274 642126 511308 642160
rect 511274 642058 511308 642092
rect 511274 641990 511308 642024
rect 511274 641922 511308 641956
rect 511274 641854 511308 641888
rect 511274 641786 511308 641820
rect 511274 641718 511308 641752
rect 511274 641650 511308 641684
rect 511274 641582 511308 641616
rect 511274 641514 511308 641548
rect 511274 641446 511308 641480
rect 511732 642330 511766 642364
rect 511732 642262 511766 642296
rect 511732 642194 511766 642228
rect 511732 642126 511766 642160
rect 511732 642058 511766 642092
rect 511732 641990 511766 642024
rect 511732 641922 511766 641956
rect 511732 641854 511766 641888
rect 511732 641786 511766 641820
rect 511732 641718 511766 641752
rect 511732 641650 511766 641684
rect 511732 641582 511766 641616
rect 511732 641514 511766 641548
rect 511732 641446 511766 641480
rect 512190 642330 512224 642364
rect 512190 642262 512224 642296
rect 512190 642194 512224 642228
rect 512190 642126 512224 642160
rect 512190 642058 512224 642092
rect 512190 641990 512224 642024
rect 512190 641922 512224 641956
rect 512190 641854 512224 641888
rect 512190 641786 512224 641820
rect 512190 641718 512224 641752
rect 512190 641650 512224 641684
rect 512190 641582 512224 641616
rect 512190 641514 512224 641548
rect 512190 641446 512224 641480
rect 512648 642330 512682 642364
rect 512648 642262 512682 642296
rect 512648 642194 512682 642228
rect 512648 642126 512682 642160
rect 512648 642058 512682 642092
rect 512648 641990 512682 642024
rect 512648 641922 512682 641956
rect 512648 641854 512682 641888
rect 512648 641786 512682 641820
rect 512648 641718 512682 641752
rect 512648 641650 512682 641684
rect 512648 641582 512682 641616
rect 512648 641514 512682 641548
rect 512648 641446 512682 641480
rect 513106 642330 513140 642364
rect 513106 642262 513140 642296
rect 513106 642194 513140 642228
rect 513106 642126 513140 642160
rect 513106 642058 513140 642092
rect 513106 641990 513140 642024
rect 513106 641922 513140 641956
rect 513106 641854 513140 641888
rect 513106 641786 513140 641820
rect 513106 641718 513140 641752
rect 513106 641650 513140 641684
rect 513106 641582 513140 641616
rect 513106 641514 513140 641548
rect 513106 641446 513140 641480
rect 513564 642330 513598 642364
rect 513564 642262 513598 642296
rect 513564 642194 513598 642228
rect 513564 642126 513598 642160
rect 513564 642058 513598 642092
rect 513564 641990 513598 642024
rect 513564 641922 513598 641956
rect 513564 641854 513598 641888
rect 513564 641786 513598 641820
rect 513564 641718 513598 641752
rect 513564 641650 513598 641684
rect 513564 641582 513598 641616
rect 513564 641514 513598 641548
rect 513564 641446 513598 641480
rect 514022 642330 514056 642364
rect 514022 642262 514056 642296
rect 514022 642194 514056 642228
rect 514022 642126 514056 642160
rect 514022 642058 514056 642092
rect 514022 641990 514056 642024
rect 514022 641922 514056 641956
rect 514022 641854 514056 641888
rect 514022 641786 514056 641820
rect 514022 641718 514056 641752
rect 514022 641650 514056 641684
rect 514022 641582 514056 641616
rect 514022 641514 514056 641548
rect 514022 641446 514056 641480
rect 514480 642330 514514 642364
rect 514480 642262 514514 642296
rect 514480 642194 514514 642228
rect 514480 642126 514514 642160
rect 514480 642058 514514 642092
rect 514480 641990 514514 642024
rect 514480 641922 514514 641956
rect 514480 641854 514514 641888
rect 514480 641786 514514 641820
rect 514480 641718 514514 641752
rect 514480 641650 514514 641684
rect 514480 641582 514514 641616
rect 514480 641514 514514 641548
rect 514480 641446 514514 641480
rect 514938 642330 514972 642364
rect 514938 642262 514972 642296
rect 514938 642194 514972 642228
rect 514938 642126 514972 642160
rect 514938 642058 514972 642092
rect 514938 641990 514972 642024
rect 514938 641922 514972 641956
rect 514938 641854 514972 641888
rect 514938 641786 514972 641820
rect 514938 641718 514972 641752
rect 514938 641650 514972 641684
rect 514938 641582 514972 641616
rect 514938 641514 514972 641548
rect 514938 641446 514972 641480
rect 515396 642330 515430 642364
rect 515396 642262 515430 642296
rect 515396 642194 515430 642228
rect 515396 642126 515430 642160
rect 515396 642058 515430 642092
rect 515396 641990 515430 642024
rect 515396 641922 515430 641956
rect 515396 641854 515430 641888
rect 515396 641786 515430 641820
rect 515396 641718 515430 641752
rect 515396 641650 515430 641684
rect 515396 641582 515430 641616
rect 515396 641514 515430 641548
rect 515396 641446 515430 641480
rect 508068 641168 508102 641202
rect 508068 641100 508102 641134
rect 508068 641032 508102 641066
rect 508068 640964 508102 640998
rect 508068 640896 508102 640930
rect 508068 640828 508102 640862
rect 508068 640760 508102 640794
rect 508068 640692 508102 640726
rect 508068 640624 508102 640658
rect 508068 640556 508102 640590
rect 508068 640488 508102 640522
rect 508068 640420 508102 640454
rect 508068 640352 508102 640386
rect 508068 640284 508102 640318
rect 508526 641168 508560 641202
rect 508526 641100 508560 641134
rect 508526 641032 508560 641066
rect 508526 640964 508560 640998
rect 508526 640896 508560 640930
rect 508526 640828 508560 640862
rect 508526 640760 508560 640794
rect 508526 640692 508560 640726
rect 508526 640624 508560 640658
rect 508526 640556 508560 640590
rect 508526 640488 508560 640522
rect 508526 640420 508560 640454
rect 508526 640352 508560 640386
rect 508526 640284 508560 640318
rect 508984 641168 509018 641202
rect 508984 641100 509018 641134
rect 508984 641032 509018 641066
rect 508984 640964 509018 640998
rect 508984 640896 509018 640930
rect 508984 640828 509018 640862
rect 508984 640760 509018 640794
rect 508984 640692 509018 640726
rect 508984 640624 509018 640658
rect 508984 640556 509018 640590
rect 508984 640488 509018 640522
rect 508984 640420 509018 640454
rect 508984 640352 509018 640386
rect 508984 640284 509018 640318
rect 509442 641168 509476 641202
rect 509442 641100 509476 641134
rect 509442 641032 509476 641066
rect 509442 640964 509476 640998
rect 509442 640896 509476 640930
rect 509442 640828 509476 640862
rect 509442 640760 509476 640794
rect 509442 640692 509476 640726
rect 509442 640624 509476 640658
rect 509442 640556 509476 640590
rect 509442 640488 509476 640522
rect 509442 640420 509476 640454
rect 509442 640352 509476 640386
rect 509442 640284 509476 640318
rect 509900 641168 509934 641202
rect 509900 641100 509934 641134
rect 509900 641032 509934 641066
rect 509900 640964 509934 640998
rect 509900 640896 509934 640930
rect 509900 640828 509934 640862
rect 509900 640760 509934 640794
rect 509900 640692 509934 640726
rect 509900 640624 509934 640658
rect 509900 640556 509934 640590
rect 509900 640488 509934 640522
rect 509900 640420 509934 640454
rect 509900 640352 509934 640386
rect 509900 640284 509934 640318
rect 510358 641168 510392 641202
rect 510358 641100 510392 641134
rect 510358 641032 510392 641066
rect 510358 640964 510392 640998
rect 510358 640896 510392 640930
rect 510358 640828 510392 640862
rect 510358 640760 510392 640794
rect 510358 640692 510392 640726
rect 510358 640624 510392 640658
rect 510358 640556 510392 640590
rect 510358 640488 510392 640522
rect 510358 640420 510392 640454
rect 510358 640352 510392 640386
rect 510358 640284 510392 640318
rect 510816 641168 510850 641202
rect 510816 641100 510850 641134
rect 510816 641032 510850 641066
rect 510816 640964 510850 640998
rect 510816 640896 510850 640930
rect 510816 640828 510850 640862
rect 510816 640760 510850 640794
rect 510816 640692 510850 640726
rect 510816 640624 510850 640658
rect 510816 640556 510850 640590
rect 510816 640488 510850 640522
rect 510816 640420 510850 640454
rect 510816 640352 510850 640386
rect 510816 640284 510850 640318
rect 511274 641168 511308 641202
rect 511274 641100 511308 641134
rect 511274 641032 511308 641066
rect 511274 640964 511308 640998
rect 511274 640896 511308 640930
rect 511274 640828 511308 640862
rect 511274 640760 511308 640794
rect 511274 640692 511308 640726
rect 511274 640624 511308 640658
rect 511274 640556 511308 640590
rect 511274 640488 511308 640522
rect 511274 640420 511308 640454
rect 511274 640352 511308 640386
rect 511274 640284 511308 640318
rect 511732 641168 511766 641202
rect 511732 641100 511766 641134
rect 511732 641032 511766 641066
rect 511732 640964 511766 640998
rect 511732 640896 511766 640930
rect 511732 640828 511766 640862
rect 511732 640760 511766 640794
rect 511732 640692 511766 640726
rect 511732 640624 511766 640658
rect 511732 640556 511766 640590
rect 511732 640488 511766 640522
rect 511732 640420 511766 640454
rect 511732 640352 511766 640386
rect 511732 640284 511766 640318
rect 512190 641168 512224 641202
rect 512190 641100 512224 641134
rect 512190 641032 512224 641066
rect 512190 640964 512224 640998
rect 512190 640896 512224 640930
rect 512190 640828 512224 640862
rect 512190 640760 512224 640794
rect 512190 640692 512224 640726
rect 512190 640624 512224 640658
rect 512190 640556 512224 640590
rect 512190 640488 512224 640522
rect 512190 640420 512224 640454
rect 512190 640352 512224 640386
rect 512190 640284 512224 640318
rect 512648 641168 512682 641202
rect 512648 641100 512682 641134
rect 512648 641032 512682 641066
rect 512648 640964 512682 640998
rect 512648 640896 512682 640930
rect 512648 640828 512682 640862
rect 512648 640760 512682 640794
rect 512648 640692 512682 640726
rect 512648 640624 512682 640658
rect 512648 640556 512682 640590
rect 512648 640488 512682 640522
rect 512648 640420 512682 640454
rect 512648 640352 512682 640386
rect 512648 640284 512682 640318
rect 513106 641168 513140 641202
rect 513106 641100 513140 641134
rect 513106 641032 513140 641066
rect 513106 640964 513140 640998
rect 513106 640896 513140 640930
rect 513106 640828 513140 640862
rect 513106 640760 513140 640794
rect 513106 640692 513140 640726
rect 513106 640624 513140 640658
rect 513106 640556 513140 640590
rect 513106 640488 513140 640522
rect 513106 640420 513140 640454
rect 513106 640352 513140 640386
rect 513106 640284 513140 640318
rect 513564 641168 513598 641202
rect 513564 641100 513598 641134
rect 513564 641032 513598 641066
rect 513564 640964 513598 640998
rect 513564 640896 513598 640930
rect 513564 640828 513598 640862
rect 513564 640760 513598 640794
rect 513564 640692 513598 640726
rect 513564 640624 513598 640658
rect 513564 640556 513598 640590
rect 513564 640488 513598 640522
rect 513564 640420 513598 640454
rect 513564 640352 513598 640386
rect 513564 640284 513598 640318
rect 514022 641168 514056 641202
rect 514022 641100 514056 641134
rect 514022 641032 514056 641066
rect 514022 640964 514056 640998
rect 514022 640896 514056 640930
rect 514022 640828 514056 640862
rect 514022 640760 514056 640794
rect 514022 640692 514056 640726
rect 514022 640624 514056 640658
rect 514022 640556 514056 640590
rect 514022 640488 514056 640522
rect 514022 640420 514056 640454
rect 514022 640352 514056 640386
rect 514022 640284 514056 640318
rect 514480 641168 514514 641202
rect 514480 641100 514514 641134
rect 514480 641032 514514 641066
rect 514480 640964 514514 640998
rect 514480 640896 514514 640930
rect 514480 640828 514514 640862
rect 514480 640760 514514 640794
rect 514480 640692 514514 640726
rect 514480 640624 514514 640658
rect 514480 640556 514514 640590
rect 514480 640488 514514 640522
rect 514480 640420 514514 640454
rect 514480 640352 514514 640386
rect 514480 640284 514514 640318
rect 514938 641168 514972 641202
rect 514938 641100 514972 641134
rect 514938 641032 514972 641066
rect 514938 640964 514972 640998
rect 514938 640896 514972 640930
rect 514938 640828 514972 640862
rect 514938 640760 514972 640794
rect 514938 640692 514972 640726
rect 514938 640624 514972 640658
rect 514938 640556 514972 640590
rect 514938 640488 514972 640522
rect 514938 640420 514972 640454
rect 514938 640352 514972 640386
rect 514938 640284 514972 640318
rect 515396 641168 515430 641202
rect 515396 641100 515430 641134
rect 515396 641032 515430 641066
rect 515396 640964 515430 640998
rect 515396 640896 515430 640930
rect 515396 640828 515430 640862
rect 515396 640760 515430 640794
rect 515396 640692 515430 640726
rect 515396 640624 515430 640658
rect 515396 640556 515430 640590
rect 515396 640488 515430 640522
rect 515396 640420 515430 640454
rect 515396 640352 515430 640386
rect 515396 640284 515430 640318
rect 515772 642330 515806 642364
rect 515772 642262 515806 642296
rect 515772 642194 515806 642228
rect 515772 642126 515806 642160
rect 515772 642058 515806 642092
rect 515772 641990 515806 642024
rect 515772 641922 515806 641956
rect 515772 641854 515806 641888
rect 515772 641786 515806 641820
rect 515772 641718 515806 641752
rect 515772 641650 515806 641684
rect 515772 641582 515806 641616
rect 515772 641514 515806 641548
rect 515772 641446 515806 641480
rect 516230 642330 516264 642364
rect 516230 642262 516264 642296
rect 516230 642194 516264 642228
rect 516230 642126 516264 642160
rect 516230 642058 516264 642092
rect 516230 641990 516264 642024
rect 516230 641922 516264 641956
rect 516230 641854 516264 641888
rect 516230 641786 516264 641820
rect 516230 641718 516264 641752
rect 516230 641650 516264 641684
rect 516230 641582 516264 641616
rect 516230 641514 516264 641548
rect 516230 641446 516264 641480
rect 516688 642330 516722 642364
rect 516688 642262 516722 642296
rect 516688 642194 516722 642228
rect 516688 642126 516722 642160
rect 516688 642058 516722 642092
rect 516688 641990 516722 642024
rect 516688 641922 516722 641956
rect 516688 641854 516722 641888
rect 516688 641786 516722 641820
rect 516688 641718 516722 641752
rect 516688 641650 516722 641684
rect 516688 641582 516722 641616
rect 516688 641514 516722 641548
rect 516688 641446 516722 641480
<< mvpdiffc >>
rect 508068 645428 508102 645462
rect 508068 645360 508102 645394
rect 508068 645292 508102 645326
rect 508068 645224 508102 645258
rect 508068 645156 508102 645190
rect 508068 645088 508102 645122
rect 508068 645020 508102 645054
rect 508068 644952 508102 644986
rect 508068 644884 508102 644918
rect 508068 644816 508102 644850
rect 508068 644748 508102 644782
rect 508068 644680 508102 644714
rect 508068 644612 508102 644646
rect 508068 644544 508102 644578
rect 508526 645428 508560 645462
rect 508526 645360 508560 645394
rect 508526 645292 508560 645326
rect 508526 645224 508560 645258
rect 508526 645156 508560 645190
rect 508526 645088 508560 645122
rect 508526 645020 508560 645054
rect 508526 644952 508560 644986
rect 508526 644884 508560 644918
rect 508526 644816 508560 644850
rect 508526 644748 508560 644782
rect 508526 644680 508560 644714
rect 508526 644612 508560 644646
rect 508526 644544 508560 644578
rect 508984 645428 509018 645462
rect 508984 645360 509018 645394
rect 508984 645292 509018 645326
rect 508984 645224 509018 645258
rect 508984 645156 509018 645190
rect 508984 645088 509018 645122
rect 508984 645020 509018 645054
rect 508984 644952 509018 644986
rect 508984 644884 509018 644918
rect 508984 644816 509018 644850
rect 508984 644748 509018 644782
rect 508984 644680 509018 644714
rect 508984 644612 509018 644646
rect 508984 644544 509018 644578
rect 509442 645428 509476 645462
rect 509442 645360 509476 645394
rect 509442 645292 509476 645326
rect 509442 645224 509476 645258
rect 509442 645156 509476 645190
rect 509442 645088 509476 645122
rect 509442 645020 509476 645054
rect 509442 644952 509476 644986
rect 509442 644884 509476 644918
rect 509442 644816 509476 644850
rect 509442 644748 509476 644782
rect 509442 644680 509476 644714
rect 509442 644612 509476 644646
rect 509442 644544 509476 644578
rect 509900 645428 509934 645462
rect 509900 645360 509934 645394
rect 509900 645292 509934 645326
rect 509900 645224 509934 645258
rect 509900 645156 509934 645190
rect 509900 645088 509934 645122
rect 509900 645020 509934 645054
rect 509900 644952 509934 644986
rect 509900 644884 509934 644918
rect 509900 644816 509934 644850
rect 509900 644748 509934 644782
rect 509900 644680 509934 644714
rect 509900 644612 509934 644646
rect 509900 644544 509934 644578
rect 510358 645428 510392 645462
rect 510358 645360 510392 645394
rect 510358 645292 510392 645326
rect 510358 645224 510392 645258
rect 510358 645156 510392 645190
rect 510358 645088 510392 645122
rect 510358 645020 510392 645054
rect 510358 644952 510392 644986
rect 510358 644884 510392 644918
rect 510358 644816 510392 644850
rect 510358 644748 510392 644782
rect 510358 644680 510392 644714
rect 510358 644612 510392 644646
rect 510358 644544 510392 644578
rect 510816 645428 510850 645462
rect 510816 645360 510850 645394
rect 510816 645292 510850 645326
rect 510816 645224 510850 645258
rect 510816 645156 510850 645190
rect 510816 645088 510850 645122
rect 510816 645020 510850 645054
rect 510816 644952 510850 644986
rect 510816 644884 510850 644918
rect 510816 644816 510850 644850
rect 510816 644748 510850 644782
rect 510816 644680 510850 644714
rect 510816 644612 510850 644646
rect 510816 644544 510850 644578
rect 511274 645428 511308 645462
rect 511274 645360 511308 645394
rect 511274 645292 511308 645326
rect 511274 645224 511308 645258
rect 511274 645156 511308 645190
rect 511274 645088 511308 645122
rect 511274 645020 511308 645054
rect 511274 644952 511308 644986
rect 511274 644884 511308 644918
rect 511274 644816 511308 644850
rect 511274 644748 511308 644782
rect 511274 644680 511308 644714
rect 511274 644612 511308 644646
rect 511274 644544 511308 644578
rect 511732 645428 511766 645462
rect 511732 645360 511766 645394
rect 511732 645292 511766 645326
rect 511732 645224 511766 645258
rect 511732 645156 511766 645190
rect 511732 645088 511766 645122
rect 511732 645020 511766 645054
rect 511732 644952 511766 644986
rect 511732 644884 511766 644918
rect 511732 644816 511766 644850
rect 511732 644748 511766 644782
rect 511732 644680 511766 644714
rect 511732 644612 511766 644646
rect 511732 644544 511766 644578
rect 512190 645428 512224 645462
rect 512190 645360 512224 645394
rect 512190 645292 512224 645326
rect 512190 645224 512224 645258
rect 512190 645156 512224 645190
rect 512190 645088 512224 645122
rect 512190 645020 512224 645054
rect 512190 644952 512224 644986
rect 512190 644884 512224 644918
rect 512190 644816 512224 644850
rect 512190 644748 512224 644782
rect 512190 644680 512224 644714
rect 512190 644612 512224 644646
rect 512190 644544 512224 644578
rect 512648 645428 512682 645462
rect 512648 645360 512682 645394
rect 512648 645292 512682 645326
rect 512648 645224 512682 645258
rect 512648 645156 512682 645190
rect 512648 645088 512682 645122
rect 512648 645020 512682 645054
rect 512648 644952 512682 644986
rect 512648 644884 512682 644918
rect 512648 644816 512682 644850
rect 512648 644748 512682 644782
rect 512648 644680 512682 644714
rect 512648 644612 512682 644646
rect 512648 644544 512682 644578
rect 513106 645428 513140 645462
rect 513106 645360 513140 645394
rect 513106 645292 513140 645326
rect 513106 645224 513140 645258
rect 513106 645156 513140 645190
rect 513106 645088 513140 645122
rect 513106 645020 513140 645054
rect 513106 644952 513140 644986
rect 513106 644884 513140 644918
rect 513106 644816 513140 644850
rect 513106 644748 513140 644782
rect 513106 644680 513140 644714
rect 513106 644612 513140 644646
rect 513106 644544 513140 644578
rect 513564 645428 513598 645462
rect 513564 645360 513598 645394
rect 513564 645292 513598 645326
rect 513564 645224 513598 645258
rect 513564 645156 513598 645190
rect 513564 645088 513598 645122
rect 513564 645020 513598 645054
rect 513564 644952 513598 644986
rect 513564 644884 513598 644918
rect 513564 644816 513598 644850
rect 513564 644748 513598 644782
rect 513564 644680 513598 644714
rect 513564 644612 513598 644646
rect 513564 644544 513598 644578
rect 514022 645428 514056 645462
rect 514022 645360 514056 645394
rect 514022 645292 514056 645326
rect 514022 645224 514056 645258
rect 514022 645156 514056 645190
rect 514022 645088 514056 645122
rect 514022 645020 514056 645054
rect 514022 644952 514056 644986
rect 514022 644884 514056 644918
rect 514022 644816 514056 644850
rect 514022 644748 514056 644782
rect 514022 644680 514056 644714
rect 514022 644612 514056 644646
rect 514022 644544 514056 644578
rect 514480 645428 514514 645462
rect 514480 645360 514514 645394
rect 514480 645292 514514 645326
rect 514480 645224 514514 645258
rect 514480 645156 514514 645190
rect 514480 645088 514514 645122
rect 514480 645020 514514 645054
rect 514480 644952 514514 644986
rect 514480 644884 514514 644918
rect 514480 644816 514514 644850
rect 514480 644748 514514 644782
rect 514480 644680 514514 644714
rect 514480 644612 514514 644646
rect 514480 644544 514514 644578
rect 514938 645428 514972 645462
rect 514938 645360 514972 645394
rect 514938 645292 514972 645326
rect 514938 645224 514972 645258
rect 514938 645156 514972 645190
rect 514938 645088 514972 645122
rect 514938 645020 514972 645054
rect 514938 644952 514972 644986
rect 514938 644884 514972 644918
rect 514938 644816 514972 644850
rect 514938 644748 514972 644782
rect 514938 644680 514972 644714
rect 514938 644612 514972 644646
rect 514938 644544 514972 644578
rect 515396 645428 515430 645462
rect 515396 645360 515430 645394
rect 515396 645292 515430 645326
rect 515396 645224 515430 645258
rect 515396 645156 515430 645190
rect 515396 645088 515430 645122
rect 515396 645020 515430 645054
rect 515396 644952 515430 644986
rect 515396 644884 515430 644918
rect 515396 644816 515430 644850
rect 515396 644748 515430 644782
rect 515396 644680 515430 644714
rect 515396 644612 515430 644646
rect 515396 644544 515430 644578
rect 508068 644262 508102 644296
rect 508068 644194 508102 644228
rect 508068 644126 508102 644160
rect 508068 644058 508102 644092
rect 508068 643990 508102 644024
rect 508068 643922 508102 643956
rect 508068 643854 508102 643888
rect 508068 643786 508102 643820
rect 508068 643718 508102 643752
rect 508068 643650 508102 643684
rect 508068 643582 508102 643616
rect 508068 643514 508102 643548
rect 508068 643446 508102 643480
rect 508068 643378 508102 643412
rect 508526 644262 508560 644296
rect 508526 644194 508560 644228
rect 508526 644126 508560 644160
rect 508526 644058 508560 644092
rect 508526 643990 508560 644024
rect 508526 643922 508560 643956
rect 508526 643854 508560 643888
rect 508526 643786 508560 643820
rect 508526 643718 508560 643752
rect 508526 643650 508560 643684
rect 508526 643582 508560 643616
rect 508526 643514 508560 643548
rect 508526 643446 508560 643480
rect 508526 643378 508560 643412
rect 508984 644262 509018 644296
rect 508984 644194 509018 644228
rect 508984 644126 509018 644160
rect 508984 644058 509018 644092
rect 508984 643990 509018 644024
rect 508984 643922 509018 643956
rect 508984 643854 509018 643888
rect 508984 643786 509018 643820
rect 508984 643718 509018 643752
rect 508984 643650 509018 643684
rect 508984 643582 509018 643616
rect 508984 643514 509018 643548
rect 508984 643446 509018 643480
rect 508984 643378 509018 643412
rect 509442 644262 509476 644296
rect 509442 644194 509476 644228
rect 509442 644126 509476 644160
rect 509442 644058 509476 644092
rect 509442 643990 509476 644024
rect 509442 643922 509476 643956
rect 509442 643854 509476 643888
rect 509442 643786 509476 643820
rect 509442 643718 509476 643752
rect 509442 643650 509476 643684
rect 509442 643582 509476 643616
rect 509442 643514 509476 643548
rect 509442 643446 509476 643480
rect 509442 643378 509476 643412
rect 509900 644262 509934 644296
rect 509900 644194 509934 644228
rect 509900 644126 509934 644160
rect 509900 644058 509934 644092
rect 509900 643990 509934 644024
rect 509900 643922 509934 643956
rect 509900 643854 509934 643888
rect 509900 643786 509934 643820
rect 509900 643718 509934 643752
rect 509900 643650 509934 643684
rect 509900 643582 509934 643616
rect 509900 643514 509934 643548
rect 509900 643446 509934 643480
rect 509900 643378 509934 643412
rect 510358 644262 510392 644296
rect 510358 644194 510392 644228
rect 510358 644126 510392 644160
rect 510358 644058 510392 644092
rect 510358 643990 510392 644024
rect 510358 643922 510392 643956
rect 510358 643854 510392 643888
rect 510358 643786 510392 643820
rect 510358 643718 510392 643752
rect 510358 643650 510392 643684
rect 510358 643582 510392 643616
rect 510358 643514 510392 643548
rect 510358 643446 510392 643480
rect 510358 643378 510392 643412
rect 510816 644262 510850 644296
rect 510816 644194 510850 644228
rect 510816 644126 510850 644160
rect 510816 644058 510850 644092
rect 510816 643990 510850 644024
rect 510816 643922 510850 643956
rect 510816 643854 510850 643888
rect 510816 643786 510850 643820
rect 510816 643718 510850 643752
rect 510816 643650 510850 643684
rect 510816 643582 510850 643616
rect 510816 643514 510850 643548
rect 510816 643446 510850 643480
rect 510816 643378 510850 643412
rect 511274 644262 511308 644296
rect 511274 644194 511308 644228
rect 511274 644126 511308 644160
rect 511274 644058 511308 644092
rect 511274 643990 511308 644024
rect 511274 643922 511308 643956
rect 511274 643854 511308 643888
rect 511274 643786 511308 643820
rect 511274 643718 511308 643752
rect 511274 643650 511308 643684
rect 511274 643582 511308 643616
rect 511274 643514 511308 643548
rect 511274 643446 511308 643480
rect 511274 643378 511308 643412
rect 511732 644262 511766 644296
rect 511732 644194 511766 644228
rect 511732 644126 511766 644160
rect 511732 644058 511766 644092
rect 511732 643990 511766 644024
rect 511732 643922 511766 643956
rect 511732 643854 511766 643888
rect 511732 643786 511766 643820
rect 511732 643718 511766 643752
rect 511732 643650 511766 643684
rect 511732 643582 511766 643616
rect 511732 643514 511766 643548
rect 511732 643446 511766 643480
rect 511732 643378 511766 643412
rect 512190 644262 512224 644296
rect 512190 644194 512224 644228
rect 512190 644126 512224 644160
rect 512190 644058 512224 644092
rect 512190 643990 512224 644024
rect 512190 643922 512224 643956
rect 512190 643854 512224 643888
rect 512190 643786 512224 643820
rect 512190 643718 512224 643752
rect 512190 643650 512224 643684
rect 512190 643582 512224 643616
rect 512190 643514 512224 643548
rect 512190 643446 512224 643480
rect 512190 643378 512224 643412
rect 512648 644262 512682 644296
rect 512648 644194 512682 644228
rect 512648 644126 512682 644160
rect 512648 644058 512682 644092
rect 512648 643990 512682 644024
rect 512648 643922 512682 643956
rect 512648 643854 512682 643888
rect 512648 643786 512682 643820
rect 512648 643718 512682 643752
rect 512648 643650 512682 643684
rect 512648 643582 512682 643616
rect 512648 643514 512682 643548
rect 512648 643446 512682 643480
rect 512648 643378 512682 643412
rect 513106 644262 513140 644296
rect 513106 644194 513140 644228
rect 513106 644126 513140 644160
rect 513106 644058 513140 644092
rect 513106 643990 513140 644024
rect 513106 643922 513140 643956
rect 513106 643854 513140 643888
rect 513106 643786 513140 643820
rect 513106 643718 513140 643752
rect 513106 643650 513140 643684
rect 513106 643582 513140 643616
rect 513106 643514 513140 643548
rect 513106 643446 513140 643480
rect 513106 643378 513140 643412
rect 513564 644262 513598 644296
rect 513564 644194 513598 644228
rect 513564 644126 513598 644160
rect 513564 644058 513598 644092
rect 513564 643990 513598 644024
rect 513564 643922 513598 643956
rect 513564 643854 513598 643888
rect 513564 643786 513598 643820
rect 513564 643718 513598 643752
rect 513564 643650 513598 643684
rect 513564 643582 513598 643616
rect 513564 643514 513598 643548
rect 513564 643446 513598 643480
rect 513564 643378 513598 643412
rect 514022 644262 514056 644296
rect 514022 644194 514056 644228
rect 514022 644126 514056 644160
rect 514022 644058 514056 644092
rect 514022 643990 514056 644024
rect 514022 643922 514056 643956
rect 514022 643854 514056 643888
rect 514022 643786 514056 643820
rect 514022 643718 514056 643752
rect 514022 643650 514056 643684
rect 514022 643582 514056 643616
rect 514022 643514 514056 643548
rect 514022 643446 514056 643480
rect 514022 643378 514056 643412
rect 514480 644262 514514 644296
rect 514480 644194 514514 644228
rect 514480 644126 514514 644160
rect 514480 644058 514514 644092
rect 514480 643990 514514 644024
rect 514480 643922 514514 643956
rect 514480 643854 514514 643888
rect 514480 643786 514514 643820
rect 514480 643718 514514 643752
rect 514480 643650 514514 643684
rect 514480 643582 514514 643616
rect 514480 643514 514514 643548
rect 514480 643446 514514 643480
rect 514480 643378 514514 643412
rect 514938 644262 514972 644296
rect 514938 644194 514972 644228
rect 514938 644126 514972 644160
rect 514938 644058 514972 644092
rect 514938 643990 514972 644024
rect 514938 643922 514972 643956
rect 514938 643854 514972 643888
rect 514938 643786 514972 643820
rect 514938 643718 514972 643752
rect 514938 643650 514972 643684
rect 514938 643582 514972 643616
rect 514938 643514 514972 643548
rect 514938 643446 514972 643480
rect 514938 643378 514972 643412
rect 515396 644262 515430 644296
rect 515396 644194 515430 644228
rect 515396 644126 515430 644160
rect 515396 644058 515430 644092
rect 515396 643990 515430 644024
rect 515396 643922 515430 643956
rect 515396 643854 515430 643888
rect 515396 643786 515430 643820
rect 515396 643718 515430 643752
rect 515396 643650 515430 643684
rect 515396 643582 515430 643616
rect 515396 643514 515430 643548
rect 515396 643446 515430 643480
rect 515396 643378 515430 643412
rect 515772 645272 515806 645306
rect 515772 645204 515806 645238
rect 515772 645136 515806 645170
rect 515772 645068 515806 645102
rect 515772 645000 515806 645034
rect 515772 644932 515806 644966
rect 515772 644864 515806 644898
rect 515772 644796 515806 644830
rect 515772 644728 515806 644762
rect 515772 644660 515806 644694
rect 515772 644592 515806 644626
rect 515772 644524 515806 644558
rect 515772 644456 515806 644490
rect 515772 644388 515806 644422
rect 515772 644320 515806 644354
rect 515772 644252 515806 644286
rect 515772 644184 515806 644218
rect 515772 644116 515806 644150
rect 515772 644048 515806 644082
rect 515772 643980 515806 644014
rect 515772 643912 515806 643946
rect 515772 643844 515806 643878
rect 515772 643776 515806 643810
rect 515772 643708 515806 643742
rect 515772 643640 515806 643674
rect 515772 643572 515806 643606
rect 515772 643504 515806 643538
rect 515772 643436 515806 643470
rect 515772 643368 515806 643402
rect 516230 645272 516264 645306
rect 516230 645204 516264 645238
rect 516230 645136 516264 645170
rect 516230 645068 516264 645102
rect 516230 645000 516264 645034
rect 516230 644932 516264 644966
rect 516230 644864 516264 644898
rect 516230 644796 516264 644830
rect 516230 644728 516264 644762
rect 516230 644660 516264 644694
rect 516230 644592 516264 644626
rect 516230 644524 516264 644558
rect 516230 644456 516264 644490
rect 516230 644388 516264 644422
rect 516230 644320 516264 644354
rect 516230 644252 516264 644286
rect 516230 644184 516264 644218
rect 516230 644116 516264 644150
rect 516230 644048 516264 644082
rect 516230 643980 516264 644014
rect 516230 643912 516264 643946
rect 516230 643844 516264 643878
rect 516230 643776 516264 643810
rect 516230 643708 516264 643742
rect 516230 643640 516264 643674
rect 516230 643572 516264 643606
rect 516230 643504 516264 643538
rect 516230 643436 516264 643470
rect 516230 643368 516264 643402
rect 516688 645272 516722 645306
rect 516688 645204 516722 645238
rect 516688 645136 516722 645170
rect 516688 645068 516722 645102
rect 516688 645000 516722 645034
rect 516688 644932 516722 644966
rect 516688 644864 516722 644898
rect 516688 644796 516722 644830
rect 516688 644728 516722 644762
rect 516688 644660 516722 644694
rect 516688 644592 516722 644626
rect 516688 644524 516722 644558
rect 516688 644456 516722 644490
rect 516688 644388 516722 644422
rect 516688 644320 516722 644354
rect 516688 644252 516722 644286
rect 516688 644184 516722 644218
rect 516688 644116 516722 644150
rect 516688 644048 516722 644082
rect 516688 643980 516722 644014
rect 516688 643912 516722 643946
rect 516688 643844 516722 643878
rect 516688 643776 516722 643810
rect 516688 643708 516722 643742
rect 516688 643640 516722 643674
rect 516688 643572 516722 643606
rect 516688 643504 516722 643538
rect 516688 643436 516722 643470
rect 516688 643368 516722 643402
<< mvpsubdiff >>
rect 507820 642702 516974 642728
rect 507820 642600 507846 642702
rect 507948 642600 507992 642702
rect 515506 642600 515550 642702
rect 515652 642600 515722 642702
rect 516776 642600 516846 642702
rect 516948 642600 516974 642702
rect 507820 642574 516974 642600
rect 507820 642528 507974 642574
rect 507820 640182 507846 642528
rect 507948 640182 507974 642528
rect 515524 642528 515678 642574
rect 507820 640136 507974 640182
rect 515524 640182 515550 642528
rect 515652 641288 515678 642528
rect 516820 642528 516974 642574
rect 516820 641288 516846 642528
rect 515652 641262 516846 641288
rect 515652 641160 515722 641262
rect 516776 641160 516846 641262
rect 515652 641094 516846 641160
rect 515652 640182 515722 641094
rect 515524 640176 515722 640182
rect 516776 640182 516846 641094
rect 516948 640182 516974 642528
rect 516776 640176 516974 640182
rect 515524 640136 516974 640176
rect 507820 640110 516974 640136
rect 507820 640008 507846 640110
rect 507948 640008 507994 640110
rect 516800 640008 516846 640110
rect 516948 640008 516974 640110
rect 507820 639982 516974 640008
<< mvnsubdiff >>
rect 507820 645725 516974 645751
rect 507820 645623 507846 645725
rect 507948 645623 507992 645725
rect 515506 645623 515550 645725
rect 515652 645623 515722 645725
rect 516776 645623 516846 645725
rect 516948 645623 516974 645725
rect 507820 645597 516974 645623
rect 507820 645551 507974 645597
rect 507820 643205 507846 645551
rect 507948 643205 507974 645551
rect 515524 645581 516974 645597
rect 515524 645551 515722 645581
rect 507820 643159 507974 643205
rect 515524 643205 515550 645551
rect 515652 645479 515722 645551
rect 516776 645551 516974 645581
rect 516776 645479 516846 645551
rect 515652 645453 516846 645479
rect 515652 643205 515678 645453
rect 515524 643159 515678 643205
rect 516820 643205 516846 645453
rect 516948 643205 516974 645551
rect 516820 643159 516974 643205
rect 507820 643133 516974 643159
rect 507820 643031 507846 643133
rect 507948 643031 507992 643133
rect 515506 643031 515550 643133
rect 515652 643031 515722 643133
rect 516776 643031 516846 643133
rect 516948 643031 516974 643133
rect 507820 643005 516974 643031
<< mvpsubdiffcont >>
rect 507846 642600 507948 642702
rect 507992 642600 515506 642702
rect 515550 642600 515652 642702
rect 515722 642600 516776 642702
rect 516846 642600 516948 642702
rect 507846 640182 507948 642528
rect 515550 640182 515652 642528
rect 515722 641160 516776 641262
rect 515722 640176 516776 641094
rect 516846 640182 516948 642528
rect 507846 640008 507948 640110
rect 507994 640008 516800 640110
rect 516846 640008 516948 640110
<< mvnsubdiffcont >>
rect 507846 645623 507948 645725
rect 507992 645623 515506 645725
rect 515550 645623 515652 645725
rect 515722 645623 516776 645725
rect 516846 645623 516948 645725
rect 507846 643205 507948 645551
rect 515550 643205 515652 645551
rect 515722 645479 516776 645581
rect 516846 643205 516948 645551
rect 507846 643031 507948 643133
rect 507992 643031 515506 643133
rect 515550 643031 515652 643133
rect 515722 643031 516776 643133
rect 516846 643031 516948 643133
<< poly >>
rect 508114 645503 508514 645529
rect 508572 645503 508972 645529
rect 509030 645503 509430 645529
rect 509488 645503 509888 645529
rect 509946 645503 510346 645529
rect 510404 645503 510804 645529
rect 510862 645503 511262 645529
rect 511320 645503 511720 645529
rect 511778 645503 512178 645529
rect 512236 645503 512636 645529
rect 512694 645503 513094 645529
rect 513152 645503 513552 645529
rect 513610 645503 514010 645529
rect 514068 645503 514468 645529
rect 514526 645503 514926 645529
rect 514984 645503 515384 645529
rect 508114 644456 508514 644503
rect 508114 644422 508161 644456
rect 508195 644422 508229 644456
rect 508263 644422 508297 644456
rect 508331 644422 508365 644456
rect 508399 644422 508433 644456
rect 508467 644422 508514 644456
rect 508114 644406 508514 644422
rect 508572 644456 508972 644503
rect 508572 644422 508619 644456
rect 508653 644422 508687 644456
rect 508721 644422 508755 644456
rect 508789 644422 508823 644456
rect 508857 644422 508891 644456
rect 508925 644422 508972 644456
rect 508572 644406 508972 644422
rect 509030 644456 509430 644503
rect 509030 644422 509077 644456
rect 509111 644422 509145 644456
rect 509179 644422 509213 644456
rect 509247 644422 509281 644456
rect 509315 644422 509349 644456
rect 509383 644422 509430 644456
rect 509030 644406 509430 644422
rect 509488 644456 509888 644503
rect 509488 644422 509535 644456
rect 509569 644422 509603 644456
rect 509637 644422 509671 644456
rect 509705 644422 509739 644456
rect 509773 644422 509807 644456
rect 509841 644422 509888 644456
rect 509488 644406 509888 644422
rect 509946 644456 510346 644503
rect 509946 644422 509993 644456
rect 510027 644422 510061 644456
rect 510095 644422 510129 644456
rect 510163 644422 510197 644456
rect 510231 644422 510265 644456
rect 510299 644422 510346 644456
rect 509946 644406 510346 644422
rect 510404 644456 510804 644503
rect 510404 644422 510451 644456
rect 510485 644422 510519 644456
rect 510553 644422 510587 644456
rect 510621 644422 510655 644456
rect 510689 644422 510723 644456
rect 510757 644422 510804 644456
rect 510404 644406 510804 644422
rect 510862 644456 511262 644503
rect 510862 644422 510909 644456
rect 510943 644422 510977 644456
rect 511011 644422 511045 644456
rect 511079 644422 511113 644456
rect 511147 644422 511181 644456
rect 511215 644422 511262 644456
rect 510862 644406 511262 644422
rect 511320 644456 511720 644503
rect 511320 644422 511367 644456
rect 511401 644422 511435 644456
rect 511469 644422 511503 644456
rect 511537 644422 511571 644456
rect 511605 644422 511639 644456
rect 511673 644422 511720 644456
rect 511320 644406 511720 644422
rect 511778 644456 512178 644503
rect 511778 644422 511825 644456
rect 511859 644422 511893 644456
rect 511927 644422 511961 644456
rect 511995 644422 512029 644456
rect 512063 644422 512097 644456
rect 512131 644422 512178 644456
rect 511778 644406 512178 644422
rect 512236 644456 512636 644503
rect 512236 644422 512283 644456
rect 512317 644422 512351 644456
rect 512385 644422 512419 644456
rect 512453 644422 512487 644456
rect 512521 644422 512555 644456
rect 512589 644422 512636 644456
rect 512236 644406 512636 644422
rect 512694 644456 513094 644503
rect 512694 644422 512741 644456
rect 512775 644422 512809 644456
rect 512843 644422 512877 644456
rect 512911 644422 512945 644456
rect 512979 644422 513013 644456
rect 513047 644422 513094 644456
rect 512694 644406 513094 644422
rect 513152 644456 513552 644503
rect 513152 644422 513199 644456
rect 513233 644422 513267 644456
rect 513301 644422 513335 644456
rect 513369 644422 513403 644456
rect 513437 644422 513471 644456
rect 513505 644422 513552 644456
rect 513152 644406 513552 644422
rect 513610 644456 514010 644503
rect 513610 644422 513657 644456
rect 513691 644422 513725 644456
rect 513759 644422 513793 644456
rect 513827 644422 513861 644456
rect 513895 644422 513929 644456
rect 513963 644422 514010 644456
rect 513610 644406 514010 644422
rect 514068 644456 514468 644503
rect 514068 644422 514115 644456
rect 514149 644422 514183 644456
rect 514217 644422 514251 644456
rect 514285 644422 514319 644456
rect 514353 644422 514387 644456
rect 514421 644422 514468 644456
rect 514068 644406 514468 644422
rect 514526 644456 514926 644503
rect 514526 644422 514573 644456
rect 514607 644422 514641 644456
rect 514675 644422 514709 644456
rect 514743 644422 514777 644456
rect 514811 644422 514845 644456
rect 514879 644422 514926 644456
rect 514526 644406 514926 644422
rect 514984 644456 515384 644503
rect 514984 644422 515031 644456
rect 515065 644422 515099 644456
rect 515133 644422 515167 644456
rect 515201 644422 515235 644456
rect 515269 644422 515303 644456
rect 515337 644422 515384 644456
rect 514984 644406 515384 644422
rect 508114 644337 508514 644363
rect 508572 644337 508972 644363
rect 509030 644337 509430 644363
rect 509488 644337 509888 644363
rect 509946 644337 510346 644363
rect 510404 644337 510804 644363
rect 510862 644337 511262 644363
rect 511320 644337 511720 644363
rect 511778 644337 512178 644363
rect 512236 644337 512636 644363
rect 512694 644337 513094 644363
rect 513152 644337 513552 644363
rect 513610 644337 514010 644363
rect 514068 644337 514468 644363
rect 514526 644337 514926 644363
rect 514984 644337 515384 644363
rect 508114 643290 508514 643337
rect 508114 643256 508161 643290
rect 508195 643256 508229 643290
rect 508263 643256 508297 643290
rect 508331 643256 508365 643290
rect 508399 643256 508433 643290
rect 508467 643256 508514 643290
rect 508114 643240 508514 643256
rect 508572 643290 508972 643337
rect 508572 643256 508619 643290
rect 508653 643256 508687 643290
rect 508721 643256 508755 643290
rect 508789 643256 508823 643290
rect 508857 643256 508891 643290
rect 508925 643256 508972 643290
rect 508572 643240 508972 643256
rect 509030 643290 509430 643337
rect 509030 643256 509077 643290
rect 509111 643256 509145 643290
rect 509179 643256 509213 643290
rect 509247 643256 509281 643290
rect 509315 643256 509349 643290
rect 509383 643256 509430 643290
rect 509030 643240 509430 643256
rect 509488 643290 509888 643337
rect 509488 643256 509535 643290
rect 509569 643256 509603 643290
rect 509637 643256 509671 643290
rect 509705 643256 509739 643290
rect 509773 643256 509807 643290
rect 509841 643256 509888 643290
rect 509488 643240 509888 643256
rect 509946 643290 510346 643337
rect 509946 643256 509993 643290
rect 510027 643256 510061 643290
rect 510095 643256 510129 643290
rect 510163 643256 510197 643290
rect 510231 643256 510265 643290
rect 510299 643256 510346 643290
rect 509946 643240 510346 643256
rect 510404 643290 510804 643337
rect 510404 643256 510451 643290
rect 510485 643256 510519 643290
rect 510553 643256 510587 643290
rect 510621 643256 510655 643290
rect 510689 643256 510723 643290
rect 510757 643256 510804 643290
rect 510404 643240 510804 643256
rect 510862 643290 511262 643337
rect 510862 643256 510909 643290
rect 510943 643256 510977 643290
rect 511011 643256 511045 643290
rect 511079 643256 511113 643290
rect 511147 643256 511181 643290
rect 511215 643256 511262 643290
rect 510862 643240 511262 643256
rect 511320 643290 511720 643337
rect 511320 643256 511367 643290
rect 511401 643256 511435 643290
rect 511469 643256 511503 643290
rect 511537 643256 511571 643290
rect 511605 643256 511639 643290
rect 511673 643256 511720 643290
rect 511320 643240 511720 643256
rect 511778 643290 512178 643337
rect 511778 643256 511825 643290
rect 511859 643256 511893 643290
rect 511927 643256 511961 643290
rect 511995 643256 512029 643290
rect 512063 643256 512097 643290
rect 512131 643256 512178 643290
rect 511778 643240 512178 643256
rect 512236 643290 512636 643337
rect 512236 643256 512283 643290
rect 512317 643256 512351 643290
rect 512385 643256 512419 643290
rect 512453 643256 512487 643290
rect 512521 643256 512555 643290
rect 512589 643256 512636 643290
rect 512236 643240 512636 643256
rect 512694 643290 513094 643337
rect 512694 643256 512741 643290
rect 512775 643256 512809 643290
rect 512843 643256 512877 643290
rect 512911 643256 512945 643290
rect 512979 643256 513013 643290
rect 513047 643256 513094 643290
rect 512694 643240 513094 643256
rect 513152 643290 513552 643337
rect 513152 643256 513199 643290
rect 513233 643256 513267 643290
rect 513301 643256 513335 643290
rect 513369 643256 513403 643290
rect 513437 643256 513471 643290
rect 513505 643256 513552 643290
rect 513152 643240 513552 643256
rect 513610 643290 514010 643337
rect 513610 643256 513657 643290
rect 513691 643256 513725 643290
rect 513759 643256 513793 643290
rect 513827 643256 513861 643290
rect 513895 643256 513929 643290
rect 513963 643256 514010 643290
rect 513610 643240 514010 643256
rect 514068 643290 514468 643337
rect 514068 643256 514115 643290
rect 514149 643256 514183 643290
rect 514217 643256 514251 643290
rect 514285 643256 514319 643290
rect 514353 643256 514387 643290
rect 514421 643256 514468 643290
rect 514068 643240 514468 643256
rect 514526 643290 514926 643337
rect 514526 643256 514573 643290
rect 514607 643256 514641 643290
rect 514675 643256 514709 643290
rect 514743 643256 514777 643290
rect 514811 643256 514845 643290
rect 514879 643256 514926 643290
rect 514526 643240 514926 643256
rect 514984 643290 515384 643337
rect 514984 643256 515031 643290
rect 515065 643256 515099 643290
rect 515133 643256 515167 643290
rect 515201 643256 515235 643290
rect 515269 643256 515303 643290
rect 515337 643256 515384 643290
rect 514984 643240 515384 643256
rect 515818 645337 516218 645363
rect 516276 645337 516676 645363
rect 515818 643290 516218 643337
rect 515818 643256 515865 643290
rect 515899 643256 515933 643290
rect 515967 643256 516001 643290
rect 516035 643256 516069 643290
rect 516103 643256 516137 643290
rect 516171 643256 516218 643290
rect 515818 643240 516218 643256
rect 516276 643290 516676 643337
rect 516276 643256 516323 643290
rect 516357 643256 516391 643290
rect 516425 643256 516459 643290
rect 516493 643256 516527 643290
rect 516561 643256 516595 643290
rect 516629 643256 516676 643290
rect 516276 643240 516676 643256
rect 508114 642477 508514 642493
rect 508114 642443 508161 642477
rect 508195 642443 508229 642477
rect 508263 642443 508297 642477
rect 508331 642443 508365 642477
rect 508399 642443 508433 642477
rect 508467 642443 508514 642477
rect 508114 642405 508514 642443
rect 508572 642477 508972 642493
rect 508572 642443 508619 642477
rect 508653 642443 508687 642477
rect 508721 642443 508755 642477
rect 508789 642443 508823 642477
rect 508857 642443 508891 642477
rect 508925 642443 508972 642477
rect 508572 642405 508972 642443
rect 509030 642477 509430 642493
rect 509030 642443 509077 642477
rect 509111 642443 509145 642477
rect 509179 642443 509213 642477
rect 509247 642443 509281 642477
rect 509315 642443 509349 642477
rect 509383 642443 509430 642477
rect 509030 642405 509430 642443
rect 509488 642477 509888 642493
rect 509488 642443 509535 642477
rect 509569 642443 509603 642477
rect 509637 642443 509671 642477
rect 509705 642443 509739 642477
rect 509773 642443 509807 642477
rect 509841 642443 509888 642477
rect 509488 642405 509888 642443
rect 509946 642477 510346 642493
rect 509946 642443 509993 642477
rect 510027 642443 510061 642477
rect 510095 642443 510129 642477
rect 510163 642443 510197 642477
rect 510231 642443 510265 642477
rect 510299 642443 510346 642477
rect 509946 642405 510346 642443
rect 510404 642477 510804 642493
rect 510404 642443 510451 642477
rect 510485 642443 510519 642477
rect 510553 642443 510587 642477
rect 510621 642443 510655 642477
rect 510689 642443 510723 642477
rect 510757 642443 510804 642477
rect 510404 642405 510804 642443
rect 510862 642477 511262 642493
rect 510862 642443 510909 642477
rect 510943 642443 510977 642477
rect 511011 642443 511045 642477
rect 511079 642443 511113 642477
rect 511147 642443 511181 642477
rect 511215 642443 511262 642477
rect 510862 642405 511262 642443
rect 511320 642477 511720 642493
rect 511320 642443 511367 642477
rect 511401 642443 511435 642477
rect 511469 642443 511503 642477
rect 511537 642443 511571 642477
rect 511605 642443 511639 642477
rect 511673 642443 511720 642477
rect 511320 642405 511720 642443
rect 511778 642477 512178 642493
rect 511778 642443 511825 642477
rect 511859 642443 511893 642477
rect 511927 642443 511961 642477
rect 511995 642443 512029 642477
rect 512063 642443 512097 642477
rect 512131 642443 512178 642477
rect 511778 642405 512178 642443
rect 512236 642477 512636 642493
rect 512236 642443 512283 642477
rect 512317 642443 512351 642477
rect 512385 642443 512419 642477
rect 512453 642443 512487 642477
rect 512521 642443 512555 642477
rect 512589 642443 512636 642477
rect 512236 642405 512636 642443
rect 512694 642477 513094 642493
rect 512694 642443 512741 642477
rect 512775 642443 512809 642477
rect 512843 642443 512877 642477
rect 512911 642443 512945 642477
rect 512979 642443 513013 642477
rect 513047 642443 513094 642477
rect 512694 642405 513094 642443
rect 513152 642477 513552 642493
rect 513152 642443 513199 642477
rect 513233 642443 513267 642477
rect 513301 642443 513335 642477
rect 513369 642443 513403 642477
rect 513437 642443 513471 642477
rect 513505 642443 513552 642477
rect 513152 642405 513552 642443
rect 513610 642477 514010 642493
rect 513610 642443 513657 642477
rect 513691 642443 513725 642477
rect 513759 642443 513793 642477
rect 513827 642443 513861 642477
rect 513895 642443 513929 642477
rect 513963 642443 514010 642477
rect 513610 642405 514010 642443
rect 514068 642477 514468 642493
rect 514068 642443 514115 642477
rect 514149 642443 514183 642477
rect 514217 642443 514251 642477
rect 514285 642443 514319 642477
rect 514353 642443 514387 642477
rect 514421 642443 514468 642477
rect 514068 642405 514468 642443
rect 514526 642477 514926 642493
rect 514526 642443 514573 642477
rect 514607 642443 514641 642477
rect 514675 642443 514709 642477
rect 514743 642443 514777 642477
rect 514811 642443 514845 642477
rect 514879 642443 514926 642477
rect 514526 642405 514926 642443
rect 514984 642477 515384 642493
rect 514984 642443 515031 642477
rect 515065 642443 515099 642477
rect 515133 642443 515167 642477
rect 515201 642443 515235 642477
rect 515269 642443 515303 642477
rect 515337 642443 515384 642477
rect 514984 642405 515384 642443
rect 508114 641379 508514 641405
rect 508572 641379 508972 641405
rect 509030 641379 509430 641405
rect 509488 641379 509888 641405
rect 509946 641379 510346 641405
rect 510404 641379 510804 641405
rect 510862 641379 511262 641405
rect 511320 641379 511720 641405
rect 511778 641379 512178 641405
rect 512236 641379 512636 641405
rect 512694 641379 513094 641405
rect 513152 641379 513552 641405
rect 513610 641379 514010 641405
rect 514068 641379 514468 641405
rect 514526 641379 514926 641405
rect 514984 641379 515384 641405
rect 508114 641315 508514 641331
rect 508114 641281 508161 641315
rect 508195 641281 508229 641315
rect 508263 641281 508297 641315
rect 508331 641281 508365 641315
rect 508399 641281 508433 641315
rect 508467 641281 508514 641315
rect 508114 641243 508514 641281
rect 508572 641315 508972 641331
rect 508572 641281 508619 641315
rect 508653 641281 508687 641315
rect 508721 641281 508755 641315
rect 508789 641281 508823 641315
rect 508857 641281 508891 641315
rect 508925 641281 508972 641315
rect 508572 641243 508972 641281
rect 509030 641315 509430 641331
rect 509030 641281 509077 641315
rect 509111 641281 509145 641315
rect 509179 641281 509213 641315
rect 509247 641281 509281 641315
rect 509315 641281 509349 641315
rect 509383 641281 509430 641315
rect 509030 641243 509430 641281
rect 509488 641315 509888 641331
rect 509488 641281 509535 641315
rect 509569 641281 509603 641315
rect 509637 641281 509671 641315
rect 509705 641281 509739 641315
rect 509773 641281 509807 641315
rect 509841 641281 509888 641315
rect 509488 641243 509888 641281
rect 509946 641315 510346 641331
rect 509946 641281 509993 641315
rect 510027 641281 510061 641315
rect 510095 641281 510129 641315
rect 510163 641281 510197 641315
rect 510231 641281 510265 641315
rect 510299 641281 510346 641315
rect 509946 641243 510346 641281
rect 510404 641315 510804 641331
rect 510404 641281 510451 641315
rect 510485 641281 510519 641315
rect 510553 641281 510587 641315
rect 510621 641281 510655 641315
rect 510689 641281 510723 641315
rect 510757 641281 510804 641315
rect 510404 641243 510804 641281
rect 510862 641315 511262 641331
rect 510862 641281 510909 641315
rect 510943 641281 510977 641315
rect 511011 641281 511045 641315
rect 511079 641281 511113 641315
rect 511147 641281 511181 641315
rect 511215 641281 511262 641315
rect 510862 641243 511262 641281
rect 511320 641315 511720 641331
rect 511320 641281 511367 641315
rect 511401 641281 511435 641315
rect 511469 641281 511503 641315
rect 511537 641281 511571 641315
rect 511605 641281 511639 641315
rect 511673 641281 511720 641315
rect 511320 641243 511720 641281
rect 511778 641315 512178 641331
rect 511778 641281 511825 641315
rect 511859 641281 511893 641315
rect 511927 641281 511961 641315
rect 511995 641281 512029 641315
rect 512063 641281 512097 641315
rect 512131 641281 512178 641315
rect 511778 641243 512178 641281
rect 512236 641315 512636 641331
rect 512236 641281 512283 641315
rect 512317 641281 512351 641315
rect 512385 641281 512419 641315
rect 512453 641281 512487 641315
rect 512521 641281 512555 641315
rect 512589 641281 512636 641315
rect 512236 641243 512636 641281
rect 512694 641315 513094 641331
rect 512694 641281 512741 641315
rect 512775 641281 512809 641315
rect 512843 641281 512877 641315
rect 512911 641281 512945 641315
rect 512979 641281 513013 641315
rect 513047 641281 513094 641315
rect 512694 641243 513094 641281
rect 513152 641315 513552 641331
rect 513152 641281 513199 641315
rect 513233 641281 513267 641315
rect 513301 641281 513335 641315
rect 513369 641281 513403 641315
rect 513437 641281 513471 641315
rect 513505 641281 513552 641315
rect 513152 641243 513552 641281
rect 513610 641315 514010 641331
rect 513610 641281 513657 641315
rect 513691 641281 513725 641315
rect 513759 641281 513793 641315
rect 513827 641281 513861 641315
rect 513895 641281 513929 641315
rect 513963 641281 514010 641315
rect 513610 641243 514010 641281
rect 514068 641315 514468 641331
rect 514068 641281 514115 641315
rect 514149 641281 514183 641315
rect 514217 641281 514251 641315
rect 514285 641281 514319 641315
rect 514353 641281 514387 641315
rect 514421 641281 514468 641315
rect 514068 641243 514468 641281
rect 514526 641315 514926 641331
rect 514526 641281 514573 641315
rect 514607 641281 514641 641315
rect 514675 641281 514709 641315
rect 514743 641281 514777 641315
rect 514811 641281 514845 641315
rect 514879 641281 514926 641315
rect 514526 641243 514926 641281
rect 514984 641315 515384 641331
rect 514984 641281 515031 641315
rect 515065 641281 515099 641315
rect 515133 641281 515167 641315
rect 515201 641281 515235 641315
rect 515269 641281 515303 641315
rect 515337 641281 515384 641315
rect 514984 641243 515384 641281
rect 508114 640217 508514 640243
rect 508572 640217 508972 640243
rect 509030 640217 509430 640243
rect 509488 640217 509888 640243
rect 509946 640217 510346 640243
rect 510404 640217 510804 640243
rect 510862 640217 511262 640243
rect 511320 640217 511720 640243
rect 511778 640217 512178 640243
rect 512236 640217 512636 640243
rect 512694 640217 513094 640243
rect 513152 640217 513552 640243
rect 513610 640217 514010 640243
rect 514068 640217 514468 640243
rect 514526 640217 514926 640243
rect 514984 640217 515384 640243
rect 515818 642477 516218 642493
rect 515818 642443 515865 642477
rect 515899 642443 515933 642477
rect 515967 642443 516001 642477
rect 516035 642443 516069 642477
rect 516103 642443 516137 642477
rect 516171 642443 516218 642477
rect 515818 642405 516218 642443
rect 516276 642477 516676 642493
rect 516276 642443 516323 642477
rect 516357 642443 516391 642477
rect 516425 642443 516459 642477
rect 516493 642443 516527 642477
rect 516561 642443 516595 642477
rect 516629 642443 516676 642477
rect 516276 642405 516676 642443
rect 515818 641379 516218 641405
rect 516276 641379 516676 641405
<< polycont >>
rect 508161 644422 508195 644456
rect 508229 644422 508263 644456
rect 508297 644422 508331 644456
rect 508365 644422 508399 644456
rect 508433 644422 508467 644456
rect 508619 644422 508653 644456
rect 508687 644422 508721 644456
rect 508755 644422 508789 644456
rect 508823 644422 508857 644456
rect 508891 644422 508925 644456
rect 509077 644422 509111 644456
rect 509145 644422 509179 644456
rect 509213 644422 509247 644456
rect 509281 644422 509315 644456
rect 509349 644422 509383 644456
rect 509535 644422 509569 644456
rect 509603 644422 509637 644456
rect 509671 644422 509705 644456
rect 509739 644422 509773 644456
rect 509807 644422 509841 644456
rect 509993 644422 510027 644456
rect 510061 644422 510095 644456
rect 510129 644422 510163 644456
rect 510197 644422 510231 644456
rect 510265 644422 510299 644456
rect 510451 644422 510485 644456
rect 510519 644422 510553 644456
rect 510587 644422 510621 644456
rect 510655 644422 510689 644456
rect 510723 644422 510757 644456
rect 510909 644422 510943 644456
rect 510977 644422 511011 644456
rect 511045 644422 511079 644456
rect 511113 644422 511147 644456
rect 511181 644422 511215 644456
rect 511367 644422 511401 644456
rect 511435 644422 511469 644456
rect 511503 644422 511537 644456
rect 511571 644422 511605 644456
rect 511639 644422 511673 644456
rect 511825 644422 511859 644456
rect 511893 644422 511927 644456
rect 511961 644422 511995 644456
rect 512029 644422 512063 644456
rect 512097 644422 512131 644456
rect 512283 644422 512317 644456
rect 512351 644422 512385 644456
rect 512419 644422 512453 644456
rect 512487 644422 512521 644456
rect 512555 644422 512589 644456
rect 512741 644422 512775 644456
rect 512809 644422 512843 644456
rect 512877 644422 512911 644456
rect 512945 644422 512979 644456
rect 513013 644422 513047 644456
rect 513199 644422 513233 644456
rect 513267 644422 513301 644456
rect 513335 644422 513369 644456
rect 513403 644422 513437 644456
rect 513471 644422 513505 644456
rect 513657 644422 513691 644456
rect 513725 644422 513759 644456
rect 513793 644422 513827 644456
rect 513861 644422 513895 644456
rect 513929 644422 513963 644456
rect 514115 644422 514149 644456
rect 514183 644422 514217 644456
rect 514251 644422 514285 644456
rect 514319 644422 514353 644456
rect 514387 644422 514421 644456
rect 514573 644422 514607 644456
rect 514641 644422 514675 644456
rect 514709 644422 514743 644456
rect 514777 644422 514811 644456
rect 514845 644422 514879 644456
rect 515031 644422 515065 644456
rect 515099 644422 515133 644456
rect 515167 644422 515201 644456
rect 515235 644422 515269 644456
rect 515303 644422 515337 644456
rect 508161 643256 508195 643290
rect 508229 643256 508263 643290
rect 508297 643256 508331 643290
rect 508365 643256 508399 643290
rect 508433 643256 508467 643290
rect 508619 643256 508653 643290
rect 508687 643256 508721 643290
rect 508755 643256 508789 643290
rect 508823 643256 508857 643290
rect 508891 643256 508925 643290
rect 509077 643256 509111 643290
rect 509145 643256 509179 643290
rect 509213 643256 509247 643290
rect 509281 643256 509315 643290
rect 509349 643256 509383 643290
rect 509535 643256 509569 643290
rect 509603 643256 509637 643290
rect 509671 643256 509705 643290
rect 509739 643256 509773 643290
rect 509807 643256 509841 643290
rect 509993 643256 510027 643290
rect 510061 643256 510095 643290
rect 510129 643256 510163 643290
rect 510197 643256 510231 643290
rect 510265 643256 510299 643290
rect 510451 643256 510485 643290
rect 510519 643256 510553 643290
rect 510587 643256 510621 643290
rect 510655 643256 510689 643290
rect 510723 643256 510757 643290
rect 510909 643256 510943 643290
rect 510977 643256 511011 643290
rect 511045 643256 511079 643290
rect 511113 643256 511147 643290
rect 511181 643256 511215 643290
rect 511367 643256 511401 643290
rect 511435 643256 511469 643290
rect 511503 643256 511537 643290
rect 511571 643256 511605 643290
rect 511639 643256 511673 643290
rect 511825 643256 511859 643290
rect 511893 643256 511927 643290
rect 511961 643256 511995 643290
rect 512029 643256 512063 643290
rect 512097 643256 512131 643290
rect 512283 643256 512317 643290
rect 512351 643256 512385 643290
rect 512419 643256 512453 643290
rect 512487 643256 512521 643290
rect 512555 643256 512589 643290
rect 512741 643256 512775 643290
rect 512809 643256 512843 643290
rect 512877 643256 512911 643290
rect 512945 643256 512979 643290
rect 513013 643256 513047 643290
rect 513199 643256 513233 643290
rect 513267 643256 513301 643290
rect 513335 643256 513369 643290
rect 513403 643256 513437 643290
rect 513471 643256 513505 643290
rect 513657 643256 513691 643290
rect 513725 643256 513759 643290
rect 513793 643256 513827 643290
rect 513861 643256 513895 643290
rect 513929 643256 513963 643290
rect 514115 643256 514149 643290
rect 514183 643256 514217 643290
rect 514251 643256 514285 643290
rect 514319 643256 514353 643290
rect 514387 643256 514421 643290
rect 514573 643256 514607 643290
rect 514641 643256 514675 643290
rect 514709 643256 514743 643290
rect 514777 643256 514811 643290
rect 514845 643256 514879 643290
rect 515031 643256 515065 643290
rect 515099 643256 515133 643290
rect 515167 643256 515201 643290
rect 515235 643256 515269 643290
rect 515303 643256 515337 643290
rect 515865 643256 515899 643290
rect 515933 643256 515967 643290
rect 516001 643256 516035 643290
rect 516069 643256 516103 643290
rect 516137 643256 516171 643290
rect 516323 643256 516357 643290
rect 516391 643256 516425 643290
rect 516459 643256 516493 643290
rect 516527 643256 516561 643290
rect 516595 643256 516629 643290
rect 508161 642443 508195 642477
rect 508229 642443 508263 642477
rect 508297 642443 508331 642477
rect 508365 642443 508399 642477
rect 508433 642443 508467 642477
rect 508619 642443 508653 642477
rect 508687 642443 508721 642477
rect 508755 642443 508789 642477
rect 508823 642443 508857 642477
rect 508891 642443 508925 642477
rect 509077 642443 509111 642477
rect 509145 642443 509179 642477
rect 509213 642443 509247 642477
rect 509281 642443 509315 642477
rect 509349 642443 509383 642477
rect 509535 642443 509569 642477
rect 509603 642443 509637 642477
rect 509671 642443 509705 642477
rect 509739 642443 509773 642477
rect 509807 642443 509841 642477
rect 509993 642443 510027 642477
rect 510061 642443 510095 642477
rect 510129 642443 510163 642477
rect 510197 642443 510231 642477
rect 510265 642443 510299 642477
rect 510451 642443 510485 642477
rect 510519 642443 510553 642477
rect 510587 642443 510621 642477
rect 510655 642443 510689 642477
rect 510723 642443 510757 642477
rect 510909 642443 510943 642477
rect 510977 642443 511011 642477
rect 511045 642443 511079 642477
rect 511113 642443 511147 642477
rect 511181 642443 511215 642477
rect 511367 642443 511401 642477
rect 511435 642443 511469 642477
rect 511503 642443 511537 642477
rect 511571 642443 511605 642477
rect 511639 642443 511673 642477
rect 511825 642443 511859 642477
rect 511893 642443 511927 642477
rect 511961 642443 511995 642477
rect 512029 642443 512063 642477
rect 512097 642443 512131 642477
rect 512283 642443 512317 642477
rect 512351 642443 512385 642477
rect 512419 642443 512453 642477
rect 512487 642443 512521 642477
rect 512555 642443 512589 642477
rect 512741 642443 512775 642477
rect 512809 642443 512843 642477
rect 512877 642443 512911 642477
rect 512945 642443 512979 642477
rect 513013 642443 513047 642477
rect 513199 642443 513233 642477
rect 513267 642443 513301 642477
rect 513335 642443 513369 642477
rect 513403 642443 513437 642477
rect 513471 642443 513505 642477
rect 513657 642443 513691 642477
rect 513725 642443 513759 642477
rect 513793 642443 513827 642477
rect 513861 642443 513895 642477
rect 513929 642443 513963 642477
rect 514115 642443 514149 642477
rect 514183 642443 514217 642477
rect 514251 642443 514285 642477
rect 514319 642443 514353 642477
rect 514387 642443 514421 642477
rect 514573 642443 514607 642477
rect 514641 642443 514675 642477
rect 514709 642443 514743 642477
rect 514777 642443 514811 642477
rect 514845 642443 514879 642477
rect 515031 642443 515065 642477
rect 515099 642443 515133 642477
rect 515167 642443 515201 642477
rect 515235 642443 515269 642477
rect 515303 642443 515337 642477
rect 508161 641281 508195 641315
rect 508229 641281 508263 641315
rect 508297 641281 508331 641315
rect 508365 641281 508399 641315
rect 508433 641281 508467 641315
rect 508619 641281 508653 641315
rect 508687 641281 508721 641315
rect 508755 641281 508789 641315
rect 508823 641281 508857 641315
rect 508891 641281 508925 641315
rect 509077 641281 509111 641315
rect 509145 641281 509179 641315
rect 509213 641281 509247 641315
rect 509281 641281 509315 641315
rect 509349 641281 509383 641315
rect 509535 641281 509569 641315
rect 509603 641281 509637 641315
rect 509671 641281 509705 641315
rect 509739 641281 509773 641315
rect 509807 641281 509841 641315
rect 509993 641281 510027 641315
rect 510061 641281 510095 641315
rect 510129 641281 510163 641315
rect 510197 641281 510231 641315
rect 510265 641281 510299 641315
rect 510451 641281 510485 641315
rect 510519 641281 510553 641315
rect 510587 641281 510621 641315
rect 510655 641281 510689 641315
rect 510723 641281 510757 641315
rect 510909 641281 510943 641315
rect 510977 641281 511011 641315
rect 511045 641281 511079 641315
rect 511113 641281 511147 641315
rect 511181 641281 511215 641315
rect 511367 641281 511401 641315
rect 511435 641281 511469 641315
rect 511503 641281 511537 641315
rect 511571 641281 511605 641315
rect 511639 641281 511673 641315
rect 511825 641281 511859 641315
rect 511893 641281 511927 641315
rect 511961 641281 511995 641315
rect 512029 641281 512063 641315
rect 512097 641281 512131 641315
rect 512283 641281 512317 641315
rect 512351 641281 512385 641315
rect 512419 641281 512453 641315
rect 512487 641281 512521 641315
rect 512555 641281 512589 641315
rect 512741 641281 512775 641315
rect 512809 641281 512843 641315
rect 512877 641281 512911 641315
rect 512945 641281 512979 641315
rect 513013 641281 513047 641315
rect 513199 641281 513233 641315
rect 513267 641281 513301 641315
rect 513335 641281 513369 641315
rect 513403 641281 513437 641315
rect 513471 641281 513505 641315
rect 513657 641281 513691 641315
rect 513725 641281 513759 641315
rect 513793 641281 513827 641315
rect 513861 641281 513895 641315
rect 513929 641281 513963 641315
rect 514115 641281 514149 641315
rect 514183 641281 514217 641315
rect 514251 641281 514285 641315
rect 514319 641281 514353 641315
rect 514387 641281 514421 641315
rect 514573 641281 514607 641315
rect 514641 641281 514675 641315
rect 514709 641281 514743 641315
rect 514777 641281 514811 641315
rect 514845 641281 514879 641315
rect 515031 641281 515065 641315
rect 515099 641281 515133 641315
rect 515167 641281 515201 641315
rect 515235 641281 515269 641315
rect 515303 641281 515337 641315
rect 515865 642443 515899 642477
rect 515933 642443 515967 642477
rect 516001 642443 516035 642477
rect 516069 642443 516103 642477
rect 516137 642443 516171 642477
rect 516323 642443 516357 642477
rect 516391 642443 516425 642477
rect 516459 642443 516493 642477
rect 516527 642443 516561 642477
rect 516595 642443 516629 642477
<< locali >>
rect 507828 645725 516966 645743
rect 507828 645623 507846 645725
rect 507948 645623 507992 645725
rect 515506 645623 515550 645725
rect 515652 645623 515722 645725
rect 516776 645623 516846 645725
rect 516948 645623 516966 645725
rect 507828 645605 516966 645623
rect 507828 645551 507966 645605
rect 507828 643205 507846 645551
rect 507948 643205 507966 645551
rect 515532 645581 516966 645605
rect 515532 645551 515722 645581
rect 508068 645488 508102 645507
rect 508068 645416 508102 645428
rect 508068 645344 508102 645360
rect 508068 645272 508102 645292
rect 508068 645200 508102 645224
rect 508068 645128 508102 645156
rect 508068 645056 508102 645088
rect 508068 644986 508102 645020
rect 508068 644918 508102 644950
rect 508068 644850 508102 644878
rect 508068 644782 508102 644806
rect 508068 644714 508102 644734
rect 508068 644646 508102 644662
rect 508068 644578 508102 644590
rect 508068 644499 508102 644518
rect 508526 645488 508560 645507
rect 508526 645416 508560 645428
rect 508526 645344 508560 645360
rect 508526 645272 508560 645292
rect 508526 645200 508560 645224
rect 508526 645128 508560 645156
rect 508526 645056 508560 645088
rect 508526 644986 508560 645020
rect 508526 644918 508560 644950
rect 508526 644850 508560 644878
rect 508526 644782 508560 644806
rect 508526 644714 508560 644734
rect 508526 644646 508560 644662
rect 508526 644578 508560 644590
rect 508526 644499 508560 644518
rect 508984 645488 509018 645507
rect 508984 645416 509018 645428
rect 508984 645344 509018 645360
rect 508984 645272 509018 645292
rect 508984 645200 509018 645224
rect 508984 645128 509018 645156
rect 508984 645056 509018 645088
rect 508984 644986 509018 645020
rect 508984 644918 509018 644950
rect 508984 644850 509018 644878
rect 508984 644782 509018 644806
rect 508984 644714 509018 644734
rect 508984 644646 509018 644662
rect 508984 644578 509018 644590
rect 508984 644499 509018 644518
rect 509442 645488 509476 645507
rect 509442 645416 509476 645428
rect 509442 645344 509476 645360
rect 509442 645272 509476 645292
rect 509442 645200 509476 645224
rect 509442 645128 509476 645156
rect 509442 645056 509476 645088
rect 509442 644986 509476 645020
rect 509442 644918 509476 644950
rect 509442 644850 509476 644878
rect 509442 644782 509476 644806
rect 509442 644714 509476 644734
rect 509442 644646 509476 644662
rect 509442 644578 509476 644590
rect 509442 644499 509476 644518
rect 509900 645488 509934 645507
rect 509900 645416 509934 645428
rect 509900 645344 509934 645360
rect 509900 645272 509934 645292
rect 509900 645200 509934 645224
rect 509900 645128 509934 645156
rect 509900 645056 509934 645088
rect 509900 644986 509934 645020
rect 509900 644918 509934 644950
rect 509900 644850 509934 644878
rect 509900 644782 509934 644806
rect 509900 644714 509934 644734
rect 509900 644646 509934 644662
rect 509900 644578 509934 644590
rect 509900 644499 509934 644518
rect 510358 645488 510392 645507
rect 510358 645416 510392 645428
rect 510358 645344 510392 645360
rect 510358 645272 510392 645292
rect 510358 645200 510392 645224
rect 510358 645128 510392 645156
rect 510358 645056 510392 645088
rect 510358 644986 510392 645020
rect 510358 644918 510392 644950
rect 510358 644850 510392 644878
rect 510358 644782 510392 644806
rect 510358 644714 510392 644734
rect 510358 644646 510392 644662
rect 510358 644578 510392 644590
rect 510358 644499 510392 644518
rect 510816 645488 510850 645507
rect 510816 645416 510850 645428
rect 510816 645344 510850 645360
rect 510816 645272 510850 645292
rect 510816 645200 510850 645224
rect 510816 645128 510850 645156
rect 510816 645056 510850 645088
rect 510816 644986 510850 645020
rect 510816 644918 510850 644950
rect 510816 644850 510850 644878
rect 510816 644782 510850 644806
rect 510816 644714 510850 644734
rect 510816 644646 510850 644662
rect 510816 644578 510850 644590
rect 510816 644499 510850 644518
rect 511274 645488 511308 645507
rect 511274 645416 511308 645428
rect 511274 645344 511308 645360
rect 511274 645272 511308 645292
rect 511274 645200 511308 645224
rect 511274 645128 511308 645156
rect 511274 645056 511308 645088
rect 511274 644986 511308 645020
rect 511274 644918 511308 644950
rect 511274 644850 511308 644878
rect 511274 644782 511308 644806
rect 511274 644714 511308 644734
rect 511274 644646 511308 644662
rect 511274 644578 511308 644590
rect 511274 644499 511308 644518
rect 511732 645488 511766 645507
rect 511732 645416 511766 645428
rect 511732 645344 511766 645360
rect 511732 645272 511766 645292
rect 511732 645200 511766 645224
rect 511732 645128 511766 645156
rect 511732 645056 511766 645088
rect 511732 644986 511766 645020
rect 511732 644918 511766 644950
rect 511732 644850 511766 644878
rect 511732 644782 511766 644806
rect 511732 644714 511766 644734
rect 511732 644646 511766 644662
rect 511732 644578 511766 644590
rect 511732 644499 511766 644518
rect 512190 645488 512224 645507
rect 512190 645416 512224 645428
rect 512190 645344 512224 645360
rect 512190 645272 512224 645292
rect 512190 645200 512224 645224
rect 512190 645128 512224 645156
rect 512190 645056 512224 645088
rect 512190 644986 512224 645020
rect 512190 644918 512224 644950
rect 512190 644850 512224 644878
rect 512190 644782 512224 644806
rect 512190 644714 512224 644734
rect 512190 644646 512224 644662
rect 512190 644578 512224 644590
rect 512190 644499 512224 644518
rect 512648 645488 512682 645507
rect 512648 645416 512682 645428
rect 512648 645344 512682 645360
rect 512648 645272 512682 645292
rect 512648 645200 512682 645224
rect 512648 645128 512682 645156
rect 512648 645056 512682 645088
rect 512648 644986 512682 645020
rect 512648 644918 512682 644950
rect 512648 644850 512682 644878
rect 512648 644782 512682 644806
rect 512648 644714 512682 644734
rect 512648 644646 512682 644662
rect 512648 644578 512682 644590
rect 512648 644499 512682 644518
rect 513106 645488 513140 645507
rect 513106 645416 513140 645428
rect 513106 645344 513140 645360
rect 513106 645272 513140 645292
rect 513106 645200 513140 645224
rect 513106 645128 513140 645156
rect 513106 645056 513140 645088
rect 513106 644986 513140 645020
rect 513106 644918 513140 644950
rect 513106 644850 513140 644878
rect 513106 644782 513140 644806
rect 513106 644714 513140 644734
rect 513106 644646 513140 644662
rect 513106 644578 513140 644590
rect 513106 644499 513140 644518
rect 513564 645488 513598 645507
rect 513564 645416 513598 645428
rect 513564 645344 513598 645360
rect 513564 645272 513598 645292
rect 513564 645200 513598 645224
rect 513564 645128 513598 645156
rect 513564 645056 513598 645088
rect 513564 644986 513598 645020
rect 513564 644918 513598 644950
rect 513564 644850 513598 644878
rect 513564 644782 513598 644806
rect 513564 644714 513598 644734
rect 513564 644646 513598 644662
rect 513564 644578 513598 644590
rect 513564 644499 513598 644518
rect 514022 645488 514056 645507
rect 514022 645416 514056 645428
rect 514022 645344 514056 645360
rect 514022 645272 514056 645292
rect 514022 645200 514056 645224
rect 514022 645128 514056 645156
rect 514022 645056 514056 645088
rect 514022 644986 514056 645020
rect 514022 644918 514056 644950
rect 514022 644850 514056 644878
rect 514022 644782 514056 644806
rect 514022 644714 514056 644734
rect 514022 644646 514056 644662
rect 514022 644578 514056 644590
rect 514022 644499 514056 644518
rect 514480 645488 514514 645507
rect 514480 645416 514514 645428
rect 514480 645344 514514 645360
rect 514480 645272 514514 645292
rect 514480 645200 514514 645224
rect 514480 645128 514514 645156
rect 514480 645056 514514 645088
rect 514480 644986 514514 645020
rect 514480 644918 514514 644950
rect 514480 644850 514514 644878
rect 514480 644782 514514 644806
rect 514480 644714 514514 644734
rect 514480 644646 514514 644662
rect 514480 644578 514514 644590
rect 514480 644499 514514 644518
rect 514938 645488 514972 645507
rect 514938 645416 514972 645428
rect 514938 645344 514972 645360
rect 514938 645272 514972 645292
rect 514938 645200 514972 645224
rect 514938 645128 514972 645156
rect 514938 645056 514972 645088
rect 514938 644986 514972 645020
rect 514938 644918 514972 644950
rect 514938 644850 514972 644878
rect 514938 644782 514972 644806
rect 514938 644714 514972 644734
rect 514938 644646 514972 644662
rect 514938 644578 514972 644590
rect 514938 644499 514972 644518
rect 515396 645488 515430 645507
rect 515396 645416 515430 645428
rect 515396 645344 515430 645360
rect 515396 645272 515430 645292
rect 515396 645200 515430 645224
rect 515396 645128 515430 645156
rect 515396 645056 515430 645088
rect 515396 644986 515430 645020
rect 515396 644918 515430 644950
rect 515396 644850 515430 644878
rect 515396 644782 515430 644806
rect 515396 644714 515430 644734
rect 515396 644646 515430 644662
rect 515396 644578 515430 644590
rect 515396 644499 515430 644518
rect 508114 644422 508153 644456
rect 508195 644422 508225 644456
rect 508263 644422 508297 644456
rect 508331 644422 508365 644456
rect 508403 644422 508433 644456
rect 508475 644422 508514 644456
rect 508572 644422 508611 644456
rect 508653 644422 508683 644456
rect 508721 644422 508755 644456
rect 508789 644422 508823 644456
rect 508861 644422 508891 644456
rect 508933 644422 508972 644456
rect 509030 644422 509069 644456
rect 509111 644422 509141 644456
rect 509179 644422 509213 644456
rect 509247 644422 509281 644456
rect 509319 644422 509349 644456
rect 509391 644422 509430 644456
rect 509488 644422 509527 644456
rect 509569 644422 509599 644456
rect 509637 644422 509671 644456
rect 509705 644422 509739 644456
rect 509777 644422 509807 644456
rect 509849 644422 509888 644456
rect 509946 644422 509985 644456
rect 510027 644422 510057 644456
rect 510095 644422 510129 644456
rect 510163 644422 510197 644456
rect 510235 644422 510265 644456
rect 510307 644422 510346 644456
rect 510404 644422 510443 644456
rect 510485 644422 510515 644456
rect 510553 644422 510587 644456
rect 510621 644422 510655 644456
rect 510693 644422 510723 644456
rect 510765 644422 510804 644456
rect 510862 644422 510901 644456
rect 510943 644422 510973 644456
rect 511011 644422 511045 644456
rect 511079 644422 511113 644456
rect 511151 644422 511181 644456
rect 511223 644422 511262 644456
rect 511320 644422 511359 644456
rect 511401 644422 511431 644456
rect 511469 644422 511503 644456
rect 511537 644422 511571 644456
rect 511609 644422 511639 644456
rect 511681 644422 511720 644456
rect 511778 644422 511817 644456
rect 511859 644422 511889 644456
rect 511927 644422 511961 644456
rect 511995 644422 512029 644456
rect 512067 644422 512097 644456
rect 512139 644422 512178 644456
rect 512236 644422 512275 644456
rect 512317 644422 512347 644456
rect 512385 644422 512419 644456
rect 512453 644422 512487 644456
rect 512525 644422 512555 644456
rect 512597 644422 512636 644456
rect 512694 644422 512733 644456
rect 512775 644422 512805 644456
rect 512843 644422 512877 644456
rect 512911 644422 512945 644456
rect 512983 644422 513013 644456
rect 513055 644422 513094 644456
rect 513152 644422 513191 644456
rect 513233 644422 513263 644456
rect 513301 644422 513335 644456
rect 513369 644422 513403 644456
rect 513441 644422 513471 644456
rect 513513 644422 513552 644456
rect 513610 644422 513649 644456
rect 513691 644422 513721 644456
rect 513759 644422 513793 644456
rect 513827 644422 513861 644456
rect 513899 644422 513929 644456
rect 513971 644422 514010 644456
rect 514068 644422 514107 644456
rect 514149 644422 514179 644456
rect 514217 644422 514251 644456
rect 514285 644422 514319 644456
rect 514357 644422 514387 644456
rect 514429 644422 514468 644456
rect 514526 644422 514565 644456
rect 514607 644422 514637 644456
rect 514675 644422 514709 644456
rect 514743 644422 514777 644456
rect 514815 644422 514845 644456
rect 514887 644422 514926 644456
rect 514984 644422 515023 644456
rect 515065 644422 515095 644456
rect 515133 644422 515167 644456
rect 515201 644422 515235 644456
rect 515273 644422 515303 644456
rect 515345 644422 515384 644456
rect 508068 644322 508102 644341
rect 508068 644250 508102 644262
rect 508068 644178 508102 644194
rect 508068 644106 508102 644126
rect 508068 644034 508102 644058
rect 508068 643962 508102 643990
rect 508068 643890 508102 643922
rect 508068 643820 508102 643854
rect 508068 643752 508102 643784
rect 508068 643684 508102 643712
rect 508068 643616 508102 643640
rect 508068 643548 508102 643568
rect 508068 643480 508102 643496
rect 508068 643412 508102 643424
rect 508068 643333 508102 643352
rect 508526 644322 508560 644341
rect 508526 644250 508560 644262
rect 508526 644178 508560 644194
rect 508526 644106 508560 644126
rect 508526 644034 508560 644058
rect 508526 643962 508560 643990
rect 508526 643890 508560 643922
rect 508526 643820 508560 643854
rect 508526 643752 508560 643784
rect 508526 643684 508560 643712
rect 508526 643616 508560 643640
rect 508526 643548 508560 643568
rect 508526 643480 508560 643496
rect 508526 643412 508560 643424
rect 508526 643333 508560 643352
rect 508984 644322 509018 644341
rect 508984 644250 509018 644262
rect 508984 644178 509018 644194
rect 508984 644106 509018 644126
rect 508984 644034 509018 644058
rect 508984 643962 509018 643990
rect 508984 643890 509018 643922
rect 508984 643820 509018 643854
rect 508984 643752 509018 643784
rect 508984 643684 509018 643712
rect 508984 643616 509018 643640
rect 508984 643548 509018 643568
rect 508984 643480 509018 643496
rect 508984 643412 509018 643424
rect 508984 643333 509018 643352
rect 509442 644322 509476 644341
rect 509442 644250 509476 644262
rect 509442 644178 509476 644194
rect 509442 644106 509476 644126
rect 509442 644034 509476 644058
rect 509442 643962 509476 643990
rect 509442 643890 509476 643922
rect 509442 643820 509476 643854
rect 509442 643752 509476 643784
rect 509442 643684 509476 643712
rect 509442 643616 509476 643640
rect 509442 643548 509476 643568
rect 509442 643480 509476 643496
rect 509442 643412 509476 643424
rect 509442 643333 509476 643352
rect 509900 644322 509934 644341
rect 509900 644250 509934 644262
rect 509900 644178 509934 644194
rect 509900 644106 509934 644126
rect 509900 644034 509934 644058
rect 509900 643962 509934 643990
rect 509900 643890 509934 643922
rect 509900 643820 509934 643854
rect 509900 643752 509934 643784
rect 509900 643684 509934 643712
rect 509900 643616 509934 643640
rect 509900 643548 509934 643568
rect 509900 643480 509934 643496
rect 509900 643412 509934 643424
rect 509900 643333 509934 643352
rect 510358 644322 510392 644341
rect 510358 644250 510392 644262
rect 510358 644178 510392 644194
rect 510358 644106 510392 644126
rect 510358 644034 510392 644058
rect 510358 643962 510392 643990
rect 510358 643890 510392 643922
rect 510358 643820 510392 643854
rect 510358 643752 510392 643784
rect 510358 643684 510392 643712
rect 510358 643616 510392 643640
rect 510358 643548 510392 643568
rect 510358 643480 510392 643496
rect 510358 643412 510392 643424
rect 510358 643333 510392 643352
rect 510816 644322 510850 644341
rect 510816 644250 510850 644262
rect 510816 644178 510850 644194
rect 510816 644106 510850 644126
rect 510816 644034 510850 644058
rect 510816 643962 510850 643990
rect 510816 643890 510850 643922
rect 510816 643820 510850 643854
rect 510816 643752 510850 643784
rect 510816 643684 510850 643712
rect 510816 643616 510850 643640
rect 510816 643548 510850 643568
rect 510816 643480 510850 643496
rect 510816 643412 510850 643424
rect 510816 643333 510850 643352
rect 511274 644322 511308 644341
rect 511274 644250 511308 644262
rect 511274 644178 511308 644194
rect 511274 644106 511308 644126
rect 511274 644034 511308 644058
rect 511274 643962 511308 643990
rect 511274 643890 511308 643922
rect 511274 643820 511308 643854
rect 511274 643752 511308 643784
rect 511274 643684 511308 643712
rect 511274 643616 511308 643640
rect 511274 643548 511308 643568
rect 511274 643480 511308 643496
rect 511274 643412 511308 643424
rect 511274 643333 511308 643352
rect 511732 644322 511766 644341
rect 511732 644250 511766 644262
rect 511732 644178 511766 644194
rect 511732 644106 511766 644126
rect 511732 644034 511766 644058
rect 511732 643962 511766 643990
rect 511732 643890 511766 643922
rect 511732 643820 511766 643854
rect 511732 643752 511766 643784
rect 511732 643684 511766 643712
rect 511732 643616 511766 643640
rect 511732 643548 511766 643568
rect 511732 643480 511766 643496
rect 511732 643412 511766 643424
rect 511732 643333 511766 643352
rect 512190 644322 512224 644341
rect 512190 644250 512224 644262
rect 512190 644178 512224 644194
rect 512190 644106 512224 644126
rect 512190 644034 512224 644058
rect 512190 643962 512224 643990
rect 512190 643890 512224 643922
rect 512190 643820 512224 643854
rect 512190 643752 512224 643784
rect 512190 643684 512224 643712
rect 512190 643616 512224 643640
rect 512190 643548 512224 643568
rect 512190 643480 512224 643496
rect 512190 643412 512224 643424
rect 512190 643333 512224 643352
rect 512648 644322 512682 644341
rect 512648 644250 512682 644262
rect 512648 644178 512682 644194
rect 512648 644106 512682 644126
rect 512648 644034 512682 644058
rect 512648 643962 512682 643990
rect 512648 643890 512682 643922
rect 512648 643820 512682 643854
rect 512648 643752 512682 643784
rect 512648 643684 512682 643712
rect 512648 643616 512682 643640
rect 512648 643548 512682 643568
rect 512648 643480 512682 643496
rect 512648 643412 512682 643424
rect 512648 643333 512682 643352
rect 513106 644322 513140 644341
rect 513106 644250 513140 644262
rect 513106 644178 513140 644194
rect 513106 644106 513140 644126
rect 513106 644034 513140 644058
rect 513106 643962 513140 643990
rect 513106 643890 513140 643922
rect 513106 643820 513140 643854
rect 513106 643752 513140 643784
rect 513106 643684 513140 643712
rect 513106 643616 513140 643640
rect 513106 643548 513140 643568
rect 513106 643480 513140 643496
rect 513106 643412 513140 643424
rect 513106 643333 513140 643352
rect 513564 644322 513598 644341
rect 513564 644250 513598 644262
rect 513564 644178 513598 644194
rect 513564 644106 513598 644126
rect 513564 644034 513598 644058
rect 513564 643962 513598 643990
rect 513564 643890 513598 643922
rect 513564 643820 513598 643854
rect 513564 643752 513598 643784
rect 513564 643684 513598 643712
rect 513564 643616 513598 643640
rect 513564 643548 513598 643568
rect 513564 643480 513598 643496
rect 513564 643412 513598 643424
rect 513564 643333 513598 643352
rect 514022 644322 514056 644341
rect 514022 644250 514056 644262
rect 514022 644178 514056 644194
rect 514022 644106 514056 644126
rect 514022 644034 514056 644058
rect 514022 643962 514056 643990
rect 514022 643890 514056 643922
rect 514022 643820 514056 643854
rect 514022 643752 514056 643784
rect 514022 643684 514056 643712
rect 514022 643616 514056 643640
rect 514022 643548 514056 643568
rect 514022 643480 514056 643496
rect 514022 643412 514056 643424
rect 514022 643333 514056 643352
rect 514480 644322 514514 644341
rect 514480 644250 514514 644262
rect 514480 644178 514514 644194
rect 514480 644106 514514 644126
rect 514480 644034 514514 644058
rect 514480 643962 514514 643990
rect 514480 643890 514514 643922
rect 514480 643820 514514 643854
rect 514480 643752 514514 643784
rect 514480 643684 514514 643712
rect 514480 643616 514514 643640
rect 514480 643548 514514 643568
rect 514480 643480 514514 643496
rect 514480 643412 514514 643424
rect 514480 643333 514514 643352
rect 514938 644322 514972 644341
rect 514938 644250 514972 644262
rect 514938 644178 514972 644194
rect 514938 644106 514972 644126
rect 514938 644034 514972 644058
rect 514938 643962 514972 643990
rect 514938 643890 514972 643922
rect 514938 643820 514972 643854
rect 514938 643752 514972 643784
rect 514938 643684 514972 643712
rect 514938 643616 514972 643640
rect 514938 643548 514972 643568
rect 514938 643480 514972 643496
rect 514938 643412 514972 643424
rect 514938 643333 514972 643352
rect 515396 644322 515430 644341
rect 515396 644250 515430 644262
rect 515396 644178 515430 644194
rect 515396 644106 515430 644126
rect 515396 644034 515430 644058
rect 515396 643962 515430 643990
rect 515396 643890 515430 643922
rect 515396 643820 515430 643854
rect 515396 643752 515430 643784
rect 515396 643684 515430 643712
rect 515396 643616 515430 643640
rect 515396 643548 515430 643568
rect 515396 643480 515430 643496
rect 515396 643412 515430 643424
rect 515396 643333 515430 643352
rect 508114 643256 508153 643290
rect 508195 643256 508225 643290
rect 508263 643256 508297 643290
rect 508331 643256 508365 643290
rect 508403 643256 508433 643290
rect 508475 643256 508514 643290
rect 508572 643256 508611 643290
rect 508653 643256 508683 643290
rect 508721 643256 508755 643290
rect 508789 643256 508823 643290
rect 508861 643256 508891 643290
rect 508933 643256 508972 643290
rect 509030 643256 509069 643290
rect 509111 643256 509141 643290
rect 509179 643256 509213 643290
rect 509247 643256 509281 643290
rect 509319 643256 509349 643290
rect 509391 643256 509430 643290
rect 509488 643256 509527 643290
rect 509569 643256 509599 643290
rect 509637 643256 509671 643290
rect 509705 643256 509739 643290
rect 509777 643256 509807 643290
rect 509849 643256 509888 643290
rect 509946 643256 509985 643290
rect 510027 643256 510057 643290
rect 510095 643256 510129 643290
rect 510163 643256 510197 643290
rect 510235 643256 510265 643290
rect 510307 643256 510346 643290
rect 510404 643256 510443 643290
rect 510485 643256 510515 643290
rect 510553 643256 510587 643290
rect 510621 643256 510655 643290
rect 510693 643256 510723 643290
rect 510765 643256 510804 643290
rect 510862 643256 510901 643290
rect 510943 643256 510973 643290
rect 511011 643256 511045 643290
rect 511079 643256 511113 643290
rect 511151 643256 511181 643290
rect 511223 643256 511262 643290
rect 511320 643256 511359 643290
rect 511401 643256 511431 643290
rect 511469 643256 511503 643290
rect 511537 643256 511571 643290
rect 511609 643256 511639 643290
rect 511681 643256 511720 643290
rect 511778 643256 511817 643290
rect 511859 643256 511889 643290
rect 511927 643256 511961 643290
rect 511995 643256 512029 643290
rect 512067 643256 512097 643290
rect 512139 643256 512178 643290
rect 512236 643256 512275 643290
rect 512317 643256 512347 643290
rect 512385 643256 512419 643290
rect 512453 643256 512487 643290
rect 512525 643256 512555 643290
rect 512597 643256 512636 643290
rect 512694 643256 512733 643290
rect 512775 643256 512805 643290
rect 512843 643256 512877 643290
rect 512911 643256 512945 643290
rect 512983 643256 513013 643290
rect 513055 643256 513094 643290
rect 513152 643256 513191 643290
rect 513233 643256 513263 643290
rect 513301 643256 513335 643290
rect 513369 643256 513403 643290
rect 513441 643256 513471 643290
rect 513513 643256 513552 643290
rect 513610 643256 513649 643290
rect 513691 643256 513721 643290
rect 513759 643256 513793 643290
rect 513827 643256 513861 643290
rect 513899 643256 513929 643290
rect 513971 643256 514010 643290
rect 514068 643256 514107 643290
rect 514149 643256 514179 643290
rect 514217 643256 514251 643290
rect 514285 643256 514319 643290
rect 514357 643256 514387 643290
rect 514429 643256 514468 643290
rect 514526 643256 514565 643290
rect 514607 643256 514637 643290
rect 514675 643256 514709 643290
rect 514743 643256 514777 643290
rect 514815 643256 514845 643290
rect 514887 643256 514926 643290
rect 514984 643256 515023 643290
rect 515065 643256 515095 643290
rect 515133 643256 515167 643290
rect 515201 643256 515235 643290
rect 515273 643256 515303 643290
rect 515345 643256 515384 643290
rect 507828 643151 507966 643205
rect 515532 643205 515550 645551
rect 515652 645479 515722 645551
rect 516776 645551 516966 645581
rect 516776 645479 516846 645551
rect 515652 645461 516846 645479
rect 515652 643205 515670 645461
rect 515772 645306 515806 645341
rect 515772 645238 515806 645256
rect 515772 645170 515806 645184
rect 515772 645102 515806 645112
rect 515772 645034 515806 645040
rect 515772 644966 515806 644968
rect 515772 644930 515806 644932
rect 515772 644858 515806 644864
rect 515772 644786 515806 644796
rect 515772 644714 515806 644728
rect 515772 644642 515806 644660
rect 515772 644570 515806 644592
rect 515772 644498 515806 644524
rect 515772 644426 515806 644456
rect 515772 644354 515806 644388
rect 515772 644286 515806 644320
rect 515772 644218 515806 644248
rect 515772 644150 515806 644176
rect 515772 644082 515806 644104
rect 515772 644014 515806 644032
rect 515772 643946 515806 643960
rect 515772 643878 515806 643888
rect 515772 643810 515806 643816
rect 515772 643742 515806 643744
rect 515772 643706 515806 643708
rect 515772 643634 515806 643640
rect 515772 643562 515806 643572
rect 515772 643490 515806 643504
rect 515772 643418 515806 643436
rect 515772 643333 515806 643368
rect 516230 645306 516264 645341
rect 516230 645238 516264 645256
rect 516230 645170 516264 645184
rect 516230 645102 516264 645112
rect 516230 645034 516264 645040
rect 516230 644966 516264 644968
rect 516230 644930 516264 644932
rect 516230 644858 516264 644864
rect 516230 644786 516264 644796
rect 516230 644714 516264 644728
rect 516230 644642 516264 644660
rect 516230 644570 516264 644592
rect 516230 644498 516264 644524
rect 516230 644426 516264 644456
rect 516230 644354 516264 644388
rect 516230 644286 516264 644320
rect 516230 644218 516264 644248
rect 516230 644150 516264 644176
rect 516230 644082 516264 644104
rect 516230 644014 516264 644032
rect 516230 643946 516264 643960
rect 516230 643878 516264 643888
rect 516230 643810 516264 643816
rect 516230 643742 516264 643744
rect 516230 643706 516264 643708
rect 516230 643634 516264 643640
rect 516230 643562 516264 643572
rect 516230 643490 516264 643504
rect 516230 643418 516264 643436
rect 516230 643333 516264 643368
rect 516688 645306 516722 645341
rect 516688 645238 516722 645256
rect 516688 645170 516722 645184
rect 516688 645102 516722 645112
rect 516688 645034 516722 645040
rect 516688 644966 516722 644968
rect 516688 644930 516722 644932
rect 516688 644858 516722 644864
rect 516688 644786 516722 644796
rect 516688 644714 516722 644728
rect 516688 644642 516722 644660
rect 516688 644570 516722 644592
rect 516688 644498 516722 644524
rect 516688 644426 516722 644456
rect 516688 644354 516722 644388
rect 516688 644286 516722 644320
rect 516688 644218 516722 644248
rect 516688 644150 516722 644176
rect 516688 644082 516722 644104
rect 516688 644014 516722 644032
rect 516688 643946 516722 643960
rect 516688 643878 516722 643888
rect 516688 643810 516722 643816
rect 516688 643742 516722 643744
rect 516688 643706 516722 643708
rect 516688 643634 516722 643640
rect 516688 643562 516722 643572
rect 516688 643490 516722 643504
rect 516688 643418 516722 643436
rect 516688 643333 516722 643368
rect 515818 643256 515857 643290
rect 515899 643256 515929 643290
rect 515967 643256 516001 643290
rect 516035 643256 516069 643290
rect 516107 643256 516137 643290
rect 516179 643256 516218 643290
rect 516276 643256 516315 643290
rect 516357 643256 516387 643290
rect 516425 643256 516459 643290
rect 516493 643256 516527 643290
rect 516565 643256 516595 643290
rect 516637 643256 516676 643290
rect 515532 643151 515670 643205
rect 516828 643205 516846 645461
rect 516948 643205 516966 645551
rect 516828 643151 516966 643205
rect 507828 643133 516966 643151
rect 507828 643031 507846 643133
rect 507948 643031 507992 643133
rect 515506 643031 515550 643133
rect 515652 643031 515722 643133
rect 516776 643031 516846 643133
rect 516948 643031 516966 643133
rect 507828 643013 516966 643031
rect 507828 642702 516966 642720
rect 507828 642600 507846 642702
rect 507948 642600 507992 642702
rect 515506 642600 515550 642702
rect 515652 642600 515722 642702
rect 516776 642600 516846 642702
rect 516948 642600 516966 642702
rect 507828 642582 516966 642600
rect 507828 642528 507966 642582
rect 507828 640182 507846 642528
rect 507948 640182 507966 642528
rect 515532 642528 515670 642582
rect 508114 642443 508153 642477
rect 508195 642443 508225 642477
rect 508263 642443 508297 642477
rect 508331 642443 508365 642477
rect 508403 642443 508433 642477
rect 508475 642443 508514 642477
rect 508572 642443 508611 642477
rect 508653 642443 508683 642477
rect 508721 642443 508755 642477
rect 508789 642443 508823 642477
rect 508861 642443 508891 642477
rect 508933 642443 508972 642477
rect 509030 642443 509069 642477
rect 509111 642443 509141 642477
rect 509179 642443 509213 642477
rect 509247 642443 509281 642477
rect 509319 642443 509349 642477
rect 509391 642443 509430 642477
rect 509488 642443 509527 642477
rect 509569 642443 509599 642477
rect 509637 642443 509671 642477
rect 509705 642443 509739 642477
rect 509777 642443 509807 642477
rect 509849 642443 509888 642477
rect 509946 642443 509985 642477
rect 510027 642443 510057 642477
rect 510095 642443 510129 642477
rect 510163 642443 510197 642477
rect 510235 642443 510265 642477
rect 510307 642443 510346 642477
rect 510404 642443 510443 642477
rect 510485 642443 510515 642477
rect 510553 642443 510587 642477
rect 510621 642443 510655 642477
rect 510693 642443 510723 642477
rect 510765 642443 510804 642477
rect 510862 642443 510901 642477
rect 510943 642443 510973 642477
rect 511011 642443 511045 642477
rect 511079 642443 511113 642477
rect 511151 642443 511181 642477
rect 511223 642443 511262 642477
rect 511320 642443 511359 642477
rect 511401 642443 511431 642477
rect 511469 642443 511503 642477
rect 511537 642443 511571 642477
rect 511609 642443 511639 642477
rect 511681 642443 511720 642477
rect 511778 642443 511817 642477
rect 511859 642443 511889 642477
rect 511927 642443 511961 642477
rect 511995 642443 512029 642477
rect 512067 642443 512097 642477
rect 512139 642443 512178 642477
rect 512236 642443 512275 642477
rect 512317 642443 512347 642477
rect 512385 642443 512419 642477
rect 512453 642443 512487 642477
rect 512525 642443 512555 642477
rect 512597 642443 512636 642477
rect 512694 642443 512733 642477
rect 512775 642443 512805 642477
rect 512843 642443 512877 642477
rect 512911 642443 512945 642477
rect 512983 642443 513013 642477
rect 513055 642443 513094 642477
rect 513152 642443 513191 642477
rect 513233 642443 513263 642477
rect 513301 642443 513335 642477
rect 513369 642443 513403 642477
rect 513441 642443 513471 642477
rect 513513 642443 513552 642477
rect 513610 642443 513649 642477
rect 513691 642443 513721 642477
rect 513759 642443 513793 642477
rect 513827 642443 513861 642477
rect 513899 642443 513929 642477
rect 513971 642443 514010 642477
rect 514068 642443 514107 642477
rect 514149 642443 514179 642477
rect 514217 642443 514251 642477
rect 514285 642443 514319 642477
rect 514357 642443 514387 642477
rect 514429 642443 514468 642477
rect 514526 642443 514565 642477
rect 514607 642443 514637 642477
rect 514675 642443 514709 642477
rect 514743 642443 514777 642477
rect 514815 642443 514845 642477
rect 514887 642443 514926 642477
rect 514984 642443 515023 642477
rect 515065 642443 515095 642477
rect 515133 642443 515167 642477
rect 515201 642443 515235 642477
rect 515273 642443 515303 642477
rect 515345 642443 515384 642477
rect 508068 642390 508102 642409
rect 508068 642318 508102 642330
rect 508068 642246 508102 642262
rect 508068 642174 508102 642194
rect 508068 642102 508102 642126
rect 508068 642030 508102 642058
rect 508068 641958 508102 641990
rect 508068 641888 508102 641922
rect 508068 641820 508102 641852
rect 508068 641752 508102 641780
rect 508068 641684 508102 641708
rect 508068 641616 508102 641636
rect 508068 641548 508102 641564
rect 508068 641480 508102 641492
rect 508068 641401 508102 641420
rect 508526 642390 508560 642409
rect 508526 642318 508560 642330
rect 508526 642246 508560 642262
rect 508526 642174 508560 642194
rect 508526 642102 508560 642126
rect 508526 642030 508560 642058
rect 508526 641958 508560 641990
rect 508526 641888 508560 641922
rect 508526 641820 508560 641852
rect 508526 641752 508560 641780
rect 508526 641684 508560 641708
rect 508526 641616 508560 641636
rect 508526 641548 508560 641564
rect 508526 641480 508560 641492
rect 508526 641401 508560 641420
rect 508984 642390 509018 642409
rect 508984 642318 509018 642330
rect 508984 642246 509018 642262
rect 508984 642174 509018 642194
rect 508984 642102 509018 642126
rect 508984 642030 509018 642058
rect 508984 641958 509018 641990
rect 508984 641888 509018 641922
rect 508984 641820 509018 641852
rect 508984 641752 509018 641780
rect 508984 641684 509018 641708
rect 508984 641616 509018 641636
rect 508984 641548 509018 641564
rect 508984 641480 509018 641492
rect 508984 641401 509018 641420
rect 509442 642390 509476 642409
rect 509442 642318 509476 642330
rect 509442 642246 509476 642262
rect 509442 642174 509476 642194
rect 509442 642102 509476 642126
rect 509442 642030 509476 642058
rect 509442 641958 509476 641990
rect 509442 641888 509476 641922
rect 509442 641820 509476 641852
rect 509442 641752 509476 641780
rect 509442 641684 509476 641708
rect 509442 641616 509476 641636
rect 509442 641548 509476 641564
rect 509442 641480 509476 641492
rect 509442 641401 509476 641420
rect 509900 642390 509934 642409
rect 509900 642318 509934 642330
rect 509900 642246 509934 642262
rect 509900 642174 509934 642194
rect 509900 642102 509934 642126
rect 509900 642030 509934 642058
rect 509900 641958 509934 641990
rect 509900 641888 509934 641922
rect 509900 641820 509934 641852
rect 509900 641752 509934 641780
rect 509900 641684 509934 641708
rect 509900 641616 509934 641636
rect 509900 641548 509934 641564
rect 509900 641480 509934 641492
rect 509900 641401 509934 641420
rect 510358 642390 510392 642409
rect 510358 642318 510392 642330
rect 510358 642246 510392 642262
rect 510358 642174 510392 642194
rect 510358 642102 510392 642126
rect 510358 642030 510392 642058
rect 510358 641958 510392 641990
rect 510358 641888 510392 641922
rect 510358 641820 510392 641852
rect 510358 641752 510392 641780
rect 510358 641684 510392 641708
rect 510358 641616 510392 641636
rect 510358 641548 510392 641564
rect 510358 641480 510392 641492
rect 510358 641401 510392 641420
rect 510816 642390 510850 642409
rect 510816 642318 510850 642330
rect 510816 642246 510850 642262
rect 510816 642174 510850 642194
rect 510816 642102 510850 642126
rect 510816 642030 510850 642058
rect 510816 641958 510850 641990
rect 510816 641888 510850 641922
rect 510816 641820 510850 641852
rect 510816 641752 510850 641780
rect 510816 641684 510850 641708
rect 510816 641616 510850 641636
rect 510816 641548 510850 641564
rect 510816 641480 510850 641492
rect 510816 641401 510850 641420
rect 511274 642390 511308 642409
rect 511274 642318 511308 642330
rect 511274 642246 511308 642262
rect 511274 642174 511308 642194
rect 511274 642102 511308 642126
rect 511274 642030 511308 642058
rect 511274 641958 511308 641990
rect 511274 641888 511308 641922
rect 511274 641820 511308 641852
rect 511274 641752 511308 641780
rect 511274 641684 511308 641708
rect 511274 641616 511308 641636
rect 511274 641548 511308 641564
rect 511274 641480 511308 641492
rect 511274 641401 511308 641420
rect 511732 642390 511766 642409
rect 511732 642318 511766 642330
rect 511732 642246 511766 642262
rect 511732 642174 511766 642194
rect 511732 642102 511766 642126
rect 511732 642030 511766 642058
rect 511732 641958 511766 641990
rect 511732 641888 511766 641922
rect 511732 641820 511766 641852
rect 511732 641752 511766 641780
rect 511732 641684 511766 641708
rect 511732 641616 511766 641636
rect 511732 641548 511766 641564
rect 511732 641480 511766 641492
rect 511732 641401 511766 641420
rect 512190 642390 512224 642409
rect 512190 642318 512224 642330
rect 512190 642246 512224 642262
rect 512190 642174 512224 642194
rect 512190 642102 512224 642126
rect 512190 642030 512224 642058
rect 512190 641958 512224 641990
rect 512190 641888 512224 641922
rect 512190 641820 512224 641852
rect 512190 641752 512224 641780
rect 512190 641684 512224 641708
rect 512190 641616 512224 641636
rect 512190 641548 512224 641564
rect 512190 641480 512224 641492
rect 512190 641401 512224 641420
rect 512648 642390 512682 642409
rect 512648 642318 512682 642330
rect 512648 642246 512682 642262
rect 512648 642174 512682 642194
rect 512648 642102 512682 642126
rect 512648 642030 512682 642058
rect 512648 641958 512682 641990
rect 512648 641888 512682 641922
rect 512648 641820 512682 641852
rect 512648 641752 512682 641780
rect 512648 641684 512682 641708
rect 512648 641616 512682 641636
rect 512648 641548 512682 641564
rect 512648 641480 512682 641492
rect 512648 641401 512682 641420
rect 513106 642390 513140 642409
rect 513106 642318 513140 642330
rect 513106 642246 513140 642262
rect 513106 642174 513140 642194
rect 513106 642102 513140 642126
rect 513106 642030 513140 642058
rect 513106 641958 513140 641990
rect 513106 641888 513140 641922
rect 513106 641820 513140 641852
rect 513106 641752 513140 641780
rect 513106 641684 513140 641708
rect 513106 641616 513140 641636
rect 513106 641548 513140 641564
rect 513106 641480 513140 641492
rect 513106 641401 513140 641420
rect 513564 642390 513598 642409
rect 513564 642318 513598 642330
rect 513564 642246 513598 642262
rect 513564 642174 513598 642194
rect 513564 642102 513598 642126
rect 513564 642030 513598 642058
rect 513564 641958 513598 641990
rect 513564 641888 513598 641922
rect 513564 641820 513598 641852
rect 513564 641752 513598 641780
rect 513564 641684 513598 641708
rect 513564 641616 513598 641636
rect 513564 641548 513598 641564
rect 513564 641480 513598 641492
rect 513564 641401 513598 641420
rect 514022 642390 514056 642409
rect 514022 642318 514056 642330
rect 514022 642246 514056 642262
rect 514022 642174 514056 642194
rect 514022 642102 514056 642126
rect 514022 642030 514056 642058
rect 514022 641958 514056 641990
rect 514022 641888 514056 641922
rect 514022 641820 514056 641852
rect 514022 641752 514056 641780
rect 514022 641684 514056 641708
rect 514022 641616 514056 641636
rect 514022 641548 514056 641564
rect 514022 641480 514056 641492
rect 514022 641401 514056 641420
rect 514480 642390 514514 642409
rect 514480 642318 514514 642330
rect 514480 642246 514514 642262
rect 514480 642174 514514 642194
rect 514480 642102 514514 642126
rect 514480 642030 514514 642058
rect 514480 641958 514514 641990
rect 514480 641888 514514 641922
rect 514480 641820 514514 641852
rect 514480 641752 514514 641780
rect 514480 641684 514514 641708
rect 514480 641616 514514 641636
rect 514480 641548 514514 641564
rect 514480 641480 514514 641492
rect 514480 641401 514514 641420
rect 514938 642390 514972 642409
rect 514938 642318 514972 642330
rect 514938 642246 514972 642262
rect 514938 642174 514972 642194
rect 514938 642102 514972 642126
rect 514938 642030 514972 642058
rect 514938 641958 514972 641990
rect 514938 641888 514972 641922
rect 514938 641820 514972 641852
rect 514938 641752 514972 641780
rect 514938 641684 514972 641708
rect 514938 641616 514972 641636
rect 514938 641548 514972 641564
rect 514938 641480 514972 641492
rect 514938 641401 514972 641420
rect 515396 642390 515430 642409
rect 515396 642318 515430 642330
rect 515396 642246 515430 642262
rect 515396 642174 515430 642194
rect 515396 642102 515430 642126
rect 515396 642030 515430 642058
rect 515396 641958 515430 641990
rect 515396 641888 515430 641922
rect 515396 641820 515430 641852
rect 515396 641752 515430 641780
rect 515396 641684 515430 641708
rect 515396 641616 515430 641636
rect 515396 641548 515430 641564
rect 515396 641480 515430 641492
rect 515396 641401 515430 641420
rect 508114 641281 508153 641315
rect 508195 641281 508225 641315
rect 508263 641281 508297 641315
rect 508331 641281 508365 641315
rect 508403 641281 508433 641315
rect 508475 641281 508514 641315
rect 508572 641281 508611 641315
rect 508653 641281 508683 641315
rect 508721 641281 508755 641315
rect 508789 641281 508823 641315
rect 508861 641281 508891 641315
rect 508933 641281 508972 641315
rect 509030 641281 509069 641315
rect 509111 641281 509141 641315
rect 509179 641281 509213 641315
rect 509247 641281 509281 641315
rect 509319 641281 509349 641315
rect 509391 641281 509430 641315
rect 509488 641281 509527 641315
rect 509569 641281 509599 641315
rect 509637 641281 509671 641315
rect 509705 641281 509739 641315
rect 509777 641281 509807 641315
rect 509849 641281 509888 641315
rect 509946 641281 509985 641315
rect 510027 641281 510057 641315
rect 510095 641281 510129 641315
rect 510163 641281 510197 641315
rect 510235 641281 510265 641315
rect 510307 641281 510346 641315
rect 510404 641281 510443 641315
rect 510485 641281 510515 641315
rect 510553 641281 510587 641315
rect 510621 641281 510655 641315
rect 510693 641281 510723 641315
rect 510765 641281 510804 641315
rect 510862 641281 510901 641315
rect 510943 641281 510973 641315
rect 511011 641281 511045 641315
rect 511079 641281 511113 641315
rect 511151 641281 511181 641315
rect 511223 641281 511262 641315
rect 511320 641281 511359 641315
rect 511401 641281 511431 641315
rect 511469 641281 511503 641315
rect 511537 641281 511571 641315
rect 511609 641281 511639 641315
rect 511681 641281 511720 641315
rect 511778 641281 511817 641315
rect 511859 641281 511889 641315
rect 511927 641281 511961 641315
rect 511995 641281 512029 641315
rect 512067 641281 512097 641315
rect 512139 641281 512178 641315
rect 512236 641281 512275 641315
rect 512317 641281 512347 641315
rect 512385 641281 512419 641315
rect 512453 641281 512487 641315
rect 512525 641281 512555 641315
rect 512597 641281 512636 641315
rect 512694 641281 512733 641315
rect 512775 641281 512805 641315
rect 512843 641281 512877 641315
rect 512911 641281 512945 641315
rect 512983 641281 513013 641315
rect 513055 641281 513094 641315
rect 513152 641281 513191 641315
rect 513233 641281 513263 641315
rect 513301 641281 513335 641315
rect 513369 641281 513403 641315
rect 513441 641281 513471 641315
rect 513513 641281 513552 641315
rect 513610 641281 513649 641315
rect 513691 641281 513721 641315
rect 513759 641281 513793 641315
rect 513827 641281 513861 641315
rect 513899 641281 513929 641315
rect 513971 641281 514010 641315
rect 514068 641281 514107 641315
rect 514149 641281 514179 641315
rect 514217 641281 514251 641315
rect 514285 641281 514319 641315
rect 514357 641281 514387 641315
rect 514429 641281 514468 641315
rect 514526 641281 514565 641315
rect 514607 641281 514637 641315
rect 514675 641281 514709 641315
rect 514743 641281 514777 641315
rect 514815 641281 514845 641315
rect 514887 641281 514926 641315
rect 514984 641281 515023 641315
rect 515065 641281 515095 641315
rect 515133 641281 515167 641315
rect 515201 641281 515235 641315
rect 515273 641281 515303 641315
rect 515345 641281 515384 641315
rect 508068 641228 508102 641247
rect 508068 641156 508102 641168
rect 508068 641084 508102 641100
rect 508068 641012 508102 641032
rect 508068 640940 508102 640964
rect 508068 640868 508102 640896
rect 508068 640796 508102 640828
rect 508068 640726 508102 640760
rect 508068 640658 508102 640690
rect 508068 640590 508102 640618
rect 508068 640522 508102 640546
rect 508068 640454 508102 640474
rect 508068 640386 508102 640402
rect 508068 640318 508102 640330
rect 508068 640239 508102 640258
rect 508526 641228 508560 641247
rect 508526 641156 508560 641168
rect 508526 641084 508560 641100
rect 508526 641012 508560 641032
rect 508526 640940 508560 640964
rect 508526 640868 508560 640896
rect 508526 640796 508560 640828
rect 508526 640726 508560 640760
rect 508526 640658 508560 640690
rect 508526 640590 508560 640618
rect 508526 640522 508560 640546
rect 508526 640454 508560 640474
rect 508526 640386 508560 640402
rect 508526 640318 508560 640330
rect 508526 640239 508560 640258
rect 508984 641228 509018 641247
rect 508984 641156 509018 641168
rect 508984 641084 509018 641100
rect 508984 641012 509018 641032
rect 508984 640940 509018 640964
rect 508984 640868 509018 640896
rect 508984 640796 509018 640828
rect 508984 640726 509018 640760
rect 508984 640658 509018 640690
rect 508984 640590 509018 640618
rect 508984 640522 509018 640546
rect 508984 640454 509018 640474
rect 508984 640386 509018 640402
rect 508984 640318 509018 640330
rect 508984 640239 509018 640258
rect 509442 641228 509476 641247
rect 509442 641156 509476 641168
rect 509442 641084 509476 641100
rect 509442 641012 509476 641032
rect 509442 640940 509476 640964
rect 509442 640868 509476 640896
rect 509442 640796 509476 640828
rect 509442 640726 509476 640760
rect 509442 640658 509476 640690
rect 509442 640590 509476 640618
rect 509442 640522 509476 640546
rect 509442 640454 509476 640474
rect 509442 640386 509476 640402
rect 509442 640318 509476 640330
rect 509442 640239 509476 640258
rect 509900 641228 509934 641247
rect 509900 641156 509934 641168
rect 509900 641084 509934 641100
rect 509900 641012 509934 641032
rect 509900 640940 509934 640964
rect 509900 640868 509934 640896
rect 509900 640796 509934 640828
rect 509900 640726 509934 640760
rect 509900 640658 509934 640690
rect 509900 640590 509934 640618
rect 509900 640522 509934 640546
rect 509900 640454 509934 640474
rect 509900 640386 509934 640402
rect 509900 640318 509934 640330
rect 509900 640239 509934 640258
rect 510358 641228 510392 641247
rect 510358 641156 510392 641168
rect 510358 641084 510392 641100
rect 510358 641012 510392 641032
rect 510358 640940 510392 640964
rect 510358 640868 510392 640896
rect 510358 640796 510392 640828
rect 510358 640726 510392 640760
rect 510358 640658 510392 640690
rect 510358 640590 510392 640618
rect 510358 640522 510392 640546
rect 510358 640454 510392 640474
rect 510358 640386 510392 640402
rect 510358 640318 510392 640330
rect 510358 640239 510392 640258
rect 510816 641228 510850 641247
rect 510816 641156 510850 641168
rect 510816 641084 510850 641100
rect 510816 641012 510850 641032
rect 510816 640940 510850 640964
rect 510816 640868 510850 640896
rect 510816 640796 510850 640828
rect 510816 640726 510850 640760
rect 510816 640658 510850 640690
rect 510816 640590 510850 640618
rect 510816 640522 510850 640546
rect 510816 640454 510850 640474
rect 510816 640386 510850 640402
rect 510816 640318 510850 640330
rect 510816 640239 510850 640258
rect 511274 641228 511308 641247
rect 511274 641156 511308 641168
rect 511274 641084 511308 641100
rect 511274 641012 511308 641032
rect 511274 640940 511308 640964
rect 511274 640868 511308 640896
rect 511274 640796 511308 640828
rect 511274 640726 511308 640760
rect 511274 640658 511308 640690
rect 511274 640590 511308 640618
rect 511274 640522 511308 640546
rect 511274 640454 511308 640474
rect 511274 640386 511308 640402
rect 511274 640318 511308 640330
rect 511274 640239 511308 640258
rect 511732 641228 511766 641247
rect 511732 641156 511766 641168
rect 511732 641084 511766 641100
rect 511732 641012 511766 641032
rect 511732 640940 511766 640964
rect 511732 640868 511766 640896
rect 511732 640796 511766 640828
rect 511732 640726 511766 640760
rect 511732 640658 511766 640690
rect 511732 640590 511766 640618
rect 511732 640522 511766 640546
rect 511732 640454 511766 640474
rect 511732 640386 511766 640402
rect 511732 640318 511766 640330
rect 511732 640239 511766 640258
rect 512190 641228 512224 641247
rect 512190 641156 512224 641168
rect 512190 641084 512224 641100
rect 512190 641012 512224 641032
rect 512190 640940 512224 640964
rect 512190 640868 512224 640896
rect 512190 640796 512224 640828
rect 512190 640726 512224 640760
rect 512190 640658 512224 640690
rect 512190 640590 512224 640618
rect 512190 640522 512224 640546
rect 512190 640454 512224 640474
rect 512190 640386 512224 640402
rect 512190 640318 512224 640330
rect 512190 640239 512224 640258
rect 512648 641228 512682 641247
rect 512648 641156 512682 641168
rect 512648 641084 512682 641100
rect 512648 641012 512682 641032
rect 512648 640940 512682 640964
rect 512648 640868 512682 640896
rect 512648 640796 512682 640828
rect 512648 640726 512682 640760
rect 512648 640658 512682 640690
rect 512648 640590 512682 640618
rect 512648 640522 512682 640546
rect 512648 640454 512682 640474
rect 512648 640386 512682 640402
rect 512648 640318 512682 640330
rect 512648 640239 512682 640258
rect 513106 641228 513140 641247
rect 513106 641156 513140 641168
rect 513106 641084 513140 641100
rect 513106 641012 513140 641032
rect 513106 640940 513140 640964
rect 513106 640868 513140 640896
rect 513106 640796 513140 640828
rect 513106 640726 513140 640760
rect 513106 640658 513140 640690
rect 513106 640590 513140 640618
rect 513106 640522 513140 640546
rect 513106 640454 513140 640474
rect 513106 640386 513140 640402
rect 513106 640318 513140 640330
rect 513106 640239 513140 640258
rect 513564 641228 513598 641247
rect 513564 641156 513598 641168
rect 513564 641084 513598 641100
rect 513564 641012 513598 641032
rect 513564 640940 513598 640964
rect 513564 640868 513598 640896
rect 513564 640796 513598 640828
rect 513564 640726 513598 640760
rect 513564 640658 513598 640690
rect 513564 640590 513598 640618
rect 513564 640522 513598 640546
rect 513564 640454 513598 640474
rect 513564 640386 513598 640402
rect 513564 640318 513598 640330
rect 513564 640239 513598 640258
rect 514022 641228 514056 641247
rect 514022 641156 514056 641168
rect 514022 641084 514056 641100
rect 514022 641012 514056 641032
rect 514022 640940 514056 640964
rect 514022 640868 514056 640896
rect 514022 640796 514056 640828
rect 514022 640726 514056 640760
rect 514022 640658 514056 640690
rect 514022 640590 514056 640618
rect 514022 640522 514056 640546
rect 514022 640454 514056 640474
rect 514022 640386 514056 640402
rect 514022 640318 514056 640330
rect 514022 640239 514056 640258
rect 514480 641228 514514 641247
rect 514480 641156 514514 641168
rect 514480 641084 514514 641100
rect 514480 641012 514514 641032
rect 514480 640940 514514 640964
rect 514480 640868 514514 640896
rect 514480 640796 514514 640828
rect 514480 640726 514514 640760
rect 514480 640658 514514 640690
rect 514480 640590 514514 640618
rect 514480 640522 514514 640546
rect 514480 640454 514514 640474
rect 514480 640386 514514 640402
rect 514480 640318 514514 640330
rect 514480 640239 514514 640258
rect 514938 641228 514972 641247
rect 514938 641156 514972 641168
rect 514938 641084 514972 641100
rect 514938 641012 514972 641032
rect 514938 640940 514972 640964
rect 514938 640868 514972 640896
rect 514938 640796 514972 640828
rect 514938 640726 514972 640760
rect 514938 640658 514972 640690
rect 514938 640590 514972 640618
rect 514938 640522 514972 640546
rect 514938 640454 514972 640474
rect 514938 640386 514972 640402
rect 514938 640318 514972 640330
rect 514938 640239 514972 640258
rect 515396 641228 515430 641247
rect 515396 641156 515430 641168
rect 515396 641084 515430 641100
rect 515396 641012 515430 641032
rect 515396 640940 515430 640964
rect 515396 640868 515430 640896
rect 515396 640796 515430 640828
rect 515396 640726 515430 640760
rect 515396 640658 515430 640690
rect 515396 640590 515430 640618
rect 515396 640522 515430 640546
rect 515396 640454 515430 640474
rect 515396 640386 515430 640402
rect 515396 640318 515430 640330
rect 515396 640239 515430 640258
rect 507828 640128 507966 640182
rect 515532 640182 515550 642528
rect 515652 641280 515670 642528
rect 516828 642528 516966 642582
rect 515818 642443 515857 642477
rect 515899 642443 515929 642477
rect 515967 642443 516001 642477
rect 516035 642443 516069 642477
rect 516107 642443 516137 642477
rect 516179 642443 516218 642477
rect 516276 642443 516315 642477
rect 516357 642443 516387 642477
rect 516425 642443 516459 642477
rect 516493 642443 516527 642477
rect 516565 642443 516595 642477
rect 516637 642443 516676 642477
rect 515772 642390 515806 642409
rect 515772 642318 515806 642330
rect 515772 642246 515806 642262
rect 515772 642174 515806 642194
rect 515772 642102 515806 642126
rect 515772 642030 515806 642058
rect 515772 641958 515806 641990
rect 515772 641888 515806 641922
rect 515772 641820 515806 641852
rect 515772 641752 515806 641780
rect 515772 641684 515806 641708
rect 515772 641616 515806 641636
rect 515772 641548 515806 641564
rect 515772 641480 515806 641492
rect 515772 641401 515806 641420
rect 516230 642390 516264 642409
rect 516230 642318 516264 642330
rect 516230 642246 516264 642262
rect 516230 642174 516264 642194
rect 516230 642102 516264 642126
rect 516230 642030 516264 642058
rect 516230 641958 516264 641990
rect 516230 641888 516264 641922
rect 516230 641820 516264 641852
rect 516230 641752 516264 641780
rect 516230 641684 516264 641708
rect 516230 641616 516264 641636
rect 516230 641548 516264 641564
rect 516230 641480 516264 641492
rect 516230 641401 516264 641420
rect 516688 642390 516722 642409
rect 516688 642318 516722 642330
rect 516688 642246 516722 642262
rect 516688 642174 516722 642194
rect 516688 642102 516722 642126
rect 516688 642030 516722 642058
rect 516688 641958 516722 641990
rect 516688 641888 516722 641922
rect 516688 641820 516722 641852
rect 516688 641752 516722 641780
rect 516688 641684 516722 641708
rect 516688 641616 516722 641636
rect 516688 641548 516722 641564
rect 516688 641480 516722 641492
rect 516688 641401 516722 641420
rect 516828 641280 516846 642528
rect 515652 641262 516846 641280
rect 515652 641160 515722 641262
rect 516776 641160 516846 641262
rect 515652 641094 516846 641160
rect 515652 640502 515722 641094
rect 515652 640182 515722 640324
rect 515532 640176 515722 640182
rect 516776 640182 516846 641094
rect 516948 640182 516966 642528
rect 516776 640176 516966 640182
rect 515532 640128 516966 640176
rect 507828 640110 516966 640128
rect 507828 640008 507846 640110
rect 507948 640008 507994 640110
rect 516800 640008 516846 640110
rect 516948 640008 516966 640110
rect 507828 639990 516966 640008
<< viali >>
rect 507879 645376 507913 645410
rect 507879 645304 507913 645338
rect 507879 645232 507913 645266
rect 507880 643744 507914 643778
rect 507880 643672 507914 643706
rect 507880 643600 507914 643634
rect 508068 645462 508102 645488
rect 508068 645454 508102 645462
rect 508068 645394 508102 645416
rect 508068 645382 508102 645394
rect 508068 645326 508102 645344
rect 508068 645310 508102 645326
rect 508068 645258 508102 645272
rect 508068 645238 508102 645258
rect 508068 645190 508102 645200
rect 508068 645166 508102 645190
rect 508068 645122 508102 645128
rect 508068 645094 508102 645122
rect 508068 645054 508102 645056
rect 508068 645022 508102 645054
rect 508068 644952 508102 644984
rect 508068 644950 508102 644952
rect 508068 644884 508102 644912
rect 508068 644878 508102 644884
rect 508068 644816 508102 644840
rect 508068 644806 508102 644816
rect 508068 644748 508102 644768
rect 508068 644734 508102 644748
rect 508068 644680 508102 644696
rect 508068 644662 508102 644680
rect 508068 644612 508102 644624
rect 508068 644590 508102 644612
rect 508068 644544 508102 644552
rect 508068 644518 508102 644544
rect 508526 645462 508560 645488
rect 508526 645454 508560 645462
rect 508526 645394 508560 645416
rect 508526 645382 508560 645394
rect 508526 645326 508560 645344
rect 508526 645310 508560 645326
rect 508526 645258 508560 645272
rect 508526 645238 508560 645258
rect 508526 645190 508560 645200
rect 508526 645166 508560 645190
rect 508526 645122 508560 645128
rect 508526 645094 508560 645122
rect 508526 645054 508560 645056
rect 508526 645022 508560 645054
rect 508526 644952 508560 644984
rect 508526 644950 508560 644952
rect 508526 644884 508560 644912
rect 508526 644878 508560 644884
rect 508526 644816 508560 644840
rect 508526 644806 508560 644816
rect 508526 644748 508560 644768
rect 508526 644734 508560 644748
rect 508526 644680 508560 644696
rect 508526 644662 508560 644680
rect 508526 644612 508560 644624
rect 508526 644590 508560 644612
rect 508526 644544 508560 644552
rect 508526 644518 508560 644544
rect 508984 645462 509018 645488
rect 508984 645454 509018 645462
rect 508984 645394 509018 645416
rect 508984 645382 509018 645394
rect 508984 645326 509018 645344
rect 508984 645310 509018 645326
rect 508984 645258 509018 645272
rect 508984 645238 509018 645258
rect 508984 645190 509018 645200
rect 508984 645166 509018 645190
rect 508984 645122 509018 645128
rect 508984 645094 509018 645122
rect 508984 645054 509018 645056
rect 508984 645022 509018 645054
rect 508984 644952 509018 644984
rect 508984 644950 509018 644952
rect 508984 644884 509018 644912
rect 508984 644878 509018 644884
rect 508984 644816 509018 644840
rect 508984 644806 509018 644816
rect 508984 644748 509018 644768
rect 508984 644734 509018 644748
rect 508984 644680 509018 644696
rect 508984 644662 509018 644680
rect 508984 644612 509018 644624
rect 508984 644590 509018 644612
rect 508984 644544 509018 644552
rect 508984 644518 509018 644544
rect 509442 645462 509476 645488
rect 509442 645454 509476 645462
rect 509442 645394 509476 645416
rect 509442 645382 509476 645394
rect 509442 645326 509476 645344
rect 509442 645310 509476 645326
rect 509442 645258 509476 645272
rect 509442 645238 509476 645258
rect 509442 645190 509476 645200
rect 509442 645166 509476 645190
rect 509442 645122 509476 645128
rect 509442 645094 509476 645122
rect 509442 645054 509476 645056
rect 509442 645022 509476 645054
rect 509442 644952 509476 644984
rect 509442 644950 509476 644952
rect 509442 644884 509476 644912
rect 509442 644878 509476 644884
rect 509442 644816 509476 644840
rect 509442 644806 509476 644816
rect 509442 644748 509476 644768
rect 509442 644734 509476 644748
rect 509442 644680 509476 644696
rect 509442 644662 509476 644680
rect 509442 644612 509476 644624
rect 509442 644590 509476 644612
rect 509442 644544 509476 644552
rect 509442 644518 509476 644544
rect 509900 645462 509934 645488
rect 509900 645454 509934 645462
rect 509900 645394 509934 645416
rect 509900 645382 509934 645394
rect 509900 645326 509934 645344
rect 509900 645310 509934 645326
rect 509900 645258 509934 645272
rect 509900 645238 509934 645258
rect 509900 645190 509934 645200
rect 509900 645166 509934 645190
rect 509900 645122 509934 645128
rect 509900 645094 509934 645122
rect 509900 645054 509934 645056
rect 509900 645022 509934 645054
rect 509900 644952 509934 644984
rect 509900 644950 509934 644952
rect 509900 644884 509934 644912
rect 509900 644878 509934 644884
rect 509900 644816 509934 644840
rect 509900 644806 509934 644816
rect 509900 644748 509934 644768
rect 509900 644734 509934 644748
rect 509900 644680 509934 644696
rect 509900 644662 509934 644680
rect 509900 644612 509934 644624
rect 509900 644590 509934 644612
rect 509900 644544 509934 644552
rect 509900 644518 509934 644544
rect 510358 645462 510392 645488
rect 510358 645454 510392 645462
rect 510358 645394 510392 645416
rect 510358 645382 510392 645394
rect 510358 645326 510392 645344
rect 510358 645310 510392 645326
rect 510358 645258 510392 645272
rect 510358 645238 510392 645258
rect 510358 645190 510392 645200
rect 510358 645166 510392 645190
rect 510358 645122 510392 645128
rect 510358 645094 510392 645122
rect 510358 645054 510392 645056
rect 510358 645022 510392 645054
rect 510358 644952 510392 644984
rect 510358 644950 510392 644952
rect 510358 644884 510392 644912
rect 510358 644878 510392 644884
rect 510358 644816 510392 644840
rect 510358 644806 510392 644816
rect 510358 644748 510392 644768
rect 510358 644734 510392 644748
rect 510358 644680 510392 644696
rect 510358 644662 510392 644680
rect 510358 644612 510392 644624
rect 510358 644590 510392 644612
rect 510358 644544 510392 644552
rect 510358 644518 510392 644544
rect 510816 645462 510850 645488
rect 510816 645454 510850 645462
rect 510816 645394 510850 645416
rect 510816 645382 510850 645394
rect 510816 645326 510850 645344
rect 510816 645310 510850 645326
rect 510816 645258 510850 645272
rect 510816 645238 510850 645258
rect 510816 645190 510850 645200
rect 510816 645166 510850 645190
rect 510816 645122 510850 645128
rect 510816 645094 510850 645122
rect 510816 645054 510850 645056
rect 510816 645022 510850 645054
rect 510816 644952 510850 644984
rect 510816 644950 510850 644952
rect 510816 644884 510850 644912
rect 510816 644878 510850 644884
rect 510816 644816 510850 644840
rect 510816 644806 510850 644816
rect 510816 644748 510850 644768
rect 510816 644734 510850 644748
rect 510816 644680 510850 644696
rect 510816 644662 510850 644680
rect 510816 644612 510850 644624
rect 510816 644590 510850 644612
rect 510816 644544 510850 644552
rect 510816 644518 510850 644544
rect 511274 645462 511308 645488
rect 511274 645454 511308 645462
rect 511274 645394 511308 645416
rect 511274 645382 511308 645394
rect 511274 645326 511308 645344
rect 511274 645310 511308 645326
rect 511274 645258 511308 645272
rect 511274 645238 511308 645258
rect 511274 645190 511308 645200
rect 511274 645166 511308 645190
rect 511274 645122 511308 645128
rect 511274 645094 511308 645122
rect 511274 645054 511308 645056
rect 511274 645022 511308 645054
rect 511274 644952 511308 644984
rect 511274 644950 511308 644952
rect 511274 644884 511308 644912
rect 511274 644878 511308 644884
rect 511274 644816 511308 644840
rect 511274 644806 511308 644816
rect 511274 644748 511308 644768
rect 511274 644734 511308 644748
rect 511274 644680 511308 644696
rect 511274 644662 511308 644680
rect 511274 644612 511308 644624
rect 511274 644590 511308 644612
rect 511274 644544 511308 644552
rect 511274 644518 511308 644544
rect 511732 645462 511766 645488
rect 511732 645454 511766 645462
rect 511732 645394 511766 645416
rect 511732 645382 511766 645394
rect 511732 645326 511766 645344
rect 511732 645310 511766 645326
rect 511732 645258 511766 645272
rect 511732 645238 511766 645258
rect 511732 645190 511766 645200
rect 511732 645166 511766 645190
rect 511732 645122 511766 645128
rect 511732 645094 511766 645122
rect 511732 645054 511766 645056
rect 511732 645022 511766 645054
rect 511732 644952 511766 644984
rect 511732 644950 511766 644952
rect 511732 644884 511766 644912
rect 511732 644878 511766 644884
rect 511732 644816 511766 644840
rect 511732 644806 511766 644816
rect 511732 644748 511766 644768
rect 511732 644734 511766 644748
rect 511732 644680 511766 644696
rect 511732 644662 511766 644680
rect 511732 644612 511766 644624
rect 511732 644590 511766 644612
rect 511732 644544 511766 644552
rect 511732 644518 511766 644544
rect 512190 645462 512224 645488
rect 512190 645454 512224 645462
rect 512190 645394 512224 645416
rect 512190 645382 512224 645394
rect 512190 645326 512224 645344
rect 512190 645310 512224 645326
rect 512190 645258 512224 645272
rect 512190 645238 512224 645258
rect 512190 645190 512224 645200
rect 512190 645166 512224 645190
rect 512190 645122 512224 645128
rect 512190 645094 512224 645122
rect 512190 645054 512224 645056
rect 512190 645022 512224 645054
rect 512190 644952 512224 644984
rect 512190 644950 512224 644952
rect 512190 644884 512224 644912
rect 512190 644878 512224 644884
rect 512190 644816 512224 644840
rect 512190 644806 512224 644816
rect 512190 644748 512224 644768
rect 512190 644734 512224 644748
rect 512190 644680 512224 644696
rect 512190 644662 512224 644680
rect 512190 644612 512224 644624
rect 512190 644590 512224 644612
rect 512190 644544 512224 644552
rect 512190 644518 512224 644544
rect 512648 645462 512682 645488
rect 512648 645454 512682 645462
rect 512648 645394 512682 645416
rect 512648 645382 512682 645394
rect 512648 645326 512682 645344
rect 512648 645310 512682 645326
rect 512648 645258 512682 645272
rect 512648 645238 512682 645258
rect 512648 645190 512682 645200
rect 512648 645166 512682 645190
rect 512648 645122 512682 645128
rect 512648 645094 512682 645122
rect 512648 645054 512682 645056
rect 512648 645022 512682 645054
rect 512648 644952 512682 644984
rect 512648 644950 512682 644952
rect 512648 644884 512682 644912
rect 512648 644878 512682 644884
rect 512648 644816 512682 644840
rect 512648 644806 512682 644816
rect 512648 644748 512682 644768
rect 512648 644734 512682 644748
rect 512648 644680 512682 644696
rect 512648 644662 512682 644680
rect 512648 644612 512682 644624
rect 512648 644590 512682 644612
rect 512648 644544 512682 644552
rect 512648 644518 512682 644544
rect 513106 645462 513140 645488
rect 513106 645454 513140 645462
rect 513106 645394 513140 645416
rect 513106 645382 513140 645394
rect 513106 645326 513140 645344
rect 513106 645310 513140 645326
rect 513106 645258 513140 645272
rect 513106 645238 513140 645258
rect 513106 645190 513140 645200
rect 513106 645166 513140 645190
rect 513106 645122 513140 645128
rect 513106 645094 513140 645122
rect 513106 645054 513140 645056
rect 513106 645022 513140 645054
rect 513106 644952 513140 644984
rect 513106 644950 513140 644952
rect 513106 644884 513140 644912
rect 513106 644878 513140 644884
rect 513106 644816 513140 644840
rect 513106 644806 513140 644816
rect 513106 644748 513140 644768
rect 513106 644734 513140 644748
rect 513106 644680 513140 644696
rect 513106 644662 513140 644680
rect 513106 644612 513140 644624
rect 513106 644590 513140 644612
rect 513106 644544 513140 644552
rect 513106 644518 513140 644544
rect 513564 645462 513598 645488
rect 513564 645454 513598 645462
rect 513564 645394 513598 645416
rect 513564 645382 513598 645394
rect 513564 645326 513598 645344
rect 513564 645310 513598 645326
rect 513564 645258 513598 645272
rect 513564 645238 513598 645258
rect 513564 645190 513598 645200
rect 513564 645166 513598 645190
rect 513564 645122 513598 645128
rect 513564 645094 513598 645122
rect 513564 645054 513598 645056
rect 513564 645022 513598 645054
rect 513564 644952 513598 644984
rect 513564 644950 513598 644952
rect 513564 644884 513598 644912
rect 513564 644878 513598 644884
rect 513564 644816 513598 644840
rect 513564 644806 513598 644816
rect 513564 644748 513598 644768
rect 513564 644734 513598 644748
rect 513564 644680 513598 644696
rect 513564 644662 513598 644680
rect 513564 644612 513598 644624
rect 513564 644590 513598 644612
rect 513564 644544 513598 644552
rect 513564 644518 513598 644544
rect 514022 645462 514056 645488
rect 514022 645454 514056 645462
rect 514022 645394 514056 645416
rect 514022 645382 514056 645394
rect 514022 645326 514056 645344
rect 514022 645310 514056 645326
rect 514022 645258 514056 645272
rect 514022 645238 514056 645258
rect 514022 645190 514056 645200
rect 514022 645166 514056 645190
rect 514022 645122 514056 645128
rect 514022 645094 514056 645122
rect 514022 645054 514056 645056
rect 514022 645022 514056 645054
rect 514022 644952 514056 644984
rect 514022 644950 514056 644952
rect 514022 644884 514056 644912
rect 514022 644878 514056 644884
rect 514022 644816 514056 644840
rect 514022 644806 514056 644816
rect 514022 644748 514056 644768
rect 514022 644734 514056 644748
rect 514022 644680 514056 644696
rect 514022 644662 514056 644680
rect 514022 644612 514056 644624
rect 514022 644590 514056 644612
rect 514022 644544 514056 644552
rect 514022 644518 514056 644544
rect 514480 645462 514514 645488
rect 514480 645454 514514 645462
rect 514480 645394 514514 645416
rect 514480 645382 514514 645394
rect 514480 645326 514514 645344
rect 514480 645310 514514 645326
rect 514480 645258 514514 645272
rect 514480 645238 514514 645258
rect 514480 645190 514514 645200
rect 514480 645166 514514 645190
rect 514480 645122 514514 645128
rect 514480 645094 514514 645122
rect 514480 645054 514514 645056
rect 514480 645022 514514 645054
rect 514480 644952 514514 644984
rect 514480 644950 514514 644952
rect 514480 644884 514514 644912
rect 514480 644878 514514 644884
rect 514480 644816 514514 644840
rect 514480 644806 514514 644816
rect 514480 644748 514514 644768
rect 514480 644734 514514 644748
rect 514480 644680 514514 644696
rect 514480 644662 514514 644680
rect 514480 644612 514514 644624
rect 514480 644590 514514 644612
rect 514480 644544 514514 644552
rect 514480 644518 514514 644544
rect 514938 645462 514972 645488
rect 514938 645454 514972 645462
rect 514938 645394 514972 645416
rect 514938 645382 514972 645394
rect 514938 645326 514972 645344
rect 514938 645310 514972 645326
rect 514938 645258 514972 645272
rect 514938 645238 514972 645258
rect 514938 645190 514972 645200
rect 514938 645166 514972 645190
rect 514938 645122 514972 645128
rect 514938 645094 514972 645122
rect 514938 645054 514972 645056
rect 514938 645022 514972 645054
rect 514938 644952 514972 644984
rect 514938 644950 514972 644952
rect 514938 644884 514972 644912
rect 514938 644878 514972 644884
rect 514938 644816 514972 644840
rect 514938 644806 514972 644816
rect 514938 644748 514972 644768
rect 514938 644734 514972 644748
rect 514938 644680 514972 644696
rect 514938 644662 514972 644680
rect 514938 644612 514972 644624
rect 514938 644590 514972 644612
rect 514938 644544 514972 644552
rect 514938 644518 514972 644544
rect 515396 645462 515430 645488
rect 515396 645454 515430 645462
rect 515396 645394 515430 645416
rect 515396 645382 515430 645394
rect 515396 645326 515430 645344
rect 515396 645310 515430 645326
rect 515396 645258 515430 645272
rect 515396 645238 515430 645258
rect 515396 645190 515430 645200
rect 515396 645166 515430 645190
rect 515396 645122 515430 645128
rect 515396 645094 515430 645122
rect 515396 645054 515430 645056
rect 515396 645022 515430 645054
rect 515396 644952 515430 644984
rect 515396 644950 515430 644952
rect 515396 644884 515430 644912
rect 515396 644878 515430 644884
rect 515396 644816 515430 644840
rect 515396 644806 515430 644816
rect 515396 644748 515430 644768
rect 515396 644734 515430 644748
rect 515396 644680 515430 644696
rect 515396 644662 515430 644680
rect 515396 644612 515430 644624
rect 515396 644590 515430 644612
rect 515396 644544 515430 644552
rect 515396 644518 515430 644544
rect 508153 644422 508161 644456
rect 508161 644422 508187 644456
rect 508225 644422 508229 644456
rect 508229 644422 508259 644456
rect 508297 644422 508331 644456
rect 508369 644422 508399 644456
rect 508399 644422 508403 644456
rect 508441 644422 508467 644456
rect 508467 644422 508475 644456
rect 508611 644422 508619 644456
rect 508619 644422 508645 644456
rect 508683 644422 508687 644456
rect 508687 644422 508717 644456
rect 508755 644422 508789 644456
rect 508827 644422 508857 644456
rect 508857 644422 508861 644456
rect 508899 644422 508925 644456
rect 508925 644422 508933 644456
rect 509069 644422 509077 644456
rect 509077 644422 509103 644456
rect 509141 644422 509145 644456
rect 509145 644422 509175 644456
rect 509213 644422 509247 644456
rect 509285 644422 509315 644456
rect 509315 644422 509319 644456
rect 509357 644422 509383 644456
rect 509383 644422 509391 644456
rect 509527 644422 509535 644456
rect 509535 644422 509561 644456
rect 509599 644422 509603 644456
rect 509603 644422 509633 644456
rect 509671 644422 509705 644456
rect 509743 644422 509773 644456
rect 509773 644422 509777 644456
rect 509815 644422 509841 644456
rect 509841 644422 509849 644456
rect 509985 644422 509993 644456
rect 509993 644422 510019 644456
rect 510057 644422 510061 644456
rect 510061 644422 510091 644456
rect 510129 644422 510163 644456
rect 510201 644422 510231 644456
rect 510231 644422 510235 644456
rect 510273 644422 510299 644456
rect 510299 644422 510307 644456
rect 510443 644422 510451 644456
rect 510451 644422 510477 644456
rect 510515 644422 510519 644456
rect 510519 644422 510549 644456
rect 510587 644422 510621 644456
rect 510659 644422 510689 644456
rect 510689 644422 510693 644456
rect 510731 644422 510757 644456
rect 510757 644422 510765 644456
rect 510901 644422 510909 644456
rect 510909 644422 510935 644456
rect 510973 644422 510977 644456
rect 510977 644422 511007 644456
rect 511045 644422 511079 644456
rect 511117 644422 511147 644456
rect 511147 644422 511151 644456
rect 511189 644422 511215 644456
rect 511215 644422 511223 644456
rect 511359 644422 511367 644456
rect 511367 644422 511393 644456
rect 511431 644422 511435 644456
rect 511435 644422 511465 644456
rect 511503 644422 511537 644456
rect 511575 644422 511605 644456
rect 511605 644422 511609 644456
rect 511647 644422 511673 644456
rect 511673 644422 511681 644456
rect 511817 644422 511825 644456
rect 511825 644422 511851 644456
rect 511889 644422 511893 644456
rect 511893 644422 511923 644456
rect 511961 644422 511995 644456
rect 512033 644422 512063 644456
rect 512063 644422 512067 644456
rect 512105 644422 512131 644456
rect 512131 644422 512139 644456
rect 512275 644422 512283 644456
rect 512283 644422 512309 644456
rect 512347 644422 512351 644456
rect 512351 644422 512381 644456
rect 512419 644422 512453 644456
rect 512491 644422 512521 644456
rect 512521 644422 512525 644456
rect 512563 644422 512589 644456
rect 512589 644422 512597 644456
rect 512733 644422 512741 644456
rect 512741 644422 512767 644456
rect 512805 644422 512809 644456
rect 512809 644422 512839 644456
rect 512877 644422 512911 644456
rect 512949 644422 512979 644456
rect 512979 644422 512983 644456
rect 513021 644422 513047 644456
rect 513047 644422 513055 644456
rect 513191 644422 513199 644456
rect 513199 644422 513225 644456
rect 513263 644422 513267 644456
rect 513267 644422 513297 644456
rect 513335 644422 513369 644456
rect 513407 644422 513437 644456
rect 513437 644422 513441 644456
rect 513479 644422 513505 644456
rect 513505 644422 513513 644456
rect 513649 644422 513657 644456
rect 513657 644422 513683 644456
rect 513721 644422 513725 644456
rect 513725 644422 513755 644456
rect 513793 644422 513827 644456
rect 513865 644422 513895 644456
rect 513895 644422 513899 644456
rect 513937 644422 513963 644456
rect 513963 644422 513971 644456
rect 514107 644422 514115 644456
rect 514115 644422 514141 644456
rect 514179 644422 514183 644456
rect 514183 644422 514213 644456
rect 514251 644422 514285 644456
rect 514323 644422 514353 644456
rect 514353 644422 514357 644456
rect 514395 644422 514421 644456
rect 514421 644422 514429 644456
rect 514565 644422 514573 644456
rect 514573 644422 514599 644456
rect 514637 644422 514641 644456
rect 514641 644422 514671 644456
rect 514709 644422 514743 644456
rect 514781 644422 514811 644456
rect 514811 644422 514815 644456
rect 514853 644422 514879 644456
rect 514879 644422 514887 644456
rect 515023 644422 515031 644456
rect 515031 644422 515057 644456
rect 515095 644422 515099 644456
rect 515099 644422 515129 644456
rect 515167 644422 515201 644456
rect 515239 644422 515269 644456
rect 515269 644422 515273 644456
rect 515311 644422 515337 644456
rect 515337 644422 515345 644456
rect 508068 644296 508102 644322
rect 508068 644288 508102 644296
rect 508068 644228 508102 644250
rect 508068 644216 508102 644228
rect 508068 644160 508102 644178
rect 508068 644144 508102 644160
rect 508068 644092 508102 644106
rect 508068 644072 508102 644092
rect 508068 644024 508102 644034
rect 508068 644000 508102 644024
rect 508068 643956 508102 643962
rect 508068 643928 508102 643956
rect 508068 643888 508102 643890
rect 508068 643856 508102 643888
rect 508068 643786 508102 643818
rect 508068 643784 508102 643786
rect 508068 643718 508102 643746
rect 508068 643712 508102 643718
rect 508068 643650 508102 643674
rect 508068 643640 508102 643650
rect 508068 643582 508102 643602
rect 508068 643568 508102 643582
rect 508068 643514 508102 643530
rect 508068 643496 508102 643514
rect 508068 643446 508102 643458
rect 508068 643424 508102 643446
rect 508068 643378 508102 643386
rect 508068 643352 508102 643378
rect 508526 644296 508560 644322
rect 508526 644288 508560 644296
rect 508526 644228 508560 644250
rect 508526 644216 508560 644228
rect 508526 644160 508560 644178
rect 508526 644144 508560 644160
rect 508526 644092 508560 644106
rect 508526 644072 508560 644092
rect 508526 644024 508560 644034
rect 508526 644000 508560 644024
rect 508526 643956 508560 643962
rect 508526 643928 508560 643956
rect 508526 643888 508560 643890
rect 508526 643856 508560 643888
rect 508526 643786 508560 643818
rect 508526 643784 508560 643786
rect 508526 643718 508560 643746
rect 508526 643712 508560 643718
rect 508526 643650 508560 643674
rect 508526 643640 508560 643650
rect 508526 643582 508560 643602
rect 508526 643568 508560 643582
rect 508526 643514 508560 643530
rect 508526 643496 508560 643514
rect 508526 643446 508560 643458
rect 508526 643424 508560 643446
rect 508526 643378 508560 643386
rect 508526 643352 508560 643378
rect 508984 644296 509018 644322
rect 508984 644288 509018 644296
rect 508984 644228 509018 644250
rect 508984 644216 509018 644228
rect 508984 644160 509018 644178
rect 508984 644144 509018 644160
rect 508984 644092 509018 644106
rect 508984 644072 509018 644092
rect 508984 644024 509018 644034
rect 508984 644000 509018 644024
rect 508984 643956 509018 643962
rect 508984 643928 509018 643956
rect 508984 643888 509018 643890
rect 508984 643856 509018 643888
rect 508984 643786 509018 643818
rect 508984 643784 509018 643786
rect 508984 643718 509018 643746
rect 508984 643712 509018 643718
rect 508984 643650 509018 643674
rect 508984 643640 509018 643650
rect 508984 643582 509018 643602
rect 508984 643568 509018 643582
rect 508984 643514 509018 643530
rect 508984 643496 509018 643514
rect 508984 643446 509018 643458
rect 508984 643424 509018 643446
rect 508984 643378 509018 643386
rect 508984 643352 509018 643378
rect 509442 644296 509476 644322
rect 509442 644288 509476 644296
rect 509442 644228 509476 644250
rect 509442 644216 509476 644228
rect 509442 644160 509476 644178
rect 509442 644144 509476 644160
rect 509442 644092 509476 644106
rect 509442 644072 509476 644092
rect 509442 644024 509476 644034
rect 509442 644000 509476 644024
rect 509442 643956 509476 643962
rect 509442 643928 509476 643956
rect 509442 643888 509476 643890
rect 509442 643856 509476 643888
rect 509442 643786 509476 643818
rect 509442 643784 509476 643786
rect 509442 643718 509476 643746
rect 509442 643712 509476 643718
rect 509442 643650 509476 643674
rect 509442 643640 509476 643650
rect 509442 643582 509476 643602
rect 509442 643568 509476 643582
rect 509442 643514 509476 643530
rect 509442 643496 509476 643514
rect 509442 643446 509476 643458
rect 509442 643424 509476 643446
rect 509442 643378 509476 643386
rect 509442 643352 509476 643378
rect 509900 644296 509934 644322
rect 509900 644288 509934 644296
rect 509900 644228 509934 644250
rect 509900 644216 509934 644228
rect 509900 644160 509934 644178
rect 509900 644144 509934 644160
rect 509900 644092 509934 644106
rect 509900 644072 509934 644092
rect 509900 644024 509934 644034
rect 509900 644000 509934 644024
rect 509900 643956 509934 643962
rect 509900 643928 509934 643956
rect 509900 643888 509934 643890
rect 509900 643856 509934 643888
rect 509900 643786 509934 643818
rect 509900 643784 509934 643786
rect 509900 643718 509934 643746
rect 509900 643712 509934 643718
rect 509900 643650 509934 643674
rect 509900 643640 509934 643650
rect 509900 643582 509934 643602
rect 509900 643568 509934 643582
rect 509900 643514 509934 643530
rect 509900 643496 509934 643514
rect 509900 643446 509934 643458
rect 509900 643424 509934 643446
rect 509900 643378 509934 643386
rect 509900 643352 509934 643378
rect 510358 644296 510392 644322
rect 510358 644288 510392 644296
rect 510358 644228 510392 644250
rect 510358 644216 510392 644228
rect 510358 644160 510392 644178
rect 510358 644144 510392 644160
rect 510358 644092 510392 644106
rect 510358 644072 510392 644092
rect 510358 644024 510392 644034
rect 510358 644000 510392 644024
rect 510358 643956 510392 643962
rect 510358 643928 510392 643956
rect 510358 643888 510392 643890
rect 510358 643856 510392 643888
rect 510358 643786 510392 643818
rect 510358 643784 510392 643786
rect 510358 643718 510392 643746
rect 510358 643712 510392 643718
rect 510358 643650 510392 643674
rect 510358 643640 510392 643650
rect 510358 643582 510392 643602
rect 510358 643568 510392 643582
rect 510358 643514 510392 643530
rect 510358 643496 510392 643514
rect 510358 643446 510392 643458
rect 510358 643424 510392 643446
rect 510358 643378 510392 643386
rect 510358 643352 510392 643378
rect 510816 644296 510850 644322
rect 510816 644288 510850 644296
rect 510816 644228 510850 644250
rect 510816 644216 510850 644228
rect 510816 644160 510850 644178
rect 510816 644144 510850 644160
rect 510816 644092 510850 644106
rect 510816 644072 510850 644092
rect 510816 644024 510850 644034
rect 510816 644000 510850 644024
rect 510816 643956 510850 643962
rect 510816 643928 510850 643956
rect 510816 643888 510850 643890
rect 510816 643856 510850 643888
rect 510816 643786 510850 643818
rect 510816 643784 510850 643786
rect 510816 643718 510850 643746
rect 510816 643712 510850 643718
rect 510816 643650 510850 643674
rect 510816 643640 510850 643650
rect 510816 643582 510850 643602
rect 510816 643568 510850 643582
rect 510816 643514 510850 643530
rect 510816 643496 510850 643514
rect 510816 643446 510850 643458
rect 510816 643424 510850 643446
rect 510816 643378 510850 643386
rect 510816 643352 510850 643378
rect 511274 644296 511308 644322
rect 511274 644288 511308 644296
rect 511274 644228 511308 644250
rect 511274 644216 511308 644228
rect 511274 644160 511308 644178
rect 511274 644144 511308 644160
rect 511274 644092 511308 644106
rect 511274 644072 511308 644092
rect 511274 644024 511308 644034
rect 511274 644000 511308 644024
rect 511274 643956 511308 643962
rect 511274 643928 511308 643956
rect 511274 643888 511308 643890
rect 511274 643856 511308 643888
rect 511274 643786 511308 643818
rect 511274 643784 511308 643786
rect 511274 643718 511308 643746
rect 511274 643712 511308 643718
rect 511274 643650 511308 643674
rect 511274 643640 511308 643650
rect 511274 643582 511308 643602
rect 511274 643568 511308 643582
rect 511274 643514 511308 643530
rect 511274 643496 511308 643514
rect 511274 643446 511308 643458
rect 511274 643424 511308 643446
rect 511274 643378 511308 643386
rect 511274 643352 511308 643378
rect 511732 644296 511766 644322
rect 511732 644288 511766 644296
rect 511732 644228 511766 644250
rect 511732 644216 511766 644228
rect 511732 644160 511766 644178
rect 511732 644144 511766 644160
rect 511732 644092 511766 644106
rect 511732 644072 511766 644092
rect 511732 644024 511766 644034
rect 511732 644000 511766 644024
rect 511732 643956 511766 643962
rect 511732 643928 511766 643956
rect 511732 643888 511766 643890
rect 511732 643856 511766 643888
rect 511732 643786 511766 643818
rect 511732 643784 511766 643786
rect 511732 643718 511766 643746
rect 511732 643712 511766 643718
rect 511732 643650 511766 643674
rect 511732 643640 511766 643650
rect 511732 643582 511766 643602
rect 511732 643568 511766 643582
rect 511732 643514 511766 643530
rect 511732 643496 511766 643514
rect 511732 643446 511766 643458
rect 511732 643424 511766 643446
rect 511732 643378 511766 643386
rect 511732 643352 511766 643378
rect 512190 644296 512224 644322
rect 512190 644288 512224 644296
rect 512190 644228 512224 644250
rect 512190 644216 512224 644228
rect 512190 644160 512224 644178
rect 512190 644144 512224 644160
rect 512190 644092 512224 644106
rect 512190 644072 512224 644092
rect 512190 644024 512224 644034
rect 512190 644000 512224 644024
rect 512190 643956 512224 643962
rect 512190 643928 512224 643956
rect 512190 643888 512224 643890
rect 512190 643856 512224 643888
rect 512190 643786 512224 643818
rect 512190 643784 512224 643786
rect 512190 643718 512224 643746
rect 512190 643712 512224 643718
rect 512190 643650 512224 643674
rect 512190 643640 512224 643650
rect 512190 643582 512224 643602
rect 512190 643568 512224 643582
rect 512190 643514 512224 643530
rect 512190 643496 512224 643514
rect 512190 643446 512224 643458
rect 512190 643424 512224 643446
rect 512190 643378 512224 643386
rect 512190 643352 512224 643378
rect 512648 644296 512682 644322
rect 512648 644288 512682 644296
rect 512648 644228 512682 644250
rect 512648 644216 512682 644228
rect 512648 644160 512682 644178
rect 512648 644144 512682 644160
rect 512648 644092 512682 644106
rect 512648 644072 512682 644092
rect 512648 644024 512682 644034
rect 512648 644000 512682 644024
rect 512648 643956 512682 643962
rect 512648 643928 512682 643956
rect 512648 643888 512682 643890
rect 512648 643856 512682 643888
rect 512648 643786 512682 643818
rect 512648 643784 512682 643786
rect 512648 643718 512682 643746
rect 512648 643712 512682 643718
rect 512648 643650 512682 643674
rect 512648 643640 512682 643650
rect 512648 643582 512682 643602
rect 512648 643568 512682 643582
rect 512648 643514 512682 643530
rect 512648 643496 512682 643514
rect 512648 643446 512682 643458
rect 512648 643424 512682 643446
rect 512648 643378 512682 643386
rect 512648 643352 512682 643378
rect 513106 644296 513140 644322
rect 513106 644288 513140 644296
rect 513106 644228 513140 644250
rect 513106 644216 513140 644228
rect 513106 644160 513140 644178
rect 513106 644144 513140 644160
rect 513106 644092 513140 644106
rect 513106 644072 513140 644092
rect 513106 644024 513140 644034
rect 513106 644000 513140 644024
rect 513106 643956 513140 643962
rect 513106 643928 513140 643956
rect 513106 643888 513140 643890
rect 513106 643856 513140 643888
rect 513106 643786 513140 643818
rect 513106 643784 513140 643786
rect 513106 643718 513140 643746
rect 513106 643712 513140 643718
rect 513106 643650 513140 643674
rect 513106 643640 513140 643650
rect 513106 643582 513140 643602
rect 513106 643568 513140 643582
rect 513106 643514 513140 643530
rect 513106 643496 513140 643514
rect 513106 643446 513140 643458
rect 513106 643424 513140 643446
rect 513106 643378 513140 643386
rect 513106 643352 513140 643378
rect 513564 644296 513598 644322
rect 513564 644288 513598 644296
rect 513564 644228 513598 644250
rect 513564 644216 513598 644228
rect 513564 644160 513598 644178
rect 513564 644144 513598 644160
rect 513564 644092 513598 644106
rect 513564 644072 513598 644092
rect 513564 644024 513598 644034
rect 513564 644000 513598 644024
rect 513564 643956 513598 643962
rect 513564 643928 513598 643956
rect 513564 643888 513598 643890
rect 513564 643856 513598 643888
rect 513564 643786 513598 643818
rect 513564 643784 513598 643786
rect 513564 643718 513598 643746
rect 513564 643712 513598 643718
rect 513564 643650 513598 643674
rect 513564 643640 513598 643650
rect 513564 643582 513598 643602
rect 513564 643568 513598 643582
rect 513564 643514 513598 643530
rect 513564 643496 513598 643514
rect 513564 643446 513598 643458
rect 513564 643424 513598 643446
rect 513564 643378 513598 643386
rect 513564 643352 513598 643378
rect 514022 644296 514056 644322
rect 514022 644288 514056 644296
rect 514022 644228 514056 644250
rect 514022 644216 514056 644228
rect 514022 644160 514056 644178
rect 514022 644144 514056 644160
rect 514022 644092 514056 644106
rect 514022 644072 514056 644092
rect 514022 644024 514056 644034
rect 514022 644000 514056 644024
rect 514022 643956 514056 643962
rect 514022 643928 514056 643956
rect 514022 643888 514056 643890
rect 514022 643856 514056 643888
rect 514022 643786 514056 643818
rect 514022 643784 514056 643786
rect 514022 643718 514056 643746
rect 514022 643712 514056 643718
rect 514022 643650 514056 643674
rect 514022 643640 514056 643650
rect 514022 643582 514056 643602
rect 514022 643568 514056 643582
rect 514022 643514 514056 643530
rect 514022 643496 514056 643514
rect 514022 643446 514056 643458
rect 514022 643424 514056 643446
rect 514022 643378 514056 643386
rect 514022 643352 514056 643378
rect 514480 644296 514514 644322
rect 514480 644288 514514 644296
rect 514480 644228 514514 644250
rect 514480 644216 514514 644228
rect 514480 644160 514514 644178
rect 514480 644144 514514 644160
rect 514480 644092 514514 644106
rect 514480 644072 514514 644092
rect 514480 644024 514514 644034
rect 514480 644000 514514 644024
rect 514480 643956 514514 643962
rect 514480 643928 514514 643956
rect 514480 643888 514514 643890
rect 514480 643856 514514 643888
rect 514480 643786 514514 643818
rect 514480 643784 514514 643786
rect 514480 643718 514514 643746
rect 514480 643712 514514 643718
rect 514480 643650 514514 643674
rect 514480 643640 514514 643650
rect 514480 643582 514514 643602
rect 514480 643568 514514 643582
rect 514480 643514 514514 643530
rect 514480 643496 514514 643514
rect 514480 643446 514514 643458
rect 514480 643424 514514 643446
rect 514480 643378 514514 643386
rect 514480 643352 514514 643378
rect 514938 644296 514972 644322
rect 514938 644288 514972 644296
rect 514938 644228 514972 644250
rect 514938 644216 514972 644228
rect 514938 644160 514972 644178
rect 514938 644144 514972 644160
rect 514938 644092 514972 644106
rect 514938 644072 514972 644092
rect 514938 644024 514972 644034
rect 514938 644000 514972 644024
rect 514938 643956 514972 643962
rect 514938 643928 514972 643956
rect 514938 643888 514972 643890
rect 514938 643856 514972 643888
rect 514938 643786 514972 643818
rect 514938 643784 514972 643786
rect 514938 643718 514972 643746
rect 514938 643712 514972 643718
rect 514938 643650 514972 643674
rect 514938 643640 514972 643650
rect 514938 643582 514972 643602
rect 514938 643568 514972 643582
rect 514938 643514 514972 643530
rect 514938 643496 514972 643514
rect 514938 643446 514972 643458
rect 514938 643424 514972 643446
rect 514938 643378 514972 643386
rect 514938 643352 514972 643378
rect 515396 644296 515430 644322
rect 515396 644288 515430 644296
rect 515396 644228 515430 644250
rect 515396 644216 515430 644228
rect 515396 644160 515430 644178
rect 515396 644144 515430 644160
rect 515396 644092 515430 644106
rect 515396 644072 515430 644092
rect 515396 644024 515430 644034
rect 515396 644000 515430 644024
rect 515396 643956 515430 643962
rect 515396 643928 515430 643956
rect 515396 643888 515430 643890
rect 515396 643856 515430 643888
rect 515396 643786 515430 643818
rect 515396 643784 515430 643786
rect 515396 643718 515430 643746
rect 515396 643712 515430 643718
rect 515396 643650 515430 643674
rect 515396 643640 515430 643650
rect 515396 643582 515430 643602
rect 515396 643568 515430 643582
rect 515396 643514 515430 643530
rect 515396 643496 515430 643514
rect 515396 643446 515430 643458
rect 515396 643424 515430 643446
rect 515396 643378 515430 643386
rect 515396 643352 515430 643378
rect 508153 643256 508161 643290
rect 508161 643256 508187 643290
rect 508225 643256 508229 643290
rect 508229 643256 508259 643290
rect 508297 643256 508331 643290
rect 508369 643256 508399 643290
rect 508399 643256 508403 643290
rect 508441 643256 508467 643290
rect 508467 643256 508475 643290
rect 508611 643256 508619 643290
rect 508619 643256 508645 643290
rect 508683 643256 508687 643290
rect 508687 643256 508717 643290
rect 508755 643256 508789 643290
rect 508827 643256 508857 643290
rect 508857 643256 508861 643290
rect 508899 643256 508925 643290
rect 508925 643256 508933 643290
rect 509069 643256 509077 643290
rect 509077 643256 509103 643290
rect 509141 643256 509145 643290
rect 509145 643256 509175 643290
rect 509213 643256 509247 643290
rect 509285 643256 509315 643290
rect 509315 643256 509319 643290
rect 509357 643256 509383 643290
rect 509383 643256 509391 643290
rect 509527 643256 509535 643290
rect 509535 643256 509561 643290
rect 509599 643256 509603 643290
rect 509603 643256 509633 643290
rect 509671 643256 509705 643290
rect 509743 643256 509773 643290
rect 509773 643256 509777 643290
rect 509815 643256 509841 643290
rect 509841 643256 509849 643290
rect 509985 643256 509993 643290
rect 509993 643256 510019 643290
rect 510057 643256 510061 643290
rect 510061 643256 510091 643290
rect 510129 643256 510163 643290
rect 510201 643256 510231 643290
rect 510231 643256 510235 643290
rect 510273 643256 510299 643290
rect 510299 643256 510307 643290
rect 510443 643256 510451 643290
rect 510451 643256 510477 643290
rect 510515 643256 510519 643290
rect 510519 643256 510549 643290
rect 510587 643256 510621 643290
rect 510659 643256 510689 643290
rect 510689 643256 510693 643290
rect 510731 643256 510757 643290
rect 510757 643256 510765 643290
rect 510901 643256 510909 643290
rect 510909 643256 510935 643290
rect 510973 643256 510977 643290
rect 510977 643256 511007 643290
rect 511045 643256 511079 643290
rect 511117 643256 511147 643290
rect 511147 643256 511151 643290
rect 511189 643256 511215 643290
rect 511215 643256 511223 643290
rect 511359 643256 511367 643290
rect 511367 643256 511393 643290
rect 511431 643256 511435 643290
rect 511435 643256 511465 643290
rect 511503 643256 511537 643290
rect 511575 643256 511605 643290
rect 511605 643256 511609 643290
rect 511647 643256 511673 643290
rect 511673 643256 511681 643290
rect 511817 643256 511825 643290
rect 511825 643256 511851 643290
rect 511889 643256 511893 643290
rect 511893 643256 511923 643290
rect 511961 643256 511995 643290
rect 512033 643256 512063 643290
rect 512063 643256 512067 643290
rect 512105 643256 512131 643290
rect 512131 643256 512139 643290
rect 512275 643256 512283 643290
rect 512283 643256 512309 643290
rect 512347 643256 512351 643290
rect 512351 643256 512381 643290
rect 512419 643256 512453 643290
rect 512491 643256 512521 643290
rect 512521 643256 512525 643290
rect 512563 643256 512589 643290
rect 512589 643256 512597 643290
rect 512733 643256 512741 643290
rect 512741 643256 512767 643290
rect 512805 643256 512809 643290
rect 512809 643256 512839 643290
rect 512877 643256 512911 643290
rect 512949 643256 512979 643290
rect 512979 643256 512983 643290
rect 513021 643256 513047 643290
rect 513047 643256 513055 643290
rect 513191 643256 513199 643290
rect 513199 643256 513225 643290
rect 513263 643256 513267 643290
rect 513267 643256 513297 643290
rect 513335 643256 513369 643290
rect 513407 643256 513437 643290
rect 513437 643256 513441 643290
rect 513479 643256 513505 643290
rect 513505 643256 513513 643290
rect 513649 643256 513657 643290
rect 513657 643256 513683 643290
rect 513721 643256 513725 643290
rect 513725 643256 513755 643290
rect 513793 643256 513827 643290
rect 513865 643256 513895 643290
rect 513895 643256 513899 643290
rect 513937 643256 513963 643290
rect 513963 643256 513971 643290
rect 514107 643256 514115 643290
rect 514115 643256 514141 643290
rect 514179 643256 514183 643290
rect 514183 643256 514213 643290
rect 514251 643256 514285 643290
rect 514323 643256 514353 643290
rect 514353 643256 514357 643290
rect 514395 643256 514421 643290
rect 514421 643256 514429 643290
rect 514565 643256 514573 643290
rect 514573 643256 514599 643290
rect 514637 643256 514641 643290
rect 514641 643256 514671 643290
rect 514709 643256 514743 643290
rect 514781 643256 514811 643290
rect 514811 643256 514815 643290
rect 514853 643256 514879 643290
rect 514879 643256 514887 643290
rect 515023 643256 515031 643290
rect 515031 643256 515057 643290
rect 515095 643256 515099 643290
rect 515099 643256 515129 643290
rect 515167 643256 515201 643290
rect 515239 643256 515269 643290
rect 515269 643256 515273 643290
rect 515311 643256 515337 643290
rect 515337 643256 515345 643290
rect 515585 645376 515619 645410
rect 515585 645304 515619 645338
rect 515585 645232 515619 645266
rect 515584 643744 515618 643778
rect 515584 643672 515618 643706
rect 515584 643600 515618 643634
rect 515772 645272 515806 645290
rect 515772 645256 515806 645272
rect 515772 645204 515806 645218
rect 515772 645184 515806 645204
rect 515772 645136 515806 645146
rect 515772 645112 515806 645136
rect 515772 645068 515806 645074
rect 515772 645040 515806 645068
rect 515772 645000 515806 645002
rect 515772 644968 515806 645000
rect 515772 644898 515806 644930
rect 515772 644896 515806 644898
rect 515772 644830 515806 644858
rect 515772 644824 515806 644830
rect 515772 644762 515806 644786
rect 515772 644752 515806 644762
rect 515772 644694 515806 644714
rect 515772 644680 515806 644694
rect 515772 644626 515806 644642
rect 515772 644608 515806 644626
rect 515772 644558 515806 644570
rect 515772 644536 515806 644558
rect 515772 644490 515806 644498
rect 515772 644464 515806 644490
rect 515772 644422 515806 644426
rect 515772 644392 515806 644422
rect 515772 644320 515806 644354
rect 515772 644252 515806 644282
rect 515772 644248 515806 644252
rect 515772 644184 515806 644210
rect 515772 644176 515806 644184
rect 515772 644116 515806 644138
rect 515772 644104 515806 644116
rect 515772 644048 515806 644066
rect 515772 644032 515806 644048
rect 515772 643980 515806 643994
rect 515772 643960 515806 643980
rect 515772 643912 515806 643922
rect 515772 643888 515806 643912
rect 515772 643844 515806 643850
rect 515772 643816 515806 643844
rect 515772 643776 515806 643778
rect 515772 643744 515806 643776
rect 515772 643674 515806 643706
rect 515772 643672 515806 643674
rect 515772 643606 515806 643634
rect 515772 643600 515806 643606
rect 515772 643538 515806 643562
rect 515772 643528 515806 643538
rect 515772 643470 515806 643490
rect 515772 643456 515806 643470
rect 515772 643402 515806 643418
rect 515772 643384 515806 643402
rect 516230 645272 516264 645290
rect 516230 645256 516264 645272
rect 516230 645204 516264 645218
rect 516230 645184 516264 645204
rect 516230 645136 516264 645146
rect 516230 645112 516264 645136
rect 516230 645068 516264 645074
rect 516230 645040 516264 645068
rect 516230 645000 516264 645002
rect 516230 644968 516264 645000
rect 516230 644898 516264 644930
rect 516230 644896 516264 644898
rect 516230 644830 516264 644858
rect 516230 644824 516264 644830
rect 516230 644762 516264 644786
rect 516230 644752 516264 644762
rect 516230 644694 516264 644714
rect 516230 644680 516264 644694
rect 516230 644626 516264 644642
rect 516230 644608 516264 644626
rect 516230 644558 516264 644570
rect 516230 644536 516264 644558
rect 516230 644490 516264 644498
rect 516230 644464 516264 644490
rect 516230 644422 516264 644426
rect 516230 644392 516264 644422
rect 516230 644320 516264 644354
rect 516230 644252 516264 644282
rect 516230 644248 516264 644252
rect 516230 644184 516264 644210
rect 516230 644176 516264 644184
rect 516230 644116 516264 644138
rect 516230 644104 516264 644116
rect 516230 644048 516264 644066
rect 516230 644032 516264 644048
rect 516230 643980 516264 643994
rect 516230 643960 516264 643980
rect 516230 643912 516264 643922
rect 516230 643888 516264 643912
rect 516230 643844 516264 643850
rect 516230 643816 516264 643844
rect 516230 643776 516264 643778
rect 516230 643744 516264 643776
rect 516230 643674 516264 643706
rect 516230 643672 516264 643674
rect 516230 643606 516264 643634
rect 516230 643600 516264 643606
rect 516230 643538 516264 643562
rect 516230 643528 516264 643538
rect 516230 643470 516264 643490
rect 516230 643456 516264 643470
rect 516230 643402 516264 643418
rect 516230 643384 516264 643402
rect 516688 645272 516722 645290
rect 516688 645256 516722 645272
rect 516688 645204 516722 645218
rect 516688 645184 516722 645204
rect 516688 645136 516722 645146
rect 516688 645112 516722 645136
rect 516688 645068 516722 645074
rect 516688 645040 516722 645068
rect 516688 645000 516722 645002
rect 516688 644968 516722 645000
rect 516688 644898 516722 644930
rect 516688 644896 516722 644898
rect 516688 644830 516722 644858
rect 516688 644824 516722 644830
rect 516688 644762 516722 644786
rect 516688 644752 516722 644762
rect 516688 644694 516722 644714
rect 516688 644680 516722 644694
rect 516688 644626 516722 644642
rect 516688 644608 516722 644626
rect 516688 644558 516722 644570
rect 516688 644536 516722 644558
rect 516688 644490 516722 644498
rect 516688 644464 516722 644490
rect 516688 644422 516722 644426
rect 516688 644392 516722 644422
rect 516688 644320 516722 644354
rect 516688 644252 516722 644282
rect 516688 644248 516722 644252
rect 516688 644184 516722 644210
rect 516688 644176 516722 644184
rect 516688 644116 516722 644138
rect 516688 644104 516722 644116
rect 516688 644048 516722 644066
rect 516688 644032 516722 644048
rect 516688 643980 516722 643994
rect 516688 643960 516722 643980
rect 516688 643912 516722 643922
rect 516688 643888 516722 643912
rect 516688 643844 516722 643850
rect 516688 643816 516722 643844
rect 516688 643776 516722 643778
rect 516688 643744 516722 643776
rect 516688 643674 516722 643706
rect 516688 643672 516722 643674
rect 516688 643606 516722 643634
rect 516688 643600 516722 643606
rect 516688 643538 516722 643562
rect 516688 643528 516722 643538
rect 516688 643470 516722 643490
rect 516688 643456 516722 643470
rect 516688 643402 516722 643418
rect 516688 643384 516722 643402
rect 515857 643256 515865 643290
rect 515865 643256 515891 643290
rect 515929 643256 515933 643290
rect 515933 643256 515963 643290
rect 516001 643256 516035 643290
rect 516073 643256 516103 643290
rect 516103 643256 516107 643290
rect 516145 643256 516171 643290
rect 516171 643256 516179 643290
rect 516315 643256 516323 643290
rect 516323 643256 516349 643290
rect 516387 643256 516391 643290
rect 516391 643256 516421 643290
rect 516459 643256 516493 643290
rect 516531 643256 516561 643290
rect 516561 643256 516565 643290
rect 516603 643256 516629 643290
rect 516629 643256 516637 643290
rect 516880 645376 516914 645410
rect 516880 645304 516914 645338
rect 516880 645232 516914 645266
rect 507880 642108 507914 642142
rect 507880 642036 507914 642070
rect 507880 641964 507914 641998
rect 507879 640468 507913 640502
rect 507879 640396 507913 640430
rect 507879 640324 507913 640358
rect 508153 642443 508161 642477
rect 508161 642443 508187 642477
rect 508225 642443 508229 642477
rect 508229 642443 508259 642477
rect 508297 642443 508331 642477
rect 508369 642443 508399 642477
rect 508399 642443 508403 642477
rect 508441 642443 508467 642477
rect 508467 642443 508475 642477
rect 508611 642443 508619 642477
rect 508619 642443 508645 642477
rect 508683 642443 508687 642477
rect 508687 642443 508717 642477
rect 508755 642443 508789 642477
rect 508827 642443 508857 642477
rect 508857 642443 508861 642477
rect 508899 642443 508925 642477
rect 508925 642443 508933 642477
rect 509069 642443 509077 642477
rect 509077 642443 509103 642477
rect 509141 642443 509145 642477
rect 509145 642443 509175 642477
rect 509213 642443 509247 642477
rect 509285 642443 509315 642477
rect 509315 642443 509319 642477
rect 509357 642443 509383 642477
rect 509383 642443 509391 642477
rect 509527 642443 509535 642477
rect 509535 642443 509561 642477
rect 509599 642443 509603 642477
rect 509603 642443 509633 642477
rect 509671 642443 509705 642477
rect 509743 642443 509773 642477
rect 509773 642443 509777 642477
rect 509815 642443 509841 642477
rect 509841 642443 509849 642477
rect 509985 642443 509993 642477
rect 509993 642443 510019 642477
rect 510057 642443 510061 642477
rect 510061 642443 510091 642477
rect 510129 642443 510163 642477
rect 510201 642443 510231 642477
rect 510231 642443 510235 642477
rect 510273 642443 510299 642477
rect 510299 642443 510307 642477
rect 510443 642443 510451 642477
rect 510451 642443 510477 642477
rect 510515 642443 510519 642477
rect 510519 642443 510549 642477
rect 510587 642443 510621 642477
rect 510659 642443 510689 642477
rect 510689 642443 510693 642477
rect 510731 642443 510757 642477
rect 510757 642443 510765 642477
rect 510901 642443 510909 642477
rect 510909 642443 510935 642477
rect 510973 642443 510977 642477
rect 510977 642443 511007 642477
rect 511045 642443 511079 642477
rect 511117 642443 511147 642477
rect 511147 642443 511151 642477
rect 511189 642443 511215 642477
rect 511215 642443 511223 642477
rect 511359 642443 511367 642477
rect 511367 642443 511393 642477
rect 511431 642443 511435 642477
rect 511435 642443 511465 642477
rect 511503 642443 511537 642477
rect 511575 642443 511605 642477
rect 511605 642443 511609 642477
rect 511647 642443 511673 642477
rect 511673 642443 511681 642477
rect 511817 642443 511825 642477
rect 511825 642443 511851 642477
rect 511889 642443 511893 642477
rect 511893 642443 511923 642477
rect 511961 642443 511995 642477
rect 512033 642443 512063 642477
rect 512063 642443 512067 642477
rect 512105 642443 512131 642477
rect 512131 642443 512139 642477
rect 512275 642443 512283 642477
rect 512283 642443 512309 642477
rect 512347 642443 512351 642477
rect 512351 642443 512381 642477
rect 512419 642443 512453 642477
rect 512491 642443 512521 642477
rect 512521 642443 512525 642477
rect 512563 642443 512589 642477
rect 512589 642443 512597 642477
rect 512733 642443 512741 642477
rect 512741 642443 512767 642477
rect 512805 642443 512809 642477
rect 512809 642443 512839 642477
rect 512877 642443 512911 642477
rect 512949 642443 512979 642477
rect 512979 642443 512983 642477
rect 513021 642443 513047 642477
rect 513047 642443 513055 642477
rect 513191 642443 513199 642477
rect 513199 642443 513225 642477
rect 513263 642443 513267 642477
rect 513267 642443 513297 642477
rect 513335 642443 513369 642477
rect 513407 642443 513437 642477
rect 513437 642443 513441 642477
rect 513479 642443 513505 642477
rect 513505 642443 513513 642477
rect 513649 642443 513657 642477
rect 513657 642443 513683 642477
rect 513721 642443 513725 642477
rect 513725 642443 513755 642477
rect 513793 642443 513827 642477
rect 513865 642443 513895 642477
rect 513895 642443 513899 642477
rect 513937 642443 513963 642477
rect 513963 642443 513971 642477
rect 514107 642443 514115 642477
rect 514115 642443 514141 642477
rect 514179 642443 514183 642477
rect 514183 642443 514213 642477
rect 514251 642443 514285 642477
rect 514323 642443 514353 642477
rect 514353 642443 514357 642477
rect 514395 642443 514421 642477
rect 514421 642443 514429 642477
rect 514565 642443 514573 642477
rect 514573 642443 514599 642477
rect 514637 642443 514641 642477
rect 514641 642443 514671 642477
rect 514709 642443 514743 642477
rect 514781 642443 514811 642477
rect 514811 642443 514815 642477
rect 514853 642443 514879 642477
rect 514879 642443 514887 642477
rect 515023 642443 515031 642477
rect 515031 642443 515057 642477
rect 515095 642443 515099 642477
rect 515099 642443 515129 642477
rect 515167 642443 515201 642477
rect 515239 642443 515269 642477
rect 515269 642443 515273 642477
rect 515311 642443 515337 642477
rect 515337 642443 515345 642477
rect 508068 642364 508102 642390
rect 508068 642356 508102 642364
rect 508068 642296 508102 642318
rect 508068 642284 508102 642296
rect 508068 642228 508102 642246
rect 508068 642212 508102 642228
rect 508068 642160 508102 642174
rect 508068 642140 508102 642160
rect 508068 642092 508102 642102
rect 508068 642068 508102 642092
rect 508068 642024 508102 642030
rect 508068 641996 508102 642024
rect 508068 641956 508102 641958
rect 508068 641924 508102 641956
rect 508068 641854 508102 641886
rect 508068 641852 508102 641854
rect 508068 641786 508102 641814
rect 508068 641780 508102 641786
rect 508068 641718 508102 641742
rect 508068 641708 508102 641718
rect 508068 641650 508102 641670
rect 508068 641636 508102 641650
rect 508068 641582 508102 641598
rect 508068 641564 508102 641582
rect 508068 641514 508102 641526
rect 508068 641492 508102 641514
rect 508068 641446 508102 641454
rect 508068 641420 508102 641446
rect 508526 642364 508560 642390
rect 508526 642356 508560 642364
rect 508526 642296 508560 642318
rect 508526 642284 508560 642296
rect 508526 642228 508560 642246
rect 508526 642212 508560 642228
rect 508526 642160 508560 642174
rect 508526 642140 508560 642160
rect 508526 642092 508560 642102
rect 508526 642068 508560 642092
rect 508526 642024 508560 642030
rect 508526 641996 508560 642024
rect 508526 641956 508560 641958
rect 508526 641924 508560 641956
rect 508526 641854 508560 641886
rect 508526 641852 508560 641854
rect 508526 641786 508560 641814
rect 508526 641780 508560 641786
rect 508526 641718 508560 641742
rect 508526 641708 508560 641718
rect 508526 641650 508560 641670
rect 508526 641636 508560 641650
rect 508526 641582 508560 641598
rect 508526 641564 508560 641582
rect 508526 641514 508560 641526
rect 508526 641492 508560 641514
rect 508526 641446 508560 641454
rect 508526 641420 508560 641446
rect 508984 642364 509018 642390
rect 508984 642356 509018 642364
rect 508984 642296 509018 642318
rect 508984 642284 509018 642296
rect 508984 642228 509018 642246
rect 508984 642212 509018 642228
rect 508984 642160 509018 642174
rect 508984 642140 509018 642160
rect 508984 642092 509018 642102
rect 508984 642068 509018 642092
rect 508984 642024 509018 642030
rect 508984 641996 509018 642024
rect 508984 641956 509018 641958
rect 508984 641924 509018 641956
rect 508984 641854 509018 641886
rect 508984 641852 509018 641854
rect 508984 641786 509018 641814
rect 508984 641780 509018 641786
rect 508984 641718 509018 641742
rect 508984 641708 509018 641718
rect 508984 641650 509018 641670
rect 508984 641636 509018 641650
rect 508984 641582 509018 641598
rect 508984 641564 509018 641582
rect 508984 641514 509018 641526
rect 508984 641492 509018 641514
rect 508984 641446 509018 641454
rect 508984 641420 509018 641446
rect 509442 642364 509476 642390
rect 509442 642356 509476 642364
rect 509442 642296 509476 642318
rect 509442 642284 509476 642296
rect 509442 642228 509476 642246
rect 509442 642212 509476 642228
rect 509442 642160 509476 642174
rect 509442 642140 509476 642160
rect 509442 642092 509476 642102
rect 509442 642068 509476 642092
rect 509442 642024 509476 642030
rect 509442 641996 509476 642024
rect 509442 641956 509476 641958
rect 509442 641924 509476 641956
rect 509442 641854 509476 641886
rect 509442 641852 509476 641854
rect 509442 641786 509476 641814
rect 509442 641780 509476 641786
rect 509442 641718 509476 641742
rect 509442 641708 509476 641718
rect 509442 641650 509476 641670
rect 509442 641636 509476 641650
rect 509442 641582 509476 641598
rect 509442 641564 509476 641582
rect 509442 641514 509476 641526
rect 509442 641492 509476 641514
rect 509442 641446 509476 641454
rect 509442 641420 509476 641446
rect 509900 642364 509934 642390
rect 509900 642356 509934 642364
rect 509900 642296 509934 642318
rect 509900 642284 509934 642296
rect 509900 642228 509934 642246
rect 509900 642212 509934 642228
rect 509900 642160 509934 642174
rect 509900 642140 509934 642160
rect 509900 642092 509934 642102
rect 509900 642068 509934 642092
rect 509900 642024 509934 642030
rect 509900 641996 509934 642024
rect 509900 641956 509934 641958
rect 509900 641924 509934 641956
rect 509900 641854 509934 641886
rect 509900 641852 509934 641854
rect 509900 641786 509934 641814
rect 509900 641780 509934 641786
rect 509900 641718 509934 641742
rect 509900 641708 509934 641718
rect 509900 641650 509934 641670
rect 509900 641636 509934 641650
rect 509900 641582 509934 641598
rect 509900 641564 509934 641582
rect 509900 641514 509934 641526
rect 509900 641492 509934 641514
rect 509900 641446 509934 641454
rect 509900 641420 509934 641446
rect 510358 642364 510392 642390
rect 510358 642356 510392 642364
rect 510358 642296 510392 642318
rect 510358 642284 510392 642296
rect 510358 642228 510392 642246
rect 510358 642212 510392 642228
rect 510358 642160 510392 642174
rect 510358 642140 510392 642160
rect 510358 642092 510392 642102
rect 510358 642068 510392 642092
rect 510358 642024 510392 642030
rect 510358 641996 510392 642024
rect 510358 641956 510392 641958
rect 510358 641924 510392 641956
rect 510358 641854 510392 641886
rect 510358 641852 510392 641854
rect 510358 641786 510392 641814
rect 510358 641780 510392 641786
rect 510358 641718 510392 641742
rect 510358 641708 510392 641718
rect 510358 641650 510392 641670
rect 510358 641636 510392 641650
rect 510358 641582 510392 641598
rect 510358 641564 510392 641582
rect 510358 641514 510392 641526
rect 510358 641492 510392 641514
rect 510358 641446 510392 641454
rect 510358 641420 510392 641446
rect 510816 642364 510850 642390
rect 510816 642356 510850 642364
rect 510816 642296 510850 642318
rect 510816 642284 510850 642296
rect 510816 642228 510850 642246
rect 510816 642212 510850 642228
rect 510816 642160 510850 642174
rect 510816 642140 510850 642160
rect 510816 642092 510850 642102
rect 510816 642068 510850 642092
rect 510816 642024 510850 642030
rect 510816 641996 510850 642024
rect 510816 641956 510850 641958
rect 510816 641924 510850 641956
rect 510816 641854 510850 641886
rect 510816 641852 510850 641854
rect 510816 641786 510850 641814
rect 510816 641780 510850 641786
rect 510816 641718 510850 641742
rect 510816 641708 510850 641718
rect 510816 641650 510850 641670
rect 510816 641636 510850 641650
rect 510816 641582 510850 641598
rect 510816 641564 510850 641582
rect 510816 641514 510850 641526
rect 510816 641492 510850 641514
rect 510816 641446 510850 641454
rect 510816 641420 510850 641446
rect 511274 642364 511308 642390
rect 511274 642356 511308 642364
rect 511274 642296 511308 642318
rect 511274 642284 511308 642296
rect 511274 642228 511308 642246
rect 511274 642212 511308 642228
rect 511274 642160 511308 642174
rect 511274 642140 511308 642160
rect 511274 642092 511308 642102
rect 511274 642068 511308 642092
rect 511274 642024 511308 642030
rect 511274 641996 511308 642024
rect 511274 641956 511308 641958
rect 511274 641924 511308 641956
rect 511274 641854 511308 641886
rect 511274 641852 511308 641854
rect 511274 641786 511308 641814
rect 511274 641780 511308 641786
rect 511274 641718 511308 641742
rect 511274 641708 511308 641718
rect 511274 641650 511308 641670
rect 511274 641636 511308 641650
rect 511274 641582 511308 641598
rect 511274 641564 511308 641582
rect 511274 641514 511308 641526
rect 511274 641492 511308 641514
rect 511274 641446 511308 641454
rect 511274 641420 511308 641446
rect 511732 642364 511766 642390
rect 511732 642356 511766 642364
rect 511732 642296 511766 642318
rect 511732 642284 511766 642296
rect 511732 642228 511766 642246
rect 511732 642212 511766 642228
rect 511732 642160 511766 642174
rect 511732 642140 511766 642160
rect 511732 642092 511766 642102
rect 511732 642068 511766 642092
rect 511732 642024 511766 642030
rect 511732 641996 511766 642024
rect 511732 641956 511766 641958
rect 511732 641924 511766 641956
rect 511732 641854 511766 641886
rect 511732 641852 511766 641854
rect 511732 641786 511766 641814
rect 511732 641780 511766 641786
rect 511732 641718 511766 641742
rect 511732 641708 511766 641718
rect 511732 641650 511766 641670
rect 511732 641636 511766 641650
rect 511732 641582 511766 641598
rect 511732 641564 511766 641582
rect 511732 641514 511766 641526
rect 511732 641492 511766 641514
rect 511732 641446 511766 641454
rect 511732 641420 511766 641446
rect 512190 642364 512224 642390
rect 512190 642356 512224 642364
rect 512190 642296 512224 642318
rect 512190 642284 512224 642296
rect 512190 642228 512224 642246
rect 512190 642212 512224 642228
rect 512190 642160 512224 642174
rect 512190 642140 512224 642160
rect 512190 642092 512224 642102
rect 512190 642068 512224 642092
rect 512190 642024 512224 642030
rect 512190 641996 512224 642024
rect 512190 641956 512224 641958
rect 512190 641924 512224 641956
rect 512190 641854 512224 641886
rect 512190 641852 512224 641854
rect 512190 641786 512224 641814
rect 512190 641780 512224 641786
rect 512190 641718 512224 641742
rect 512190 641708 512224 641718
rect 512190 641650 512224 641670
rect 512190 641636 512224 641650
rect 512190 641582 512224 641598
rect 512190 641564 512224 641582
rect 512190 641514 512224 641526
rect 512190 641492 512224 641514
rect 512190 641446 512224 641454
rect 512190 641420 512224 641446
rect 512648 642364 512682 642390
rect 512648 642356 512682 642364
rect 512648 642296 512682 642318
rect 512648 642284 512682 642296
rect 512648 642228 512682 642246
rect 512648 642212 512682 642228
rect 512648 642160 512682 642174
rect 512648 642140 512682 642160
rect 512648 642092 512682 642102
rect 512648 642068 512682 642092
rect 512648 642024 512682 642030
rect 512648 641996 512682 642024
rect 512648 641956 512682 641958
rect 512648 641924 512682 641956
rect 512648 641854 512682 641886
rect 512648 641852 512682 641854
rect 512648 641786 512682 641814
rect 512648 641780 512682 641786
rect 512648 641718 512682 641742
rect 512648 641708 512682 641718
rect 512648 641650 512682 641670
rect 512648 641636 512682 641650
rect 512648 641582 512682 641598
rect 512648 641564 512682 641582
rect 512648 641514 512682 641526
rect 512648 641492 512682 641514
rect 512648 641446 512682 641454
rect 512648 641420 512682 641446
rect 513106 642364 513140 642390
rect 513106 642356 513140 642364
rect 513106 642296 513140 642318
rect 513106 642284 513140 642296
rect 513106 642228 513140 642246
rect 513106 642212 513140 642228
rect 513106 642160 513140 642174
rect 513106 642140 513140 642160
rect 513106 642092 513140 642102
rect 513106 642068 513140 642092
rect 513106 642024 513140 642030
rect 513106 641996 513140 642024
rect 513106 641956 513140 641958
rect 513106 641924 513140 641956
rect 513106 641854 513140 641886
rect 513106 641852 513140 641854
rect 513106 641786 513140 641814
rect 513106 641780 513140 641786
rect 513106 641718 513140 641742
rect 513106 641708 513140 641718
rect 513106 641650 513140 641670
rect 513106 641636 513140 641650
rect 513106 641582 513140 641598
rect 513106 641564 513140 641582
rect 513106 641514 513140 641526
rect 513106 641492 513140 641514
rect 513106 641446 513140 641454
rect 513106 641420 513140 641446
rect 513564 642364 513598 642390
rect 513564 642356 513598 642364
rect 513564 642296 513598 642318
rect 513564 642284 513598 642296
rect 513564 642228 513598 642246
rect 513564 642212 513598 642228
rect 513564 642160 513598 642174
rect 513564 642140 513598 642160
rect 513564 642092 513598 642102
rect 513564 642068 513598 642092
rect 513564 642024 513598 642030
rect 513564 641996 513598 642024
rect 513564 641956 513598 641958
rect 513564 641924 513598 641956
rect 513564 641854 513598 641886
rect 513564 641852 513598 641854
rect 513564 641786 513598 641814
rect 513564 641780 513598 641786
rect 513564 641718 513598 641742
rect 513564 641708 513598 641718
rect 513564 641650 513598 641670
rect 513564 641636 513598 641650
rect 513564 641582 513598 641598
rect 513564 641564 513598 641582
rect 513564 641514 513598 641526
rect 513564 641492 513598 641514
rect 513564 641446 513598 641454
rect 513564 641420 513598 641446
rect 514022 642364 514056 642390
rect 514022 642356 514056 642364
rect 514022 642296 514056 642318
rect 514022 642284 514056 642296
rect 514022 642228 514056 642246
rect 514022 642212 514056 642228
rect 514022 642160 514056 642174
rect 514022 642140 514056 642160
rect 514022 642092 514056 642102
rect 514022 642068 514056 642092
rect 514022 642024 514056 642030
rect 514022 641996 514056 642024
rect 514022 641956 514056 641958
rect 514022 641924 514056 641956
rect 514022 641854 514056 641886
rect 514022 641852 514056 641854
rect 514022 641786 514056 641814
rect 514022 641780 514056 641786
rect 514022 641718 514056 641742
rect 514022 641708 514056 641718
rect 514022 641650 514056 641670
rect 514022 641636 514056 641650
rect 514022 641582 514056 641598
rect 514022 641564 514056 641582
rect 514022 641514 514056 641526
rect 514022 641492 514056 641514
rect 514022 641446 514056 641454
rect 514022 641420 514056 641446
rect 514480 642364 514514 642390
rect 514480 642356 514514 642364
rect 514480 642296 514514 642318
rect 514480 642284 514514 642296
rect 514480 642228 514514 642246
rect 514480 642212 514514 642228
rect 514480 642160 514514 642174
rect 514480 642140 514514 642160
rect 514480 642092 514514 642102
rect 514480 642068 514514 642092
rect 514480 642024 514514 642030
rect 514480 641996 514514 642024
rect 514480 641956 514514 641958
rect 514480 641924 514514 641956
rect 514480 641854 514514 641886
rect 514480 641852 514514 641854
rect 514480 641786 514514 641814
rect 514480 641780 514514 641786
rect 514480 641718 514514 641742
rect 514480 641708 514514 641718
rect 514480 641650 514514 641670
rect 514480 641636 514514 641650
rect 514480 641582 514514 641598
rect 514480 641564 514514 641582
rect 514480 641514 514514 641526
rect 514480 641492 514514 641514
rect 514480 641446 514514 641454
rect 514480 641420 514514 641446
rect 514938 642364 514972 642390
rect 514938 642356 514972 642364
rect 514938 642296 514972 642318
rect 514938 642284 514972 642296
rect 514938 642228 514972 642246
rect 514938 642212 514972 642228
rect 514938 642160 514972 642174
rect 514938 642140 514972 642160
rect 514938 642092 514972 642102
rect 514938 642068 514972 642092
rect 514938 642024 514972 642030
rect 514938 641996 514972 642024
rect 514938 641956 514972 641958
rect 514938 641924 514972 641956
rect 514938 641854 514972 641886
rect 514938 641852 514972 641854
rect 514938 641786 514972 641814
rect 514938 641780 514972 641786
rect 514938 641718 514972 641742
rect 514938 641708 514972 641718
rect 514938 641650 514972 641670
rect 514938 641636 514972 641650
rect 514938 641582 514972 641598
rect 514938 641564 514972 641582
rect 514938 641514 514972 641526
rect 514938 641492 514972 641514
rect 514938 641446 514972 641454
rect 514938 641420 514972 641446
rect 515396 642364 515430 642390
rect 515396 642356 515430 642364
rect 515396 642296 515430 642318
rect 515396 642284 515430 642296
rect 515396 642228 515430 642246
rect 515396 642212 515430 642228
rect 515396 642160 515430 642174
rect 515396 642140 515430 642160
rect 515396 642092 515430 642102
rect 515396 642068 515430 642092
rect 515396 642024 515430 642030
rect 515396 641996 515430 642024
rect 515396 641956 515430 641958
rect 515396 641924 515430 641956
rect 515396 641854 515430 641886
rect 515396 641852 515430 641854
rect 515396 641786 515430 641814
rect 515396 641780 515430 641786
rect 515396 641718 515430 641742
rect 515396 641708 515430 641718
rect 515396 641650 515430 641670
rect 515396 641636 515430 641650
rect 515396 641582 515430 641598
rect 515396 641564 515430 641582
rect 515396 641514 515430 641526
rect 515396 641492 515430 641514
rect 515396 641446 515430 641454
rect 515396 641420 515430 641446
rect 508153 641281 508161 641315
rect 508161 641281 508187 641315
rect 508225 641281 508229 641315
rect 508229 641281 508259 641315
rect 508297 641281 508331 641315
rect 508369 641281 508399 641315
rect 508399 641281 508403 641315
rect 508441 641281 508467 641315
rect 508467 641281 508475 641315
rect 508611 641281 508619 641315
rect 508619 641281 508645 641315
rect 508683 641281 508687 641315
rect 508687 641281 508717 641315
rect 508755 641281 508789 641315
rect 508827 641281 508857 641315
rect 508857 641281 508861 641315
rect 508899 641281 508925 641315
rect 508925 641281 508933 641315
rect 509069 641281 509077 641315
rect 509077 641281 509103 641315
rect 509141 641281 509145 641315
rect 509145 641281 509175 641315
rect 509213 641281 509247 641315
rect 509285 641281 509315 641315
rect 509315 641281 509319 641315
rect 509357 641281 509383 641315
rect 509383 641281 509391 641315
rect 509527 641281 509535 641315
rect 509535 641281 509561 641315
rect 509599 641281 509603 641315
rect 509603 641281 509633 641315
rect 509671 641281 509705 641315
rect 509743 641281 509773 641315
rect 509773 641281 509777 641315
rect 509815 641281 509841 641315
rect 509841 641281 509849 641315
rect 509985 641281 509993 641315
rect 509993 641281 510019 641315
rect 510057 641281 510061 641315
rect 510061 641281 510091 641315
rect 510129 641281 510163 641315
rect 510201 641281 510231 641315
rect 510231 641281 510235 641315
rect 510273 641281 510299 641315
rect 510299 641281 510307 641315
rect 510443 641281 510451 641315
rect 510451 641281 510477 641315
rect 510515 641281 510519 641315
rect 510519 641281 510549 641315
rect 510587 641281 510621 641315
rect 510659 641281 510689 641315
rect 510689 641281 510693 641315
rect 510731 641281 510757 641315
rect 510757 641281 510765 641315
rect 510901 641281 510909 641315
rect 510909 641281 510935 641315
rect 510973 641281 510977 641315
rect 510977 641281 511007 641315
rect 511045 641281 511079 641315
rect 511117 641281 511147 641315
rect 511147 641281 511151 641315
rect 511189 641281 511215 641315
rect 511215 641281 511223 641315
rect 511359 641281 511367 641315
rect 511367 641281 511393 641315
rect 511431 641281 511435 641315
rect 511435 641281 511465 641315
rect 511503 641281 511537 641315
rect 511575 641281 511605 641315
rect 511605 641281 511609 641315
rect 511647 641281 511673 641315
rect 511673 641281 511681 641315
rect 511817 641281 511825 641315
rect 511825 641281 511851 641315
rect 511889 641281 511893 641315
rect 511893 641281 511923 641315
rect 511961 641281 511995 641315
rect 512033 641281 512063 641315
rect 512063 641281 512067 641315
rect 512105 641281 512131 641315
rect 512131 641281 512139 641315
rect 512275 641281 512283 641315
rect 512283 641281 512309 641315
rect 512347 641281 512351 641315
rect 512351 641281 512381 641315
rect 512419 641281 512453 641315
rect 512491 641281 512521 641315
rect 512521 641281 512525 641315
rect 512563 641281 512589 641315
rect 512589 641281 512597 641315
rect 512733 641281 512741 641315
rect 512741 641281 512767 641315
rect 512805 641281 512809 641315
rect 512809 641281 512839 641315
rect 512877 641281 512911 641315
rect 512949 641281 512979 641315
rect 512979 641281 512983 641315
rect 513021 641281 513047 641315
rect 513047 641281 513055 641315
rect 513191 641281 513199 641315
rect 513199 641281 513225 641315
rect 513263 641281 513267 641315
rect 513267 641281 513297 641315
rect 513335 641281 513369 641315
rect 513407 641281 513437 641315
rect 513437 641281 513441 641315
rect 513479 641281 513505 641315
rect 513505 641281 513513 641315
rect 513649 641281 513657 641315
rect 513657 641281 513683 641315
rect 513721 641281 513725 641315
rect 513725 641281 513755 641315
rect 513793 641281 513827 641315
rect 513865 641281 513895 641315
rect 513895 641281 513899 641315
rect 513937 641281 513963 641315
rect 513963 641281 513971 641315
rect 514107 641281 514115 641315
rect 514115 641281 514141 641315
rect 514179 641281 514183 641315
rect 514183 641281 514213 641315
rect 514251 641281 514285 641315
rect 514323 641281 514353 641315
rect 514353 641281 514357 641315
rect 514395 641281 514421 641315
rect 514421 641281 514429 641315
rect 514565 641281 514573 641315
rect 514573 641281 514599 641315
rect 514637 641281 514641 641315
rect 514641 641281 514671 641315
rect 514709 641281 514743 641315
rect 514781 641281 514811 641315
rect 514811 641281 514815 641315
rect 514853 641281 514879 641315
rect 514879 641281 514887 641315
rect 515023 641281 515031 641315
rect 515031 641281 515057 641315
rect 515095 641281 515099 641315
rect 515099 641281 515129 641315
rect 515167 641281 515201 641315
rect 515239 641281 515269 641315
rect 515269 641281 515273 641315
rect 515311 641281 515337 641315
rect 515337 641281 515345 641315
rect 508068 641202 508102 641228
rect 508068 641194 508102 641202
rect 508068 641134 508102 641156
rect 508068 641122 508102 641134
rect 508068 641066 508102 641084
rect 508068 641050 508102 641066
rect 508068 640998 508102 641012
rect 508068 640978 508102 640998
rect 508068 640930 508102 640940
rect 508068 640906 508102 640930
rect 508068 640862 508102 640868
rect 508068 640834 508102 640862
rect 508068 640794 508102 640796
rect 508068 640762 508102 640794
rect 508068 640692 508102 640724
rect 508068 640690 508102 640692
rect 508068 640624 508102 640652
rect 508068 640618 508102 640624
rect 508068 640556 508102 640580
rect 508068 640546 508102 640556
rect 508068 640488 508102 640508
rect 508068 640474 508102 640488
rect 508068 640420 508102 640436
rect 508068 640402 508102 640420
rect 508068 640352 508102 640364
rect 508068 640330 508102 640352
rect 508068 640284 508102 640292
rect 508068 640258 508102 640284
rect 508526 641202 508560 641228
rect 508526 641194 508560 641202
rect 508526 641134 508560 641156
rect 508526 641122 508560 641134
rect 508526 641066 508560 641084
rect 508526 641050 508560 641066
rect 508526 640998 508560 641012
rect 508526 640978 508560 640998
rect 508526 640930 508560 640940
rect 508526 640906 508560 640930
rect 508526 640862 508560 640868
rect 508526 640834 508560 640862
rect 508526 640794 508560 640796
rect 508526 640762 508560 640794
rect 508526 640692 508560 640724
rect 508526 640690 508560 640692
rect 508526 640624 508560 640652
rect 508526 640618 508560 640624
rect 508526 640556 508560 640580
rect 508526 640546 508560 640556
rect 508526 640488 508560 640508
rect 508526 640474 508560 640488
rect 508526 640420 508560 640436
rect 508526 640402 508560 640420
rect 508526 640352 508560 640364
rect 508526 640330 508560 640352
rect 508526 640284 508560 640292
rect 508526 640258 508560 640284
rect 508984 641202 509018 641228
rect 508984 641194 509018 641202
rect 508984 641134 509018 641156
rect 508984 641122 509018 641134
rect 508984 641066 509018 641084
rect 508984 641050 509018 641066
rect 508984 640998 509018 641012
rect 508984 640978 509018 640998
rect 508984 640930 509018 640940
rect 508984 640906 509018 640930
rect 508984 640862 509018 640868
rect 508984 640834 509018 640862
rect 508984 640794 509018 640796
rect 508984 640762 509018 640794
rect 508984 640692 509018 640724
rect 508984 640690 509018 640692
rect 508984 640624 509018 640652
rect 508984 640618 509018 640624
rect 508984 640556 509018 640580
rect 508984 640546 509018 640556
rect 508984 640488 509018 640508
rect 508984 640474 509018 640488
rect 508984 640420 509018 640436
rect 508984 640402 509018 640420
rect 508984 640352 509018 640364
rect 508984 640330 509018 640352
rect 508984 640284 509018 640292
rect 508984 640258 509018 640284
rect 509442 641202 509476 641228
rect 509442 641194 509476 641202
rect 509442 641134 509476 641156
rect 509442 641122 509476 641134
rect 509442 641066 509476 641084
rect 509442 641050 509476 641066
rect 509442 640998 509476 641012
rect 509442 640978 509476 640998
rect 509442 640930 509476 640940
rect 509442 640906 509476 640930
rect 509442 640862 509476 640868
rect 509442 640834 509476 640862
rect 509442 640794 509476 640796
rect 509442 640762 509476 640794
rect 509442 640692 509476 640724
rect 509442 640690 509476 640692
rect 509442 640624 509476 640652
rect 509442 640618 509476 640624
rect 509442 640556 509476 640580
rect 509442 640546 509476 640556
rect 509442 640488 509476 640508
rect 509442 640474 509476 640488
rect 509442 640420 509476 640436
rect 509442 640402 509476 640420
rect 509442 640352 509476 640364
rect 509442 640330 509476 640352
rect 509442 640284 509476 640292
rect 509442 640258 509476 640284
rect 509900 641202 509934 641228
rect 509900 641194 509934 641202
rect 509900 641134 509934 641156
rect 509900 641122 509934 641134
rect 509900 641066 509934 641084
rect 509900 641050 509934 641066
rect 509900 640998 509934 641012
rect 509900 640978 509934 640998
rect 509900 640930 509934 640940
rect 509900 640906 509934 640930
rect 509900 640862 509934 640868
rect 509900 640834 509934 640862
rect 509900 640794 509934 640796
rect 509900 640762 509934 640794
rect 509900 640692 509934 640724
rect 509900 640690 509934 640692
rect 509900 640624 509934 640652
rect 509900 640618 509934 640624
rect 509900 640556 509934 640580
rect 509900 640546 509934 640556
rect 509900 640488 509934 640508
rect 509900 640474 509934 640488
rect 509900 640420 509934 640436
rect 509900 640402 509934 640420
rect 509900 640352 509934 640364
rect 509900 640330 509934 640352
rect 509900 640284 509934 640292
rect 509900 640258 509934 640284
rect 510358 641202 510392 641228
rect 510358 641194 510392 641202
rect 510358 641134 510392 641156
rect 510358 641122 510392 641134
rect 510358 641066 510392 641084
rect 510358 641050 510392 641066
rect 510358 640998 510392 641012
rect 510358 640978 510392 640998
rect 510358 640930 510392 640940
rect 510358 640906 510392 640930
rect 510358 640862 510392 640868
rect 510358 640834 510392 640862
rect 510358 640794 510392 640796
rect 510358 640762 510392 640794
rect 510358 640692 510392 640724
rect 510358 640690 510392 640692
rect 510358 640624 510392 640652
rect 510358 640618 510392 640624
rect 510358 640556 510392 640580
rect 510358 640546 510392 640556
rect 510358 640488 510392 640508
rect 510358 640474 510392 640488
rect 510358 640420 510392 640436
rect 510358 640402 510392 640420
rect 510358 640352 510392 640364
rect 510358 640330 510392 640352
rect 510358 640284 510392 640292
rect 510358 640258 510392 640284
rect 510816 641202 510850 641228
rect 510816 641194 510850 641202
rect 510816 641134 510850 641156
rect 510816 641122 510850 641134
rect 510816 641066 510850 641084
rect 510816 641050 510850 641066
rect 510816 640998 510850 641012
rect 510816 640978 510850 640998
rect 510816 640930 510850 640940
rect 510816 640906 510850 640930
rect 510816 640862 510850 640868
rect 510816 640834 510850 640862
rect 510816 640794 510850 640796
rect 510816 640762 510850 640794
rect 510816 640692 510850 640724
rect 510816 640690 510850 640692
rect 510816 640624 510850 640652
rect 510816 640618 510850 640624
rect 510816 640556 510850 640580
rect 510816 640546 510850 640556
rect 510816 640488 510850 640508
rect 510816 640474 510850 640488
rect 510816 640420 510850 640436
rect 510816 640402 510850 640420
rect 510816 640352 510850 640364
rect 510816 640330 510850 640352
rect 510816 640284 510850 640292
rect 510816 640258 510850 640284
rect 511274 641202 511308 641228
rect 511274 641194 511308 641202
rect 511274 641134 511308 641156
rect 511274 641122 511308 641134
rect 511274 641066 511308 641084
rect 511274 641050 511308 641066
rect 511274 640998 511308 641012
rect 511274 640978 511308 640998
rect 511274 640930 511308 640940
rect 511274 640906 511308 640930
rect 511274 640862 511308 640868
rect 511274 640834 511308 640862
rect 511274 640794 511308 640796
rect 511274 640762 511308 640794
rect 511274 640692 511308 640724
rect 511274 640690 511308 640692
rect 511274 640624 511308 640652
rect 511274 640618 511308 640624
rect 511274 640556 511308 640580
rect 511274 640546 511308 640556
rect 511274 640488 511308 640508
rect 511274 640474 511308 640488
rect 511274 640420 511308 640436
rect 511274 640402 511308 640420
rect 511274 640352 511308 640364
rect 511274 640330 511308 640352
rect 511274 640284 511308 640292
rect 511274 640258 511308 640284
rect 511732 641202 511766 641228
rect 511732 641194 511766 641202
rect 511732 641134 511766 641156
rect 511732 641122 511766 641134
rect 511732 641066 511766 641084
rect 511732 641050 511766 641066
rect 511732 640998 511766 641012
rect 511732 640978 511766 640998
rect 511732 640930 511766 640940
rect 511732 640906 511766 640930
rect 511732 640862 511766 640868
rect 511732 640834 511766 640862
rect 511732 640794 511766 640796
rect 511732 640762 511766 640794
rect 511732 640692 511766 640724
rect 511732 640690 511766 640692
rect 511732 640624 511766 640652
rect 511732 640618 511766 640624
rect 511732 640556 511766 640580
rect 511732 640546 511766 640556
rect 511732 640488 511766 640508
rect 511732 640474 511766 640488
rect 511732 640420 511766 640436
rect 511732 640402 511766 640420
rect 511732 640352 511766 640364
rect 511732 640330 511766 640352
rect 511732 640284 511766 640292
rect 511732 640258 511766 640284
rect 512190 641202 512224 641228
rect 512190 641194 512224 641202
rect 512190 641134 512224 641156
rect 512190 641122 512224 641134
rect 512190 641066 512224 641084
rect 512190 641050 512224 641066
rect 512190 640998 512224 641012
rect 512190 640978 512224 640998
rect 512190 640930 512224 640940
rect 512190 640906 512224 640930
rect 512190 640862 512224 640868
rect 512190 640834 512224 640862
rect 512190 640794 512224 640796
rect 512190 640762 512224 640794
rect 512190 640692 512224 640724
rect 512190 640690 512224 640692
rect 512190 640624 512224 640652
rect 512190 640618 512224 640624
rect 512190 640556 512224 640580
rect 512190 640546 512224 640556
rect 512190 640488 512224 640508
rect 512190 640474 512224 640488
rect 512190 640420 512224 640436
rect 512190 640402 512224 640420
rect 512190 640352 512224 640364
rect 512190 640330 512224 640352
rect 512190 640284 512224 640292
rect 512190 640258 512224 640284
rect 512648 641202 512682 641228
rect 512648 641194 512682 641202
rect 512648 641134 512682 641156
rect 512648 641122 512682 641134
rect 512648 641066 512682 641084
rect 512648 641050 512682 641066
rect 512648 640998 512682 641012
rect 512648 640978 512682 640998
rect 512648 640930 512682 640940
rect 512648 640906 512682 640930
rect 512648 640862 512682 640868
rect 512648 640834 512682 640862
rect 512648 640794 512682 640796
rect 512648 640762 512682 640794
rect 512648 640692 512682 640724
rect 512648 640690 512682 640692
rect 512648 640624 512682 640652
rect 512648 640618 512682 640624
rect 512648 640556 512682 640580
rect 512648 640546 512682 640556
rect 512648 640488 512682 640508
rect 512648 640474 512682 640488
rect 512648 640420 512682 640436
rect 512648 640402 512682 640420
rect 512648 640352 512682 640364
rect 512648 640330 512682 640352
rect 512648 640284 512682 640292
rect 512648 640258 512682 640284
rect 513106 641202 513140 641228
rect 513106 641194 513140 641202
rect 513106 641134 513140 641156
rect 513106 641122 513140 641134
rect 513106 641066 513140 641084
rect 513106 641050 513140 641066
rect 513106 640998 513140 641012
rect 513106 640978 513140 640998
rect 513106 640930 513140 640940
rect 513106 640906 513140 640930
rect 513106 640862 513140 640868
rect 513106 640834 513140 640862
rect 513106 640794 513140 640796
rect 513106 640762 513140 640794
rect 513106 640692 513140 640724
rect 513106 640690 513140 640692
rect 513106 640624 513140 640652
rect 513106 640618 513140 640624
rect 513106 640556 513140 640580
rect 513106 640546 513140 640556
rect 513106 640488 513140 640508
rect 513106 640474 513140 640488
rect 513106 640420 513140 640436
rect 513106 640402 513140 640420
rect 513106 640352 513140 640364
rect 513106 640330 513140 640352
rect 513106 640284 513140 640292
rect 513106 640258 513140 640284
rect 513564 641202 513598 641228
rect 513564 641194 513598 641202
rect 513564 641134 513598 641156
rect 513564 641122 513598 641134
rect 513564 641066 513598 641084
rect 513564 641050 513598 641066
rect 513564 640998 513598 641012
rect 513564 640978 513598 640998
rect 513564 640930 513598 640940
rect 513564 640906 513598 640930
rect 513564 640862 513598 640868
rect 513564 640834 513598 640862
rect 513564 640794 513598 640796
rect 513564 640762 513598 640794
rect 513564 640692 513598 640724
rect 513564 640690 513598 640692
rect 513564 640624 513598 640652
rect 513564 640618 513598 640624
rect 513564 640556 513598 640580
rect 513564 640546 513598 640556
rect 513564 640488 513598 640508
rect 513564 640474 513598 640488
rect 513564 640420 513598 640436
rect 513564 640402 513598 640420
rect 513564 640352 513598 640364
rect 513564 640330 513598 640352
rect 513564 640284 513598 640292
rect 513564 640258 513598 640284
rect 514022 641202 514056 641228
rect 514022 641194 514056 641202
rect 514022 641134 514056 641156
rect 514022 641122 514056 641134
rect 514022 641066 514056 641084
rect 514022 641050 514056 641066
rect 514022 640998 514056 641012
rect 514022 640978 514056 640998
rect 514022 640930 514056 640940
rect 514022 640906 514056 640930
rect 514022 640862 514056 640868
rect 514022 640834 514056 640862
rect 514022 640794 514056 640796
rect 514022 640762 514056 640794
rect 514022 640692 514056 640724
rect 514022 640690 514056 640692
rect 514022 640624 514056 640652
rect 514022 640618 514056 640624
rect 514022 640556 514056 640580
rect 514022 640546 514056 640556
rect 514022 640488 514056 640508
rect 514022 640474 514056 640488
rect 514022 640420 514056 640436
rect 514022 640402 514056 640420
rect 514022 640352 514056 640364
rect 514022 640330 514056 640352
rect 514022 640284 514056 640292
rect 514022 640258 514056 640284
rect 514480 641202 514514 641228
rect 514480 641194 514514 641202
rect 514480 641134 514514 641156
rect 514480 641122 514514 641134
rect 514480 641066 514514 641084
rect 514480 641050 514514 641066
rect 514480 640998 514514 641012
rect 514480 640978 514514 640998
rect 514480 640930 514514 640940
rect 514480 640906 514514 640930
rect 514480 640862 514514 640868
rect 514480 640834 514514 640862
rect 514480 640794 514514 640796
rect 514480 640762 514514 640794
rect 514480 640692 514514 640724
rect 514480 640690 514514 640692
rect 514480 640624 514514 640652
rect 514480 640618 514514 640624
rect 514480 640556 514514 640580
rect 514480 640546 514514 640556
rect 514480 640488 514514 640508
rect 514480 640474 514514 640488
rect 514480 640420 514514 640436
rect 514480 640402 514514 640420
rect 514480 640352 514514 640364
rect 514480 640330 514514 640352
rect 514480 640284 514514 640292
rect 514480 640258 514514 640284
rect 514938 641202 514972 641228
rect 514938 641194 514972 641202
rect 514938 641134 514972 641156
rect 514938 641122 514972 641134
rect 514938 641066 514972 641084
rect 514938 641050 514972 641066
rect 514938 640998 514972 641012
rect 514938 640978 514972 640998
rect 514938 640930 514972 640940
rect 514938 640906 514972 640930
rect 514938 640862 514972 640868
rect 514938 640834 514972 640862
rect 514938 640794 514972 640796
rect 514938 640762 514972 640794
rect 514938 640692 514972 640724
rect 514938 640690 514972 640692
rect 514938 640624 514972 640652
rect 514938 640618 514972 640624
rect 514938 640556 514972 640580
rect 514938 640546 514972 640556
rect 514938 640488 514972 640508
rect 514938 640474 514972 640488
rect 514938 640420 514972 640436
rect 514938 640402 514972 640420
rect 514938 640352 514972 640364
rect 514938 640330 514972 640352
rect 514938 640284 514972 640292
rect 514938 640258 514972 640284
rect 515396 641202 515430 641228
rect 515396 641194 515430 641202
rect 515396 641134 515430 641156
rect 515396 641122 515430 641134
rect 515396 641066 515430 641084
rect 515396 641050 515430 641066
rect 515396 640998 515430 641012
rect 515396 640978 515430 640998
rect 515396 640930 515430 640940
rect 515396 640906 515430 640930
rect 515396 640862 515430 640868
rect 515396 640834 515430 640862
rect 515396 640794 515430 640796
rect 515396 640762 515430 640794
rect 515396 640692 515430 640724
rect 515396 640690 515430 640692
rect 515396 640624 515430 640652
rect 515396 640618 515430 640624
rect 515396 640556 515430 640580
rect 515396 640546 515430 640556
rect 515396 640488 515430 640508
rect 515396 640474 515430 640488
rect 515396 640420 515430 640436
rect 515396 640402 515430 640420
rect 515396 640352 515430 640364
rect 515396 640330 515430 640352
rect 515396 640284 515430 640292
rect 515396 640258 515430 640284
rect 515584 642108 515618 642142
rect 515584 642036 515618 642070
rect 515584 641964 515618 641998
rect 515857 642443 515865 642477
rect 515865 642443 515891 642477
rect 515929 642443 515933 642477
rect 515933 642443 515963 642477
rect 516001 642443 516035 642477
rect 516073 642443 516103 642477
rect 516103 642443 516107 642477
rect 516145 642443 516171 642477
rect 516171 642443 516179 642477
rect 516315 642443 516323 642477
rect 516323 642443 516349 642477
rect 516387 642443 516391 642477
rect 516391 642443 516421 642477
rect 516459 642443 516493 642477
rect 516531 642443 516561 642477
rect 516561 642443 516565 642477
rect 516603 642443 516629 642477
rect 516629 642443 516637 642477
rect 515772 642364 515806 642390
rect 515772 642356 515806 642364
rect 515772 642296 515806 642318
rect 515772 642284 515806 642296
rect 515772 642228 515806 642246
rect 515772 642212 515806 642228
rect 515772 642160 515806 642174
rect 515772 642140 515806 642160
rect 515772 642092 515806 642102
rect 515772 642068 515806 642092
rect 515772 642024 515806 642030
rect 515772 641996 515806 642024
rect 515772 641956 515806 641958
rect 515772 641924 515806 641956
rect 515772 641854 515806 641886
rect 515772 641852 515806 641854
rect 515772 641786 515806 641814
rect 515772 641780 515806 641786
rect 515772 641718 515806 641742
rect 515772 641708 515806 641718
rect 515772 641650 515806 641670
rect 515772 641636 515806 641650
rect 515772 641582 515806 641598
rect 515772 641564 515806 641582
rect 515772 641514 515806 641526
rect 515772 641492 515806 641514
rect 515772 641446 515806 641454
rect 515772 641420 515806 641446
rect 516230 642364 516264 642390
rect 516230 642356 516264 642364
rect 516230 642296 516264 642318
rect 516230 642284 516264 642296
rect 516230 642228 516264 642246
rect 516230 642212 516264 642228
rect 516230 642160 516264 642174
rect 516230 642140 516264 642160
rect 516230 642092 516264 642102
rect 516230 642068 516264 642092
rect 516230 642024 516264 642030
rect 516230 641996 516264 642024
rect 516230 641956 516264 641958
rect 516230 641924 516264 641956
rect 516230 641854 516264 641886
rect 516230 641852 516264 641854
rect 516230 641786 516264 641814
rect 516230 641780 516264 641786
rect 516230 641718 516264 641742
rect 516230 641708 516264 641718
rect 516230 641650 516264 641670
rect 516230 641636 516264 641650
rect 516230 641582 516264 641598
rect 516230 641564 516264 641582
rect 516230 641514 516264 641526
rect 516230 641492 516264 641514
rect 516230 641446 516264 641454
rect 516230 641420 516264 641446
rect 516688 642364 516722 642390
rect 516688 642356 516722 642364
rect 516688 642296 516722 642318
rect 516688 642284 516722 642296
rect 516688 642228 516722 642246
rect 516688 642212 516722 642228
rect 516688 642160 516722 642174
rect 516688 642140 516722 642160
rect 516688 642092 516722 642102
rect 516688 642068 516722 642092
rect 516688 642024 516722 642030
rect 516688 641996 516722 642024
rect 516688 641956 516722 641958
rect 516688 641924 516722 641956
rect 516688 641854 516722 641886
rect 516688 641852 516722 641854
rect 516688 641786 516722 641814
rect 516688 641780 516722 641786
rect 516688 641718 516722 641742
rect 516688 641708 516722 641718
rect 516688 641650 516722 641670
rect 516688 641636 516722 641650
rect 516688 641582 516722 641598
rect 516688 641564 516722 641582
rect 516688 641514 516722 641526
rect 516688 641492 516722 641514
rect 516688 641446 516722 641454
rect 516688 641420 516722 641446
rect 515650 640324 515652 640502
rect 515652 640324 515722 640502
rect 515722 640324 516044 640502
<< metal1 >>
rect 508062 645488 508108 645503
rect 508062 645454 508068 645488
rect 508102 645454 508108 645488
rect 507867 645417 507925 645422
rect 508062 645417 508108 645454
rect 508520 645488 508566 645503
rect 508520 645454 508526 645488
rect 508560 645454 508566 645488
rect 508520 645417 508566 645454
rect 508978 645488 509024 645503
rect 508978 645454 508984 645488
rect 509018 645454 509024 645488
rect 508978 645417 509024 645454
rect 509436 645488 509482 645503
rect 509436 645454 509442 645488
rect 509476 645454 509482 645488
rect 507864 645411 507928 645417
rect 507864 645359 507870 645411
rect 507922 645359 507928 645411
rect 507864 645347 507928 645359
rect 507864 645295 507870 645347
rect 507922 645295 507928 645347
rect 507864 645283 507928 645295
rect 507864 645231 507870 645283
rect 507922 645231 507928 645283
rect 507864 645225 507928 645231
rect 508053 645416 508117 645417
rect 508053 645411 508068 645416
rect 508102 645411 508117 645416
rect 508053 645359 508059 645411
rect 508111 645359 508117 645411
rect 508053 645347 508117 645359
rect 508053 645295 508059 645347
rect 508111 645295 508117 645347
rect 508053 645283 508117 645295
rect 508053 645231 508059 645283
rect 508111 645231 508117 645283
rect 508053 645225 508117 645231
rect 508511 645416 508575 645417
rect 508511 645411 508526 645416
rect 508560 645411 508575 645416
rect 508511 645359 508517 645411
rect 508569 645359 508575 645411
rect 508511 645347 508575 645359
rect 508511 645295 508517 645347
rect 508569 645295 508575 645347
rect 508511 645283 508575 645295
rect 508511 645231 508517 645283
rect 508569 645231 508575 645283
rect 508511 645225 508575 645231
rect 508969 645416 509033 645417
rect 508969 645411 508984 645416
rect 509018 645411 509033 645416
rect 508969 645359 508975 645411
rect 509027 645359 509033 645411
rect 508969 645347 509033 645359
rect 508969 645295 508975 645347
rect 509027 645295 509033 645347
rect 508969 645283 509033 645295
rect 508969 645231 508975 645283
rect 509027 645231 509033 645283
rect 508969 645225 509033 645231
rect 509436 645416 509482 645454
rect 509894 645488 509940 645503
rect 509894 645454 509900 645488
rect 509934 645454 509940 645488
rect 509894 645417 509940 645454
rect 510352 645488 510398 645503
rect 510352 645454 510358 645488
rect 510392 645454 510398 645488
rect 509436 645382 509442 645416
rect 509476 645382 509482 645416
rect 509436 645344 509482 645382
rect 509436 645310 509442 645344
rect 509476 645310 509482 645344
rect 509436 645272 509482 645310
rect 509436 645238 509442 645272
rect 509476 645238 509482 645272
rect 507867 645220 507925 645225
rect 508062 645200 508108 645225
rect 508062 645166 508068 645200
rect 508102 645166 508108 645200
rect 508062 645128 508108 645166
rect 508062 645094 508068 645128
rect 508102 645094 508108 645128
rect 508062 645056 508108 645094
rect 508062 645022 508068 645056
rect 508102 645022 508108 645056
rect 508062 644984 508108 645022
rect 508062 644950 508068 644984
rect 508102 644950 508108 644984
rect 508062 644912 508108 644950
rect 508062 644878 508068 644912
rect 508102 644878 508108 644912
rect 508062 644840 508108 644878
rect 508062 644806 508068 644840
rect 508102 644806 508108 644840
rect 508062 644768 508108 644806
rect 508062 644734 508068 644768
rect 508102 644734 508108 644768
rect 508062 644696 508108 644734
rect 508062 644662 508068 644696
rect 508102 644662 508108 644696
rect 508062 644624 508108 644662
rect 508062 644590 508068 644624
rect 508102 644590 508108 644624
rect 508062 644552 508108 644590
rect 508062 644518 508068 644552
rect 508102 644518 508108 644552
rect 508062 644503 508108 644518
rect 508520 645200 508566 645225
rect 508520 645166 508526 645200
rect 508560 645166 508566 645200
rect 508520 645128 508566 645166
rect 508520 645094 508526 645128
rect 508560 645094 508566 645128
rect 508520 645056 508566 645094
rect 508520 645022 508526 645056
rect 508560 645022 508566 645056
rect 508520 644984 508566 645022
rect 508520 644950 508526 644984
rect 508560 644950 508566 644984
rect 508520 644912 508566 644950
rect 508520 644878 508526 644912
rect 508560 644878 508566 644912
rect 508520 644840 508566 644878
rect 508520 644806 508526 644840
rect 508560 644806 508566 644840
rect 508520 644768 508566 644806
rect 508520 644734 508526 644768
rect 508560 644734 508566 644768
rect 508520 644696 508566 644734
rect 508520 644662 508526 644696
rect 508560 644662 508566 644696
rect 508520 644624 508566 644662
rect 508520 644590 508526 644624
rect 508560 644590 508566 644624
rect 508520 644552 508566 644590
rect 508520 644518 508526 644552
rect 508560 644518 508566 644552
rect 508520 644462 508566 644518
rect 508978 645200 509024 645225
rect 508978 645166 508984 645200
rect 509018 645166 509024 645200
rect 508978 645128 509024 645166
rect 508978 645094 508984 645128
rect 509018 645094 509024 645128
rect 508978 645056 509024 645094
rect 508978 645022 508984 645056
rect 509018 645022 509024 645056
rect 508978 644984 509024 645022
rect 508978 644950 508984 644984
rect 509018 644950 509024 644984
rect 508978 644912 509024 644950
rect 508978 644878 508984 644912
rect 509018 644878 509024 644912
rect 508978 644840 509024 644878
rect 508978 644806 508984 644840
rect 509018 644806 509024 644840
rect 508978 644768 509024 644806
rect 509436 645200 509482 645238
rect 509885 645416 509949 645417
rect 509885 645411 509900 645416
rect 509934 645411 509949 645416
rect 509885 645359 509891 645411
rect 509943 645359 509949 645411
rect 509885 645347 509949 645359
rect 509885 645295 509891 645347
rect 509943 645295 509949 645347
rect 509885 645283 509949 645295
rect 509885 645231 509891 645283
rect 509943 645231 509949 645283
rect 509885 645225 509949 645231
rect 510352 645416 510398 645454
rect 510810 645488 510856 645503
rect 510810 645454 510816 645488
rect 510850 645454 510856 645488
rect 510810 645417 510856 645454
rect 511268 645488 511314 645503
rect 511268 645454 511274 645488
rect 511308 645454 511314 645488
rect 510352 645382 510358 645416
rect 510392 645382 510398 645416
rect 510352 645344 510398 645382
rect 510352 645310 510358 645344
rect 510392 645310 510398 645344
rect 510352 645272 510398 645310
rect 510352 645238 510358 645272
rect 510392 645238 510398 645272
rect 509436 645166 509442 645200
rect 509476 645166 509482 645200
rect 509436 645128 509482 645166
rect 509436 645094 509442 645128
rect 509476 645094 509482 645128
rect 509436 645056 509482 645094
rect 509436 645022 509442 645056
rect 509476 645022 509482 645056
rect 509436 644984 509482 645022
rect 509436 644950 509442 644984
rect 509476 644950 509482 644984
rect 509436 644912 509482 644950
rect 509436 644878 509442 644912
rect 509476 644878 509482 644912
rect 509436 644840 509482 644878
rect 509436 644806 509442 644840
rect 509476 644806 509482 644840
rect 509436 644782 509482 644806
rect 509894 645200 509940 645225
rect 509894 645166 509900 645200
rect 509934 645166 509940 645200
rect 509894 645128 509940 645166
rect 509894 645094 509900 645128
rect 509934 645094 509940 645128
rect 509894 645056 509940 645094
rect 509894 645022 509900 645056
rect 509934 645022 509940 645056
rect 509894 644984 509940 645022
rect 509894 644950 509900 644984
rect 509934 644950 509940 644984
rect 509894 644912 509940 644950
rect 509894 644878 509900 644912
rect 509934 644878 509940 644912
rect 509894 644840 509940 644878
rect 509894 644806 509900 644840
rect 509934 644806 509940 644840
rect 508978 644734 508984 644768
rect 509018 644734 509024 644768
rect 508978 644696 509024 644734
rect 508978 644662 508984 644696
rect 509018 644662 509024 644696
rect 508978 644624 509024 644662
rect 508978 644590 508984 644624
rect 509018 644590 509024 644624
rect 509427 644776 509491 644782
rect 509427 644724 509433 644776
rect 509485 644724 509491 644776
rect 509427 644712 509491 644724
rect 509427 644660 509433 644712
rect 509485 644660 509491 644712
rect 509427 644648 509491 644660
rect 509427 644596 509433 644648
rect 509485 644596 509491 644648
rect 509427 644590 509442 644596
rect 509476 644590 509491 644596
rect 509894 644768 509940 644806
rect 510352 645200 510398 645238
rect 510801 645416 510865 645417
rect 510801 645411 510816 645416
rect 510850 645411 510865 645416
rect 510801 645359 510807 645411
rect 510859 645359 510865 645411
rect 510801 645347 510865 645359
rect 510801 645295 510807 645347
rect 510859 645295 510865 645347
rect 510801 645283 510865 645295
rect 510801 645231 510807 645283
rect 510859 645231 510865 645283
rect 510801 645225 510865 645231
rect 511268 645416 511314 645454
rect 511726 645488 511772 645503
rect 511726 645454 511732 645488
rect 511766 645454 511772 645488
rect 511726 645417 511772 645454
rect 512184 645488 512230 645503
rect 512184 645454 512190 645488
rect 512224 645454 512230 645488
rect 511268 645382 511274 645416
rect 511308 645382 511314 645416
rect 511268 645344 511314 645382
rect 511268 645310 511274 645344
rect 511308 645310 511314 645344
rect 511268 645272 511314 645310
rect 511268 645238 511274 645272
rect 511308 645238 511314 645272
rect 510352 645166 510358 645200
rect 510392 645166 510398 645200
rect 510352 645128 510398 645166
rect 510352 645094 510358 645128
rect 510392 645094 510398 645128
rect 510352 645056 510398 645094
rect 510352 645022 510358 645056
rect 510392 645022 510398 645056
rect 510352 644984 510398 645022
rect 510352 644950 510358 644984
rect 510392 644950 510398 644984
rect 510352 644912 510398 644950
rect 510352 644878 510358 644912
rect 510392 644878 510398 644912
rect 510352 644840 510398 644878
rect 510352 644806 510358 644840
rect 510392 644806 510398 644840
rect 510352 644782 510398 644806
rect 510810 645200 510856 645225
rect 510810 645166 510816 645200
rect 510850 645166 510856 645200
rect 510810 645128 510856 645166
rect 510810 645094 510816 645128
rect 510850 645094 510856 645128
rect 511268 645200 511314 645238
rect 511717 645416 511781 645417
rect 511717 645411 511732 645416
rect 511766 645411 511781 645416
rect 511717 645359 511723 645411
rect 511775 645359 511781 645411
rect 511717 645347 511781 645359
rect 511717 645295 511723 645347
rect 511775 645295 511781 645347
rect 511717 645283 511781 645295
rect 511717 645231 511723 645283
rect 511775 645231 511781 645283
rect 511717 645225 511781 645231
rect 512184 645416 512230 645454
rect 512642 645488 512688 645503
rect 512642 645454 512648 645488
rect 512682 645454 512688 645488
rect 512642 645417 512688 645454
rect 513100 645488 513146 645503
rect 513100 645454 513106 645488
rect 513140 645454 513146 645488
rect 512184 645382 512190 645416
rect 512224 645382 512230 645416
rect 512184 645344 512230 645382
rect 512184 645310 512190 645344
rect 512224 645310 512230 645344
rect 512184 645272 512230 645310
rect 512184 645238 512190 645272
rect 512224 645238 512230 645272
rect 511268 645166 511274 645200
rect 511308 645166 511314 645200
rect 511268 645128 511314 645166
rect 511268 645094 511274 645128
rect 511308 645094 511314 645128
rect 511726 645200 511772 645225
rect 511726 645166 511732 645200
rect 511766 645166 511772 645200
rect 511726 645128 511772 645166
rect 511726 645094 511732 645128
rect 511766 645094 511772 645128
rect 512184 645200 512230 645238
rect 512633 645416 512697 645417
rect 512633 645411 512648 645416
rect 512682 645411 512697 645416
rect 512633 645359 512639 645411
rect 512691 645359 512697 645411
rect 512633 645347 512697 645359
rect 512633 645295 512639 645347
rect 512691 645295 512697 645347
rect 512633 645283 512697 645295
rect 512633 645231 512639 645283
rect 512691 645231 512697 645283
rect 512633 645225 512697 645231
rect 513100 645416 513146 645454
rect 513558 645488 513604 645503
rect 513558 645454 513564 645488
rect 513598 645454 513604 645488
rect 513558 645417 513604 645454
rect 514016 645488 514062 645503
rect 514016 645454 514022 645488
rect 514056 645454 514062 645488
rect 513100 645382 513106 645416
rect 513140 645382 513146 645416
rect 513100 645344 513146 645382
rect 513100 645310 513106 645344
rect 513140 645310 513146 645344
rect 513100 645272 513146 645310
rect 513100 645238 513106 645272
rect 513140 645238 513146 645272
rect 512184 645166 512190 645200
rect 512224 645166 512230 645200
rect 512184 645128 512230 645166
rect 512184 645094 512190 645128
rect 512224 645094 512230 645128
rect 512642 645200 512688 645225
rect 512642 645166 512648 645200
rect 512682 645166 512688 645200
rect 512642 645128 512688 645166
rect 512642 645094 512648 645128
rect 512682 645094 512688 645128
rect 510810 645056 510856 645094
rect 510810 645022 510816 645056
rect 510850 645022 510856 645056
rect 510810 644984 510856 645022
rect 510810 644950 510816 644984
rect 510850 644950 510856 644984
rect 510810 644912 510856 644950
rect 510810 644878 510816 644912
rect 510850 644878 510856 644912
rect 511259 645088 511323 645094
rect 511259 645036 511265 645088
rect 511317 645036 511323 645088
rect 511259 645024 511274 645036
rect 511308 645024 511323 645036
rect 511259 644972 511265 645024
rect 511317 644972 511323 645024
rect 511259 644960 511274 644972
rect 511308 644960 511323 644972
rect 511259 644908 511265 644960
rect 511317 644908 511323 644960
rect 511259 644902 511274 644908
rect 510810 644840 510856 644878
rect 510810 644806 510816 644840
rect 510850 644806 510856 644840
rect 509894 644734 509900 644768
rect 509934 644734 509940 644768
rect 509894 644696 509940 644734
rect 509894 644662 509900 644696
rect 509934 644662 509940 644696
rect 509894 644624 509940 644662
rect 509894 644590 509900 644624
rect 509934 644590 509940 644624
rect 510343 644776 510407 644782
rect 510343 644724 510349 644776
rect 510401 644724 510407 644776
rect 510343 644712 510407 644724
rect 510343 644660 510349 644712
rect 510401 644660 510407 644712
rect 510343 644648 510407 644660
rect 510343 644596 510349 644648
rect 510401 644596 510407 644648
rect 510343 644590 510358 644596
rect 510392 644590 510407 644596
rect 510810 644768 510856 644806
rect 510810 644734 510816 644768
rect 510850 644734 510856 644768
rect 510810 644696 510856 644734
rect 510810 644662 510816 644696
rect 510850 644662 510856 644696
rect 510810 644624 510856 644662
rect 510810 644590 510816 644624
rect 510850 644590 510856 644624
rect 508978 644552 509024 644590
rect 508978 644518 508984 644552
rect 509018 644518 509024 644552
rect 508978 644503 509024 644518
rect 509436 644552 509482 644590
rect 509436 644518 509442 644552
rect 509476 644518 509482 644552
rect 509436 644503 509482 644518
rect 509894 644552 509940 644590
rect 509894 644518 509900 644552
rect 509934 644518 509940 644552
rect 509894 644503 509940 644518
rect 510352 644552 510398 644590
rect 510352 644518 510358 644552
rect 510392 644518 510398 644552
rect 510352 644462 510398 644518
rect 510810 644552 510856 644590
rect 510810 644518 510816 644552
rect 510850 644518 510856 644552
rect 510810 644503 510856 644518
rect 511268 644878 511274 644902
rect 511308 644902 511323 644908
rect 511726 645056 511772 645094
rect 511726 645022 511732 645056
rect 511766 645022 511772 645056
rect 511726 644984 511772 645022
rect 511726 644950 511732 644984
rect 511766 644950 511772 644984
rect 511726 644912 511772 644950
rect 511308 644878 511314 644902
rect 511268 644840 511314 644878
rect 511268 644806 511274 644840
rect 511308 644806 511314 644840
rect 511268 644768 511314 644806
rect 511268 644734 511274 644768
rect 511308 644734 511314 644768
rect 511268 644696 511314 644734
rect 511268 644662 511274 644696
rect 511308 644662 511314 644696
rect 511268 644624 511314 644662
rect 511268 644590 511274 644624
rect 511308 644590 511314 644624
rect 511268 644552 511314 644590
rect 511268 644518 511274 644552
rect 511308 644518 511314 644552
rect 511268 644462 511314 644518
rect 511726 644878 511732 644912
rect 511766 644878 511772 644912
rect 512175 645088 512239 645094
rect 512175 645036 512181 645088
rect 512233 645036 512239 645088
rect 512175 645024 512190 645036
rect 512224 645024 512239 645036
rect 512175 644972 512181 645024
rect 512233 644972 512239 645024
rect 512175 644960 512190 644972
rect 512224 644960 512239 644972
rect 512175 644908 512181 644960
rect 512233 644908 512239 644960
rect 512175 644902 512190 644908
rect 511726 644840 511772 644878
rect 511726 644806 511732 644840
rect 511766 644806 511772 644840
rect 511726 644768 511772 644806
rect 511726 644734 511732 644768
rect 511766 644734 511772 644768
rect 511726 644696 511772 644734
rect 511726 644662 511732 644696
rect 511766 644662 511772 644696
rect 511726 644624 511772 644662
rect 511726 644590 511732 644624
rect 511766 644590 511772 644624
rect 511726 644552 511772 644590
rect 511726 644518 511732 644552
rect 511766 644518 511772 644552
rect 511726 644503 511772 644518
rect 512184 644878 512190 644902
rect 512224 644902 512239 644908
rect 512642 645056 512688 645094
rect 512642 645022 512648 645056
rect 512682 645022 512688 645056
rect 512642 644984 512688 645022
rect 512642 644950 512648 644984
rect 512682 644950 512688 644984
rect 512642 644912 512688 644950
rect 512224 644878 512230 644902
rect 512184 644840 512230 644878
rect 512184 644806 512190 644840
rect 512224 644806 512230 644840
rect 512184 644768 512230 644806
rect 512184 644734 512190 644768
rect 512224 644734 512230 644768
rect 512184 644696 512230 644734
rect 512184 644662 512190 644696
rect 512224 644662 512230 644696
rect 512184 644624 512230 644662
rect 512184 644590 512190 644624
rect 512224 644590 512230 644624
rect 512184 644552 512230 644590
rect 512184 644518 512190 644552
rect 512224 644518 512230 644552
rect 512184 644503 512230 644518
rect 512642 644878 512648 644912
rect 512682 644878 512688 644912
rect 512642 644840 512688 644878
rect 512642 644806 512648 644840
rect 512682 644806 512688 644840
rect 512642 644768 512688 644806
rect 513100 645200 513146 645238
rect 513549 645416 513613 645417
rect 513549 645411 513564 645416
rect 513598 645411 513613 645416
rect 513549 645359 513555 645411
rect 513607 645359 513613 645411
rect 513549 645347 513613 645359
rect 513549 645295 513555 645347
rect 513607 645295 513613 645347
rect 513549 645283 513613 645295
rect 513549 645231 513555 645283
rect 513607 645231 513613 645283
rect 513549 645225 513613 645231
rect 514016 645416 514062 645454
rect 514474 645488 514520 645503
rect 514474 645454 514480 645488
rect 514514 645454 514520 645488
rect 514474 645417 514520 645454
rect 514932 645488 514978 645503
rect 514932 645454 514938 645488
rect 514972 645454 514978 645488
rect 514932 645417 514978 645454
rect 515390 645488 515436 645503
rect 515390 645454 515396 645488
rect 515430 645454 515436 645488
rect 515390 645417 515436 645454
rect 515573 645417 515631 645422
rect 516868 645417 516926 645422
rect 514016 645382 514022 645416
rect 514056 645382 514062 645416
rect 514016 645344 514062 645382
rect 514016 645310 514022 645344
rect 514056 645310 514062 645344
rect 514016 645272 514062 645310
rect 514016 645238 514022 645272
rect 514056 645238 514062 645272
rect 513100 645166 513106 645200
rect 513140 645166 513146 645200
rect 513100 645128 513146 645166
rect 513100 645094 513106 645128
rect 513140 645094 513146 645128
rect 513100 645056 513146 645094
rect 513100 645022 513106 645056
rect 513140 645022 513146 645056
rect 513100 644984 513146 645022
rect 513100 644950 513106 644984
rect 513140 644950 513146 644984
rect 513100 644912 513146 644950
rect 513100 644878 513106 644912
rect 513140 644878 513146 644912
rect 513100 644840 513146 644878
rect 513100 644806 513106 644840
rect 513140 644806 513146 644840
rect 513100 644782 513146 644806
rect 513558 645200 513604 645225
rect 513558 645166 513564 645200
rect 513598 645166 513604 645200
rect 513558 645128 513604 645166
rect 513558 645094 513564 645128
rect 513598 645094 513604 645128
rect 513558 645056 513604 645094
rect 513558 645022 513564 645056
rect 513598 645022 513604 645056
rect 513558 644984 513604 645022
rect 513558 644950 513564 644984
rect 513598 644950 513604 644984
rect 513558 644912 513604 644950
rect 513558 644878 513564 644912
rect 513598 644878 513604 644912
rect 513558 644840 513604 644878
rect 513558 644806 513564 644840
rect 513598 644806 513604 644840
rect 512642 644734 512648 644768
rect 512682 644734 512688 644768
rect 512642 644696 512688 644734
rect 512642 644662 512648 644696
rect 512682 644662 512688 644696
rect 512642 644624 512688 644662
rect 512642 644590 512648 644624
rect 512682 644590 512688 644624
rect 513091 644776 513155 644782
rect 513091 644724 513097 644776
rect 513149 644724 513155 644776
rect 513091 644712 513155 644724
rect 513091 644660 513097 644712
rect 513149 644660 513155 644712
rect 513091 644648 513155 644660
rect 513091 644596 513097 644648
rect 513149 644596 513155 644648
rect 513091 644590 513106 644596
rect 513140 644590 513155 644596
rect 513558 644768 513604 644806
rect 514016 645200 514062 645238
rect 514465 645416 514529 645417
rect 514465 645411 514480 645416
rect 514514 645411 514529 645416
rect 514465 645359 514471 645411
rect 514523 645359 514529 645411
rect 514465 645347 514529 645359
rect 514465 645295 514471 645347
rect 514523 645295 514529 645347
rect 514465 645283 514529 645295
rect 514465 645231 514471 645283
rect 514523 645231 514529 645283
rect 514465 645225 514529 645231
rect 514923 645416 514987 645417
rect 514923 645411 514938 645416
rect 514972 645411 514987 645416
rect 514923 645359 514929 645411
rect 514981 645359 514987 645411
rect 514923 645347 514987 645359
rect 514923 645295 514929 645347
rect 514981 645295 514987 645347
rect 514923 645283 514987 645295
rect 514923 645231 514929 645283
rect 514981 645231 514987 645283
rect 514923 645225 514987 645231
rect 515381 645416 515445 645417
rect 515381 645411 515396 645416
rect 515430 645411 515445 645416
rect 515381 645359 515387 645411
rect 515439 645359 515445 645411
rect 515381 645347 515445 645359
rect 515381 645295 515387 645347
rect 515439 645295 515445 645347
rect 515381 645283 515445 645295
rect 515381 645231 515387 645283
rect 515439 645231 515445 645283
rect 515381 645225 515445 645231
rect 515570 645411 515634 645417
rect 515570 645359 515576 645411
rect 515628 645359 515634 645411
rect 515570 645347 515634 645359
rect 515570 645295 515576 645347
rect 515628 645295 515634 645347
rect 516865 645411 516929 645417
rect 516865 645359 516871 645411
rect 516923 645359 516929 645411
rect 516865 645347 516929 645359
rect 515570 645283 515634 645295
rect 515570 645231 515576 645283
rect 515628 645231 515634 645283
rect 515570 645225 515634 645231
rect 515766 645290 515812 645337
rect 515766 645256 515772 645290
rect 515806 645256 515812 645290
rect 514016 645166 514022 645200
rect 514056 645166 514062 645200
rect 514016 645128 514062 645166
rect 514016 645094 514022 645128
rect 514056 645094 514062 645128
rect 514016 645056 514062 645094
rect 514016 645022 514022 645056
rect 514056 645022 514062 645056
rect 514016 644984 514062 645022
rect 514016 644950 514022 644984
rect 514056 644950 514062 644984
rect 514016 644912 514062 644950
rect 514016 644878 514022 644912
rect 514056 644878 514062 644912
rect 514016 644840 514062 644878
rect 514016 644806 514022 644840
rect 514056 644806 514062 644840
rect 514016 644782 514062 644806
rect 514474 645200 514520 645225
rect 514474 645166 514480 645200
rect 514514 645166 514520 645200
rect 514474 645128 514520 645166
rect 514474 645094 514480 645128
rect 514514 645094 514520 645128
rect 514474 645056 514520 645094
rect 514474 645022 514480 645056
rect 514514 645022 514520 645056
rect 514474 644984 514520 645022
rect 514474 644950 514480 644984
rect 514514 644950 514520 644984
rect 514474 644912 514520 644950
rect 514474 644878 514480 644912
rect 514514 644878 514520 644912
rect 514474 644840 514520 644878
rect 514474 644806 514480 644840
rect 514514 644806 514520 644840
rect 513558 644734 513564 644768
rect 513598 644734 513604 644768
rect 513558 644696 513604 644734
rect 513558 644662 513564 644696
rect 513598 644662 513604 644696
rect 513558 644624 513604 644662
rect 513558 644590 513564 644624
rect 513598 644590 513604 644624
rect 514007 644776 514071 644782
rect 514007 644724 514013 644776
rect 514065 644724 514071 644776
rect 514007 644712 514071 644724
rect 514007 644660 514013 644712
rect 514065 644660 514071 644712
rect 514007 644648 514071 644660
rect 514007 644596 514013 644648
rect 514065 644596 514071 644648
rect 514007 644590 514022 644596
rect 514056 644590 514071 644596
rect 514474 644768 514520 644806
rect 514474 644734 514480 644768
rect 514514 644734 514520 644768
rect 514474 644696 514520 644734
rect 514474 644662 514480 644696
rect 514514 644662 514520 644696
rect 514474 644624 514520 644662
rect 514474 644590 514480 644624
rect 514514 644590 514520 644624
rect 512642 644552 512688 644590
rect 512642 644518 512648 644552
rect 512682 644518 512688 644552
rect 512642 644503 512688 644518
rect 513100 644552 513146 644590
rect 513100 644518 513106 644552
rect 513140 644518 513146 644552
rect 513100 644462 513146 644518
rect 513558 644552 513604 644590
rect 513558 644518 513564 644552
rect 513598 644518 513604 644552
rect 513558 644503 513604 644518
rect 514016 644552 514062 644590
rect 514016 644518 514022 644552
rect 514056 644518 514062 644552
rect 514016 644503 514062 644518
rect 514474 644552 514520 644590
rect 514474 644518 514480 644552
rect 514514 644518 514520 644552
rect 514474 644503 514520 644518
rect 514932 645200 514978 645225
rect 514932 645166 514938 645200
rect 514972 645166 514978 645200
rect 514932 645128 514978 645166
rect 514932 645094 514938 645128
rect 514972 645094 514978 645128
rect 514932 645056 514978 645094
rect 514932 645022 514938 645056
rect 514972 645022 514978 645056
rect 514932 644984 514978 645022
rect 514932 644950 514938 644984
rect 514972 644950 514978 644984
rect 514932 644912 514978 644950
rect 514932 644878 514938 644912
rect 514972 644878 514978 644912
rect 514932 644840 514978 644878
rect 514932 644806 514938 644840
rect 514972 644806 514978 644840
rect 514932 644768 514978 644806
rect 514932 644734 514938 644768
rect 514972 644734 514978 644768
rect 514932 644696 514978 644734
rect 514932 644662 514938 644696
rect 514972 644662 514978 644696
rect 514932 644624 514978 644662
rect 514932 644590 514938 644624
rect 514972 644590 514978 644624
rect 514932 644552 514978 644590
rect 514932 644518 514938 644552
rect 514972 644518 514978 644552
rect 514932 644462 514978 644518
rect 515390 645200 515436 645225
rect 515573 645220 515631 645225
rect 515390 645166 515396 645200
rect 515430 645166 515436 645200
rect 515390 645128 515436 645166
rect 515390 645094 515396 645128
rect 515430 645094 515436 645128
rect 515390 645056 515436 645094
rect 515390 645022 515396 645056
rect 515430 645022 515436 645056
rect 515390 644984 515436 645022
rect 515390 644950 515396 644984
rect 515430 644950 515436 644984
rect 515390 644912 515436 644950
rect 515390 644878 515396 644912
rect 515430 644878 515436 644912
rect 515390 644840 515436 644878
rect 515390 644806 515396 644840
rect 515430 644806 515436 644840
rect 515390 644768 515436 644806
rect 515390 644734 515396 644768
rect 515430 644734 515436 644768
rect 515390 644696 515436 644734
rect 515390 644662 515396 644696
rect 515430 644662 515436 644696
rect 515390 644624 515436 644662
rect 515390 644590 515396 644624
rect 515430 644590 515436 644624
rect 515390 644552 515436 644590
rect 515766 645218 515812 645256
rect 516224 645290 516270 645337
rect 516224 645256 516230 645290
rect 516264 645256 516270 645290
rect 516224 645255 516270 645256
rect 516682 645290 516728 645337
rect 516682 645256 516688 645290
rect 516722 645256 516728 645290
rect 515766 645184 515772 645218
rect 515806 645184 515812 645218
rect 515766 645146 515812 645184
rect 515766 645112 515772 645146
rect 515806 645112 515812 645146
rect 515766 645074 515812 645112
rect 515766 645040 515772 645074
rect 515806 645040 515812 645074
rect 515766 645002 515812 645040
rect 515766 644968 515772 645002
rect 515806 644968 515812 645002
rect 515766 644930 515812 644968
rect 515766 644896 515772 644930
rect 515806 644896 515812 644930
rect 515766 644858 515812 644896
rect 516215 645249 516279 645255
rect 516215 645197 516221 645249
rect 516273 645197 516279 645249
rect 516215 645185 516230 645197
rect 516264 645185 516279 645197
rect 516215 645133 516221 645185
rect 516273 645133 516279 645185
rect 516215 645121 516230 645133
rect 516264 645121 516279 645133
rect 516215 645069 516221 645121
rect 516273 645069 516279 645121
rect 516215 645057 516230 645069
rect 516264 645057 516279 645069
rect 516215 645005 516221 645057
rect 516273 645005 516279 645057
rect 516215 645002 516279 645005
rect 516215 644993 516230 645002
rect 516264 644993 516279 645002
rect 516215 644941 516221 644993
rect 516273 644941 516279 644993
rect 516215 644930 516279 644941
rect 516215 644929 516230 644930
rect 516264 644929 516279 644930
rect 516215 644877 516221 644929
rect 516273 644877 516279 644929
rect 516215 644871 516279 644877
rect 516682 645218 516728 645256
rect 516865 645295 516871 645347
rect 516923 645295 516929 645347
rect 516865 645283 516929 645295
rect 516865 645231 516871 645283
rect 516923 645231 516929 645283
rect 516865 645225 516929 645231
rect 516868 645220 516926 645225
rect 516682 645184 516688 645218
rect 516722 645184 516728 645218
rect 516682 645146 516728 645184
rect 516682 645112 516688 645146
rect 516722 645112 516728 645146
rect 516682 645074 516728 645112
rect 516682 645040 516688 645074
rect 516722 645040 516728 645074
rect 516682 645002 516728 645040
rect 516682 644968 516688 645002
rect 516722 644968 516728 645002
rect 516682 644930 516728 644968
rect 516682 644896 516688 644930
rect 516722 644896 516728 644930
rect 515766 644824 515772 644858
rect 515806 644824 515812 644858
rect 515766 644786 515812 644824
rect 515766 644752 515772 644786
rect 515806 644752 515812 644786
rect 515766 644714 515812 644752
rect 515766 644680 515772 644714
rect 515806 644680 515812 644714
rect 515766 644642 515812 644680
rect 515766 644608 515772 644642
rect 515806 644608 515812 644642
rect 515766 644570 515812 644608
rect 515766 644565 515772 644570
rect 515390 644518 515396 644552
rect 515430 644518 515436 644552
rect 515390 644503 515436 644518
rect 515757 644559 515772 644565
rect 515806 644565 515812 644570
rect 516224 644858 516270 644871
rect 516224 644824 516230 644858
rect 516264 644824 516270 644858
rect 516224 644786 516270 644824
rect 516224 644752 516230 644786
rect 516264 644752 516270 644786
rect 516224 644714 516270 644752
rect 516224 644680 516230 644714
rect 516264 644680 516270 644714
rect 516224 644642 516270 644680
rect 516224 644608 516230 644642
rect 516264 644608 516270 644642
rect 516224 644570 516270 644608
rect 515806 644559 515821 644565
rect 515757 644507 515763 644559
rect 515815 644507 515821 644559
rect 515757 644498 515821 644507
rect 515757 644495 515772 644498
rect 515806 644495 515821 644498
rect 508118 644456 508968 644462
rect 508118 644422 508153 644456
rect 508187 644422 508225 644456
rect 508259 644422 508297 644456
rect 508331 644422 508369 644456
rect 508403 644422 508441 644456
rect 508475 644422 508611 644456
rect 508645 644422 508683 644456
rect 508717 644422 508755 644456
rect 508789 644422 508827 644456
rect 508861 644422 508899 644456
rect 508933 644422 508968 644456
rect 508118 644416 508968 644422
rect 509034 644456 510800 644462
rect 509034 644422 509069 644456
rect 509103 644422 509141 644456
rect 509175 644422 509213 644456
rect 509247 644422 509285 644456
rect 509319 644422 509357 644456
rect 509391 644422 509527 644456
rect 509561 644422 509599 644456
rect 509633 644422 509671 644456
rect 509705 644422 509743 644456
rect 509777 644422 509815 644456
rect 509849 644422 509985 644456
rect 510019 644422 510057 644456
rect 510091 644422 510129 644456
rect 510163 644422 510201 644456
rect 510235 644422 510273 644456
rect 510307 644422 510443 644456
rect 510477 644422 510515 644456
rect 510549 644422 510587 644456
rect 510621 644422 510659 644456
rect 510693 644422 510731 644456
rect 510765 644422 510800 644456
rect 509034 644416 510800 644422
rect 510866 644456 512632 644462
rect 510866 644422 510901 644456
rect 510935 644422 510973 644456
rect 511007 644422 511045 644456
rect 511079 644422 511117 644456
rect 511151 644422 511189 644456
rect 511223 644422 511359 644456
rect 511393 644422 511431 644456
rect 511465 644422 511503 644456
rect 511537 644422 511575 644456
rect 511609 644422 511647 644456
rect 511681 644422 511817 644456
rect 511851 644422 511889 644456
rect 511923 644422 511961 644456
rect 511995 644422 512033 644456
rect 512067 644422 512105 644456
rect 512139 644422 512275 644456
rect 512309 644422 512347 644456
rect 512381 644422 512419 644456
rect 512453 644422 512491 644456
rect 512525 644422 512563 644456
rect 512597 644422 512632 644456
rect 510866 644416 512632 644422
rect 512698 644456 514464 644462
rect 512698 644422 512733 644456
rect 512767 644422 512805 644456
rect 512839 644422 512877 644456
rect 512911 644422 512949 644456
rect 512983 644422 513021 644456
rect 513055 644422 513191 644456
rect 513225 644422 513263 644456
rect 513297 644422 513335 644456
rect 513369 644422 513407 644456
rect 513441 644422 513479 644456
rect 513513 644422 513649 644456
rect 513683 644422 513721 644456
rect 513755 644422 513793 644456
rect 513827 644422 513865 644456
rect 513899 644422 513937 644456
rect 513971 644422 514107 644456
rect 514141 644422 514179 644456
rect 514213 644422 514251 644456
rect 514285 644422 514323 644456
rect 514357 644422 514395 644456
rect 514429 644422 514464 644456
rect 512698 644416 514464 644422
rect 514530 644456 515380 644462
rect 514530 644422 514565 644456
rect 514599 644422 514637 644456
rect 514671 644422 514709 644456
rect 514743 644422 514781 644456
rect 514815 644422 514853 644456
rect 514887 644422 515023 644456
rect 515057 644422 515095 644456
rect 515129 644422 515167 644456
rect 515201 644422 515239 644456
rect 515273 644422 515311 644456
rect 515345 644422 515380 644456
rect 514530 644416 515380 644422
rect 515757 644443 515763 644495
rect 515815 644443 515821 644495
rect 515757 644431 515821 644443
rect 515757 644379 515763 644431
rect 515815 644379 515821 644431
rect 515757 644367 515821 644379
rect 508062 644322 508108 644337
rect 508062 644288 508068 644322
rect 508102 644288 508108 644322
rect 508062 644250 508108 644288
rect 508062 644216 508068 644250
rect 508102 644216 508108 644250
rect 508062 644178 508108 644216
rect 508062 644144 508068 644178
rect 508102 644144 508108 644178
rect 508062 644106 508108 644144
rect 508062 644072 508068 644106
rect 508102 644072 508108 644106
rect 508062 644034 508108 644072
rect 508062 644000 508068 644034
rect 508102 644000 508108 644034
rect 508062 643962 508108 644000
rect 508062 643928 508068 643962
rect 508102 643928 508108 643962
rect 508062 643890 508108 643928
rect 508062 643856 508068 643890
rect 508102 643856 508108 643890
rect 508062 643818 508108 643856
rect 507868 643785 507926 643790
rect 508062 643785 508068 643818
rect 507865 643779 507929 643785
rect 507865 643727 507871 643779
rect 507923 643727 507929 643779
rect 507865 643715 507929 643727
rect 507865 643663 507871 643715
rect 507923 643663 507929 643715
rect 507865 643651 507929 643663
rect 507865 643599 507871 643651
rect 507923 643599 507929 643651
rect 507865 643593 507929 643599
rect 508053 643784 508068 643785
rect 508102 643785 508108 643818
rect 508520 644322 508566 644337
rect 508520 644288 508526 644322
rect 508560 644288 508566 644322
rect 508520 644250 508566 644288
rect 508978 644322 509024 644337
rect 508978 644288 508984 644322
rect 509018 644288 509024 644322
rect 508978 644250 509024 644288
rect 509436 644322 509482 644337
rect 509436 644288 509442 644322
rect 509476 644288 509482 644322
rect 509436 644250 509482 644288
rect 509894 644322 509940 644337
rect 509894 644288 509900 644322
rect 509934 644288 509940 644322
rect 509894 644250 509940 644288
rect 510352 644322 510398 644337
rect 510352 644288 510358 644322
rect 510392 644288 510398 644322
rect 510352 644250 510398 644288
rect 510810 644322 510856 644337
rect 510810 644288 510816 644322
rect 510850 644288 510856 644322
rect 510810 644250 510856 644288
rect 511268 644322 511314 644337
rect 511268 644288 511274 644322
rect 511308 644288 511314 644322
rect 511268 644250 511314 644288
rect 511726 644322 511772 644337
rect 511726 644288 511732 644322
rect 511766 644288 511772 644322
rect 511726 644250 511772 644288
rect 512184 644322 512230 644337
rect 512184 644288 512190 644322
rect 512224 644288 512230 644322
rect 512184 644250 512230 644288
rect 512642 644322 512688 644337
rect 512642 644288 512648 644322
rect 512682 644288 512688 644322
rect 512642 644250 512688 644288
rect 513100 644322 513146 644337
rect 513100 644288 513106 644322
rect 513140 644288 513146 644322
rect 513100 644250 513146 644288
rect 513558 644322 513604 644337
rect 513558 644288 513564 644322
rect 513598 644288 513604 644322
rect 513558 644250 513604 644288
rect 514016 644322 514062 644337
rect 514016 644288 514022 644322
rect 514056 644288 514062 644322
rect 514016 644250 514062 644288
rect 508520 644216 508526 644250
rect 508560 644216 508566 644250
rect 508520 644178 508566 644216
rect 508520 644144 508526 644178
rect 508560 644144 508566 644178
rect 508520 644106 508566 644144
rect 508520 644072 508526 644106
rect 508560 644072 508566 644106
rect 508520 644034 508566 644072
rect 508969 644244 508984 644250
rect 509018 644244 509033 644250
rect 508969 644192 508975 644244
rect 509027 644192 509033 644244
rect 508969 644180 509033 644192
rect 508969 644128 508975 644180
rect 509027 644128 509033 644180
rect 508969 644116 509033 644128
rect 508969 644064 508975 644116
rect 509027 644064 509033 644116
rect 508969 644058 509033 644064
rect 509436 644216 509442 644250
rect 509476 644216 509482 644250
rect 509436 644178 509482 644216
rect 509436 644144 509442 644178
rect 509476 644144 509482 644178
rect 509436 644106 509482 644144
rect 509436 644072 509442 644106
rect 509476 644072 509482 644106
rect 508520 644000 508526 644034
rect 508560 644000 508566 644034
rect 508520 643962 508566 644000
rect 508520 643928 508526 643962
rect 508560 643928 508566 643962
rect 508520 643890 508566 643928
rect 508520 643856 508526 643890
rect 508560 643856 508566 643890
rect 508520 643818 508566 643856
rect 508520 643785 508526 643818
rect 508102 643784 508117 643785
rect 508053 643779 508117 643784
rect 508053 643727 508059 643779
rect 508111 643727 508117 643779
rect 508053 643715 508068 643727
rect 508102 643715 508117 643727
rect 508053 643663 508059 643715
rect 508111 643663 508117 643715
rect 508053 643651 508068 643663
rect 508102 643651 508117 643663
rect 508053 643599 508059 643651
rect 508111 643599 508117 643651
rect 508053 643593 508068 643599
rect 507868 643588 507926 643593
rect 508062 643568 508068 643593
rect 508102 643593 508117 643599
rect 508511 643784 508526 643785
rect 508560 643785 508566 643818
rect 508978 644034 509024 644058
rect 508978 644000 508984 644034
rect 509018 644000 509024 644034
rect 508978 643962 509024 644000
rect 508978 643928 508984 643962
rect 509018 643928 509024 643962
rect 508978 643890 509024 643928
rect 508978 643856 508984 643890
rect 509018 643856 509024 643890
rect 508978 643818 509024 643856
rect 508560 643784 508575 643785
rect 508511 643779 508575 643784
rect 508511 643727 508517 643779
rect 508569 643727 508575 643779
rect 508511 643715 508526 643727
rect 508560 643715 508575 643727
rect 508511 643663 508517 643715
rect 508569 643663 508575 643715
rect 508511 643651 508526 643663
rect 508560 643651 508575 643663
rect 508511 643599 508517 643651
rect 508569 643599 508575 643651
rect 508511 643593 508526 643599
rect 508102 643568 508108 643593
rect 508062 643530 508108 643568
rect 508062 643496 508068 643530
rect 508102 643496 508108 643530
rect 508062 643458 508108 643496
rect 508062 643424 508068 643458
rect 508102 643424 508108 643458
rect 508062 643386 508108 643424
rect 508062 643352 508068 643386
rect 508102 643352 508108 643386
rect 508062 643296 508108 643352
rect 508520 643568 508526 643593
rect 508560 643593 508575 643599
rect 508978 643784 508984 643818
rect 509018 643784 509024 643818
rect 509436 644034 509482 644072
rect 509885 644244 509900 644250
rect 509934 644244 509949 644250
rect 509885 644192 509891 644244
rect 509943 644192 509949 644244
rect 509885 644180 509949 644192
rect 509885 644128 509891 644180
rect 509943 644128 509949 644180
rect 509885 644116 509949 644128
rect 509885 644064 509891 644116
rect 509943 644064 509949 644116
rect 509885 644058 509949 644064
rect 510352 644216 510358 644250
rect 510392 644216 510398 644250
rect 510352 644178 510398 644216
rect 510352 644144 510358 644178
rect 510392 644144 510398 644178
rect 510352 644106 510398 644144
rect 510352 644072 510358 644106
rect 510392 644072 510398 644106
rect 509436 644000 509442 644034
rect 509476 644000 509482 644034
rect 509436 643962 509482 644000
rect 509436 643928 509442 643962
rect 509476 643928 509482 643962
rect 509436 643890 509482 643928
rect 509436 643856 509442 643890
rect 509476 643856 509482 643890
rect 509436 643818 509482 643856
rect 509436 643785 509442 643818
rect 508978 643746 509024 643784
rect 508978 643712 508984 643746
rect 509018 643712 509024 643746
rect 508978 643674 509024 643712
rect 508978 643640 508984 643674
rect 509018 643640 509024 643674
rect 508978 643602 509024 643640
rect 508560 643568 508566 643593
rect 508520 643530 508566 643568
rect 508520 643496 508526 643530
rect 508560 643496 508566 643530
rect 508520 643458 508566 643496
rect 508520 643424 508526 643458
rect 508560 643424 508566 643458
rect 508520 643386 508566 643424
rect 508520 643352 508526 643386
rect 508560 643352 508566 643386
rect 508520 643337 508566 643352
rect 508978 643568 508984 643602
rect 509018 643568 509024 643602
rect 509427 643784 509442 643785
rect 509476 643785 509482 643818
rect 509894 644034 509940 644058
rect 509894 644000 509900 644034
rect 509934 644000 509940 644034
rect 509894 643962 509940 644000
rect 509894 643928 509900 643962
rect 509934 643928 509940 643962
rect 509894 643890 509940 643928
rect 509894 643856 509900 643890
rect 509934 643856 509940 643890
rect 509894 643818 509940 643856
rect 509476 643784 509491 643785
rect 509427 643779 509491 643784
rect 509427 643727 509433 643779
rect 509485 643727 509491 643779
rect 509427 643715 509442 643727
rect 509476 643715 509491 643727
rect 509427 643663 509433 643715
rect 509485 643663 509491 643715
rect 509427 643651 509442 643663
rect 509476 643651 509491 643663
rect 509427 643599 509433 643651
rect 509485 643599 509491 643651
rect 509427 643593 509442 643599
rect 508978 643530 509024 643568
rect 508978 643496 508984 643530
rect 509018 643496 509024 643530
rect 508978 643458 509024 643496
rect 508978 643424 508984 643458
rect 509018 643424 509024 643458
rect 508978 643386 509024 643424
rect 508978 643352 508984 643386
rect 509018 643352 509024 643386
rect 508978 643337 509024 643352
rect 509436 643568 509442 643593
rect 509476 643593 509491 643599
rect 509894 643784 509900 643818
rect 509934 643784 509940 643818
rect 510352 644034 510398 644072
rect 510801 644244 510816 644250
rect 510850 644244 510865 644250
rect 510801 644192 510807 644244
rect 510859 644192 510865 644244
rect 510801 644180 510865 644192
rect 510801 644128 510807 644180
rect 510859 644128 510865 644180
rect 510801 644116 510865 644128
rect 510801 644064 510807 644116
rect 510859 644064 510865 644116
rect 510801 644058 510865 644064
rect 511268 644216 511274 644250
rect 511308 644216 511314 644250
rect 511268 644178 511314 644216
rect 511268 644144 511274 644178
rect 511308 644144 511314 644178
rect 511268 644106 511314 644144
rect 511268 644072 511274 644106
rect 511308 644072 511314 644106
rect 510352 644000 510358 644034
rect 510392 644000 510398 644034
rect 510352 643962 510398 644000
rect 510352 643928 510358 643962
rect 510392 643928 510398 643962
rect 510352 643890 510398 643928
rect 510352 643856 510358 643890
rect 510392 643856 510398 643890
rect 510352 643818 510398 643856
rect 510352 643785 510358 643818
rect 509894 643746 509940 643784
rect 509894 643712 509900 643746
rect 509934 643712 509940 643746
rect 509894 643674 509940 643712
rect 509894 643640 509900 643674
rect 509934 643640 509940 643674
rect 509894 643602 509940 643640
rect 509476 643568 509482 643593
rect 509436 643530 509482 643568
rect 509436 643496 509442 643530
rect 509476 643496 509482 643530
rect 509436 643458 509482 643496
rect 509436 643424 509442 643458
rect 509476 643424 509482 643458
rect 509436 643386 509482 643424
rect 509436 643352 509442 643386
rect 509476 643383 509482 643386
rect 509894 643568 509900 643602
rect 509934 643568 509940 643602
rect 510343 643784 510358 643785
rect 510392 643785 510398 643818
rect 510810 644034 510856 644058
rect 510810 644000 510816 644034
rect 510850 644000 510856 644034
rect 510810 643962 510856 644000
rect 510810 643928 510816 643962
rect 510850 643928 510856 643962
rect 510810 643890 510856 643928
rect 510810 643856 510816 643890
rect 510850 643856 510856 643890
rect 510810 643818 510856 643856
rect 510392 643784 510407 643785
rect 510343 643779 510407 643784
rect 510343 643727 510349 643779
rect 510401 643727 510407 643779
rect 510343 643715 510358 643727
rect 510392 643715 510407 643727
rect 510343 643663 510349 643715
rect 510401 643663 510407 643715
rect 510343 643651 510358 643663
rect 510392 643651 510407 643663
rect 510343 643599 510349 643651
rect 510401 643599 510407 643651
rect 510343 643593 510358 643599
rect 509894 643530 509940 643568
rect 509894 643496 509900 643530
rect 509934 643496 509940 643530
rect 509894 643458 509940 643496
rect 509894 643424 509900 643458
rect 509934 643424 509940 643458
rect 509894 643386 509940 643424
rect 509476 643352 509538 643383
rect 509436 643337 509538 643352
rect 509894 643352 509900 643386
rect 509934 643352 509940 643386
rect 509894 643337 509940 643352
rect 510352 643568 510358 643593
rect 510392 643593 510407 643599
rect 510810 643784 510816 643818
rect 510850 643784 510856 643818
rect 511268 644034 511314 644072
rect 511717 644244 511732 644250
rect 511766 644244 511781 644250
rect 511717 644192 511723 644244
rect 511775 644192 511781 644244
rect 511717 644180 511781 644192
rect 511717 644128 511723 644180
rect 511775 644128 511781 644180
rect 511717 644116 511781 644128
rect 511717 644064 511723 644116
rect 511775 644064 511781 644116
rect 511717 644058 511781 644064
rect 512184 644216 512190 644250
rect 512224 644216 512230 644250
rect 512184 644178 512230 644216
rect 512184 644144 512190 644178
rect 512224 644144 512230 644178
rect 512184 644106 512230 644144
rect 512184 644072 512190 644106
rect 512224 644072 512230 644106
rect 511268 644000 511274 644034
rect 511308 644000 511314 644034
rect 511268 643962 511314 644000
rect 511268 643928 511274 643962
rect 511308 643928 511314 643962
rect 511268 643890 511314 643928
rect 511268 643856 511274 643890
rect 511308 643856 511314 643890
rect 511268 643818 511314 643856
rect 511268 643785 511274 643818
rect 510810 643746 510856 643784
rect 510810 643712 510816 643746
rect 510850 643712 510856 643746
rect 510810 643674 510856 643712
rect 510810 643640 510816 643674
rect 510850 643640 510856 643674
rect 510810 643602 510856 643640
rect 510392 643568 510398 643593
rect 510352 643530 510398 643568
rect 510352 643496 510358 643530
rect 510392 643496 510398 643530
rect 510352 643458 510398 643496
rect 510352 643424 510358 643458
rect 510392 643424 510398 643458
rect 510352 643386 510398 643424
rect 510352 643352 510358 643386
rect 510392 643352 510398 643386
rect 510352 643337 510398 643352
rect 510810 643568 510816 643602
rect 510850 643568 510856 643602
rect 511259 643784 511274 643785
rect 511308 643785 511314 643818
rect 511726 644034 511772 644058
rect 511726 644000 511732 644034
rect 511766 644000 511772 644034
rect 511726 643962 511772 644000
rect 511726 643928 511732 643962
rect 511766 643928 511772 643962
rect 511726 643890 511772 643928
rect 511726 643856 511732 643890
rect 511766 643856 511772 643890
rect 511726 643818 511772 643856
rect 511308 643784 511323 643785
rect 511259 643779 511323 643784
rect 511259 643727 511265 643779
rect 511317 643727 511323 643779
rect 511259 643715 511274 643727
rect 511308 643715 511323 643727
rect 511259 643663 511265 643715
rect 511317 643663 511323 643715
rect 511259 643651 511274 643663
rect 511308 643651 511323 643663
rect 511259 643599 511265 643651
rect 511317 643599 511323 643651
rect 511259 643593 511274 643599
rect 510810 643530 510856 643568
rect 510810 643496 510816 643530
rect 510850 643496 510856 643530
rect 510810 643458 510856 643496
rect 510810 643424 510816 643458
rect 510850 643424 510856 643458
rect 510810 643386 510856 643424
rect 510810 643352 510816 643386
rect 510850 643352 510856 643386
rect 510810 643337 510856 643352
rect 511268 643568 511274 643593
rect 511308 643593 511323 643599
rect 511726 643784 511732 643818
rect 511766 643784 511772 643818
rect 512184 644034 512230 644072
rect 512633 644244 512648 644250
rect 512682 644244 512697 644250
rect 512633 644192 512639 644244
rect 512691 644192 512697 644244
rect 512633 644180 512697 644192
rect 512633 644128 512639 644180
rect 512691 644128 512697 644180
rect 512633 644116 512697 644128
rect 512633 644064 512639 644116
rect 512691 644064 512697 644116
rect 512633 644058 512697 644064
rect 513100 644216 513106 644250
rect 513140 644216 513146 644250
rect 513100 644178 513146 644216
rect 513100 644144 513106 644178
rect 513140 644144 513146 644178
rect 513100 644106 513146 644144
rect 513100 644072 513106 644106
rect 513140 644072 513146 644106
rect 512184 644000 512190 644034
rect 512224 644000 512230 644034
rect 512184 643962 512230 644000
rect 512184 643928 512190 643962
rect 512224 643928 512230 643962
rect 512184 643890 512230 643928
rect 512184 643856 512190 643890
rect 512224 643856 512230 643890
rect 512184 643818 512230 643856
rect 512184 643785 512190 643818
rect 511726 643746 511772 643784
rect 511726 643712 511732 643746
rect 511766 643712 511772 643746
rect 511726 643674 511772 643712
rect 511726 643640 511732 643674
rect 511766 643640 511772 643674
rect 511726 643602 511772 643640
rect 511308 643568 511314 643593
rect 511268 643530 511314 643568
rect 511268 643496 511274 643530
rect 511308 643496 511314 643530
rect 511268 643458 511314 643496
rect 511268 643424 511274 643458
rect 511308 643424 511314 643458
rect 511268 643386 511314 643424
rect 511268 643352 511274 643386
rect 511308 643352 511314 643386
rect 511268 643337 511314 643352
rect 511726 643568 511732 643602
rect 511766 643568 511772 643602
rect 512175 643784 512190 643785
rect 512224 643785 512230 643818
rect 512642 644034 512688 644058
rect 512642 644000 512648 644034
rect 512682 644000 512688 644034
rect 512642 643962 512688 644000
rect 512642 643928 512648 643962
rect 512682 643928 512688 643962
rect 512642 643890 512688 643928
rect 512642 643856 512648 643890
rect 512682 643856 512688 643890
rect 512642 643818 512688 643856
rect 512224 643784 512239 643785
rect 512175 643779 512239 643784
rect 512175 643727 512181 643779
rect 512233 643727 512239 643779
rect 512175 643715 512190 643727
rect 512224 643715 512239 643727
rect 512175 643663 512181 643715
rect 512233 643663 512239 643715
rect 512175 643651 512190 643663
rect 512224 643651 512239 643663
rect 512175 643599 512181 643651
rect 512233 643599 512239 643651
rect 512175 643593 512190 643599
rect 511726 643530 511772 643568
rect 511726 643496 511732 643530
rect 511766 643496 511772 643530
rect 511726 643458 511772 643496
rect 511726 643424 511732 643458
rect 511766 643424 511772 643458
rect 511726 643386 511772 643424
rect 511726 643352 511732 643386
rect 511766 643352 511772 643386
rect 511726 643337 511772 643352
rect 512184 643568 512190 643593
rect 512224 643593 512239 643599
rect 512642 643784 512648 643818
rect 512682 643784 512688 643818
rect 513100 644034 513146 644072
rect 513549 644244 513564 644250
rect 513598 644244 513613 644250
rect 513549 644192 513555 644244
rect 513607 644192 513613 644244
rect 513549 644180 513613 644192
rect 513549 644128 513555 644180
rect 513607 644128 513613 644180
rect 513549 644116 513613 644128
rect 513549 644064 513555 644116
rect 513607 644064 513613 644116
rect 513549 644058 513613 644064
rect 514016 644216 514022 644250
rect 514056 644216 514062 644250
rect 514016 644178 514062 644216
rect 514016 644144 514022 644178
rect 514056 644144 514062 644178
rect 514016 644106 514062 644144
rect 514016 644072 514022 644106
rect 514056 644072 514062 644106
rect 513100 644000 513106 644034
rect 513140 644000 513146 644034
rect 513100 643962 513146 644000
rect 513100 643928 513106 643962
rect 513140 643928 513146 643962
rect 513100 643890 513146 643928
rect 513100 643856 513106 643890
rect 513140 643856 513146 643890
rect 513100 643818 513146 643856
rect 513100 643785 513106 643818
rect 512642 643746 512688 643784
rect 512642 643712 512648 643746
rect 512682 643712 512688 643746
rect 512642 643674 512688 643712
rect 512642 643640 512648 643674
rect 512682 643640 512688 643674
rect 512642 643602 512688 643640
rect 512224 643568 512230 643593
rect 512184 643530 512230 643568
rect 512184 643496 512190 643530
rect 512224 643496 512230 643530
rect 512184 643458 512230 643496
rect 512184 643424 512190 643458
rect 512224 643424 512230 643458
rect 512184 643386 512230 643424
rect 512184 643352 512190 643386
rect 512224 643352 512230 643386
rect 512184 643337 512230 643352
rect 512642 643568 512648 643602
rect 512682 643568 512688 643602
rect 513091 643784 513106 643785
rect 513140 643785 513146 643818
rect 513558 644034 513604 644058
rect 513558 644000 513564 644034
rect 513598 644000 513604 644034
rect 513558 643962 513604 644000
rect 513558 643928 513564 643962
rect 513598 643928 513604 643962
rect 513558 643890 513604 643928
rect 513558 643856 513564 643890
rect 513598 643856 513604 643890
rect 513558 643818 513604 643856
rect 513140 643784 513155 643785
rect 513091 643779 513155 643784
rect 513091 643727 513097 643779
rect 513149 643727 513155 643779
rect 513091 643715 513106 643727
rect 513140 643715 513155 643727
rect 513091 643663 513097 643715
rect 513149 643663 513155 643715
rect 513091 643651 513106 643663
rect 513140 643651 513155 643663
rect 513091 643599 513097 643651
rect 513149 643599 513155 643651
rect 513091 643593 513106 643599
rect 512642 643530 512688 643568
rect 512642 643496 512648 643530
rect 512682 643496 512688 643530
rect 512642 643458 512688 643496
rect 512642 643424 512648 643458
rect 512682 643424 512688 643458
rect 512642 643386 512688 643424
rect 512642 643352 512648 643386
rect 512682 643352 512688 643386
rect 512642 643337 512688 643352
rect 513100 643568 513106 643593
rect 513140 643593 513155 643599
rect 513558 643784 513564 643818
rect 513598 643784 513604 643818
rect 514016 644034 514062 644072
rect 514016 644000 514022 644034
rect 514056 644000 514062 644034
rect 514016 643962 514062 644000
rect 514016 643928 514022 643962
rect 514056 643928 514062 643962
rect 514016 643890 514062 643928
rect 514016 643856 514022 643890
rect 514056 643856 514062 643890
rect 514016 643818 514062 643856
rect 514016 643785 514022 643818
rect 513558 643746 513604 643784
rect 513558 643712 513564 643746
rect 513598 643712 513604 643746
rect 513558 643674 513604 643712
rect 513558 643640 513564 643674
rect 513598 643640 513604 643674
rect 513558 643602 513604 643640
rect 513140 643568 513146 643593
rect 513100 643530 513146 643568
rect 513100 643496 513106 643530
rect 513140 643496 513146 643530
rect 513100 643458 513146 643496
rect 513100 643424 513106 643458
rect 513140 643424 513146 643458
rect 513100 643386 513146 643424
rect 513100 643352 513106 643386
rect 513140 643352 513146 643386
rect 513100 643337 513146 643352
rect 513558 643568 513564 643602
rect 513598 643568 513604 643602
rect 514007 643784 514022 643785
rect 514056 643785 514062 643818
rect 514474 644322 514520 644337
rect 514474 644288 514480 644322
rect 514514 644288 514520 644322
rect 514474 644250 514520 644288
rect 514474 644216 514480 644250
rect 514514 644216 514520 644250
rect 514474 644178 514520 644216
rect 514474 644144 514480 644178
rect 514514 644144 514520 644178
rect 514474 644106 514520 644144
rect 514474 644072 514480 644106
rect 514514 644072 514520 644106
rect 514474 644034 514520 644072
rect 514474 644000 514480 644034
rect 514514 644000 514520 644034
rect 514474 643962 514520 644000
rect 514474 643928 514480 643962
rect 514514 643928 514520 643962
rect 514474 643890 514520 643928
rect 514474 643856 514480 643890
rect 514514 643856 514520 643890
rect 514474 643818 514520 643856
rect 514474 643785 514480 643818
rect 514056 643784 514071 643785
rect 514007 643779 514071 643784
rect 514007 643727 514013 643779
rect 514065 643727 514071 643779
rect 514007 643715 514022 643727
rect 514056 643715 514071 643727
rect 514007 643663 514013 643715
rect 514065 643663 514071 643715
rect 514007 643651 514022 643663
rect 514056 643651 514071 643663
rect 514007 643599 514013 643651
rect 514065 643599 514071 643651
rect 514007 643593 514022 643599
rect 513558 643530 513604 643568
rect 513558 643496 513564 643530
rect 513598 643496 513604 643530
rect 513558 643458 513604 643496
rect 513558 643424 513564 643458
rect 513598 643424 513604 643458
rect 513558 643386 513604 643424
rect 513558 643352 513564 643386
rect 513598 643352 513604 643386
rect 513558 643337 513604 643352
rect 514016 643568 514022 643593
rect 514056 643593 514071 643599
rect 514465 643784 514480 643785
rect 514514 643785 514520 643818
rect 514932 644322 514978 644337
rect 514932 644288 514938 644322
rect 514972 644288 514978 644322
rect 514932 644250 514978 644288
rect 514932 644216 514938 644250
rect 514972 644216 514978 644250
rect 514932 644178 514978 644216
rect 514932 644144 514938 644178
rect 514972 644144 514978 644178
rect 514932 644106 514978 644144
rect 514932 644072 514938 644106
rect 514972 644072 514978 644106
rect 514932 644034 514978 644072
rect 514932 644000 514938 644034
rect 514972 644000 514978 644034
rect 514932 643962 514978 644000
rect 514932 643928 514938 643962
rect 514972 643928 514978 643962
rect 514932 643890 514978 643928
rect 514932 643856 514938 643890
rect 514972 643856 514978 643890
rect 514932 643818 514978 643856
rect 514932 643785 514938 643818
rect 514514 643784 514529 643785
rect 514465 643779 514529 643784
rect 514465 643727 514471 643779
rect 514523 643727 514529 643779
rect 514465 643715 514480 643727
rect 514514 643715 514529 643727
rect 514465 643663 514471 643715
rect 514523 643663 514529 643715
rect 514465 643651 514480 643663
rect 514514 643651 514529 643663
rect 514465 643599 514471 643651
rect 514523 643599 514529 643651
rect 514465 643593 514480 643599
rect 514056 643568 514062 643593
rect 514016 643530 514062 643568
rect 514016 643496 514022 643530
rect 514056 643496 514062 643530
rect 514016 643458 514062 643496
rect 514016 643424 514022 643458
rect 514056 643424 514062 643458
rect 514016 643386 514062 643424
rect 514016 643352 514022 643386
rect 514056 643352 514062 643386
rect 509492 643296 509538 643337
rect 514016 643296 514062 643352
rect 514474 643568 514480 643593
rect 514514 643593 514529 643599
rect 514923 643784 514938 643785
rect 514972 643785 514978 643818
rect 515390 644322 515436 644337
rect 515390 644288 515396 644322
rect 515430 644288 515436 644322
rect 515390 644250 515436 644288
rect 515390 644216 515396 644250
rect 515430 644216 515436 644250
rect 515390 644178 515436 644216
rect 515757 644315 515763 644367
rect 515815 644315 515821 644367
rect 515757 644303 515821 644315
rect 515757 644251 515763 644303
rect 515815 644251 515821 644303
rect 515757 644248 515772 644251
rect 515806 644248 515821 644251
rect 515757 644239 515821 644248
rect 515757 644187 515763 644239
rect 515815 644187 515821 644239
rect 515757 644181 515772 644187
rect 515390 644144 515396 644178
rect 515430 644144 515436 644178
rect 515390 644106 515436 644144
rect 515390 644072 515396 644106
rect 515430 644072 515436 644106
rect 515390 644034 515436 644072
rect 515390 644000 515396 644034
rect 515430 644000 515436 644034
rect 515390 643962 515436 644000
rect 515390 643928 515396 643962
rect 515430 643928 515436 643962
rect 515390 643890 515436 643928
rect 515390 643856 515396 643890
rect 515430 643856 515436 643890
rect 515390 643818 515436 643856
rect 515390 643785 515396 643818
rect 514972 643784 514987 643785
rect 514923 643779 514987 643784
rect 514923 643727 514929 643779
rect 514981 643727 514987 643779
rect 514923 643715 514938 643727
rect 514972 643715 514987 643727
rect 514923 643663 514929 643715
rect 514981 643663 514987 643715
rect 514923 643651 514938 643663
rect 514972 643651 514987 643663
rect 514923 643599 514929 643651
rect 514981 643599 514987 643651
rect 514923 643593 514938 643599
rect 514514 643568 514520 643593
rect 514474 643530 514520 643568
rect 514474 643496 514480 643530
rect 514514 643496 514520 643530
rect 514474 643458 514520 643496
rect 514474 643424 514480 643458
rect 514514 643424 514520 643458
rect 514474 643386 514520 643424
rect 514474 643352 514480 643386
rect 514514 643352 514520 643386
rect 514474 643296 514520 643352
rect 514932 643568 514938 643593
rect 514972 643593 514987 643599
rect 515381 643784 515396 643785
rect 515430 643785 515436 643818
rect 515766 644176 515772 644181
rect 515806 644181 515821 644187
rect 516224 644536 516230 644570
rect 516264 644536 516270 644570
rect 516682 644858 516728 644896
rect 516682 644824 516688 644858
rect 516722 644824 516728 644858
rect 516682 644786 516728 644824
rect 516682 644752 516688 644786
rect 516722 644752 516728 644786
rect 516682 644714 516728 644752
rect 516682 644680 516688 644714
rect 516722 644680 516728 644714
rect 516682 644642 516728 644680
rect 516682 644608 516688 644642
rect 516722 644608 516728 644642
rect 516682 644570 516728 644608
rect 516682 644565 516688 644570
rect 516224 644498 516270 644536
rect 516224 644464 516230 644498
rect 516264 644464 516270 644498
rect 516224 644426 516270 644464
rect 516224 644392 516230 644426
rect 516264 644392 516270 644426
rect 516224 644354 516270 644392
rect 516224 644320 516230 644354
rect 516264 644320 516270 644354
rect 516224 644282 516270 644320
rect 516224 644248 516230 644282
rect 516264 644248 516270 644282
rect 516224 644210 516270 644248
rect 515806 644176 515812 644181
rect 515766 644138 515812 644176
rect 515766 644104 515772 644138
rect 515806 644104 515812 644138
rect 515766 644066 515812 644104
rect 515766 644032 515772 644066
rect 515806 644032 515812 644066
rect 515766 643994 515812 644032
rect 515766 643960 515772 643994
rect 515806 643960 515812 643994
rect 515766 643922 515812 643960
rect 515766 643888 515772 643922
rect 515806 643888 515812 643922
rect 515766 643850 515812 643888
rect 515766 643816 515772 643850
rect 515806 643816 515812 643850
rect 515572 643785 515630 643790
rect 515430 643784 515445 643785
rect 515381 643779 515445 643784
rect 515381 643727 515387 643779
rect 515439 643727 515445 643779
rect 515381 643715 515396 643727
rect 515430 643715 515445 643727
rect 515381 643663 515387 643715
rect 515439 643663 515445 643715
rect 515381 643651 515396 643663
rect 515430 643651 515445 643663
rect 515381 643599 515387 643651
rect 515439 643599 515445 643651
rect 515381 643593 515396 643599
rect 514972 643568 514978 643593
rect 514932 643530 514978 643568
rect 514932 643496 514938 643530
rect 514972 643496 514978 643530
rect 514932 643458 514978 643496
rect 514932 643424 514938 643458
rect 514972 643424 514978 643458
rect 514932 643386 514978 643424
rect 514932 643352 514938 643386
rect 514972 643352 514978 643386
rect 514932 643296 514978 643352
rect 515390 643568 515396 643593
rect 515430 643593 515445 643599
rect 515569 643779 515633 643785
rect 515569 643727 515575 643779
rect 515627 643727 515633 643779
rect 515569 643715 515633 643727
rect 515569 643663 515575 643715
rect 515627 643663 515633 643715
rect 515569 643651 515633 643663
rect 515569 643599 515575 643651
rect 515627 643599 515633 643651
rect 515569 643593 515633 643599
rect 515766 643778 515812 643816
rect 515766 643744 515772 643778
rect 515806 643744 515812 643778
rect 515766 643706 515812 643744
rect 515766 643672 515772 643706
rect 515806 643672 515812 643706
rect 515766 643634 515812 643672
rect 515766 643600 515772 643634
rect 515806 643600 515812 643634
rect 515430 643568 515436 643593
rect 515572 643588 515630 643593
rect 515390 643530 515436 643568
rect 515390 643496 515396 643530
rect 515430 643496 515436 643530
rect 515390 643458 515436 643496
rect 515390 643424 515396 643458
rect 515430 643424 515436 643458
rect 515390 643386 515436 643424
rect 515390 643352 515396 643386
rect 515430 643352 515436 643386
rect 515390 643337 515436 643352
rect 515766 643562 515812 643600
rect 515766 643528 515772 643562
rect 515806 643528 515812 643562
rect 515766 643490 515812 643528
rect 515766 643456 515772 643490
rect 515806 643456 515812 643490
rect 515766 643418 515812 643456
rect 515766 643384 515772 643418
rect 515806 643384 515812 643418
rect 515766 643337 515812 643384
rect 516224 644176 516230 644210
rect 516264 644176 516270 644210
rect 516673 644559 516688 644565
rect 516722 644565 516728 644570
rect 516722 644559 516737 644565
rect 516673 644507 516679 644559
rect 516731 644507 516737 644559
rect 516673 644498 516737 644507
rect 516673 644495 516688 644498
rect 516722 644495 516737 644498
rect 516673 644443 516679 644495
rect 516731 644443 516737 644495
rect 516673 644431 516737 644443
rect 516673 644379 516679 644431
rect 516731 644379 516737 644431
rect 516673 644367 516737 644379
rect 516673 644315 516679 644367
rect 516731 644315 516737 644367
rect 516673 644303 516737 644315
rect 516673 644251 516679 644303
rect 516731 644251 516737 644303
rect 516673 644248 516688 644251
rect 516722 644248 516737 644251
rect 516673 644239 516737 644248
rect 516673 644187 516679 644239
rect 516731 644187 516737 644239
rect 516673 644181 516688 644187
rect 516224 644138 516270 644176
rect 516224 644104 516230 644138
rect 516264 644104 516270 644138
rect 516224 644066 516270 644104
rect 516224 644032 516230 644066
rect 516264 644032 516270 644066
rect 516224 643994 516270 644032
rect 516224 643960 516230 643994
rect 516264 643960 516270 643994
rect 516224 643922 516270 643960
rect 516224 643888 516230 643922
rect 516264 643888 516270 643922
rect 516224 643850 516270 643888
rect 516224 643816 516230 643850
rect 516264 643816 516270 643850
rect 516224 643778 516270 643816
rect 516224 643744 516230 643778
rect 516264 643744 516270 643778
rect 516224 643706 516270 643744
rect 516224 643672 516230 643706
rect 516264 643672 516270 643706
rect 516224 643634 516270 643672
rect 516224 643600 516230 643634
rect 516264 643600 516270 643634
rect 516224 643562 516270 643600
rect 516224 643528 516230 643562
rect 516264 643528 516270 643562
rect 516224 643490 516270 643528
rect 516224 643456 516230 643490
rect 516264 643456 516270 643490
rect 516224 643418 516270 643456
rect 516224 643384 516230 643418
rect 516264 643384 516270 643418
rect 516224 643337 516270 643384
rect 516682 644176 516688 644181
rect 516722 644181 516737 644187
rect 516722 644176 516728 644181
rect 516682 644138 516728 644176
rect 516682 644104 516688 644138
rect 516722 644104 516728 644138
rect 516682 644066 516728 644104
rect 516682 644032 516688 644066
rect 516722 644032 516728 644066
rect 516682 643994 516728 644032
rect 516682 643960 516688 643994
rect 516722 643960 516728 643994
rect 516682 643922 516728 643960
rect 516682 643888 516688 643922
rect 516722 643888 516728 643922
rect 516682 643850 516728 643888
rect 516682 643816 516688 643850
rect 516722 643816 516728 643850
rect 516682 643778 516728 643816
rect 516682 643744 516688 643778
rect 516722 643744 516728 643778
rect 516682 643706 516728 643744
rect 516682 643672 516688 643706
rect 516722 643672 516728 643706
rect 516682 643634 516728 643672
rect 516682 643600 516688 643634
rect 516722 643600 516728 643634
rect 516682 643562 516728 643600
rect 516682 643528 516688 643562
rect 516722 643528 516728 643562
rect 516682 643490 516728 643528
rect 516682 643456 516688 643490
rect 516722 643456 516728 643490
rect 516682 643418 516728 643456
rect 516682 643384 516688 643418
rect 516722 643384 516728 643418
rect 516682 643337 516728 643384
rect 516348 643299 516604 643305
rect 516348 643296 516354 643299
rect 508062 643290 508510 643296
rect 508062 643256 508153 643290
rect 508187 643256 508225 643290
rect 508259 643256 508297 643290
rect 508331 643256 508369 643290
rect 508403 643256 508441 643290
rect 508475 643256 508510 643290
rect 508062 643250 508510 643256
rect 508576 643290 509426 643296
rect 508576 643256 508611 643290
rect 508645 643256 508683 643290
rect 508717 643256 508755 643290
rect 508789 643256 508827 643290
rect 508861 643256 508879 643290
rect 508933 643256 508943 643290
rect 508576 643250 508879 643256
rect 508873 643238 508879 643250
rect 508931 643238 508943 643256
rect 508995 643238 509007 643290
rect 509059 643256 509069 643290
rect 509123 643256 509141 643290
rect 509175 643256 509213 643290
rect 509247 643256 509285 643290
rect 509319 643256 509357 643290
rect 509391 643256 509426 643290
rect 509059 643238 509071 643256
rect 509123 643250 509426 643256
rect 509492 643290 509884 643296
rect 509492 643256 509527 643290
rect 509561 643256 509599 643290
rect 509633 643256 509671 643290
rect 509705 643256 509743 643290
rect 509777 643256 509815 643290
rect 509849 643256 509884 643290
rect 509492 643250 509884 643256
rect 509950 643290 511716 643296
rect 509950 643256 509985 643290
rect 510019 643256 510057 643290
rect 510091 643256 510129 643290
rect 510163 643256 510201 643290
rect 510235 643256 510273 643290
rect 510307 643256 510443 643290
rect 510477 643256 510515 643290
rect 510549 643256 510587 643290
rect 510621 643256 510659 643290
rect 510693 643256 510711 643290
rect 510765 643256 510775 643290
rect 509950 643250 510711 643256
rect 509123 643238 509129 643250
rect 508873 643232 509129 643238
rect 510705 643238 510711 643250
rect 510763 643238 510775 643256
rect 510827 643238 510839 643290
rect 510891 643256 510901 643290
rect 510955 643256 510973 643290
rect 511007 643256 511045 643290
rect 511079 643256 511117 643290
rect 511151 643256 511189 643290
rect 511223 643256 511359 643290
rect 511393 643256 511431 643290
rect 511465 643256 511503 643290
rect 511537 643256 511575 643290
rect 511609 643256 511647 643290
rect 511681 643256 511716 643290
rect 510891 643238 510903 643256
rect 510955 643250 511716 643256
rect 511782 643290 513548 643296
rect 511782 643256 511817 643290
rect 511851 643256 511889 643290
rect 511923 643256 511961 643290
rect 511995 643256 512033 643290
rect 512067 643256 512105 643290
rect 512139 643256 512275 643290
rect 512309 643256 512347 643290
rect 512381 643256 512419 643290
rect 512453 643256 512491 643290
rect 512525 643256 512543 643290
rect 512597 643256 512607 643290
rect 511782 643250 512543 643256
rect 510955 643238 510961 643250
rect 510705 643232 510961 643238
rect 512537 643238 512543 643250
rect 512595 643238 512607 643256
rect 512659 643238 512671 643290
rect 512723 643256 512733 643290
rect 512787 643256 512805 643290
rect 512839 643256 512877 643290
rect 512911 643256 512949 643290
rect 512983 643256 513021 643290
rect 513055 643256 513191 643290
rect 513225 643256 513263 643290
rect 513297 643256 513335 643290
rect 513369 643256 513407 643290
rect 513441 643256 513479 643290
rect 513513 643256 513548 643290
rect 512723 643238 512735 643256
rect 512787 643250 513548 643256
rect 513614 643290 515380 643296
rect 513614 643256 513649 643290
rect 513683 643256 513721 643290
rect 513755 643256 513793 643290
rect 513827 643256 513865 643290
rect 513899 643256 513937 643290
rect 513971 643256 514107 643290
rect 514141 643256 514179 643290
rect 514213 643256 514251 643290
rect 514285 643256 514323 643290
rect 514357 643256 514395 643290
rect 514429 643256 514565 643290
rect 514599 643256 514637 643290
rect 514671 643256 514709 643290
rect 514743 643256 514781 643290
rect 514815 643256 514853 643290
rect 514887 643256 515023 643290
rect 515057 643256 515095 643290
rect 515129 643256 515167 643290
rect 515201 643256 515239 643290
rect 515273 643256 515311 643290
rect 515345 643256 515380 643290
rect 513614 643250 515380 643256
rect 515822 643290 516214 643296
rect 515822 643256 515857 643290
rect 515891 643256 515929 643290
rect 515963 643256 516001 643290
rect 516035 643256 516073 643290
rect 516107 643256 516145 643290
rect 516179 643256 516214 643290
rect 515822 643250 516214 643256
rect 516280 643290 516354 643296
rect 516406 643290 516418 643299
rect 516470 643290 516482 643299
rect 516534 643290 516546 643299
rect 516598 643296 516604 643299
rect 516598 643290 516672 643296
rect 516280 643256 516315 643290
rect 516349 643256 516354 643290
rect 516598 643256 516603 643290
rect 516637 643256 516672 643290
rect 516280 643250 516354 643256
rect 512787 643238 512793 643250
rect 512537 643232 512793 643238
rect 515968 642914 516068 643250
rect 516348 643247 516354 643250
rect 516406 643247 516418 643256
rect 516470 643247 516482 643256
rect 516534 643247 516546 643256
rect 516598 643250 516672 643256
rect 516598 643247 516604 643250
rect 516348 643241 516604 643247
rect 515954 642908 516082 642914
rect 515954 642792 515960 642908
rect 516076 642792 516082 642908
rect 515954 642786 516082 642792
rect 508873 642495 509129 642501
rect 508873 642483 508879 642495
rect 508062 642477 508510 642483
rect 508062 642443 508153 642477
rect 508187 642443 508225 642477
rect 508259 642443 508297 642477
rect 508331 642443 508369 642477
rect 508403 642443 508441 642477
rect 508475 642443 508510 642477
rect 508062 642437 508510 642443
rect 508576 642477 508879 642483
rect 508931 642477 508943 642495
rect 508576 642443 508611 642477
rect 508645 642443 508683 642477
rect 508717 642443 508755 642477
rect 508789 642443 508827 642477
rect 508861 642443 508879 642477
rect 508933 642443 508943 642477
rect 508995 642443 509007 642495
rect 509059 642477 509071 642495
rect 509123 642483 509129 642495
rect 510705 642495 510961 642501
rect 510705 642483 510711 642495
rect 509123 642477 509426 642483
rect 509059 642443 509069 642477
rect 509123 642443 509141 642477
rect 509175 642443 509213 642477
rect 509247 642443 509285 642477
rect 509319 642443 509357 642477
rect 509391 642443 509426 642477
rect 508576 642437 509426 642443
rect 509492 642477 509884 642483
rect 509492 642443 509527 642477
rect 509561 642443 509599 642477
rect 509633 642443 509671 642477
rect 509705 642443 509743 642477
rect 509777 642443 509815 642477
rect 509849 642443 509884 642477
rect 509492 642437 509884 642443
rect 509950 642477 510711 642483
rect 510763 642477 510775 642495
rect 509950 642443 509985 642477
rect 510019 642443 510057 642477
rect 510091 642443 510129 642477
rect 510163 642443 510201 642477
rect 510235 642443 510273 642477
rect 510307 642443 510443 642477
rect 510477 642443 510515 642477
rect 510549 642443 510587 642477
rect 510621 642443 510659 642477
rect 510693 642443 510711 642477
rect 510765 642443 510775 642477
rect 510827 642443 510839 642495
rect 510891 642477 510903 642495
rect 510955 642483 510961 642495
rect 512537 642495 512793 642501
rect 512537 642483 512543 642495
rect 510955 642477 511716 642483
rect 510891 642443 510901 642477
rect 510955 642443 510973 642477
rect 511007 642443 511045 642477
rect 511079 642443 511117 642477
rect 511151 642443 511189 642477
rect 511223 642443 511359 642477
rect 511393 642443 511431 642477
rect 511465 642443 511503 642477
rect 511537 642443 511575 642477
rect 511609 642443 511647 642477
rect 511681 642443 511716 642477
rect 509950 642437 511716 642443
rect 511782 642477 512543 642483
rect 512595 642477 512607 642495
rect 511782 642443 511817 642477
rect 511851 642443 511889 642477
rect 511923 642443 511961 642477
rect 511995 642443 512033 642477
rect 512067 642443 512105 642477
rect 512139 642443 512275 642477
rect 512309 642443 512347 642477
rect 512381 642443 512419 642477
rect 512453 642443 512491 642477
rect 512525 642443 512543 642477
rect 512597 642443 512607 642477
rect 512659 642443 512671 642495
rect 512723 642477 512735 642495
rect 512787 642483 512793 642495
rect 515968 642483 516068 642786
rect 516347 642486 516603 642492
rect 516347 642483 516353 642486
rect 512787 642477 513548 642483
rect 512723 642443 512733 642477
rect 512787 642443 512805 642477
rect 512839 642443 512877 642477
rect 512911 642443 512949 642477
rect 512983 642443 513021 642477
rect 513055 642443 513191 642477
rect 513225 642443 513263 642477
rect 513297 642443 513335 642477
rect 513369 642443 513407 642477
rect 513441 642443 513479 642477
rect 513513 642443 513548 642477
rect 511782 642437 513548 642443
rect 513614 642477 515380 642483
rect 513614 642443 513649 642477
rect 513683 642443 513721 642477
rect 513755 642443 513793 642477
rect 513827 642443 513865 642477
rect 513899 642443 513937 642477
rect 513971 642443 514107 642477
rect 514141 642443 514179 642477
rect 514213 642443 514251 642477
rect 514285 642443 514323 642477
rect 514357 642443 514395 642477
rect 514429 642443 514565 642477
rect 514599 642443 514637 642477
rect 514671 642443 514709 642477
rect 514743 642443 514781 642477
rect 514815 642443 514853 642477
rect 514887 642443 515023 642477
rect 515057 642443 515095 642477
rect 515129 642443 515167 642477
rect 515201 642443 515239 642477
rect 515273 642443 515311 642477
rect 515345 642443 515380 642477
rect 513614 642437 515380 642443
rect 515822 642477 516214 642483
rect 515822 642443 515857 642477
rect 515891 642443 515929 642477
rect 515963 642443 516001 642477
rect 516035 642443 516073 642477
rect 516107 642443 516145 642477
rect 516179 642443 516214 642477
rect 515822 642437 516214 642443
rect 516280 642477 516353 642483
rect 516405 642477 516417 642486
rect 516469 642477 516481 642486
rect 516533 642477 516545 642486
rect 516597 642483 516603 642486
rect 516597 642477 516672 642483
rect 516280 642443 516315 642477
rect 516349 642443 516353 642477
rect 516597 642443 516603 642477
rect 516637 642443 516672 642477
rect 516280 642437 516353 642443
rect 508062 642390 508108 642437
rect 509492 642405 509538 642437
rect 508062 642356 508068 642390
rect 508102 642356 508108 642390
rect 508062 642318 508108 642356
rect 508062 642284 508068 642318
rect 508102 642284 508108 642318
rect 508062 642246 508108 642284
rect 508062 642212 508068 642246
rect 508102 642212 508108 642246
rect 508062 642174 508108 642212
rect 507868 642149 507926 642154
rect 508062 642149 508068 642174
rect 507865 642143 507929 642149
rect 507865 642091 507871 642143
rect 507923 642091 507929 642143
rect 507865 642079 507929 642091
rect 507865 642027 507871 642079
rect 507923 642027 507929 642079
rect 507865 642015 507929 642027
rect 507865 641963 507871 642015
rect 507923 641963 507929 642015
rect 507865 641957 507929 641963
rect 508053 642143 508068 642149
rect 508102 642149 508108 642174
rect 508520 642390 508566 642405
rect 508520 642356 508526 642390
rect 508560 642356 508566 642390
rect 508520 642318 508566 642356
rect 508520 642284 508526 642318
rect 508560 642284 508566 642318
rect 508520 642246 508566 642284
rect 508520 642212 508526 642246
rect 508560 642212 508566 642246
rect 508520 642174 508566 642212
rect 508520 642149 508526 642174
rect 508102 642143 508117 642149
rect 508053 642091 508059 642143
rect 508111 642091 508117 642143
rect 508053 642079 508068 642091
rect 508102 642079 508117 642091
rect 508053 642027 508059 642079
rect 508111 642027 508117 642079
rect 508053 642015 508068 642027
rect 508102 642015 508117 642027
rect 508053 641963 508059 642015
rect 508111 641963 508117 642015
rect 508053 641958 508117 641963
rect 508053 641957 508068 641958
rect 507868 641952 507926 641957
rect 508062 641924 508068 641957
rect 508102 641957 508117 641958
rect 508511 642143 508526 642149
rect 508560 642149 508566 642174
rect 508978 642390 509024 642405
rect 508978 642356 508984 642390
rect 509018 642356 509024 642390
rect 508978 642318 509024 642356
rect 508978 642284 508984 642318
rect 509018 642284 509024 642318
rect 508978 642246 509024 642284
rect 508978 642212 508984 642246
rect 509018 642212 509024 642246
rect 508978 642174 509024 642212
rect 508560 642143 508575 642149
rect 508511 642091 508517 642143
rect 508569 642091 508575 642143
rect 508511 642079 508526 642091
rect 508560 642079 508575 642091
rect 508511 642027 508517 642079
rect 508569 642027 508575 642079
rect 508511 642015 508526 642027
rect 508560 642015 508575 642027
rect 508511 641963 508517 642015
rect 508569 641963 508575 642015
rect 508511 641958 508575 641963
rect 508511 641957 508526 641958
rect 508102 641924 508108 641957
rect 508062 641886 508108 641924
rect 508062 641852 508068 641886
rect 508102 641852 508108 641886
rect 508062 641814 508108 641852
rect 508062 641780 508068 641814
rect 508102 641780 508108 641814
rect 508062 641742 508108 641780
rect 508062 641708 508068 641742
rect 508102 641708 508108 641742
rect 508062 641670 508108 641708
rect 508062 641636 508068 641670
rect 508102 641636 508108 641670
rect 508062 641598 508108 641636
rect 508062 641564 508068 641598
rect 508102 641564 508108 641598
rect 508062 641526 508108 641564
rect 508062 641492 508068 641526
rect 508102 641492 508108 641526
rect 508062 641454 508108 641492
rect 508062 641420 508068 641454
rect 508102 641420 508108 641454
rect 508062 641405 508108 641420
rect 508520 641924 508526 641957
rect 508560 641957 508575 641958
rect 508978 642140 508984 642174
rect 509018 642140 509024 642174
rect 509436 642390 509538 642405
rect 509436 642356 509442 642390
rect 509476 642359 509538 642390
rect 509894 642390 509940 642405
rect 509476 642356 509482 642359
rect 509436 642318 509482 642356
rect 509436 642284 509442 642318
rect 509476 642284 509482 642318
rect 509436 642246 509482 642284
rect 509436 642212 509442 642246
rect 509476 642212 509482 642246
rect 509436 642174 509482 642212
rect 509436 642149 509442 642174
rect 508978 642102 509024 642140
rect 508978 642068 508984 642102
rect 509018 642068 509024 642102
rect 508978 642030 509024 642068
rect 508978 641996 508984 642030
rect 509018 641996 509024 642030
rect 508978 641958 509024 641996
rect 508560 641924 508566 641957
rect 508520 641886 508566 641924
rect 508520 641852 508526 641886
rect 508560 641852 508566 641886
rect 508520 641814 508566 641852
rect 508520 641780 508526 641814
rect 508560 641780 508566 641814
rect 508520 641742 508566 641780
rect 508520 641708 508526 641742
rect 508560 641708 508566 641742
rect 508520 641670 508566 641708
rect 508978 641924 508984 641958
rect 509018 641924 509024 641958
rect 509427 642143 509442 642149
rect 509476 642149 509482 642174
rect 509894 642356 509900 642390
rect 509934 642356 509940 642390
rect 509894 642318 509940 642356
rect 509894 642284 509900 642318
rect 509934 642284 509940 642318
rect 509894 642246 509940 642284
rect 509894 642212 509900 642246
rect 509934 642212 509940 642246
rect 509894 642174 509940 642212
rect 509476 642143 509491 642149
rect 509427 642091 509433 642143
rect 509485 642091 509491 642143
rect 509427 642079 509442 642091
rect 509476 642079 509491 642091
rect 509427 642027 509433 642079
rect 509485 642027 509491 642079
rect 509427 642015 509442 642027
rect 509476 642015 509491 642027
rect 509427 641963 509433 642015
rect 509485 641963 509491 642015
rect 509427 641958 509491 641963
rect 509427 641957 509442 641958
rect 508978 641886 509024 641924
rect 508978 641852 508984 641886
rect 509018 641852 509024 641886
rect 508978 641814 509024 641852
rect 508978 641780 508984 641814
rect 509018 641780 509024 641814
rect 508978 641742 509024 641780
rect 508978 641708 508984 641742
rect 509018 641708 509024 641742
rect 508978 641684 509024 641708
rect 509436 641924 509442 641957
rect 509476 641957 509491 641958
rect 509894 642140 509900 642174
rect 509934 642140 509940 642174
rect 510352 642390 510398 642405
rect 510352 642356 510358 642390
rect 510392 642356 510398 642390
rect 510352 642318 510398 642356
rect 510352 642284 510358 642318
rect 510392 642284 510398 642318
rect 510352 642246 510398 642284
rect 510352 642212 510358 642246
rect 510392 642212 510398 642246
rect 510352 642174 510398 642212
rect 510352 642149 510358 642174
rect 509894 642102 509940 642140
rect 509894 642068 509900 642102
rect 509934 642068 509940 642102
rect 509894 642030 509940 642068
rect 509894 641996 509900 642030
rect 509934 641996 509940 642030
rect 509894 641958 509940 641996
rect 509476 641924 509482 641957
rect 509436 641886 509482 641924
rect 509436 641852 509442 641886
rect 509476 641852 509482 641886
rect 509436 641814 509482 641852
rect 509436 641780 509442 641814
rect 509476 641780 509482 641814
rect 509436 641742 509482 641780
rect 509436 641708 509442 641742
rect 509476 641708 509482 641742
rect 508520 641636 508526 641670
rect 508560 641636 508566 641670
rect 508520 641598 508566 641636
rect 508520 641564 508526 641598
rect 508560 641564 508566 641598
rect 508520 641526 508566 641564
rect 508520 641492 508526 641526
rect 508560 641492 508566 641526
rect 508969 641678 509033 641684
rect 508969 641626 508975 641678
rect 509027 641626 509033 641678
rect 508969 641614 509033 641626
rect 508969 641562 508975 641614
rect 509027 641562 509033 641614
rect 508969 641550 509033 641562
rect 508969 641498 508975 641550
rect 509027 641498 509033 641550
rect 508969 641492 508984 641498
rect 509018 641492 509033 641498
rect 509436 641670 509482 641708
rect 509894 641924 509900 641958
rect 509934 641924 509940 641958
rect 510343 642143 510358 642149
rect 510392 642149 510398 642174
rect 510810 642390 510856 642405
rect 510810 642356 510816 642390
rect 510850 642356 510856 642390
rect 510810 642318 510856 642356
rect 510810 642284 510816 642318
rect 510850 642284 510856 642318
rect 510810 642246 510856 642284
rect 510810 642212 510816 642246
rect 510850 642212 510856 642246
rect 510810 642174 510856 642212
rect 510392 642143 510407 642149
rect 510343 642091 510349 642143
rect 510401 642091 510407 642143
rect 510343 642079 510358 642091
rect 510392 642079 510407 642091
rect 510343 642027 510349 642079
rect 510401 642027 510407 642079
rect 510343 642015 510358 642027
rect 510392 642015 510407 642027
rect 510343 641963 510349 642015
rect 510401 641963 510407 642015
rect 510343 641958 510407 641963
rect 510343 641957 510358 641958
rect 509894 641886 509940 641924
rect 509894 641852 509900 641886
rect 509934 641852 509940 641886
rect 509894 641814 509940 641852
rect 509894 641780 509900 641814
rect 509934 641780 509940 641814
rect 509894 641742 509940 641780
rect 509894 641708 509900 641742
rect 509934 641708 509940 641742
rect 509894 641684 509940 641708
rect 510352 641924 510358 641957
rect 510392 641957 510407 641958
rect 510810 642140 510816 642174
rect 510850 642140 510856 642174
rect 511268 642390 511314 642405
rect 511268 642356 511274 642390
rect 511308 642356 511314 642390
rect 511268 642318 511314 642356
rect 511268 642284 511274 642318
rect 511308 642284 511314 642318
rect 511268 642246 511314 642284
rect 511268 642212 511274 642246
rect 511308 642212 511314 642246
rect 511268 642174 511314 642212
rect 511268 642149 511274 642174
rect 510810 642102 510856 642140
rect 510810 642068 510816 642102
rect 510850 642068 510856 642102
rect 510810 642030 510856 642068
rect 510810 641996 510816 642030
rect 510850 641996 510856 642030
rect 510810 641958 510856 641996
rect 510392 641924 510398 641957
rect 510352 641886 510398 641924
rect 510352 641852 510358 641886
rect 510392 641852 510398 641886
rect 510352 641814 510398 641852
rect 510352 641780 510358 641814
rect 510392 641780 510398 641814
rect 510352 641742 510398 641780
rect 510352 641708 510358 641742
rect 510392 641708 510398 641742
rect 509436 641636 509442 641670
rect 509476 641636 509482 641670
rect 509436 641598 509482 641636
rect 509436 641564 509442 641598
rect 509476 641564 509482 641598
rect 509436 641526 509482 641564
rect 509436 641492 509442 641526
rect 509476 641492 509482 641526
rect 509885 641678 509949 641684
rect 509885 641626 509891 641678
rect 509943 641626 509949 641678
rect 509885 641614 509949 641626
rect 509885 641562 509891 641614
rect 509943 641562 509949 641614
rect 509885 641550 509949 641562
rect 509885 641498 509891 641550
rect 509943 641498 509949 641550
rect 509885 641492 509900 641498
rect 509934 641492 509949 641498
rect 510352 641670 510398 641708
rect 510810 641924 510816 641958
rect 510850 641924 510856 641958
rect 511259 642143 511274 642149
rect 511308 642149 511314 642174
rect 511726 642390 511772 642405
rect 511726 642356 511732 642390
rect 511766 642356 511772 642390
rect 511726 642318 511772 642356
rect 511726 642284 511732 642318
rect 511766 642284 511772 642318
rect 511726 642246 511772 642284
rect 511726 642212 511732 642246
rect 511766 642212 511772 642246
rect 511726 642174 511772 642212
rect 511308 642143 511323 642149
rect 511259 642091 511265 642143
rect 511317 642091 511323 642143
rect 511259 642079 511274 642091
rect 511308 642079 511323 642091
rect 511259 642027 511265 642079
rect 511317 642027 511323 642079
rect 511259 642015 511274 642027
rect 511308 642015 511323 642027
rect 511259 641963 511265 642015
rect 511317 641963 511323 642015
rect 511259 641958 511323 641963
rect 511259 641957 511274 641958
rect 510810 641886 510856 641924
rect 510810 641852 510816 641886
rect 510850 641852 510856 641886
rect 510810 641814 510856 641852
rect 510810 641780 510816 641814
rect 510850 641780 510856 641814
rect 510810 641742 510856 641780
rect 510810 641708 510816 641742
rect 510850 641708 510856 641742
rect 510810 641684 510856 641708
rect 511268 641924 511274 641957
rect 511308 641957 511323 641958
rect 511726 642140 511732 642174
rect 511766 642140 511772 642174
rect 512184 642390 512230 642405
rect 512184 642356 512190 642390
rect 512224 642356 512230 642390
rect 512184 642318 512230 642356
rect 512184 642284 512190 642318
rect 512224 642284 512230 642318
rect 512184 642246 512230 642284
rect 512184 642212 512190 642246
rect 512224 642212 512230 642246
rect 512184 642174 512230 642212
rect 512184 642149 512190 642174
rect 511726 642102 511772 642140
rect 511726 642068 511732 642102
rect 511766 642068 511772 642102
rect 511726 642030 511772 642068
rect 511726 641996 511732 642030
rect 511766 641996 511772 642030
rect 511726 641958 511772 641996
rect 511308 641924 511314 641957
rect 511268 641886 511314 641924
rect 511268 641852 511274 641886
rect 511308 641852 511314 641886
rect 511268 641814 511314 641852
rect 511268 641780 511274 641814
rect 511308 641780 511314 641814
rect 511268 641742 511314 641780
rect 511268 641708 511274 641742
rect 511308 641708 511314 641742
rect 510352 641636 510358 641670
rect 510392 641636 510398 641670
rect 510352 641598 510398 641636
rect 510352 641564 510358 641598
rect 510392 641564 510398 641598
rect 510352 641526 510398 641564
rect 510352 641492 510358 641526
rect 510392 641492 510398 641526
rect 510801 641678 510865 641684
rect 510801 641626 510807 641678
rect 510859 641626 510865 641678
rect 510801 641614 510865 641626
rect 510801 641562 510807 641614
rect 510859 641562 510865 641614
rect 510801 641550 510865 641562
rect 510801 641498 510807 641550
rect 510859 641498 510865 641550
rect 510801 641492 510816 641498
rect 510850 641492 510865 641498
rect 511268 641670 511314 641708
rect 511726 641924 511732 641958
rect 511766 641924 511772 641958
rect 512175 642143 512190 642149
rect 512224 642149 512230 642174
rect 512642 642390 512688 642405
rect 512642 642356 512648 642390
rect 512682 642356 512688 642390
rect 512642 642318 512688 642356
rect 512642 642284 512648 642318
rect 512682 642284 512688 642318
rect 512642 642246 512688 642284
rect 512642 642212 512648 642246
rect 512682 642212 512688 642246
rect 512642 642174 512688 642212
rect 512224 642143 512239 642149
rect 512175 642091 512181 642143
rect 512233 642091 512239 642143
rect 512175 642079 512190 642091
rect 512224 642079 512239 642091
rect 512175 642027 512181 642079
rect 512233 642027 512239 642079
rect 512175 642015 512190 642027
rect 512224 642015 512239 642027
rect 512175 641963 512181 642015
rect 512233 641963 512239 642015
rect 512175 641958 512239 641963
rect 512175 641957 512190 641958
rect 511726 641886 511772 641924
rect 511726 641852 511732 641886
rect 511766 641852 511772 641886
rect 511726 641814 511772 641852
rect 511726 641780 511732 641814
rect 511766 641780 511772 641814
rect 511726 641742 511772 641780
rect 511726 641708 511732 641742
rect 511766 641708 511772 641742
rect 511726 641684 511772 641708
rect 512184 641924 512190 641957
rect 512224 641957 512239 641958
rect 512642 642140 512648 642174
rect 512682 642140 512688 642174
rect 513100 642390 513146 642405
rect 513100 642356 513106 642390
rect 513140 642356 513146 642390
rect 513100 642318 513146 642356
rect 513100 642284 513106 642318
rect 513140 642284 513146 642318
rect 513100 642246 513146 642284
rect 513100 642212 513106 642246
rect 513140 642212 513146 642246
rect 513100 642174 513146 642212
rect 513100 642149 513106 642174
rect 512642 642102 512688 642140
rect 512642 642068 512648 642102
rect 512682 642068 512688 642102
rect 512642 642030 512688 642068
rect 512642 641996 512648 642030
rect 512682 641996 512688 642030
rect 512642 641958 512688 641996
rect 512224 641924 512230 641957
rect 512184 641886 512230 641924
rect 512184 641852 512190 641886
rect 512224 641852 512230 641886
rect 512184 641814 512230 641852
rect 512184 641780 512190 641814
rect 512224 641780 512230 641814
rect 512184 641742 512230 641780
rect 512184 641708 512190 641742
rect 512224 641708 512230 641742
rect 511268 641636 511274 641670
rect 511308 641636 511314 641670
rect 511268 641598 511314 641636
rect 511268 641564 511274 641598
rect 511308 641564 511314 641598
rect 511268 641526 511314 641564
rect 511268 641492 511274 641526
rect 511308 641492 511314 641526
rect 511717 641678 511781 641684
rect 511717 641626 511723 641678
rect 511775 641626 511781 641678
rect 511717 641614 511781 641626
rect 511717 641562 511723 641614
rect 511775 641562 511781 641614
rect 511717 641550 511781 641562
rect 511717 641498 511723 641550
rect 511775 641498 511781 641550
rect 511717 641492 511732 641498
rect 511766 641492 511781 641498
rect 512184 641670 512230 641708
rect 512642 641924 512648 641958
rect 512682 641924 512688 641958
rect 513091 642143 513106 642149
rect 513140 642149 513146 642174
rect 513558 642390 513604 642405
rect 513558 642356 513564 642390
rect 513598 642356 513604 642390
rect 513558 642318 513604 642356
rect 513558 642284 513564 642318
rect 513598 642284 513604 642318
rect 513558 642246 513604 642284
rect 513558 642212 513564 642246
rect 513598 642212 513604 642246
rect 513558 642174 513604 642212
rect 513140 642143 513155 642149
rect 513091 642091 513097 642143
rect 513149 642091 513155 642143
rect 513091 642079 513106 642091
rect 513140 642079 513155 642091
rect 513091 642027 513097 642079
rect 513149 642027 513155 642079
rect 513091 642015 513106 642027
rect 513140 642015 513155 642027
rect 513091 641963 513097 642015
rect 513149 641963 513155 642015
rect 513091 641958 513155 641963
rect 513091 641957 513106 641958
rect 512642 641886 512688 641924
rect 512642 641852 512648 641886
rect 512682 641852 512688 641886
rect 512642 641814 512688 641852
rect 512642 641780 512648 641814
rect 512682 641780 512688 641814
rect 512642 641742 512688 641780
rect 512642 641708 512648 641742
rect 512682 641708 512688 641742
rect 512642 641684 512688 641708
rect 513100 641924 513106 641957
rect 513140 641957 513155 641958
rect 513558 642140 513564 642174
rect 513598 642140 513604 642174
rect 514016 642390 514062 642437
rect 514016 642356 514022 642390
rect 514056 642356 514062 642390
rect 514016 642318 514062 642356
rect 514016 642284 514022 642318
rect 514056 642284 514062 642318
rect 514016 642246 514062 642284
rect 514016 642212 514022 642246
rect 514056 642212 514062 642246
rect 514016 642174 514062 642212
rect 514016 642149 514022 642174
rect 513558 642102 513604 642140
rect 513558 642068 513564 642102
rect 513598 642068 513604 642102
rect 513558 642030 513604 642068
rect 513558 641996 513564 642030
rect 513598 641996 513604 642030
rect 513558 641958 513604 641996
rect 513140 641924 513146 641957
rect 513100 641886 513146 641924
rect 513100 641852 513106 641886
rect 513140 641852 513146 641886
rect 513100 641814 513146 641852
rect 513100 641780 513106 641814
rect 513140 641780 513146 641814
rect 513100 641742 513146 641780
rect 513100 641708 513106 641742
rect 513140 641708 513146 641742
rect 512184 641636 512190 641670
rect 512224 641636 512230 641670
rect 512184 641598 512230 641636
rect 512184 641564 512190 641598
rect 512224 641564 512230 641598
rect 512184 641526 512230 641564
rect 512184 641492 512190 641526
rect 512224 641492 512230 641526
rect 512633 641678 512697 641684
rect 512633 641626 512639 641678
rect 512691 641626 512697 641678
rect 512633 641614 512697 641626
rect 512633 641562 512639 641614
rect 512691 641562 512697 641614
rect 512633 641550 512697 641562
rect 512633 641498 512639 641550
rect 512691 641498 512697 641550
rect 512633 641492 512648 641498
rect 512682 641492 512697 641498
rect 513100 641670 513146 641708
rect 513558 641924 513564 641958
rect 513598 641924 513604 641958
rect 514007 642143 514022 642149
rect 514056 642149 514062 642174
rect 514474 642390 514520 642437
rect 514474 642356 514480 642390
rect 514514 642356 514520 642390
rect 514474 642318 514520 642356
rect 514474 642284 514480 642318
rect 514514 642284 514520 642318
rect 514474 642246 514520 642284
rect 514474 642212 514480 642246
rect 514514 642212 514520 642246
rect 514474 642174 514520 642212
rect 514474 642149 514480 642174
rect 514056 642143 514071 642149
rect 514007 642091 514013 642143
rect 514065 642091 514071 642143
rect 514007 642079 514022 642091
rect 514056 642079 514071 642091
rect 514007 642027 514013 642079
rect 514065 642027 514071 642079
rect 514007 642015 514022 642027
rect 514056 642015 514071 642027
rect 514007 641963 514013 642015
rect 514065 641963 514071 642015
rect 514007 641958 514071 641963
rect 514007 641957 514022 641958
rect 513558 641886 513604 641924
rect 513558 641852 513564 641886
rect 513598 641852 513604 641886
rect 513558 641814 513604 641852
rect 513558 641780 513564 641814
rect 513598 641780 513604 641814
rect 513558 641742 513604 641780
rect 513558 641708 513564 641742
rect 513598 641708 513604 641742
rect 513558 641684 513604 641708
rect 514016 641924 514022 641957
rect 514056 641957 514071 641958
rect 514465 642143 514480 642149
rect 514514 642149 514520 642174
rect 514932 642390 514978 642437
rect 516347 642434 516353 642437
rect 516405 642434 516417 642443
rect 516469 642434 516481 642443
rect 516533 642434 516545 642443
rect 516597 642437 516672 642443
rect 516597 642434 516603 642437
rect 516347 642428 516603 642434
rect 514932 642356 514938 642390
rect 514972 642356 514978 642390
rect 514932 642318 514978 642356
rect 514932 642284 514938 642318
rect 514972 642284 514978 642318
rect 514932 642246 514978 642284
rect 514932 642212 514938 642246
rect 514972 642212 514978 642246
rect 514932 642174 514978 642212
rect 514932 642149 514938 642174
rect 514514 642143 514529 642149
rect 514465 642091 514471 642143
rect 514523 642091 514529 642143
rect 514465 642079 514480 642091
rect 514514 642079 514529 642091
rect 514465 642027 514471 642079
rect 514523 642027 514529 642079
rect 514465 642015 514480 642027
rect 514514 642015 514529 642027
rect 514465 641963 514471 642015
rect 514523 641963 514529 642015
rect 514465 641958 514529 641963
rect 514465 641957 514480 641958
rect 514056 641924 514062 641957
rect 514016 641886 514062 641924
rect 514016 641852 514022 641886
rect 514056 641852 514062 641886
rect 514016 641814 514062 641852
rect 514016 641780 514022 641814
rect 514056 641780 514062 641814
rect 514016 641742 514062 641780
rect 514016 641708 514022 641742
rect 514056 641708 514062 641742
rect 513100 641636 513106 641670
rect 513140 641636 513146 641670
rect 513100 641598 513146 641636
rect 513100 641564 513106 641598
rect 513140 641564 513146 641598
rect 513100 641526 513146 641564
rect 513100 641492 513106 641526
rect 513140 641492 513146 641526
rect 513549 641678 513613 641684
rect 513549 641626 513555 641678
rect 513607 641626 513613 641678
rect 513549 641614 513613 641626
rect 513549 641562 513555 641614
rect 513607 641562 513613 641614
rect 513549 641550 513613 641562
rect 513549 641498 513555 641550
rect 513607 641498 513613 641550
rect 513549 641492 513564 641498
rect 513598 641492 513613 641498
rect 514016 641670 514062 641708
rect 514016 641636 514022 641670
rect 514056 641636 514062 641670
rect 514016 641598 514062 641636
rect 514016 641564 514022 641598
rect 514056 641564 514062 641598
rect 514016 641526 514062 641564
rect 514016 641492 514022 641526
rect 514056 641492 514062 641526
rect 508520 641454 508566 641492
rect 508520 641420 508526 641454
rect 508560 641420 508566 641454
rect 508520 641405 508566 641420
rect 508978 641454 509024 641492
rect 508978 641420 508984 641454
rect 509018 641420 509024 641454
rect 508978 641405 509024 641420
rect 509436 641454 509482 641492
rect 509436 641420 509442 641454
rect 509476 641420 509482 641454
rect 509436 641405 509482 641420
rect 509894 641454 509940 641492
rect 509894 641420 509900 641454
rect 509934 641420 509940 641454
rect 509894 641405 509940 641420
rect 510352 641454 510398 641492
rect 510352 641420 510358 641454
rect 510392 641420 510398 641454
rect 510352 641405 510398 641420
rect 510810 641454 510856 641492
rect 510810 641420 510816 641454
rect 510850 641420 510856 641454
rect 510810 641405 510856 641420
rect 511268 641454 511314 641492
rect 511268 641420 511274 641454
rect 511308 641420 511314 641454
rect 511268 641405 511314 641420
rect 511726 641454 511772 641492
rect 511726 641420 511732 641454
rect 511766 641420 511772 641454
rect 511726 641405 511772 641420
rect 512184 641454 512230 641492
rect 512184 641420 512190 641454
rect 512224 641420 512230 641454
rect 512184 641405 512230 641420
rect 512642 641454 512688 641492
rect 512642 641420 512648 641454
rect 512682 641420 512688 641454
rect 512642 641405 512688 641420
rect 513100 641454 513146 641492
rect 513100 641420 513106 641454
rect 513140 641420 513146 641454
rect 513100 641405 513146 641420
rect 513558 641454 513604 641492
rect 513558 641420 513564 641454
rect 513598 641420 513604 641454
rect 513558 641405 513604 641420
rect 514016 641454 514062 641492
rect 514016 641420 514022 641454
rect 514056 641420 514062 641454
rect 514016 641405 514062 641420
rect 514474 641924 514480 641957
rect 514514 641957 514529 641958
rect 514923 642143 514938 642149
rect 514972 642149 514978 642174
rect 515390 642390 515436 642405
rect 515390 642356 515396 642390
rect 515430 642356 515436 642390
rect 515390 642318 515436 642356
rect 515390 642284 515396 642318
rect 515430 642284 515436 642318
rect 515390 642246 515436 642284
rect 515766 642390 515812 642405
rect 515766 642356 515772 642390
rect 515806 642356 515812 642390
rect 515766 642318 515812 642356
rect 515766 642284 515772 642318
rect 515806 642284 515812 642318
rect 515766 642249 515812 642284
rect 516224 642390 516270 642405
rect 516224 642356 516230 642390
rect 516264 642356 516270 642390
rect 516224 642318 516270 642356
rect 516224 642284 516230 642318
rect 516264 642284 516270 642318
rect 515390 642212 515396 642246
rect 515430 642212 515436 642246
rect 515390 642174 515436 642212
rect 515390 642149 515396 642174
rect 514972 642143 514987 642149
rect 514923 642091 514929 642143
rect 514981 642091 514987 642143
rect 514923 642079 514938 642091
rect 514972 642079 514987 642091
rect 514923 642027 514929 642079
rect 514981 642027 514987 642079
rect 514923 642015 514938 642027
rect 514972 642015 514987 642027
rect 514923 641963 514929 642015
rect 514981 641963 514987 642015
rect 514923 641958 514987 641963
rect 514923 641957 514938 641958
rect 514514 641924 514520 641957
rect 514474 641886 514520 641924
rect 514474 641852 514480 641886
rect 514514 641852 514520 641886
rect 514474 641814 514520 641852
rect 514474 641780 514480 641814
rect 514514 641780 514520 641814
rect 514474 641742 514520 641780
rect 514474 641708 514480 641742
rect 514514 641708 514520 641742
rect 514474 641670 514520 641708
rect 514474 641636 514480 641670
rect 514514 641636 514520 641670
rect 514474 641598 514520 641636
rect 514474 641564 514480 641598
rect 514514 641564 514520 641598
rect 514474 641526 514520 641564
rect 514474 641492 514480 641526
rect 514514 641492 514520 641526
rect 514474 641454 514520 641492
rect 514474 641420 514480 641454
rect 514514 641420 514520 641454
rect 514474 641405 514520 641420
rect 514932 641924 514938 641957
rect 514972 641957 514987 641958
rect 515381 642143 515396 642149
rect 515430 642149 515436 642174
rect 515757 642246 515821 642249
rect 515757 642243 515772 642246
rect 515806 642243 515821 642246
rect 515757 642191 515763 642243
rect 515815 642191 515821 642243
rect 515757 642179 515821 642191
rect 515572 642149 515630 642154
rect 515430 642143 515445 642149
rect 515381 642091 515387 642143
rect 515439 642091 515445 642143
rect 515381 642079 515396 642091
rect 515430 642079 515445 642091
rect 515381 642027 515387 642079
rect 515439 642027 515445 642079
rect 515381 642015 515396 642027
rect 515430 642015 515445 642027
rect 515381 641963 515387 642015
rect 515439 641963 515445 642015
rect 515381 641958 515445 641963
rect 515381 641957 515396 641958
rect 514972 641924 514978 641957
rect 514932 641886 514978 641924
rect 514932 641852 514938 641886
rect 514972 641852 514978 641886
rect 514932 641814 514978 641852
rect 514932 641780 514938 641814
rect 514972 641780 514978 641814
rect 514932 641742 514978 641780
rect 514932 641708 514938 641742
rect 514972 641708 514978 641742
rect 514932 641670 514978 641708
rect 514932 641636 514938 641670
rect 514972 641636 514978 641670
rect 514932 641598 514978 641636
rect 514932 641564 514938 641598
rect 514972 641564 514978 641598
rect 514932 641526 514978 641564
rect 514932 641492 514938 641526
rect 514972 641492 514978 641526
rect 514932 641454 514978 641492
rect 514932 641420 514938 641454
rect 514972 641420 514978 641454
rect 514932 641405 514978 641420
rect 515390 641924 515396 641957
rect 515430 641957 515445 641958
rect 515569 642143 515633 642149
rect 515569 642091 515575 642143
rect 515627 642091 515633 642143
rect 515569 642079 515633 642091
rect 515569 642027 515575 642079
rect 515627 642027 515633 642079
rect 515569 642015 515633 642027
rect 515569 641963 515575 642015
rect 515627 641963 515633 642015
rect 515569 641957 515633 641963
rect 515757 642127 515763 642179
rect 515815 642127 515821 642179
rect 515757 642115 515821 642127
rect 515757 642063 515763 642115
rect 515815 642063 515821 642115
rect 515757 642051 515821 642063
rect 515757 641999 515763 642051
rect 515815 641999 515821 642051
rect 515757 641996 515772 641999
rect 515806 641996 515821 641999
rect 515757 641987 515821 641996
rect 515430 641924 515436 641957
rect 515572 641952 515630 641957
rect 515390 641886 515436 641924
rect 515390 641852 515396 641886
rect 515430 641852 515436 641886
rect 515757 641935 515763 641987
rect 515815 641935 515821 641987
rect 515757 641924 515772 641935
rect 515806 641924 515821 641935
rect 515757 641923 515821 641924
rect 515757 641871 515763 641923
rect 515815 641871 515821 641923
rect 515757 641865 515772 641871
rect 515390 641814 515436 641852
rect 515390 641780 515396 641814
rect 515430 641780 515436 641814
rect 515390 641742 515436 641780
rect 515390 641708 515396 641742
rect 515430 641708 515436 641742
rect 515390 641670 515436 641708
rect 515390 641636 515396 641670
rect 515430 641636 515436 641670
rect 515390 641598 515436 641636
rect 515390 641564 515396 641598
rect 515430 641564 515436 641598
rect 515390 641526 515436 641564
rect 515390 641492 515396 641526
rect 515430 641492 515436 641526
rect 515390 641454 515436 641492
rect 515390 641420 515396 641454
rect 515430 641420 515436 641454
rect 515390 641405 515436 641420
rect 515766 641852 515772 641865
rect 515806 641865 515821 641871
rect 516224 642246 516270 642284
rect 516682 642390 516728 642405
rect 516682 642356 516688 642390
rect 516722 642356 516728 642390
rect 516682 642318 516728 642356
rect 516682 642284 516688 642318
rect 516722 642284 516728 642318
rect 516682 642249 516728 642284
rect 516224 642212 516230 642246
rect 516264 642212 516270 642246
rect 516224 642174 516270 642212
rect 516224 642140 516230 642174
rect 516264 642140 516270 642174
rect 516224 642102 516270 642140
rect 516224 642068 516230 642102
rect 516264 642068 516270 642102
rect 516224 642030 516270 642068
rect 516224 641996 516230 642030
rect 516264 641996 516270 642030
rect 516224 641958 516270 641996
rect 516224 641924 516230 641958
rect 516264 641924 516270 641958
rect 516224 641886 516270 641924
rect 515806 641852 515812 641865
rect 515766 641814 515812 641852
rect 515766 641780 515772 641814
rect 515806 641780 515812 641814
rect 516224 641852 516230 641886
rect 516264 641852 516270 641886
rect 516673 642246 516737 642249
rect 516673 642243 516688 642246
rect 516722 642243 516737 642246
rect 516673 642191 516679 642243
rect 516731 642191 516737 642243
rect 516673 642179 516737 642191
rect 516673 642127 516679 642179
rect 516731 642127 516737 642179
rect 516673 642115 516737 642127
rect 516673 642063 516679 642115
rect 516731 642063 516737 642115
rect 516673 642051 516737 642063
rect 516673 641999 516679 642051
rect 516731 641999 516737 642051
rect 516673 641996 516688 641999
rect 516722 641996 516737 641999
rect 516673 641987 516737 641996
rect 516673 641935 516679 641987
rect 516731 641935 516737 641987
rect 516673 641924 516688 641935
rect 516722 641924 516737 641935
rect 516673 641923 516737 641924
rect 516673 641871 516679 641923
rect 516731 641871 516737 641923
rect 516673 641865 516688 641871
rect 516224 641814 516270 641852
rect 516224 641797 516230 641814
rect 515766 641742 515812 641780
rect 515766 641708 515772 641742
rect 515806 641708 515812 641742
rect 515766 641670 515812 641708
rect 515766 641636 515772 641670
rect 515806 641636 515812 641670
rect 515766 641598 515812 641636
rect 515766 641564 515772 641598
rect 515806 641564 515812 641598
rect 515766 641526 515812 641564
rect 515766 641492 515772 641526
rect 515806 641492 515812 641526
rect 515766 641454 515812 641492
rect 516215 641791 516230 641797
rect 516264 641797 516270 641814
rect 516682 641852 516688 641865
rect 516722 641865 516737 641871
rect 516722 641852 516728 641865
rect 516682 641814 516728 641852
rect 516264 641791 516279 641797
rect 516215 641739 516221 641791
rect 516273 641739 516279 641791
rect 516215 641727 516230 641739
rect 516264 641727 516279 641739
rect 516215 641675 516221 641727
rect 516273 641675 516279 641727
rect 516215 641670 516279 641675
rect 516215 641663 516230 641670
rect 516264 641663 516279 641670
rect 516215 641611 516221 641663
rect 516273 641611 516279 641663
rect 516215 641599 516279 641611
rect 516215 641547 516221 641599
rect 516273 641547 516279 641599
rect 516215 641535 516279 641547
rect 516215 641483 516221 641535
rect 516273 641483 516279 641535
rect 516215 641477 516279 641483
rect 516682 641780 516688 641814
rect 516722 641780 516728 641814
rect 516682 641742 516728 641780
rect 516682 641708 516688 641742
rect 516722 641708 516728 641742
rect 516682 641670 516728 641708
rect 516682 641636 516688 641670
rect 516722 641636 516728 641670
rect 516682 641598 516728 641636
rect 516682 641564 516688 641598
rect 516722 641564 516728 641598
rect 516682 641526 516728 641564
rect 516682 641492 516688 641526
rect 516722 641492 516728 641526
rect 515766 641420 515772 641454
rect 515806 641420 515812 641454
rect 515766 641405 515812 641420
rect 516224 641454 516270 641477
rect 516224 641420 516230 641454
rect 516264 641420 516270 641454
rect 516224 641405 516270 641420
rect 516682 641454 516728 641492
rect 516682 641420 516688 641454
rect 516722 641420 516728 641454
rect 516682 641405 516728 641420
rect 508118 641315 508968 641321
rect 508118 641281 508153 641315
rect 508187 641281 508225 641315
rect 508259 641281 508297 641315
rect 508331 641281 508369 641315
rect 508403 641281 508441 641315
rect 508475 641281 508611 641315
rect 508645 641281 508683 641315
rect 508717 641281 508755 641315
rect 508789 641281 508827 641315
rect 508861 641281 508899 641315
rect 508933 641281 508968 641315
rect 508118 641275 508968 641281
rect 509034 641315 510800 641321
rect 509034 641281 509069 641315
rect 509103 641281 509141 641315
rect 509175 641281 509213 641315
rect 509247 641281 509285 641315
rect 509319 641281 509357 641315
rect 509391 641281 509527 641315
rect 509561 641281 509599 641315
rect 509633 641281 509671 641315
rect 509705 641281 509743 641315
rect 509777 641281 509815 641315
rect 509849 641281 509985 641315
rect 510019 641281 510057 641315
rect 510091 641281 510129 641315
rect 510163 641281 510201 641315
rect 510235 641281 510273 641315
rect 510307 641281 510443 641315
rect 510477 641281 510515 641315
rect 510549 641281 510587 641315
rect 510621 641281 510659 641315
rect 510693 641281 510731 641315
rect 510765 641281 510800 641315
rect 509034 641275 510800 641281
rect 510866 641315 512632 641321
rect 510866 641281 510901 641315
rect 510935 641281 510973 641315
rect 511007 641281 511045 641315
rect 511079 641281 511117 641315
rect 511151 641281 511189 641315
rect 511223 641281 511359 641315
rect 511393 641281 511431 641315
rect 511465 641281 511503 641315
rect 511537 641281 511575 641315
rect 511609 641281 511647 641315
rect 511681 641281 511817 641315
rect 511851 641281 511889 641315
rect 511923 641281 511961 641315
rect 511995 641281 512033 641315
rect 512067 641281 512105 641315
rect 512139 641281 512275 641315
rect 512309 641281 512347 641315
rect 512381 641281 512419 641315
rect 512453 641281 512491 641315
rect 512525 641281 512563 641315
rect 512597 641281 512632 641315
rect 510866 641275 512632 641281
rect 512698 641315 514464 641321
rect 512698 641281 512733 641315
rect 512767 641281 512805 641315
rect 512839 641281 512877 641315
rect 512911 641281 512949 641315
rect 512983 641281 513021 641315
rect 513055 641281 513191 641315
rect 513225 641281 513263 641315
rect 513297 641281 513335 641315
rect 513369 641281 513407 641315
rect 513441 641281 513479 641315
rect 513513 641281 513649 641315
rect 513683 641281 513721 641315
rect 513755 641281 513793 641315
rect 513827 641281 513865 641315
rect 513899 641281 513937 641315
rect 513971 641281 514107 641315
rect 514141 641281 514179 641315
rect 514213 641281 514251 641315
rect 514285 641281 514323 641315
rect 514357 641281 514395 641315
rect 514429 641281 514464 641315
rect 512698 641275 514464 641281
rect 514530 641315 515380 641321
rect 514530 641281 514565 641315
rect 514599 641281 514637 641315
rect 514671 641281 514709 641315
rect 514743 641281 514781 641315
rect 514815 641281 514853 641315
rect 514887 641281 515023 641315
rect 515057 641281 515095 641315
rect 515129 641281 515167 641315
rect 515201 641281 515239 641315
rect 515273 641281 515311 641315
rect 515345 641281 515380 641315
rect 514530 641275 515380 641281
rect 508062 641228 508108 641243
rect 508062 641194 508068 641228
rect 508102 641194 508108 641228
rect 508062 641156 508108 641194
rect 508062 641122 508068 641156
rect 508102 641122 508108 641156
rect 508062 641084 508108 641122
rect 508062 641050 508068 641084
rect 508102 641050 508108 641084
rect 508062 641012 508108 641050
rect 508062 640978 508068 641012
rect 508102 640978 508108 641012
rect 508062 640940 508108 640978
rect 508062 640906 508068 640940
rect 508102 640906 508108 640940
rect 508062 640868 508108 640906
rect 508062 640834 508068 640868
rect 508102 640834 508108 640868
rect 508062 640796 508108 640834
rect 508062 640762 508068 640796
rect 508102 640762 508108 640796
rect 508062 640724 508108 640762
rect 508062 640690 508068 640724
rect 508102 640690 508108 640724
rect 508062 640652 508108 640690
rect 508062 640618 508068 640652
rect 508102 640618 508108 640652
rect 508062 640580 508108 640618
rect 508062 640546 508068 640580
rect 508102 640546 508108 640580
rect 507867 640509 507925 640514
rect 508062 640509 508108 640546
rect 508520 641228 508566 641275
rect 508520 641194 508526 641228
rect 508560 641194 508566 641228
rect 508520 641156 508566 641194
rect 508520 641122 508526 641156
rect 508560 641122 508566 641156
rect 508520 641084 508566 641122
rect 508520 641050 508526 641084
rect 508560 641050 508566 641084
rect 508520 641012 508566 641050
rect 508520 640978 508526 641012
rect 508560 640978 508566 641012
rect 508520 640940 508566 640978
rect 508520 640906 508526 640940
rect 508560 640906 508566 640940
rect 508520 640868 508566 640906
rect 508520 640834 508526 640868
rect 508560 640834 508566 640868
rect 508520 640796 508566 640834
rect 508520 640762 508526 640796
rect 508560 640762 508566 640796
rect 508520 640724 508566 640762
rect 508520 640690 508526 640724
rect 508560 640690 508566 640724
rect 508520 640652 508566 640690
rect 508520 640618 508526 640652
rect 508560 640618 508566 640652
rect 508520 640580 508566 640618
rect 508520 640546 508526 640580
rect 508560 640546 508566 640580
rect 508520 640509 508566 640546
rect 508978 641228 509024 641243
rect 508978 641194 508984 641228
rect 509018 641194 509024 641228
rect 509436 641228 509482 641243
rect 509436 641194 509442 641228
rect 509476 641194 509482 641228
rect 509894 641228 509940 641243
rect 509894 641194 509900 641228
rect 509934 641194 509940 641228
rect 510352 641228 510398 641275
rect 510352 641194 510358 641228
rect 510392 641194 510398 641228
rect 510810 641228 510856 641243
rect 510810 641194 510816 641228
rect 510850 641194 510856 641228
rect 508978 641156 509024 641194
rect 508978 641122 508984 641156
rect 509018 641122 509024 641156
rect 508978 641084 509024 641122
rect 508978 641050 508984 641084
rect 509018 641050 509024 641084
rect 508978 641012 509024 641050
rect 508978 640978 508984 641012
rect 509018 640978 509024 641012
rect 509427 641188 509491 641194
rect 509427 641136 509433 641188
rect 509485 641136 509491 641188
rect 509427 641124 509442 641136
rect 509476 641124 509491 641136
rect 509427 641072 509433 641124
rect 509485 641072 509491 641124
rect 509427 641060 509442 641072
rect 509476 641060 509491 641072
rect 509427 641008 509433 641060
rect 509485 641008 509491 641060
rect 509427 641002 509442 641008
rect 508978 640940 509024 640978
rect 508978 640906 508984 640940
rect 509018 640906 509024 640940
rect 508978 640868 509024 640906
rect 508978 640834 508984 640868
rect 509018 640834 509024 640868
rect 508978 640796 509024 640834
rect 508978 640762 508984 640796
rect 509018 640762 509024 640796
rect 508978 640724 509024 640762
rect 508978 640690 508984 640724
rect 509018 640690 509024 640724
rect 508978 640652 509024 640690
rect 508978 640618 508984 640652
rect 509018 640618 509024 640652
rect 508978 640580 509024 640618
rect 508978 640546 508984 640580
rect 509018 640546 509024 640580
rect 508978 640509 509024 640546
rect 509436 640978 509442 641002
rect 509476 641002 509491 641008
rect 509894 641156 509940 641194
rect 509894 641122 509900 641156
rect 509934 641122 509940 641156
rect 509894 641084 509940 641122
rect 509894 641050 509900 641084
rect 509934 641050 509940 641084
rect 509894 641012 509940 641050
rect 509476 640978 509482 641002
rect 509436 640940 509482 640978
rect 509436 640906 509442 640940
rect 509476 640906 509482 640940
rect 509436 640868 509482 640906
rect 509436 640834 509442 640868
rect 509476 640834 509482 640868
rect 509436 640796 509482 640834
rect 509436 640762 509442 640796
rect 509476 640762 509482 640796
rect 509436 640724 509482 640762
rect 509436 640690 509442 640724
rect 509476 640690 509482 640724
rect 509436 640652 509482 640690
rect 509436 640618 509442 640652
rect 509476 640618 509482 640652
rect 509436 640580 509482 640618
rect 509436 640546 509442 640580
rect 509476 640546 509482 640580
rect 507864 640503 507928 640509
rect 507864 640451 507870 640503
rect 507922 640451 507928 640503
rect 507864 640439 507928 640451
rect 507864 640387 507870 640439
rect 507922 640387 507928 640439
rect 507864 640375 507928 640387
rect 507864 640323 507870 640375
rect 507922 640323 507928 640375
rect 507864 640317 507928 640323
rect 508053 640508 508117 640509
rect 508053 640503 508068 640508
rect 508102 640503 508117 640508
rect 508053 640451 508059 640503
rect 508111 640451 508117 640503
rect 508053 640439 508117 640451
rect 508053 640387 508059 640439
rect 508111 640387 508117 640439
rect 508053 640375 508117 640387
rect 508053 640323 508059 640375
rect 508111 640323 508117 640375
rect 508053 640317 508117 640323
rect 508511 640508 508575 640509
rect 508511 640503 508526 640508
rect 508560 640503 508575 640508
rect 508511 640451 508517 640503
rect 508569 640451 508575 640503
rect 508511 640439 508575 640451
rect 508511 640387 508517 640439
rect 508569 640387 508575 640439
rect 508511 640375 508575 640387
rect 508511 640323 508517 640375
rect 508569 640323 508575 640375
rect 508511 640317 508575 640323
rect 508969 640508 509033 640509
rect 508969 640503 508984 640508
rect 509018 640503 509033 640508
rect 508969 640451 508975 640503
rect 509027 640451 509033 640503
rect 508969 640439 509033 640451
rect 508969 640387 508975 640439
rect 509027 640387 509033 640439
rect 508969 640375 509033 640387
rect 508969 640323 508975 640375
rect 509027 640323 509033 640375
rect 508969 640317 509033 640323
rect 509436 640508 509482 640546
rect 509894 640978 509900 641012
rect 509934 640978 509940 641012
rect 510343 641188 510407 641194
rect 510343 641136 510349 641188
rect 510401 641136 510407 641188
rect 510343 641124 510358 641136
rect 510392 641124 510407 641136
rect 510343 641072 510349 641124
rect 510401 641072 510407 641124
rect 510343 641060 510358 641072
rect 510392 641060 510407 641072
rect 510343 641008 510349 641060
rect 510401 641008 510407 641060
rect 510343 641002 510358 641008
rect 509894 640940 509940 640978
rect 509894 640906 509900 640940
rect 509934 640906 509940 640940
rect 509894 640868 509940 640906
rect 509894 640834 509900 640868
rect 509934 640834 509940 640868
rect 509894 640796 509940 640834
rect 509894 640762 509900 640796
rect 509934 640762 509940 640796
rect 509894 640724 509940 640762
rect 509894 640690 509900 640724
rect 509934 640690 509940 640724
rect 509894 640652 509940 640690
rect 509894 640618 509900 640652
rect 509934 640618 509940 640652
rect 509894 640580 509940 640618
rect 509894 640546 509900 640580
rect 509934 640546 509940 640580
rect 509894 640509 509940 640546
rect 510352 640978 510358 641002
rect 510392 641002 510407 641008
rect 510810 641156 510856 641194
rect 510810 641122 510816 641156
rect 510850 641122 510856 641156
rect 510810 641084 510856 641122
rect 510810 641050 510816 641084
rect 510850 641050 510856 641084
rect 510810 641012 510856 641050
rect 510392 640978 510398 641002
rect 510352 640940 510398 640978
rect 510352 640906 510358 640940
rect 510392 640906 510398 640940
rect 510352 640868 510398 640906
rect 510352 640834 510358 640868
rect 510392 640834 510398 640868
rect 510352 640796 510398 640834
rect 510352 640762 510358 640796
rect 510392 640762 510398 640796
rect 510352 640724 510398 640762
rect 510352 640690 510358 640724
rect 510392 640690 510398 640724
rect 510352 640652 510398 640690
rect 510352 640618 510358 640652
rect 510392 640618 510398 640652
rect 510352 640580 510398 640618
rect 510352 640546 510358 640580
rect 510392 640546 510398 640580
rect 509436 640474 509442 640508
rect 509476 640474 509482 640508
rect 509436 640436 509482 640474
rect 509436 640402 509442 640436
rect 509476 640402 509482 640436
rect 509436 640364 509482 640402
rect 509436 640330 509442 640364
rect 509476 640330 509482 640364
rect 507867 640312 507925 640317
rect 508062 640292 508108 640317
rect 508062 640258 508068 640292
rect 508102 640258 508108 640292
rect 508062 640243 508108 640258
rect 508520 640292 508566 640317
rect 508520 640258 508526 640292
rect 508560 640258 508566 640292
rect 508520 640243 508566 640258
rect 508978 640292 509024 640317
rect 508978 640258 508984 640292
rect 509018 640258 509024 640292
rect 508978 640243 509024 640258
rect 509436 640292 509482 640330
rect 509885 640508 509949 640509
rect 509885 640503 509900 640508
rect 509934 640503 509949 640508
rect 509885 640451 509891 640503
rect 509943 640451 509949 640503
rect 509885 640439 509949 640451
rect 509885 640387 509891 640439
rect 509943 640387 509949 640439
rect 509885 640375 509949 640387
rect 509885 640323 509891 640375
rect 509943 640323 509949 640375
rect 509885 640317 509949 640323
rect 510352 640508 510398 640546
rect 510810 640978 510816 641012
rect 510850 640978 510856 641012
rect 510810 640940 510856 640978
rect 510810 640906 510816 640940
rect 510850 640906 510856 640940
rect 510810 640868 510856 640906
rect 510810 640834 510816 640868
rect 510850 640834 510856 640868
rect 511268 641228 511314 641275
rect 511268 641194 511274 641228
rect 511308 641194 511314 641228
rect 511268 641156 511314 641194
rect 511268 641122 511274 641156
rect 511308 641122 511314 641156
rect 511268 641084 511314 641122
rect 511268 641050 511274 641084
rect 511308 641050 511314 641084
rect 511268 641012 511314 641050
rect 511268 640978 511274 641012
rect 511308 640978 511314 641012
rect 511268 640940 511314 640978
rect 511268 640906 511274 640940
rect 511308 640906 511314 640940
rect 511268 640868 511314 640906
rect 511268 640840 511274 640868
rect 510810 640796 510856 640834
rect 510810 640762 510816 640796
rect 510850 640762 510856 640796
rect 510810 640724 510856 640762
rect 510810 640690 510816 640724
rect 510850 640690 510856 640724
rect 510810 640652 510856 640690
rect 510810 640618 510816 640652
rect 510850 640618 510856 640652
rect 511259 640834 511274 640840
rect 511308 640840 511314 640868
rect 511726 641228 511772 641243
rect 511726 641194 511732 641228
rect 511766 641194 511772 641228
rect 511726 641156 511772 641194
rect 511726 641122 511732 641156
rect 511766 641122 511772 641156
rect 511726 641084 511772 641122
rect 511726 641050 511732 641084
rect 511766 641050 511772 641084
rect 511726 641012 511772 641050
rect 511726 640978 511732 641012
rect 511766 640978 511772 641012
rect 511726 640940 511772 640978
rect 511726 640906 511732 640940
rect 511766 640906 511772 640940
rect 511726 640868 511772 640906
rect 511308 640834 511323 640840
rect 511259 640782 511265 640834
rect 511317 640782 511323 640834
rect 511259 640770 511274 640782
rect 511308 640770 511323 640782
rect 511259 640718 511265 640770
rect 511317 640718 511323 640770
rect 511259 640706 511274 640718
rect 511308 640706 511323 640718
rect 511259 640654 511265 640706
rect 511317 640654 511323 640706
rect 511259 640652 511323 640654
rect 511259 640648 511274 640652
rect 510810 640580 510856 640618
rect 510810 640546 510816 640580
rect 510850 640546 510856 640580
rect 510810 640509 510856 640546
rect 511268 640618 511274 640648
rect 511308 640648 511323 640652
rect 511726 640834 511732 640868
rect 511766 640834 511772 640868
rect 512184 641228 512230 641243
rect 512184 641194 512190 641228
rect 512224 641194 512230 641228
rect 512184 641156 512230 641194
rect 512184 641122 512190 641156
rect 512224 641122 512230 641156
rect 512184 641084 512230 641122
rect 512184 641050 512190 641084
rect 512224 641050 512230 641084
rect 512184 641012 512230 641050
rect 512184 640978 512190 641012
rect 512224 640978 512230 641012
rect 512184 640940 512230 640978
rect 512184 640906 512190 640940
rect 512224 640906 512230 640940
rect 512184 640868 512230 640906
rect 512184 640840 512190 640868
rect 511726 640796 511772 640834
rect 511726 640762 511732 640796
rect 511766 640762 511772 640796
rect 511726 640724 511772 640762
rect 511726 640690 511732 640724
rect 511766 640690 511772 640724
rect 511726 640652 511772 640690
rect 511308 640618 511314 640648
rect 511268 640580 511314 640618
rect 511268 640546 511274 640580
rect 511308 640546 511314 640580
rect 510352 640474 510358 640508
rect 510392 640474 510398 640508
rect 510352 640436 510398 640474
rect 510352 640402 510358 640436
rect 510392 640402 510398 640436
rect 510352 640364 510398 640402
rect 510352 640330 510358 640364
rect 510392 640330 510398 640364
rect 509436 640258 509442 640292
rect 509476 640258 509482 640292
rect 509436 640243 509482 640258
rect 509894 640292 509940 640317
rect 509894 640258 509900 640292
rect 509934 640258 509940 640292
rect 509894 640243 509940 640258
rect 510352 640292 510398 640330
rect 510801 640508 510865 640509
rect 510801 640503 510816 640508
rect 510850 640503 510865 640508
rect 510801 640451 510807 640503
rect 510859 640451 510865 640503
rect 510801 640439 510865 640451
rect 510801 640387 510807 640439
rect 510859 640387 510865 640439
rect 510801 640375 510865 640387
rect 510801 640323 510807 640375
rect 510859 640323 510865 640375
rect 510801 640317 510865 640323
rect 511268 640508 511314 640546
rect 511726 640618 511732 640652
rect 511766 640618 511772 640652
rect 512175 640834 512190 640840
rect 512224 640840 512230 640868
rect 512642 641228 512688 641243
rect 512642 641194 512648 641228
rect 512682 641194 512688 641228
rect 513100 641228 513146 641275
rect 513100 641194 513106 641228
rect 513140 641194 513146 641228
rect 513558 641228 513604 641243
rect 513558 641194 513564 641228
rect 513598 641194 513604 641228
rect 514016 641228 514062 641243
rect 514016 641194 514022 641228
rect 514056 641194 514062 641228
rect 514474 641228 514520 641243
rect 514474 641194 514480 641228
rect 514514 641194 514520 641228
rect 512642 641156 512688 641194
rect 512642 641122 512648 641156
rect 512682 641122 512688 641156
rect 512642 641084 512688 641122
rect 512642 641050 512648 641084
rect 512682 641050 512688 641084
rect 512642 641012 512688 641050
rect 512642 640978 512648 641012
rect 512682 640978 512688 641012
rect 513091 641188 513155 641194
rect 513091 641136 513097 641188
rect 513149 641136 513155 641188
rect 513091 641124 513106 641136
rect 513140 641124 513155 641136
rect 513091 641072 513097 641124
rect 513149 641072 513155 641124
rect 513091 641060 513106 641072
rect 513140 641060 513155 641072
rect 513091 641008 513097 641060
rect 513149 641008 513155 641060
rect 513091 641002 513106 641008
rect 512642 640940 512688 640978
rect 512642 640906 512648 640940
rect 512682 640906 512688 640940
rect 512642 640868 512688 640906
rect 512224 640834 512239 640840
rect 512175 640782 512181 640834
rect 512233 640782 512239 640834
rect 512175 640770 512190 640782
rect 512224 640770 512239 640782
rect 512175 640718 512181 640770
rect 512233 640718 512239 640770
rect 512175 640706 512190 640718
rect 512224 640706 512239 640718
rect 512175 640654 512181 640706
rect 512233 640654 512239 640706
rect 512175 640652 512239 640654
rect 512175 640648 512190 640652
rect 511726 640580 511772 640618
rect 511726 640546 511732 640580
rect 511766 640546 511772 640580
rect 511726 640509 511772 640546
rect 512184 640618 512190 640648
rect 512224 640648 512239 640652
rect 512642 640834 512648 640868
rect 512682 640834 512688 640868
rect 512642 640796 512688 640834
rect 512642 640762 512648 640796
rect 512682 640762 512688 640796
rect 512642 640724 512688 640762
rect 512642 640690 512648 640724
rect 512682 640690 512688 640724
rect 512642 640652 512688 640690
rect 512224 640618 512230 640648
rect 512184 640580 512230 640618
rect 512184 640546 512190 640580
rect 512224 640546 512230 640580
rect 511268 640474 511274 640508
rect 511308 640474 511314 640508
rect 511268 640436 511314 640474
rect 511268 640402 511274 640436
rect 511308 640402 511314 640436
rect 511268 640364 511314 640402
rect 511268 640330 511274 640364
rect 511308 640330 511314 640364
rect 510352 640258 510358 640292
rect 510392 640258 510398 640292
rect 510352 640243 510398 640258
rect 510810 640292 510856 640317
rect 510810 640258 510816 640292
rect 510850 640258 510856 640292
rect 510810 640243 510856 640258
rect 511268 640292 511314 640330
rect 511717 640508 511781 640509
rect 511717 640503 511732 640508
rect 511766 640503 511781 640508
rect 511717 640451 511723 640503
rect 511775 640451 511781 640503
rect 511717 640439 511781 640451
rect 511717 640387 511723 640439
rect 511775 640387 511781 640439
rect 511717 640375 511781 640387
rect 511717 640323 511723 640375
rect 511775 640323 511781 640375
rect 511717 640317 511781 640323
rect 512184 640508 512230 640546
rect 512642 640618 512648 640652
rect 512682 640618 512688 640652
rect 512642 640580 512688 640618
rect 512642 640546 512648 640580
rect 512682 640546 512688 640580
rect 512642 640509 512688 640546
rect 513100 640978 513106 641002
rect 513140 641002 513155 641008
rect 513558 641156 513604 641194
rect 513558 641122 513564 641156
rect 513598 641122 513604 641156
rect 513558 641084 513604 641122
rect 513558 641050 513564 641084
rect 513598 641050 513604 641084
rect 513558 641012 513604 641050
rect 513140 640978 513146 641002
rect 513100 640940 513146 640978
rect 513100 640906 513106 640940
rect 513140 640906 513146 640940
rect 513100 640868 513146 640906
rect 513100 640834 513106 640868
rect 513140 640834 513146 640868
rect 513100 640796 513146 640834
rect 513100 640762 513106 640796
rect 513140 640762 513146 640796
rect 513100 640724 513146 640762
rect 513100 640690 513106 640724
rect 513140 640690 513146 640724
rect 513100 640652 513146 640690
rect 513100 640618 513106 640652
rect 513140 640618 513146 640652
rect 513100 640580 513146 640618
rect 513100 640546 513106 640580
rect 513140 640546 513146 640580
rect 512184 640474 512190 640508
rect 512224 640474 512230 640508
rect 512184 640436 512230 640474
rect 512184 640402 512190 640436
rect 512224 640402 512230 640436
rect 512184 640364 512230 640402
rect 512184 640330 512190 640364
rect 512224 640330 512230 640364
rect 511268 640258 511274 640292
rect 511308 640258 511314 640292
rect 511268 640243 511314 640258
rect 511726 640292 511772 640317
rect 511726 640258 511732 640292
rect 511766 640258 511772 640292
rect 511726 640243 511772 640258
rect 512184 640292 512230 640330
rect 512633 640508 512697 640509
rect 512633 640503 512648 640508
rect 512682 640503 512697 640508
rect 512633 640451 512639 640503
rect 512691 640451 512697 640503
rect 512633 640439 512697 640451
rect 512633 640387 512639 640439
rect 512691 640387 512697 640439
rect 512633 640375 512697 640387
rect 512633 640323 512639 640375
rect 512691 640323 512697 640375
rect 512633 640317 512697 640323
rect 513100 640508 513146 640546
rect 513558 640978 513564 641012
rect 513598 640978 513604 641012
rect 514007 641188 514071 641194
rect 514007 641136 514013 641188
rect 514065 641136 514071 641188
rect 514007 641124 514022 641136
rect 514056 641124 514071 641136
rect 514007 641072 514013 641124
rect 514065 641072 514071 641124
rect 514007 641060 514022 641072
rect 514056 641060 514071 641072
rect 514007 641008 514013 641060
rect 514065 641008 514071 641060
rect 514007 641002 514022 641008
rect 513558 640940 513604 640978
rect 513558 640906 513564 640940
rect 513598 640906 513604 640940
rect 513558 640868 513604 640906
rect 513558 640834 513564 640868
rect 513598 640834 513604 640868
rect 513558 640796 513604 640834
rect 513558 640762 513564 640796
rect 513598 640762 513604 640796
rect 513558 640724 513604 640762
rect 513558 640690 513564 640724
rect 513598 640690 513604 640724
rect 513558 640652 513604 640690
rect 513558 640618 513564 640652
rect 513598 640618 513604 640652
rect 513558 640580 513604 640618
rect 513558 640546 513564 640580
rect 513598 640546 513604 640580
rect 513558 640509 513604 640546
rect 514016 640978 514022 641002
rect 514056 641002 514071 641008
rect 514474 641156 514520 641194
rect 514474 641122 514480 641156
rect 514514 641122 514520 641156
rect 514474 641084 514520 641122
rect 514474 641050 514480 641084
rect 514514 641050 514520 641084
rect 514474 641012 514520 641050
rect 514056 640978 514062 641002
rect 514016 640940 514062 640978
rect 514016 640906 514022 640940
rect 514056 640906 514062 640940
rect 514016 640868 514062 640906
rect 514016 640834 514022 640868
rect 514056 640834 514062 640868
rect 514016 640796 514062 640834
rect 514016 640762 514022 640796
rect 514056 640762 514062 640796
rect 514016 640724 514062 640762
rect 514016 640690 514022 640724
rect 514056 640690 514062 640724
rect 514016 640652 514062 640690
rect 514016 640618 514022 640652
rect 514056 640618 514062 640652
rect 514016 640580 514062 640618
rect 514016 640546 514022 640580
rect 514056 640546 514062 640580
rect 513100 640474 513106 640508
rect 513140 640474 513146 640508
rect 513100 640436 513146 640474
rect 513100 640402 513106 640436
rect 513140 640402 513146 640436
rect 513100 640364 513146 640402
rect 513100 640330 513106 640364
rect 513140 640330 513146 640364
rect 512184 640258 512190 640292
rect 512224 640258 512230 640292
rect 512184 640243 512230 640258
rect 512642 640292 512688 640317
rect 512642 640258 512648 640292
rect 512682 640258 512688 640292
rect 512642 640243 512688 640258
rect 513100 640292 513146 640330
rect 513549 640508 513613 640509
rect 513549 640503 513564 640508
rect 513598 640503 513613 640508
rect 513549 640451 513555 640503
rect 513607 640451 513613 640503
rect 513549 640439 513613 640451
rect 513549 640387 513555 640439
rect 513607 640387 513613 640439
rect 513549 640375 513613 640387
rect 513549 640323 513555 640375
rect 513607 640323 513613 640375
rect 513549 640317 513613 640323
rect 514016 640508 514062 640546
rect 514474 640978 514480 641012
rect 514514 640978 514520 641012
rect 514474 640940 514520 640978
rect 514474 640906 514480 640940
rect 514514 640906 514520 640940
rect 514474 640868 514520 640906
rect 514474 640834 514480 640868
rect 514514 640834 514520 640868
rect 514474 640796 514520 640834
rect 514474 640762 514480 640796
rect 514514 640762 514520 640796
rect 514474 640724 514520 640762
rect 514474 640690 514480 640724
rect 514514 640690 514520 640724
rect 514474 640652 514520 640690
rect 514474 640618 514480 640652
rect 514514 640618 514520 640652
rect 514474 640580 514520 640618
rect 514474 640546 514480 640580
rect 514514 640546 514520 640580
rect 514474 640509 514520 640546
rect 514932 641228 514978 641275
rect 514932 641194 514938 641228
rect 514972 641194 514978 641228
rect 514932 641156 514978 641194
rect 514932 641122 514938 641156
rect 514972 641122 514978 641156
rect 514932 641084 514978 641122
rect 514932 641050 514938 641084
rect 514972 641050 514978 641084
rect 514932 641012 514978 641050
rect 514932 640978 514938 641012
rect 514972 640978 514978 641012
rect 514932 640940 514978 640978
rect 514932 640906 514938 640940
rect 514972 640906 514978 640940
rect 514932 640868 514978 640906
rect 514932 640834 514938 640868
rect 514972 640834 514978 640868
rect 514932 640796 514978 640834
rect 514932 640762 514938 640796
rect 514972 640762 514978 640796
rect 514932 640724 514978 640762
rect 514932 640690 514938 640724
rect 514972 640690 514978 640724
rect 514932 640652 514978 640690
rect 514932 640618 514938 640652
rect 514972 640618 514978 640652
rect 514932 640580 514978 640618
rect 514932 640546 514938 640580
rect 514972 640546 514978 640580
rect 514932 640509 514978 640546
rect 515390 641228 515436 641243
rect 515390 641194 515396 641228
rect 515430 641194 515436 641228
rect 515390 641156 515436 641194
rect 515390 641122 515396 641156
rect 515430 641122 515436 641156
rect 515390 641084 515436 641122
rect 515390 641050 515396 641084
rect 515430 641050 515436 641084
rect 515390 641012 515436 641050
rect 515390 640978 515396 641012
rect 515430 640978 515436 641012
rect 515390 640940 515436 640978
rect 515390 640906 515396 640940
rect 515430 640906 515436 640940
rect 515390 640868 515436 640906
rect 515390 640834 515396 640868
rect 515430 640834 515436 640868
rect 515390 640796 515436 640834
rect 515390 640762 515396 640796
rect 515430 640762 515436 640796
rect 515390 640724 515436 640762
rect 515390 640690 515396 640724
rect 515430 640690 515436 640724
rect 515390 640652 515436 640690
rect 515390 640618 515396 640652
rect 515430 640618 515436 640652
rect 515390 640580 515436 640618
rect 515390 640546 515396 640580
rect 515430 640546 515436 640580
rect 515390 640509 515436 640546
rect 514016 640474 514022 640508
rect 514056 640474 514062 640508
rect 514016 640436 514062 640474
rect 514016 640402 514022 640436
rect 514056 640402 514062 640436
rect 514016 640364 514062 640402
rect 514016 640330 514022 640364
rect 514056 640330 514062 640364
rect 513100 640258 513106 640292
rect 513140 640258 513146 640292
rect 513100 640243 513146 640258
rect 513558 640292 513604 640317
rect 513558 640258 513564 640292
rect 513598 640258 513604 640292
rect 513558 640243 513604 640258
rect 514016 640292 514062 640330
rect 514465 640508 514529 640509
rect 514465 640503 514480 640508
rect 514514 640503 514529 640508
rect 514465 640451 514471 640503
rect 514523 640451 514529 640503
rect 514465 640439 514529 640451
rect 514465 640387 514471 640439
rect 514523 640387 514529 640439
rect 514465 640375 514529 640387
rect 514465 640323 514471 640375
rect 514523 640323 514529 640375
rect 514465 640317 514529 640323
rect 514923 640508 514987 640509
rect 514923 640503 514938 640508
rect 514972 640503 514987 640508
rect 514923 640451 514929 640503
rect 514981 640451 514987 640503
rect 514923 640439 514987 640451
rect 514923 640387 514929 640439
rect 514981 640387 514987 640439
rect 514923 640375 514987 640387
rect 514923 640323 514929 640375
rect 514981 640323 514987 640375
rect 514923 640317 514987 640323
rect 515381 640508 515445 640509
rect 515381 640503 515396 640508
rect 515430 640503 515445 640508
rect 515381 640451 515387 640503
rect 515439 640451 515445 640503
rect 515381 640439 515445 640451
rect 515381 640387 515387 640439
rect 515439 640387 515445 640439
rect 515381 640375 515445 640387
rect 515381 640323 515387 640375
rect 515439 640323 515445 640375
rect 515381 640317 515445 640323
rect 515638 640503 516056 640514
rect 515638 640502 515661 640503
rect 516033 640502 516056 640503
rect 515638 640324 515650 640502
rect 516044 640324 516056 640502
rect 515638 640323 515661 640324
rect 516033 640323 516056 640324
rect 514016 640258 514022 640292
rect 514056 640258 514062 640292
rect 514016 640243 514062 640258
rect 514474 640292 514520 640317
rect 514474 640258 514480 640292
rect 514514 640258 514520 640292
rect 514474 640243 514520 640258
rect 514932 640292 514978 640317
rect 514932 640258 514938 640292
rect 514972 640258 514978 640292
rect 514932 640243 514978 640258
rect 515390 640292 515436 640317
rect 515638 640312 516056 640323
rect 515390 640258 515396 640292
rect 515430 640258 515436 640292
rect 515390 640243 515436 640258
<< via1 >>
rect 507870 645410 507922 645411
rect 507870 645376 507879 645410
rect 507879 645376 507913 645410
rect 507913 645376 507922 645410
rect 507870 645359 507922 645376
rect 507870 645338 507922 645347
rect 507870 645304 507879 645338
rect 507879 645304 507913 645338
rect 507913 645304 507922 645338
rect 507870 645295 507922 645304
rect 507870 645266 507922 645283
rect 507870 645232 507879 645266
rect 507879 645232 507913 645266
rect 507913 645232 507922 645266
rect 507870 645231 507922 645232
rect 508059 645382 508068 645411
rect 508068 645382 508102 645411
rect 508102 645382 508111 645411
rect 508059 645359 508111 645382
rect 508059 645344 508111 645347
rect 508059 645310 508068 645344
rect 508068 645310 508102 645344
rect 508102 645310 508111 645344
rect 508059 645295 508111 645310
rect 508059 645272 508111 645283
rect 508059 645238 508068 645272
rect 508068 645238 508102 645272
rect 508102 645238 508111 645272
rect 508059 645231 508111 645238
rect 508517 645382 508526 645411
rect 508526 645382 508560 645411
rect 508560 645382 508569 645411
rect 508517 645359 508569 645382
rect 508517 645344 508569 645347
rect 508517 645310 508526 645344
rect 508526 645310 508560 645344
rect 508560 645310 508569 645344
rect 508517 645295 508569 645310
rect 508517 645272 508569 645283
rect 508517 645238 508526 645272
rect 508526 645238 508560 645272
rect 508560 645238 508569 645272
rect 508517 645231 508569 645238
rect 508975 645382 508984 645411
rect 508984 645382 509018 645411
rect 509018 645382 509027 645411
rect 508975 645359 509027 645382
rect 508975 645344 509027 645347
rect 508975 645310 508984 645344
rect 508984 645310 509018 645344
rect 509018 645310 509027 645344
rect 508975 645295 509027 645310
rect 508975 645272 509027 645283
rect 508975 645238 508984 645272
rect 508984 645238 509018 645272
rect 509018 645238 509027 645272
rect 508975 645231 509027 645238
rect 509891 645382 509900 645411
rect 509900 645382 509934 645411
rect 509934 645382 509943 645411
rect 509891 645359 509943 645382
rect 509891 645344 509943 645347
rect 509891 645310 509900 645344
rect 509900 645310 509934 645344
rect 509934 645310 509943 645344
rect 509891 645295 509943 645310
rect 509891 645272 509943 645283
rect 509891 645238 509900 645272
rect 509900 645238 509934 645272
rect 509934 645238 509943 645272
rect 509891 645231 509943 645238
rect 509433 644768 509485 644776
rect 509433 644734 509442 644768
rect 509442 644734 509476 644768
rect 509476 644734 509485 644768
rect 509433 644724 509485 644734
rect 509433 644696 509485 644712
rect 509433 644662 509442 644696
rect 509442 644662 509476 644696
rect 509476 644662 509485 644696
rect 509433 644660 509485 644662
rect 509433 644624 509485 644648
rect 509433 644596 509442 644624
rect 509442 644596 509476 644624
rect 509476 644596 509485 644624
rect 510807 645382 510816 645411
rect 510816 645382 510850 645411
rect 510850 645382 510859 645411
rect 510807 645359 510859 645382
rect 510807 645344 510859 645347
rect 510807 645310 510816 645344
rect 510816 645310 510850 645344
rect 510850 645310 510859 645344
rect 510807 645295 510859 645310
rect 510807 645272 510859 645283
rect 510807 645238 510816 645272
rect 510816 645238 510850 645272
rect 510850 645238 510859 645272
rect 510807 645231 510859 645238
rect 511723 645382 511732 645411
rect 511732 645382 511766 645411
rect 511766 645382 511775 645411
rect 511723 645359 511775 645382
rect 511723 645344 511775 645347
rect 511723 645310 511732 645344
rect 511732 645310 511766 645344
rect 511766 645310 511775 645344
rect 511723 645295 511775 645310
rect 511723 645272 511775 645283
rect 511723 645238 511732 645272
rect 511732 645238 511766 645272
rect 511766 645238 511775 645272
rect 511723 645231 511775 645238
rect 512639 645382 512648 645411
rect 512648 645382 512682 645411
rect 512682 645382 512691 645411
rect 512639 645359 512691 645382
rect 512639 645344 512691 645347
rect 512639 645310 512648 645344
rect 512648 645310 512682 645344
rect 512682 645310 512691 645344
rect 512639 645295 512691 645310
rect 512639 645272 512691 645283
rect 512639 645238 512648 645272
rect 512648 645238 512682 645272
rect 512682 645238 512691 645272
rect 512639 645231 512691 645238
rect 511265 645056 511317 645088
rect 511265 645036 511274 645056
rect 511274 645036 511308 645056
rect 511308 645036 511317 645056
rect 511265 645022 511274 645024
rect 511274 645022 511308 645024
rect 511308 645022 511317 645024
rect 511265 644984 511317 645022
rect 511265 644972 511274 644984
rect 511274 644972 511308 644984
rect 511308 644972 511317 644984
rect 511265 644950 511274 644960
rect 511274 644950 511308 644960
rect 511308 644950 511317 644960
rect 511265 644912 511317 644950
rect 511265 644908 511274 644912
rect 511274 644908 511308 644912
rect 511308 644908 511317 644912
rect 510349 644768 510401 644776
rect 510349 644734 510358 644768
rect 510358 644734 510392 644768
rect 510392 644734 510401 644768
rect 510349 644724 510401 644734
rect 510349 644696 510401 644712
rect 510349 644662 510358 644696
rect 510358 644662 510392 644696
rect 510392 644662 510401 644696
rect 510349 644660 510401 644662
rect 510349 644624 510401 644648
rect 510349 644596 510358 644624
rect 510358 644596 510392 644624
rect 510392 644596 510401 644624
rect 512181 645056 512233 645088
rect 512181 645036 512190 645056
rect 512190 645036 512224 645056
rect 512224 645036 512233 645056
rect 512181 645022 512190 645024
rect 512190 645022 512224 645024
rect 512224 645022 512233 645024
rect 512181 644984 512233 645022
rect 512181 644972 512190 644984
rect 512190 644972 512224 644984
rect 512224 644972 512233 644984
rect 512181 644950 512190 644960
rect 512190 644950 512224 644960
rect 512224 644950 512233 644960
rect 512181 644912 512233 644950
rect 512181 644908 512190 644912
rect 512190 644908 512224 644912
rect 512224 644908 512233 644912
rect 513555 645382 513564 645411
rect 513564 645382 513598 645411
rect 513598 645382 513607 645411
rect 513555 645359 513607 645382
rect 513555 645344 513607 645347
rect 513555 645310 513564 645344
rect 513564 645310 513598 645344
rect 513598 645310 513607 645344
rect 513555 645295 513607 645310
rect 513555 645272 513607 645283
rect 513555 645238 513564 645272
rect 513564 645238 513598 645272
rect 513598 645238 513607 645272
rect 513555 645231 513607 645238
rect 513097 644768 513149 644776
rect 513097 644734 513106 644768
rect 513106 644734 513140 644768
rect 513140 644734 513149 644768
rect 513097 644724 513149 644734
rect 513097 644696 513149 644712
rect 513097 644662 513106 644696
rect 513106 644662 513140 644696
rect 513140 644662 513149 644696
rect 513097 644660 513149 644662
rect 513097 644624 513149 644648
rect 513097 644596 513106 644624
rect 513106 644596 513140 644624
rect 513140 644596 513149 644624
rect 514471 645382 514480 645411
rect 514480 645382 514514 645411
rect 514514 645382 514523 645411
rect 514471 645359 514523 645382
rect 514471 645344 514523 645347
rect 514471 645310 514480 645344
rect 514480 645310 514514 645344
rect 514514 645310 514523 645344
rect 514471 645295 514523 645310
rect 514471 645272 514523 645283
rect 514471 645238 514480 645272
rect 514480 645238 514514 645272
rect 514514 645238 514523 645272
rect 514471 645231 514523 645238
rect 514929 645382 514938 645411
rect 514938 645382 514972 645411
rect 514972 645382 514981 645411
rect 514929 645359 514981 645382
rect 514929 645344 514981 645347
rect 514929 645310 514938 645344
rect 514938 645310 514972 645344
rect 514972 645310 514981 645344
rect 514929 645295 514981 645310
rect 514929 645272 514981 645283
rect 514929 645238 514938 645272
rect 514938 645238 514972 645272
rect 514972 645238 514981 645272
rect 514929 645231 514981 645238
rect 515387 645382 515396 645411
rect 515396 645382 515430 645411
rect 515430 645382 515439 645411
rect 515387 645359 515439 645382
rect 515387 645344 515439 645347
rect 515387 645310 515396 645344
rect 515396 645310 515430 645344
rect 515430 645310 515439 645344
rect 515387 645295 515439 645310
rect 515387 645272 515439 645283
rect 515387 645238 515396 645272
rect 515396 645238 515430 645272
rect 515430 645238 515439 645272
rect 515387 645231 515439 645238
rect 515576 645410 515628 645411
rect 515576 645376 515585 645410
rect 515585 645376 515619 645410
rect 515619 645376 515628 645410
rect 515576 645359 515628 645376
rect 515576 645338 515628 645347
rect 515576 645304 515585 645338
rect 515585 645304 515619 645338
rect 515619 645304 515628 645338
rect 515576 645295 515628 645304
rect 516871 645410 516923 645411
rect 516871 645376 516880 645410
rect 516880 645376 516914 645410
rect 516914 645376 516923 645410
rect 516871 645359 516923 645376
rect 515576 645266 515628 645283
rect 515576 645232 515585 645266
rect 515585 645232 515619 645266
rect 515619 645232 515628 645266
rect 515576 645231 515628 645232
rect 514013 644768 514065 644776
rect 514013 644734 514022 644768
rect 514022 644734 514056 644768
rect 514056 644734 514065 644768
rect 514013 644724 514065 644734
rect 514013 644696 514065 644712
rect 514013 644662 514022 644696
rect 514022 644662 514056 644696
rect 514056 644662 514065 644696
rect 514013 644660 514065 644662
rect 514013 644624 514065 644648
rect 514013 644596 514022 644624
rect 514022 644596 514056 644624
rect 514056 644596 514065 644624
rect 516221 645218 516273 645249
rect 516221 645197 516230 645218
rect 516230 645197 516264 645218
rect 516264 645197 516273 645218
rect 516221 645184 516230 645185
rect 516230 645184 516264 645185
rect 516264 645184 516273 645185
rect 516221 645146 516273 645184
rect 516221 645133 516230 645146
rect 516230 645133 516264 645146
rect 516264 645133 516273 645146
rect 516221 645112 516230 645121
rect 516230 645112 516264 645121
rect 516264 645112 516273 645121
rect 516221 645074 516273 645112
rect 516221 645069 516230 645074
rect 516230 645069 516264 645074
rect 516264 645069 516273 645074
rect 516221 645040 516230 645057
rect 516230 645040 516264 645057
rect 516264 645040 516273 645057
rect 516221 645005 516273 645040
rect 516221 644968 516230 644993
rect 516230 644968 516264 644993
rect 516264 644968 516273 644993
rect 516221 644941 516273 644968
rect 516221 644896 516230 644929
rect 516230 644896 516264 644929
rect 516264 644896 516273 644929
rect 516221 644877 516273 644896
rect 516871 645338 516923 645347
rect 516871 645304 516880 645338
rect 516880 645304 516914 645338
rect 516914 645304 516923 645338
rect 516871 645295 516923 645304
rect 516871 645266 516923 645283
rect 516871 645232 516880 645266
rect 516880 645232 516914 645266
rect 516914 645232 516923 645266
rect 516871 645231 516923 645232
rect 515763 644536 515772 644559
rect 515772 644536 515806 644559
rect 515806 644536 515815 644559
rect 515763 644507 515815 644536
rect 515763 644464 515772 644495
rect 515772 644464 515806 644495
rect 515806 644464 515815 644495
rect 515763 644443 515815 644464
rect 515763 644426 515815 644431
rect 515763 644392 515772 644426
rect 515772 644392 515806 644426
rect 515806 644392 515815 644426
rect 515763 644379 515815 644392
rect 507871 643778 507923 643779
rect 507871 643744 507880 643778
rect 507880 643744 507914 643778
rect 507914 643744 507923 643778
rect 507871 643727 507923 643744
rect 507871 643706 507923 643715
rect 507871 643672 507880 643706
rect 507880 643672 507914 643706
rect 507914 643672 507923 643706
rect 507871 643663 507923 643672
rect 507871 643634 507923 643651
rect 507871 643600 507880 643634
rect 507880 643600 507914 643634
rect 507914 643600 507923 643634
rect 507871 643599 507923 643600
rect 508975 644216 508984 644244
rect 508984 644216 509018 644244
rect 509018 644216 509027 644244
rect 508975 644192 509027 644216
rect 508975 644178 509027 644180
rect 508975 644144 508984 644178
rect 508984 644144 509018 644178
rect 509018 644144 509027 644178
rect 508975 644128 509027 644144
rect 508975 644106 509027 644116
rect 508975 644072 508984 644106
rect 508984 644072 509018 644106
rect 509018 644072 509027 644106
rect 508975 644064 509027 644072
rect 508059 643746 508111 643779
rect 508059 643727 508068 643746
rect 508068 643727 508102 643746
rect 508102 643727 508111 643746
rect 508059 643712 508068 643715
rect 508068 643712 508102 643715
rect 508102 643712 508111 643715
rect 508059 643674 508111 643712
rect 508059 643663 508068 643674
rect 508068 643663 508102 643674
rect 508102 643663 508111 643674
rect 508059 643640 508068 643651
rect 508068 643640 508102 643651
rect 508102 643640 508111 643651
rect 508059 643602 508111 643640
rect 508059 643599 508068 643602
rect 508068 643599 508102 643602
rect 508102 643599 508111 643602
rect 508517 643746 508569 643779
rect 508517 643727 508526 643746
rect 508526 643727 508560 643746
rect 508560 643727 508569 643746
rect 508517 643712 508526 643715
rect 508526 643712 508560 643715
rect 508560 643712 508569 643715
rect 508517 643674 508569 643712
rect 508517 643663 508526 643674
rect 508526 643663 508560 643674
rect 508560 643663 508569 643674
rect 508517 643640 508526 643651
rect 508526 643640 508560 643651
rect 508560 643640 508569 643651
rect 508517 643602 508569 643640
rect 508517 643599 508526 643602
rect 508526 643599 508560 643602
rect 508560 643599 508569 643602
rect 509891 644216 509900 644244
rect 509900 644216 509934 644244
rect 509934 644216 509943 644244
rect 509891 644192 509943 644216
rect 509891 644178 509943 644180
rect 509891 644144 509900 644178
rect 509900 644144 509934 644178
rect 509934 644144 509943 644178
rect 509891 644128 509943 644144
rect 509891 644106 509943 644116
rect 509891 644072 509900 644106
rect 509900 644072 509934 644106
rect 509934 644072 509943 644106
rect 509891 644064 509943 644072
rect 509433 643746 509485 643779
rect 509433 643727 509442 643746
rect 509442 643727 509476 643746
rect 509476 643727 509485 643746
rect 509433 643712 509442 643715
rect 509442 643712 509476 643715
rect 509476 643712 509485 643715
rect 509433 643674 509485 643712
rect 509433 643663 509442 643674
rect 509442 643663 509476 643674
rect 509476 643663 509485 643674
rect 509433 643640 509442 643651
rect 509442 643640 509476 643651
rect 509476 643640 509485 643651
rect 509433 643602 509485 643640
rect 509433 643599 509442 643602
rect 509442 643599 509476 643602
rect 509476 643599 509485 643602
rect 510807 644216 510816 644244
rect 510816 644216 510850 644244
rect 510850 644216 510859 644244
rect 510807 644192 510859 644216
rect 510807 644178 510859 644180
rect 510807 644144 510816 644178
rect 510816 644144 510850 644178
rect 510850 644144 510859 644178
rect 510807 644128 510859 644144
rect 510807 644106 510859 644116
rect 510807 644072 510816 644106
rect 510816 644072 510850 644106
rect 510850 644072 510859 644106
rect 510807 644064 510859 644072
rect 510349 643746 510401 643779
rect 510349 643727 510358 643746
rect 510358 643727 510392 643746
rect 510392 643727 510401 643746
rect 510349 643712 510358 643715
rect 510358 643712 510392 643715
rect 510392 643712 510401 643715
rect 510349 643674 510401 643712
rect 510349 643663 510358 643674
rect 510358 643663 510392 643674
rect 510392 643663 510401 643674
rect 510349 643640 510358 643651
rect 510358 643640 510392 643651
rect 510392 643640 510401 643651
rect 510349 643602 510401 643640
rect 510349 643599 510358 643602
rect 510358 643599 510392 643602
rect 510392 643599 510401 643602
rect 511723 644216 511732 644244
rect 511732 644216 511766 644244
rect 511766 644216 511775 644244
rect 511723 644192 511775 644216
rect 511723 644178 511775 644180
rect 511723 644144 511732 644178
rect 511732 644144 511766 644178
rect 511766 644144 511775 644178
rect 511723 644128 511775 644144
rect 511723 644106 511775 644116
rect 511723 644072 511732 644106
rect 511732 644072 511766 644106
rect 511766 644072 511775 644106
rect 511723 644064 511775 644072
rect 511265 643746 511317 643779
rect 511265 643727 511274 643746
rect 511274 643727 511308 643746
rect 511308 643727 511317 643746
rect 511265 643712 511274 643715
rect 511274 643712 511308 643715
rect 511308 643712 511317 643715
rect 511265 643674 511317 643712
rect 511265 643663 511274 643674
rect 511274 643663 511308 643674
rect 511308 643663 511317 643674
rect 511265 643640 511274 643651
rect 511274 643640 511308 643651
rect 511308 643640 511317 643651
rect 511265 643602 511317 643640
rect 511265 643599 511274 643602
rect 511274 643599 511308 643602
rect 511308 643599 511317 643602
rect 512639 644216 512648 644244
rect 512648 644216 512682 644244
rect 512682 644216 512691 644244
rect 512639 644192 512691 644216
rect 512639 644178 512691 644180
rect 512639 644144 512648 644178
rect 512648 644144 512682 644178
rect 512682 644144 512691 644178
rect 512639 644128 512691 644144
rect 512639 644106 512691 644116
rect 512639 644072 512648 644106
rect 512648 644072 512682 644106
rect 512682 644072 512691 644106
rect 512639 644064 512691 644072
rect 512181 643746 512233 643779
rect 512181 643727 512190 643746
rect 512190 643727 512224 643746
rect 512224 643727 512233 643746
rect 512181 643712 512190 643715
rect 512190 643712 512224 643715
rect 512224 643712 512233 643715
rect 512181 643674 512233 643712
rect 512181 643663 512190 643674
rect 512190 643663 512224 643674
rect 512224 643663 512233 643674
rect 512181 643640 512190 643651
rect 512190 643640 512224 643651
rect 512224 643640 512233 643651
rect 512181 643602 512233 643640
rect 512181 643599 512190 643602
rect 512190 643599 512224 643602
rect 512224 643599 512233 643602
rect 513555 644216 513564 644244
rect 513564 644216 513598 644244
rect 513598 644216 513607 644244
rect 513555 644192 513607 644216
rect 513555 644178 513607 644180
rect 513555 644144 513564 644178
rect 513564 644144 513598 644178
rect 513598 644144 513607 644178
rect 513555 644128 513607 644144
rect 513555 644106 513607 644116
rect 513555 644072 513564 644106
rect 513564 644072 513598 644106
rect 513598 644072 513607 644106
rect 513555 644064 513607 644072
rect 513097 643746 513149 643779
rect 513097 643727 513106 643746
rect 513106 643727 513140 643746
rect 513140 643727 513149 643746
rect 513097 643712 513106 643715
rect 513106 643712 513140 643715
rect 513140 643712 513149 643715
rect 513097 643674 513149 643712
rect 513097 643663 513106 643674
rect 513106 643663 513140 643674
rect 513140 643663 513149 643674
rect 513097 643640 513106 643651
rect 513106 643640 513140 643651
rect 513140 643640 513149 643651
rect 513097 643602 513149 643640
rect 513097 643599 513106 643602
rect 513106 643599 513140 643602
rect 513140 643599 513149 643602
rect 514013 643746 514065 643779
rect 514013 643727 514022 643746
rect 514022 643727 514056 643746
rect 514056 643727 514065 643746
rect 514013 643712 514022 643715
rect 514022 643712 514056 643715
rect 514056 643712 514065 643715
rect 514013 643674 514065 643712
rect 514013 643663 514022 643674
rect 514022 643663 514056 643674
rect 514056 643663 514065 643674
rect 514013 643640 514022 643651
rect 514022 643640 514056 643651
rect 514056 643640 514065 643651
rect 514013 643602 514065 643640
rect 514013 643599 514022 643602
rect 514022 643599 514056 643602
rect 514056 643599 514065 643602
rect 514471 643746 514523 643779
rect 514471 643727 514480 643746
rect 514480 643727 514514 643746
rect 514514 643727 514523 643746
rect 514471 643712 514480 643715
rect 514480 643712 514514 643715
rect 514514 643712 514523 643715
rect 514471 643674 514523 643712
rect 514471 643663 514480 643674
rect 514480 643663 514514 643674
rect 514514 643663 514523 643674
rect 514471 643640 514480 643651
rect 514480 643640 514514 643651
rect 514514 643640 514523 643651
rect 514471 643602 514523 643640
rect 514471 643599 514480 643602
rect 514480 643599 514514 643602
rect 514514 643599 514523 643602
rect 515763 644354 515815 644367
rect 515763 644320 515772 644354
rect 515772 644320 515806 644354
rect 515806 644320 515815 644354
rect 515763 644315 515815 644320
rect 515763 644282 515815 644303
rect 515763 644251 515772 644282
rect 515772 644251 515806 644282
rect 515806 644251 515815 644282
rect 515763 644210 515815 644239
rect 515763 644187 515772 644210
rect 515772 644187 515806 644210
rect 515806 644187 515815 644210
rect 514929 643746 514981 643779
rect 514929 643727 514938 643746
rect 514938 643727 514972 643746
rect 514972 643727 514981 643746
rect 514929 643712 514938 643715
rect 514938 643712 514972 643715
rect 514972 643712 514981 643715
rect 514929 643674 514981 643712
rect 514929 643663 514938 643674
rect 514938 643663 514972 643674
rect 514972 643663 514981 643674
rect 514929 643640 514938 643651
rect 514938 643640 514972 643651
rect 514972 643640 514981 643651
rect 514929 643602 514981 643640
rect 514929 643599 514938 643602
rect 514938 643599 514972 643602
rect 514972 643599 514981 643602
rect 515387 643746 515439 643779
rect 515387 643727 515396 643746
rect 515396 643727 515430 643746
rect 515430 643727 515439 643746
rect 515387 643712 515396 643715
rect 515396 643712 515430 643715
rect 515430 643712 515439 643715
rect 515387 643674 515439 643712
rect 515387 643663 515396 643674
rect 515396 643663 515430 643674
rect 515430 643663 515439 643674
rect 515387 643640 515396 643651
rect 515396 643640 515430 643651
rect 515430 643640 515439 643651
rect 515387 643602 515439 643640
rect 515387 643599 515396 643602
rect 515396 643599 515430 643602
rect 515430 643599 515439 643602
rect 515575 643778 515627 643779
rect 515575 643744 515584 643778
rect 515584 643744 515618 643778
rect 515618 643744 515627 643778
rect 515575 643727 515627 643744
rect 515575 643706 515627 643715
rect 515575 643672 515584 643706
rect 515584 643672 515618 643706
rect 515618 643672 515627 643706
rect 515575 643663 515627 643672
rect 515575 643634 515627 643651
rect 515575 643600 515584 643634
rect 515584 643600 515618 643634
rect 515618 643600 515627 643634
rect 515575 643599 515627 643600
rect 516679 644536 516688 644559
rect 516688 644536 516722 644559
rect 516722 644536 516731 644559
rect 516679 644507 516731 644536
rect 516679 644464 516688 644495
rect 516688 644464 516722 644495
rect 516722 644464 516731 644495
rect 516679 644443 516731 644464
rect 516679 644426 516731 644431
rect 516679 644392 516688 644426
rect 516688 644392 516722 644426
rect 516722 644392 516731 644426
rect 516679 644379 516731 644392
rect 516679 644354 516731 644367
rect 516679 644320 516688 644354
rect 516688 644320 516722 644354
rect 516722 644320 516731 644354
rect 516679 644315 516731 644320
rect 516679 644282 516731 644303
rect 516679 644251 516688 644282
rect 516688 644251 516722 644282
rect 516722 644251 516731 644282
rect 516679 644210 516731 644239
rect 516679 644187 516688 644210
rect 516688 644187 516722 644210
rect 516722 644187 516731 644210
rect 508879 643256 508899 643290
rect 508899 643256 508931 643290
rect 508879 643238 508931 643256
rect 508943 643238 508995 643290
rect 509007 643238 509059 643290
rect 509071 643256 509103 643290
rect 509103 643256 509123 643290
rect 509071 643238 509123 643256
rect 510711 643256 510731 643290
rect 510731 643256 510763 643290
rect 510711 643238 510763 643256
rect 510775 643238 510827 643290
rect 510839 643238 510891 643290
rect 510903 643256 510935 643290
rect 510935 643256 510955 643290
rect 510903 643238 510955 643256
rect 512543 643256 512563 643290
rect 512563 643256 512595 643290
rect 512543 643238 512595 643256
rect 512607 643238 512659 643290
rect 512671 643238 512723 643290
rect 512735 643256 512767 643290
rect 512767 643256 512787 643290
rect 512735 643238 512787 643256
rect 516354 643290 516406 643299
rect 516418 643290 516470 643299
rect 516482 643290 516534 643299
rect 516546 643290 516598 643299
rect 516354 643256 516387 643290
rect 516387 643256 516406 643290
rect 516418 643256 516421 643290
rect 516421 643256 516459 643290
rect 516459 643256 516470 643290
rect 516482 643256 516493 643290
rect 516493 643256 516531 643290
rect 516531 643256 516534 643290
rect 516546 643256 516565 643290
rect 516565 643256 516598 643290
rect 516354 643247 516406 643256
rect 516418 643247 516470 643256
rect 516482 643247 516534 643256
rect 516546 643247 516598 643256
rect 515960 642792 516076 642908
rect 508879 642477 508931 642495
rect 508879 642443 508899 642477
rect 508899 642443 508931 642477
rect 508943 642443 508995 642495
rect 509007 642443 509059 642495
rect 509071 642477 509123 642495
rect 509071 642443 509103 642477
rect 509103 642443 509123 642477
rect 510711 642477 510763 642495
rect 510711 642443 510731 642477
rect 510731 642443 510763 642477
rect 510775 642443 510827 642495
rect 510839 642443 510891 642495
rect 510903 642477 510955 642495
rect 510903 642443 510935 642477
rect 510935 642443 510955 642477
rect 512543 642477 512595 642495
rect 512543 642443 512563 642477
rect 512563 642443 512595 642477
rect 512607 642443 512659 642495
rect 512671 642443 512723 642495
rect 512735 642477 512787 642495
rect 512735 642443 512767 642477
rect 512767 642443 512787 642477
rect 516353 642477 516405 642486
rect 516417 642477 516469 642486
rect 516481 642477 516533 642486
rect 516545 642477 516597 642486
rect 516353 642443 516387 642477
rect 516387 642443 516405 642477
rect 516417 642443 516421 642477
rect 516421 642443 516459 642477
rect 516459 642443 516469 642477
rect 516481 642443 516493 642477
rect 516493 642443 516531 642477
rect 516531 642443 516533 642477
rect 516545 642443 516565 642477
rect 516565 642443 516597 642477
rect 507871 642142 507923 642143
rect 507871 642108 507880 642142
rect 507880 642108 507914 642142
rect 507914 642108 507923 642142
rect 507871 642091 507923 642108
rect 507871 642070 507923 642079
rect 507871 642036 507880 642070
rect 507880 642036 507914 642070
rect 507914 642036 507923 642070
rect 507871 642027 507923 642036
rect 507871 641998 507923 642015
rect 507871 641964 507880 641998
rect 507880 641964 507914 641998
rect 507914 641964 507923 641998
rect 507871 641963 507923 641964
rect 508059 642140 508068 642143
rect 508068 642140 508102 642143
rect 508102 642140 508111 642143
rect 508059 642102 508111 642140
rect 508059 642091 508068 642102
rect 508068 642091 508102 642102
rect 508102 642091 508111 642102
rect 508059 642068 508068 642079
rect 508068 642068 508102 642079
rect 508102 642068 508111 642079
rect 508059 642030 508111 642068
rect 508059 642027 508068 642030
rect 508068 642027 508102 642030
rect 508102 642027 508111 642030
rect 508059 641996 508068 642015
rect 508068 641996 508102 642015
rect 508102 641996 508111 642015
rect 508059 641963 508111 641996
rect 508517 642140 508526 642143
rect 508526 642140 508560 642143
rect 508560 642140 508569 642143
rect 508517 642102 508569 642140
rect 508517 642091 508526 642102
rect 508526 642091 508560 642102
rect 508560 642091 508569 642102
rect 508517 642068 508526 642079
rect 508526 642068 508560 642079
rect 508560 642068 508569 642079
rect 508517 642030 508569 642068
rect 508517 642027 508526 642030
rect 508526 642027 508560 642030
rect 508560 642027 508569 642030
rect 508517 641996 508526 642015
rect 508526 641996 508560 642015
rect 508560 641996 508569 642015
rect 508517 641963 508569 641996
rect 509433 642140 509442 642143
rect 509442 642140 509476 642143
rect 509476 642140 509485 642143
rect 509433 642102 509485 642140
rect 509433 642091 509442 642102
rect 509442 642091 509476 642102
rect 509476 642091 509485 642102
rect 509433 642068 509442 642079
rect 509442 642068 509476 642079
rect 509476 642068 509485 642079
rect 509433 642030 509485 642068
rect 509433 642027 509442 642030
rect 509442 642027 509476 642030
rect 509476 642027 509485 642030
rect 509433 641996 509442 642015
rect 509442 641996 509476 642015
rect 509476 641996 509485 642015
rect 509433 641963 509485 641996
rect 508975 641670 509027 641678
rect 508975 641636 508984 641670
rect 508984 641636 509018 641670
rect 509018 641636 509027 641670
rect 508975 641626 509027 641636
rect 508975 641598 509027 641614
rect 508975 641564 508984 641598
rect 508984 641564 509018 641598
rect 509018 641564 509027 641598
rect 508975 641562 509027 641564
rect 508975 641526 509027 641550
rect 508975 641498 508984 641526
rect 508984 641498 509018 641526
rect 509018 641498 509027 641526
rect 510349 642140 510358 642143
rect 510358 642140 510392 642143
rect 510392 642140 510401 642143
rect 510349 642102 510401 642140
rect 510349 642091 510358 642102
rect 510358 642091 510392 642102
rect 510392 642091 510401 642102
rect 510349 642068 510358 642079
rect 510358 642068 510392 642079
rect 510392 642068 510401 642079
rect 510349 642030 510401 642068
rect 510349 642027 510358 642030
rect 510358 642027 510392 642030
rect 510392 642027 510401 642030
rect 510349 641996 510358 642015
rect 510358 641996 510392 642015
rect 510392 641996 510401 642015
rect 510349 641963 510401 641996
rect 509891 641670 509943 641678
rect 509891 641636 509900 641670
rect 509900 641636 509934 641670
rect 509934 641636 509943 641670
rect 509891 641626 509943 641636
rect 509891 641598 509943 641614
rect 509891 641564 509900 641598
rect 509900 641564 509934 641598
rect 509934 641564 509943 641598
rect 509891 641562 509943 641564
rect 509891 641526 509943 641550
rect 509891 641498 509900 641526
rect 509900 641498 509934 641526
rect 509934 641498 509943 641526
rect 511265 642140 511274 642143
rect 511274 642140 511308 642143
rect 511308 642140 511317 642143
rect 511265 642102 511317 642140
rect 511265 642091 511274 642102
rect 511274 642091 511308 642102
rect 511308 642091 511317 642102
rect 511265 642068 511274 642079
rect 511274 642068 511308 642079
rect 511308 642068 511317 642079
rect 511265 642030 511317 642068
rect 511265 642027 511274 642030
rect 511274 642027 511308 642030
rect 511308 642027 511317 642030
rect 511265 641996 511274 642015
rect 511274 641996 511308 642015
rect 511308 641996 511317 642015
rect 511265 641963 511317 641996
rect 510807 641670 510859 641678
rect 510807 641636 510816 641670
rect 510816 641636 510850 641670
rect 510850 641636 510859 641670
rect 510807 641626 510859 641636
rect 510807 641598 510859 641614
rect 510807 641564 510816 641598
rect 510816 641564 510850 641598
rect 510850 641564 510859 641598
rect 510807 641562 510859 641564
rect 510807 641526 510859 641550
rect 510807 641498 510816 641526
rect 510816 641498 510850 641526
rect 510850 641498 510859 641526
rect 512181 642140 512190 642143
rect 512190 642140 512224 642143
rect 512224 642140 512233 642143
rect 512181 642102 512233 642140
rect 512181 642091 512190 642102
rect 512190 642091 512224 642102
rect 512224 642091 512233 642102
rect 512181 642068 512190 642079
rect 512190 642068 512224 642079
rect 512224 642068 512233 642079
rect 512181 642030 512233 642068
rect 512181 642027 512190 642030
rect 512190 642027 512224 642030
rect 512224 642027 512233 642030
rect 512181 641996 512190 642015
rect 512190 641996 512224 642015
rect 512224 641996 512233 642015
rect 512181 641963 512233 641996
rect 511723 641670 511775 641678
rect 511723 641636 511732 641670
rect 511732 641636 511766 641670
rect 511766 641636 511775 641670
rect 511723 641626 511775 641636
rect 511723 641598 511775 641614
rect 511723 641564 511732 641598
rect 511732 641564 511766 641598
rect 511766 641564 511775 641598
rect 511723 641562 511775 641564
rect 511723 641526 511775 641550
rect 511723 641498 511732 641526
rect 511732 641498 511766 641526
rect 511766 641498 511775 641526
rect 513097 642140 513106 642143
rect 513106 642140 513140 642143
rect 513140 642140 513149 642143
rect 513097 642102 513149 642140
rect 513097 642091 513106 642102
rect 513106 642091 513140 642102
rect 513140 642091 513149 642102
rect 513097 642068 513106 642079
rect 513106 642068 513140 642079
rect 513140 642068 513149 642079
rect 513097 642030 513149 642068
rect 513097 642027 513106 642030
rect 513106 642027 513140 642030
rect 513140 642027 513149 642030
rect 513097 641996 513106 642015
rect 513106 641996 513140 642015
rect 513140 641996 513149 642015
rect 513097 641963 513149 641996
rect 512639 641670 512691 641678
rect 512639 641636 512648 641670
rect 512648 641636 512682 641670
rect 512682 641636 512691 641670
rect 512639 641626 512691 641636
rect 512639 641598 512691 641614
rect 512639 641564 512648 641598
rect 512648 641564 512682 641598
rect 512682 641564 512691 641598
rect 512639 641562 512691 641564
rect 512639 641526 512691 641550
rect 512639 641498 512648 641526
rect 512648 641498 512682 641526
rect 512682 641498 512691 641526
rect 514013 642140 514022 642143
rect 514022 642140 514056 642143
rect 514056 642140 514065 642143
rect 514013 642102 514065 642140
rect 514013 642091 514022 642102
rect 514022 642091 514056 642102
rect 514056 642091 514065 642102
rect 514013 642068 514022 642079
rect 514022 642068 514056 642079
rect 514056 642068 514065 642079
rect 514013 642030 514065 642068
rect 514013 642027 514022 642030
rect 514022 642027 514056 642030
rect 514056 642027 514065 642030
rect 514013 641996 514022 642015
rect 514022 641996 514056 642015
rect 514056 641996 514065 642015
rect 514013 641963 514065 641996
rect 516353 642434 516405 642443
rect 516417 642434 516469 642443
rect 516481 642434 516533 642443
rect 516545 642434 516597 642443
rect 514471 642140 514480 642143
rect 514480 642140 514514 642143
rect 514514 642140 514523 642143
rect 514471 642102 514523 642140
rect 514471 642091 514480 642102
rect 514480 642091 514514 642102
rect 514514 642091 514523 642102
rect 514471 642068 514480 642079
rect 514480 642068 514514 642079
rect 514514 642068 514523 642079
rect 514471 642030 514523 642068
rect 514471 642027 514480 642030
rect 514480 642027 514514 642030
rect 514514 642027 514523 642030
rect 514471 641996 514480 642015
rect 514480 641996 514514 642015
rect 514514 641996 514523 642015
rect 514471 641963 514523 641996
rect 513555 641670 513607 641678
rect 513555 641636 513564 641670
rect 513564 641636 513598 641670
rect 513598 641636 513607 641670
rect 513555 641626 513607 641636
rect 513555 641598 513607 641614
rect 513555 641564 513564 641598
rect 513564 641564 513598 641598
rect 513598 641564 513607 641598
rect 513555 641562 513607 641564
rect 513555 641526 513607 641550
rect 513555 641498 513564 641526
rect 513564 641498 513598 641526
rect 513598 641498 513607 641526
rect 514929 642140 514938 642143
rect 514938 642140 514972 642143
rect 514972 642140 514981 642143
rect 514929 642102 514981 642140
rect 514929 642091 514938 642102
rect 514938 642091 514972 642102
rect 514972 642091 514981 642102
rect 514929 642068 514938 642079
rect 514938 642068 514972 642079
rect 514972 642068 514981 642079
rect 514929 642030 514981 642068
rect 514929 642027 514938 642030
rect 514938 642027 514972 642030
rect 514972 642027 514981 642030
rect 514929 641996 514938 642015
rect 514938 641996 514972 642015
rect 514972 641996 514981 642015
rect 514929 641963 514981 641996
rect 515763 642212 515772 642243
rect 515772 642212 515806 642243
rect 515806 642212 515815 642243
rect 515763 642191 515815 642212
rect 515387 642140 515396 642143
rect 515396 642140 515430 642143
rect 515430 642140 515439 642143
rect 515387 642102 515439 642140
rect 515387 642091 515396 642102
rect 515396 642091 515430 642102
rect 515430 642091 515439 642102
rect 515387 642068 515396 642079
rect 515396 642068 515430 642079
rect 515430 642068 515439 642079
rect 515387 642030 515439 642068
rect 515387 642027 515396 642030
rect 515396 642027 515430 642030
rect 515430 642027 515439 642030
rect 515387 641996 515396 642015
rect 515396 641996 515430 642015
rect 515430 641996 515439 642015
rect 515387 641963 515439 641996
rect 515575 642142 515627 642143
rect 515575 642108 515584 642142
rect 515584 642108 515618 642142
rect 515618 642108 515627 642142
rect 515575 642091 515627 642108
rect 515575 642070 515627 642079
rect 515575 642036 515584 642070
rect 515584 642036 515618 642070
rect 515618 642036 515627 642070
rect 515575 642027 515627 642036
rect 515575 641998 515627 642015
rect 515575 641964 515584 641998
rect 515584 641964 515618 641998
rect 515618 641964 515627 641998
rect 515575 641963 515627 641964
rect 515763 642174 515815 642179
rect 515763 642140 515772 642174
rect 515772 642140 515806 642174
rect 515806 642140 515815 642174
rect 515763 642127 515815 642140
rect 515763 642102 515815 642115
rect 515763 642068 515772 642102
rect 515772 642068 515806 642102
rect 515806 642068 515815 642102
rect 515763 642063 515815 642068
rect 515763 642030 515815 642051
rect 515763 641999 515772 642030
rect 515772 641999 515806 642030
rect 515806 641999 515815 642030
rect 515763 641958 515815 641987
rect 515763 641935 515772 641958
rect 515772 641935 515806 641958
rect 515806 641935 515815 641958
rect 515763 641886 515815 641923
rect 515763 641871 515772 641886
rect 515772 641871 515806 641886
rect 515806 641871 515815 641886
rect 516679 642212 516688 642243
rect 516688 642212 516722 642243
rect 516722 642212 516731 642243
rect 516679 642191 516731 642212
rect 516679 642174 516731 642179
rect 516679 642140 516688 642174
rect 516688 642140 516722 642174
rect 516722 642140 516731 642174
rect 516679 642127 516731 642140
rect 516679 642102 516731 642115
rect 516679 642068 516688 642102
rect 516688 642068 516722 642102
rect 516722 642068 516731 642102
rect 516679 642063 516731 642068
rect 516679 642030 516731 642051
rect 516679 641999 516688 642030
rect 516688 641999 516722 642030
rect 516722 641999 516731 642030
rect 516679 641958 516731 641987
rect 516679 641935 516688 641958
rect 516688 641935 516722 641958
rect 516722 641935 516731 641958
rect 516679 641886 516731 641923
rect 516679 641871 516688 641886
rect 516688 641871 516722 641886
rect 516722 641871 516731 641886
rect 516221 641780 516230 641791
rect 516230 641780 516264 641791
rect 516264 641780 516273 641791
rect 516221 641742 516273 641780
rect 516221 641739 516230 641742
rect 516230 641739 516264 641742
rect 516264 641739 516273 641742
rect 516221 641708 516230 641727
rect 516230 641708 516264 641727
rect 516264 641708 516273 641727
rect 516221 641675 516273 641708
rect 516221 641636 516230 641663
rect 516230 641636 516264 641663
rect 516264 641636 516273 641663
rect 516221 641611 516273 641636
rect 516221 641598 516273 641599
rect 516221 641564 516230 641598
rect 516230 641564 516264 641598
rect 516264 641564 516273 641598
rect 516221 641547 516273 641564
rect 516221 641526 516273 641535
rect 516221 641492 516230 641526
rect 516230 641492 516264 641526
rect 516264 641492 516273 641526
rect 516221 641483 516273 641492
rect 509433 641156 509485 641188
rect 509433 641136 509442 641156
rect 509442 641136 509476 641156
rect 509476 641136 509485 641156
rect 509433 641122 509442 641124
rect 509442 641122 509476 641124
rect 509476 641122 509485 641124
rect 509433 641084 509485 641122
rect 509433 641072 509442 641084
rect 509442 641072 509476 641084
rect 509476 641072 509485 641084
rect 509433 641050 509442 641060
rect 509442 641050 509476 641060
rect 509476 641050 509485 641060
rect 509433 641012 509485 641050
rect 509433 641008 509442 641012
rect 509442 641008 509476 641012
rect 509476 641008 509485 641012
rect 507870 640502 507922 640503
rect 507870 640468 507879 640502
rect 507879 640468 507913 640502
rect 507913 640468 507922 640502
rect 507870 640451 507922 640468
rect 507870 640430 507922 640439
rect 507870 640396 507879 640430
rect 507879 640396 507913 640430
rect 507913 640396 507922 640430
rect 507870 640387 507922 640396
rect 507870 640358 507922 640375
rect 507870 640324 507879 640358
rect 507879 640324 507913 640358
rect 507913 640324 507922 640358
rect 507870 640323 507922 640324
rect 508059 640474 508068 640503
rect 508068 640474 508102 640503
rect 508102 640474 508111 640503
rect 508059 640451 508111 640474
rect 508059 640436 508111 640439
rect 508059 640402 508068 640436
rect 508068 640402 508102 640436
rect 508102 640402 508111 640436
rect 508059 640387 508111 640402
rect 508059 640364 508111 640375
rect 508059 640330 508068 640364
rect 508068 640330 508102 640364
rect 508102 640330 508111 640364
rect 508059 640323 508111 640330
rect 508517 640474 508526 640503
rect 508526 640474 508560 640503
rect 508560 640474 508569 640503
rect 508517 640451 508569 640474
rect 508517 640436 508569 640439
rect 508517 640402 508526 640436
rect 508526 640402 508560 640436
rect 508560 640402 508569 640436
rect 508517 640387 508569 640402
rect 508517 640364 508569 640375
rect 508517 640330 508526 640364
rect 508526 640330 508560 640364
rect 508560 640330 508569 640364
rect 508517 640323 508569 640330
rect 508975 640474 508984 640503
rect 508984 640474 509018 640503
rect 509018 640474 509027 640503
rect 508975 640451 509027 640474
rect 508975 640436 509027 640439
rect 508975 640402 508984 640436
rect 508984 640402 509018 640436
rect 509018 640402 509027 640436
rect 508975 640387 509027 640402
rect 508975 640364 509027 640375
rect 508975 640330 508984 640364
rect 508984 640330 509018 640364
rect 509018 640330 509027 640364
rect 508975 640323 509027 640330
rect 510349 641156 510401 641188
rect 510349 641136 510358 641156
rect 510358 641136 510392 641156
rect 510392 641136 510401 641156
rect 510349 641122 510358 641124
rect 510358 641122 510392 641124
rect 510392 641122 510401 641124
rect 510349 641084 510401 641122
rect 510349 641072 510358 641084
rect 510358 641072 510392 641084
rect 510392 641072 510401 641084
rect 510349 641050 510358 641060
rect 510358 641050 510392 641060
rect 510392 641050 510401 641060
rect 510349 641012 510401 641050
rect 510349 641008 510358 641012
rect 510358 641008 510392 641012
rect 510392 641008 510401 641012
rect 509891 640474 509900 640503
rect 509900 640474 509934 640503
rect 509934 640474 509943 640503
rect 509891 640451 509943 640474
rect 509891 640436 509943 640439
rect 509891 640402 509900 640436
rect 509900 640402 509934 640436
rect 509934 640402 509943 640436
rect 509891 640387 509943 640402
rect 509891 640364 509943 640375
rect 509891 640330 509900 640364
rect 509900 640330 509934 640364
rect 509934 640330 509943 640364
rect 509891 640323 509943 640330
rect 511265 640796 511317 640834
rect 511265 640782 511274 640796
rect 511274 640782 511308 640796
rect 511308 640782 511317 640796
rect 511265 640762 511274 640770
rect 511274 640762 511308 640770
rect 511308 640762 511317 640770
rect 511265 640724 511317 640762
rect 511265 640718 511274 640724
rect 511274 640718 511308 640724
rect 511308 640718 511317 640724
rect 511265 640690 511274 640706
rect 511274 640690 511308 640706
rect 511308 640690 511317 640706
rect 511265 640654 511317 640690
rect 510807 640474 510816 640503
rect 510816 640474 510850 640503
rect 510850 640474 510859 640503
rect 510807 640451 510859 640474
rect 510807 640436 510859 640439
rect 510807 640402 510816 640436
rect 510816 640402 510850 640436
rect 510850 640402 510859 640436
rect 510807 640387 510859 640402
rect 510807 640364 510859 640375
rect 510807 640330 510816 640364
rect 510816 640330 510850 640364
rect 510850 640330 510859 640364
rect 510807 640323 510859 640330
rect 513097 641156 513149 641188
rect 513097 641136 513106 641156
rect 513106 641136 513140 641156
rect 513140 641136 513149 641156
rect 513097 641122 513106 641124
rect 513106 641122 513140 641124
rect 513140 641122 513149 641124
rect 513097 641084 513149 641122
rect 513097 641072 513106 641084
rect 513106 641072 513140 641084
rect 513140 641072 513149 641084
rect 513097 641050 513106 641060
rect 513106 641050 513140 641060
rect 513140 641050 513149 641060
rect 513097 641012 513149 641050
rect 513097 641008 513106 641012
rect 513106 641008 513140 641012
rect 513140 641008 513149 641012
rect 512181 640796 512233 640834
rect 512181 640782 512190 640796
rect 512190 640782 512224 640796
rect 512224 640782 512233 640796
rect 512181 640762 512190 640770
rect 512190 640762 512224 640770
rect 512224 640762 512233 640770
rect 512181 640724 512233 640762
rect 512181 640718 512190 640724
rect 512190 640718 512224 640724
rect 512224 640718 512233 640724
rect 512181 640690 512190 640706
rect 512190 640690 512224 640706
rect 512224 640690 512233 640706
rect 512181 640654 512233 640690
rect 511723 640474 511732 640503
rect 511732 640474 511766 640503
rect 511766 640474 511775 640503
rect 511723 640451 511775 640474
rect 511723 640436 511775 640439
rect 511723 640402 511732 640436
rect 511732 640402 511766 640436
rect 511766 640402 511775 640436
rect 511723 640387 511775 640402
rect 511723 640364 511775 640375
rect 511723 640330 511732 640364
rect 511732 640330 511766 640364
rect 511766 640330 511775 640364
rect 511723 640323 511775 640330
rect 512639 640474 512648 640503
rect 512648 640474 512682 640503
rect 512682 640474 512691 640503
rect 512639 640451 512691 640474
rect 512639 640436 512691 640439
rect 512639 640402 512648 640436
rect 512648 640402 512682 640436
rect 512682 640402 512691 640436
rect 512639 640387 512691 640402
rect 512639 640364 512691 640375
rect 512639 640330 512648 640364
rect 512648 640330 512682 640364
rect 512682 640330 512691 640364
rect 512639 640323 512691 640330
rect 514013 641156 514065 641188
rect 514013 641136 514022 641156
rect 514022 641136 514056 641156
rect 514056 641136 514065 641156
rect 514013 641122 514022 641124
rect 514022 641122 514056 641124
rect 514056 641122 514065 641124
rect 514013 641084 514065 641122
rect 514013 641072 514022 641084
rect 514022 641072 514056 641084
rect 514056 641072 514065 641084
rect 514013 641050 514022 641060
rect 514022 641050 514056 641060
rect 514056 641050 514065 641060
rect 514013 641012 514065 641050
rect 514013 641008 514022 641012
rect 514022 641008 514056 641012
rect 514056 641008 514065 641012
rect 513555 640474 513564 640503
rect 513564 640474 513598 640503
rect 513598 640474 513607 640503
rect 513555 640451 513607 640474
rect 513555 640436 513607 640439
rect 513555 640402 513564 640436
rect 513564 640402 513598 640436
rect 513598 640402 513607 640436
rect 513555 640387 513607 640402
rect 513555 640364 513607 640375
rect 513555 640330 513564 640364
rect 513564 640330 513598 640364
rect 513598 640330 513607 640364
rect 513555 640323 513607 640330
rect 514471 640474 514480 640503
rect 514480 640474 514514 640503
rect 514514 640474 514523 640503
rect 514471 640451 514523 640474
rect 514471 640436 514523 640439
rect 514471 640402 514480 640436
rect 514480 640402 514514 640436
rect 514514 640402 514523 640436
rect 514471 640387 514523 640402
rect 514471 640364 514523 640375
rect 514471 640330 514480 640364
rect 514480 640330 514514 640364
rect 514514 640330 514523 640364
rect 514471 640323 514523 640330
rect 514929 640474 514938 640503
rect 514938 640474 514972 640503
rect 514972 640474 514981 640503
rect 514929 640451 514981 640474
rect 514929 640436 514981 640439
rect 514929 640402 514938 640436
rect 514938 640402 514972 640436
rect 514972 640402 514981 640436
rect 514929 640387 514981 640402
rect 514929 640364 514981 640375
rect 514929 640330 514938 640364
rect 514938 640330 514972 640364
rect 514972 640330 514981 640364
rect 514929 640323 514981 640330
rect 515387 640474 515396 640503
rect 515396 640474 515430 640503
rect 515430 640474 515439 640503
rect 515387 640451 515439 640474
rect 515387 640436 515439 640439
rect 515387 640402 515396 640436
rect 515396 640402 515430 640436
rect 515430 640402 515439 640436
rect 515387 640387 515439 640402
rect 515387 640364 515439 640375
rect 515387 640330 515396 640364
rect 515396 640330 515430 640364
rect 515430 640330 515439 640364
rect 515387 640323 515439 640330
rect 515661 640502 516033 640503
rect 515661 640324 516033 640502
rect 515661 640323 516033 640324
<< metal2 >>
rect 515532 645438 515670 645453
rect 507864 645411 507928 645417
rect 507864 645359 507870 645411
rect 507922 645401 507928 645411
rect 508053 645411 508117 645417
rect 508053 645401 508059 645411
rect 507922 645359 508059 645401
rect 508111 645401 508117 645411
rect 508511 645411 508575 645417
rect 508511 645401 508517 645411
rect 508111 645359 508517 645401
rect 508569 645401 508575 645411
rect 508969 645411 509033 645417
rect 508969 645401 508975 645411
rect 508569 645359 508975 645401
rect 509027 645401 509033 645411
rect 509885 645411 509949 645417
rect 509885 645401 509891 645411
rect 509027 645389 509891 645401
rect 509943 645401 509949 645411
rect 510801 645411 510865 645417
rect 510801 645401 510807 645411
rect 509943 645389 510807 645401
rect 510577 645359 510807 645389
rect 510859 645401 510865 645411
rect 511717 645411 511781 645417
rect 511717 645401 511723 645411
rect 510859 645359 511723 645401
rect 511775 645401 511781 645411
rect 512633 645411 512697 645417
rect 512633 645401 512639 645411
rect 511775 645359 512639 645401
rect 512691 645401 512697 645411
rect 513549 645411 513613 645417
rect 513549 645401 513555 645411
rect 512691 645359 513555 645401
rect 513607 645401 513613 645411
rect 514465 645411 514529 645417
rect 514465 645401 514471 645411
rect 513607 645359 514471 645401
rect 514523 645401 514529 645411
rect 514923 645411 514987 645417
rect 514923 645401 514929 645411
rect 514523 645359 514929 645401
rect 514981 645401 514987 645411
rect 515381 645411 515445 645417
rect 515381 645401 515387 645411
rect 514981 645359 515387 645401
rect 515439 645401 515445 645411
rect 515532 645401 515572 645438
rect 515439 645382 515572 645401
rect 515628 645401 515670 645438
rect 516865 645411 516929 645417
rect 516865 645401 516871 645411
rect 515439 645359 515576 645382
rect 515628 645359 516871 645401
rect 516923 645359 516929 645411
rect 507864 645347 509001 645359
rect 510577 645358 516929 645359
rect 510577 645347 515572 645358
rect 515628 645347 516929 645358
rect 507864 645295 507870 645347
rect 507922 645295 508059 645347
rect 508111 645295 508517 645347
rect 508569 645295 508975 645347
rect 510577 645295 510807 645347
rect 510859 645295 511723 645347
rect 511775 645295 512639 645347
rect 512691 645295 513555 645347
rect 513607 645295 514471 645347
rect 514523 645295 514929 645347
rect 514981 645295 515387 645347
rect 515439 645302 515572 645347
rect 515439 645295 515576 645302
rect 515628 645295 516871 645347
rect 516923 645295 516929 645347
rect 507864 645283 509001 645295
rect 510577 645283 516929 645295
rect 507864 645231 507870 645283
rect 507922 645241 508059 645283
rect 507922 645231 507928 645241
rect 507864 645225 507928 645231
rect 508053 645231 508059 645241
rect 508111 645241 508517 645283
rect 508111 645231 508117 645241
rect 508053 645225 508117 645231
rect 508511 645231 508517 645241
rect 508569 645241 508975 645283
rect 510577 645253 510807 645283
rect 508569 645231 508575 645241
rect 508511 645225 508575 645231
rect 508969 645231 508975 645241
rect 509027 645241 509891 645253
rect 509027 645231 509033 645241
rect 508969 645225 509033 645231
rect 509885 645231 509891 645241
rect 509943 645241 510807 645253
rect 509943 645231 509949 645241
rect 509885 645225 509949 645231
rect 510801 645231 510807 645241
rect 510859 645241 511723 645283
rect 510859 645231 510865 645241
rect 510801 645225 510865 645231
rect 511717 645231 511723 645241
rect 511775 645241 512639 645283
rect 511775 645231 511781 645241
rect 511717 645225 511781 645231
rect 512633 645231 512639 645241
rect 512691 645241 513555 645283
rect 512691 645231 512697 645241
rect 512633 645225 512697 645231
rect 513549 645231 513555 645241
rect 513607 645241 514471 645283
rect 513607 645231 513613 645241
rect 513549 645225 513613 645231
rect 514465 645231 514471 645241
rect 514523 645241 514929 645283
rect 514523 645231 514529 645241
rect 514465 645225 514529 645231
rect 514923 645231 514929 645241
rect 514981 645241 515387 645283
rect 514981 645231 514987 645241
rect 514923 645225 514987 645231
rect 515381 645231 515387 645241
rect 515439 645278 515576 645283
rect 515439 645241 515572 645278
rect 515439 645231 515445 645241
rect 515381 645225 515445 645231
rect 515532 645222 515572 645241
rect 515628 645249 516871 645283
rect 515628 645241 516221 645249
rect 515628 645222 515670 645241
rect 515532 645207 515670 645222
rect 516215 645197 516221 645241
rect 516273 645241 516871 645249
rect 516273 645197 516279 645241
rect 516865 645231 516871 645241
rect 516923 645231 516929 645283
rect 516865 645225 516929 645231
rect 516215 645185 516279 645197
rect 516215 645133 516221 645185
rect 516273 645133 516279 645185
rect 516215 645121 516279 645133
rect 509422 645106 509496 645115
rect 509422 645050 509431 645106
rect 509487 645050 509496 645106
rect 514002 645106 514076 645115
rect 509422 645048 509496 645050
rect 511259 645088 511323 645094
rect 511259 645048 511265 645088
rect 509422 645036 511265 645048
rect 511317 645036 511323 645088
rect 509422 645026 511323 645036
rect 509422 644970 509431 645026
rect 509487 645024 511323 645026
rect 509487 644972 511265 645024
rect 511317 644972 511323 645024
rect 509487 644970 511323 644972
rect 509422 644960 511323 644970
rect 509422 644948 511265 644960
rect 509422 644946 509496 644948
rect 509422 644890 509431 644946
rect 509487 644890 509496 644946
rect 511259 644908 511265 644948
rect 511317 644908 511323 644960
rect 511259 644902 511323 644908
rect 512175 645088 512239 645094
rect 512175 645036 512181 645088
rect 512233 645048 512239 645088
rect 514002 645050 514011 645106
rect 514067 645050 514076 645106
rect 514002 645048 514076 645050
rect 512233 645036 514076 645048
rect 512175 645026 514076 645036
rect 512175 645024 514011 645026
rect 512175 644972 512181 645024
rect 512233 644972 514011 645024
rect 512175 644970 514011 644972
rect 514067 644970 514076 645026
rect 512175 644960 514076 644970
rect 512175 644908 512181 644960
rect 512233 644948 514076 644960
rect 512233 644908 512239 644948
rect 512175 644902 512239 644908
rect 514002 644946 514076 644948
rect 509422 644881 509496 644890
rect 514002 644890 514011 644946
rect 514067 644890 514076 644946
rect 514002 644881 514076 644890
rect 516215 645069 516221 645121
rect 516273 645069 516279 645121
rect 516215 645057 516279 645069
rect 516215 645005 516221 645057
rect 516273 645005 516279 645057
rect 516215 644993 516279 645005
rect 516215 644941 516221 644993
rect 516273 644941 516279 644993
rect 516215 644929 516279 644941
rect 516215 644877 516221 644929
rect 516273 644877 516279 644929
rect 516215 644871 516279 644877
rect 509880 644794 509954 644803
rect 509427 644776 509491 644782
rect 509427 644724 509433 644776
rect 509485 644736 509491 644776
rect 509880 644738 509889 644794
rect 509945 644738 509954 644794
rect 511254 644794 511328 644803
rect 509880 644736 509954 644738
rect 509485 644724 509954 644736
rect 509427 644714 509954 644724
rect 509427 644712 509889 644714
rect 509427 644660 509433 644712
rect 509485 644660 509889 644712
rect 509427 644658 509889 644660
rect 509945 644658 509954 644714
rect 509427 644648 509954 644658
rect 509427 644596 509433 644648
rect 509485 644636 509954 644648
rect 509485 644596 509491 644636
rect 509427 644590 509491 644596
rect 509880 644634 509954 644636
rect 509880 644578 509889 644634
rect 509945 644578 509954 644634
rect 510343 644776 510407 644782
rect 510343 644724 510349 644776
rect 510401 644736 510407 644776
rect 511254 644738 511263 644794
rect 511319 644738 511328 644794
rect 511254 644736 511328 644738
rect 510401 644724 511328 644736
rect 510343 644714 511328 644724
rect 510343 644712 511263 644714
rect 510343 644660 510349 644712
rect 510401 644660 511263 644712
rect 510343 644658 511263 644660
rect 511319 644658 511328 644714
rect 510343 644648 511328 644658
rect 510343 644596 510349 644648
rect 510401 644636 511328 644648
rect 510401 644596 510407 644636
rect 510343 644590 510407 644596
rect 511254 644634 511328 644636
rect 509880 644569 509954 644578
rect 511254 644578 511263 644634
rect 511319 644578 511328 644634
rect 511254 644569 511328 644578
rect 512170 644794 512244 644803
rect 512170 644738 512179 644794
rect 512235 644738 512244 644794
rect 513544 644794 513618 644803
rect 512170 644736 512244 644738
rect 513091 644776 513155 644782
rect 513091 644736 513097 644776
rect 512170 644724 513097 644736
rect 513149 644724 513155 644776
rect 512170 644714 513155 644724
rect 512170 644658 512179 644714
rect 512235 644712 513155 644714
rect 512235 644660 513097 644712
rect 513149 644660 513155 644712
rect 512235 644658 513155 644660
rect 512170 644648 513155 644658
rect 512170 644636 513097 644648
rect 512170 644634 512244 644636
rect 512170 644578 512179 644634
rect 512235 644578 512244 644634
rect 513091 644596 513097 644636
rect 513149 644596 513155 644648
rect 513091 644590 513155 644596
rect 513544 644738 513553 644794
rect 513609 644738 513618 644794
rect 513544 644736 513618 644738
rect 514007 644776 514071 644782
rect 514007 644736 514013 644776
rect 513544 644724 514013 644736
rect 514065 644724 514071 644776
rect 513544 644714 514071 644724
rect 513544 644658 513553 644714
rect 513609 644712 514071 644714
rect 513609 644660 514013 644712
rect 514065 644660 514071 644712
rect 513609 644658 514071 644660
rect 513544 644648 514071 644658
rect 513544 644636 514013 644648
rect 513544 644634 513618 644636
rect 512170 644569 512244 644578
rect 513544 644578 513553 644634
rect 513609 644578 513618 644634
rect 514007 644596 514013 644636
rect 514065 644596 514071 644648
rect 514007 644590 514071 644596
rect 516668 644601 516742 644610
rect 513544 644569 513618 644578
rect 515757 644559 515821 644565
rect 515757 644507 515763 644559
rect 515815 644507 515821 644559
rect 515757 644495 515821 644507
rect 515757 644443 515763 644495
rect 515815 644443 515821 644495
rect 515757 644431 515821 644443
rect 515757 644379 515763 644431
rect 515815 644423 515821 644431
rect 516668 644545 516677 644601
rect 516733 644545 516742 644601
rect 516668 644521 516679 644545
rect 516731 644521 516742 644545
rect 516668 644465 516677 644521
rect 516733 644465 516742 644521
rect 516668 644443 516679 644465
rect 516731 644443 516742 644465
rect 516668 644441 516742 644443
rect 515815 644379 516526 644423
rect 515757 644367 516526 644379
rect 515757 644315 515763 644367
rect 515815 644323 516526 644367
rect 515815 644315 515821 644323
rect 515757 644303 515821 644315
rect 515757 644251 515763 644303
rect 515815 644251 515821 644303
rect 508969 644244 509033 644250
rect 508969 644192 508975 644244
rect 509027 644234 509033 644244
rect 509885 644244 509949 644250
rect 509885 644234 509891 644244
rect 509027 644192 509891 644234
rect 509943 644234 509949 644244
rect 510801 644244 510865 644250
rect 510801 644234 510807 644244
rect 509943 644192 510807 644234
rect 510859 644234 510865 644244
rect 511717 644244 511781 644250
rect 511717 644234 511723 644244
rect 510859 644192 511723 644234
rect 511775 644234 511781 644244
rect 512633 644244 512697 644250
rect 512633 644234 512639 644244
rect 511775 644192 512639 644234
rect 512691 644234 512697 644244
rect 513549 644244 513613 644250
rect 513549 644234 513555 644244
rect 512691 644192 513555 644234
rect 513607 644192 513613 644244
rect 508969 644180 513613 644192
rect 515757 644239 515821 644251
rect 515757 644187 515763 644239
rect 515815 644187 515821 644239
rect 515757 644181 515821 644187
rect 508969 644128 508975 644180
rect 509027 644128 509891 644180
rect 509943 644128 510807 644180
rect 510859 644128 511723 644180
rect 511775 644128 512639 644180
rect 512691 644128 513555 644180
rect 513607 644128 513613 644180
rect 508969 644116 513613 644128
rect 508969 644064 508975 644116
rect 509027 644074 509891 644116
rect 509027 644064 509033 644074
rect 508969 644058 509033 644064
rect 509885 644064 509891 644074
rect 509943 644074 510807 644116
rect 509943 644064 509949 644074
rect 509885 644058 509949 644064
rect 510801 644064 510807 644074
rect 510859 644074 511723 644116
rect 510859 644064 510865 644074
rect 510801 644058 510865 644064
rect 511717 644064 511723 644074
rect 511775 644074 512639 644116
rect 511775 644064 511781 644074
rect 511717 644058 511781 644064
rect 512633 644064 512639 644074
rect 512691 644074 513555 644116
rect 512691 644064 512697 644074
rect 512633 644058 512697 644064
rect 513549 644064 513555 644074
rect 513607 644064 513613 644116
rect 513549 644058 513613 644064
rect 510338 643797 510412 643806
rect 507865 643779 507929 643785
rect 507865 643727 507871 643779
rect 507923 643769 507929 643779
rect 508053 643779 508117 643785
rect 508053 643769 508059 643779
rect 507923 643757 508059 643769
rect 508111 643769 508117 643779
rect 508511 643779 508575 643785
rect 508511 643769 508517 643779
rect 508111 643757 508517 643769
rect 508569 643769 508575 643779
rect 509427 643779 509491 643785
rect 509427 643769 509433 643779
rect 508569 643757 509433 643769
rect 507923 643727 508012 643757
rect 509108 643727 509433 643757
rect 509485 643727 509491 643779
rect 507865 643715 508012 643727
rect 509108 643715 509491 643727
rect 507865 643663 507871 643715
rect 507923 643663 508012 643715
rect 509108 643663 509433 643715
rect 509485 643663 509491 643715
rect 507865 643651 508012 643663
rect 509108 643651 509491 643663
rect 507865 643599 507871 643651
rect 507923 643621 508012 643651
rect 509108 643621 509433 643651
rect 507923 643609 508059 643621
rect 507923 643599 507929 643609
rect 507865 643593 507929 643599
rect 508053 643599 508059 643609
rect 508111 643609 508517 643621
rect 508111 643599 508117 643609
rect 508053 643593 508117 643599
rect 508511 643599 508517 643609
rect 508569 643609 509433 643621
rect 508569 643599 508575 643609
rect 508511 643593 508575 643599
rect 509427 643599 509433 643609
rect 509485 643599 509491 643651
rect 509427 643593 509491 643599
rect 510338 643741 510347 643797
rect 510403 643769 510412 643797
rect 513086 643797 513160 643806
rect 511259 643779 511323 643785
rect 511259 643769 511265 643779
rect 510403 643741 511265 643769
rect 510338 643727 510349 643741
rect 510401 643727 511265 643741
rect 511317 643727 511323 643779
rect 510338 643717 511323 643727
rect 510338 643661 510347 643717
rect 510403 643715 511323 643717
rect 510403 643663 511265 643715
rect 511317 643663 511323 643715
rect 510403 643661 511323 643663
rect 510338 643651 511323 643661
rect 510338 643637 510349 643651
rect 510401 643637 511265 643651
rect 510338 643581 510347 643637
rect 510403 643609 511265 643637
rect 510403 643581 510412 643609
rect 511259 643599 511265 643609
rect 511317 643599 511323 643651
rect 511259 643593 511323 643599
rect 512175 643779 512239 643785
rect 512175 643727 512181 643779
rect 512233 643769 512239 643779
rect 513086 643769 513095 643797
rect 512233 643741 513095 643769
rect 513151 643741 513160 643797
rect 515532 643805 515670 643820
rect 512233 643727 513097 643741
rect 513149 643727 513160 643741
rect 512175 643717 513160 643727
rect 512175 643715 513095 643717
rect 512175 643663 512181 643715
rect 512233 643663 513095 643715
rect 512175 643661 513095 643663
rect 513151 643661 513160 643717
rect 512175 643651 513160 643661
rect 512175 643599 512181 643651
rect 512233 643637 513097 643651
rect 513149 643637 513160 643651
rect 512233 643609 513095 643637
rect 512233 643599 512239 643609
rect 512175 643593 512239 643599
rect 510338 643572 510412 643581
rect 513086 643581 513095 643609
rect 513151 643581 513160 643637
rect 514007 643779 514071 643785
rect 514007 643727 514013 643779
rect 514065 643769 514071 643779
rect 514465 643779 514529 643785
rect 514465 643769 514471 643779
rect 514065 643727 514471 643769
rect 514523 643769 514529 643779
rect 514923 643779 514987 643785
rect 514923 643769 514929 643779
rect 514523 643727 514929 643769
rect 514981 643769 514987 643779
rect 515381 643779 515445 643785
rect 515381 643769 515387 643779
rect 514981 643727 515387 643769
rect 515439 643769 515445 643779
rect 515532 643769 515572 643805
rect 515439 643749 515572 643769
rect 515628 643749 515670 643805
rect 515439 643727 515575 643749
rect 515627 643727 515670 643749
rect 514007 643725 515670 643727
rect 514007 643715 515572 643725
rect 514007 643663 514013 643715
rect 514065 643663 514471 643715
rect 514523 643663 514929 643715
rect 514981 643663 515387 643715
rect 515439 643669 515572 643715
rect 515628 643669 515670 643725
rect 515439 643663 515575 643669
rect 515627 643663 515670 643669
rect 514007 643651 515670 643663
rect 514007 643599 514013 643651
rect 514065 643609 514471 643651
rect 514065 643599 514071 643609
rect 514007 643593 514071 643599
rect 514465 643599 514471 643609
rect 514523 643609 514929 643651
rect 514523 643599 514529 643609
rect 514465 643593 514529 643599
rect 514923 643599 514929 643609
rect 514981 643609 515387 643651
rect 514981 643599 514987 643609
rect 514923 643593 514987 643599
rect 515381 643599 515387 643609
rect 515439 643645 515575 643651
rect 515627 643645 515670 643651
rect 515439 643609 515572 643645
rect 515439 643599 515445 643609
rect 515381 643593 515445 643599
rect 513086 643572 513160 643581
rect 515532 643589 515572 643609
rect 515628 643589 515670 643645
rect 515532 643574 515670 643589
rect 507733 643331 507887 643340
rect 507733 643195 507742 643331
rect 507878 643314 507887 643331
rect 507878 643290 509129 643314
rect 516426 643305 516526 644323
rect 516668 644385 516677 644441
rect 516733 644385 516742 644441
rect 516668 644379 516679 644385
rect 516731 644379 516742 644385
rect 516668 644367 516742 644379
rect 516668 644361 516679 644367
rect 516731 644361 516742 644367
rect 516668 644305 516677 644361
rect 516733 644305 516742 644361
rect 516668 644303 516742 644305
rect 516668 644281 516679 644303
rect 516731 644281 516742 644303
rect 516668 644225 516677 644281
rect 516733 644225 516742 644281
rect 516668 644201 516679 644225
rect 516731 644201 516742 644225
rect 516668 644145 516677 644201
rect 516733 644145 516742 644201
rect 516668 644136 516742 644145
rect 507878 643238 508879 643290
rect 508931 643238 508943 643290
rect 508995 643238 509007 643290
rect 509059 643238 509071 643290
rect 509123 643238 509129 643290
rect 507878 643214 509129 643238
rect 510676 643292 510990 643301
rect 510676 643236 510685 643292
rect 510741 643290 510765 643292
rect 510821 643290 510845 643292
rect 510901 643290 510925 643292
rect 510763 643238 510765 643290
rect 510827 643238 510839 643290
rect 510901 643238 510903 643290
rect 510741 643236 510765 643238
rect 510821 643236 510845 643238
rect 510901 643236 510925 643238
rect 510981 643236 510990 643292
rect 510676 643227 510990 643236
rect 512508 643292 512822 643301
rect 512508 643236 512517 643292
rect 512573 643290 512597 643292
rect 512653 643290 512677 643292
rect 512733 643290 512757 643292
rect 512595 643238 512597 643290
rect 512659 643238 512671 643290
rect 512733 643238 512735 643290
rect 512573 643236 512597 643238
rect 512653 643236 512677 643238
rect 512733 643236 512757 643238
rect 512813 643236 512822 643292
rect 516348 643299 516604 643305
rect 516348 643247 516354 643299
rect 516406 643247 516418 643299
rect 516470 643247 516482 643299
rect 516534 643247 516546 643299
rect 516598 643247 516604 643299
rect 516348 643241 516604 643247
rect 512508 643227 512822 643236
rect 507878 643195 507887 643214
rect 507733 643186 507887 643195
rect 512589 643058 512743 643067
rect 512589 643040 512598 643058
rect 507669 642940 512598 643040
rect 512589 642922 512598 642940
rect 512734 642922 512743 643058
rect 512589 642913 512743 642922
rect 513505 642918 513659 642927
rect 510756 642823 510910 642832
rect 510756 642805 510765 642823
rect 507669 642705 510765 642805
rect 510756 642687 510765 642705
rect 510901 642687 510910 642823
rect 513505 642782 513514 642918
rect 513650 642900 513659 642918
rect 513962 642918 514116 642927
rect 513962 642900 513971 642918
rect 513650 642800 513971 642900
rect 513650 642782 513659 642800
rect 513505 642773 513659 642782
rect 513962 642782 513971 642800
rect 514107 642900 514116 642918
rect 515954 642908 516082 642914
rect 515954 642900 515960 642908
rect 514107 642800 515960 642900
rect 514107 642782 514116 642800
rect 515954 642792 515960 642800
rect 516076 642792 516082 642908
rect 515954 642786 516082 642792
rect 513962 642773 514116 642782
rect 510756 642678 510910 642687
rect 509186 642536 509340 642545
rect 509186 642519 509195 642536
rect 507669 642495 509195 642519
rect 507669 642443 508879 642495
rect 508931 642443 508943 642495
rect 508995 642443 509007 642495
rect 509059 642443 509071 642495
rect 509123 642443 509195 642495
rect 507669 642419 509195 642443
rect 509186 642400 509195 642419
rect 509331 642400 509340 642536
rect 510676 642497 510990 642506
rect 510676 642441 510685 642497
rect 510741 642495 510765 642497
rect 510821 642495 510845 642497
rect 510901 642495 510925 642497
rect 510763 642443 510765 642495
rect 510827 642443 510839 642495
rect 510901 642443 510903 642495
rect 510741 642441 510765 642443
rect 510821 642441 510845 642443
rect 510901 642441 510925 642443
rect 510981 642441 510990 642497
rect 510676 642432 510990 642441
rect 512508 642497 512822 642506
rect 512508 642441 512517 642497
rect 512573 642495 512597 642497
rect 512653 642495 512677 642497
rect 512733 642495 512757 642497
rect 512595 642443 512597 642495
rect 512659 642443 512671 642495
rect 512733 642443 512735 642495
rect 512573 642441 512597 642443
rect 512653 642441 512677 642443
rect 512733 642441 512757 642443
rect 512813 642441 512822 642497
rect 516426 642492 516526 643241
rect 516628 642925 516782 642934
rect 516628 642789 516637 642925
rect 516773 642907 516782 642925
rect 516773 642807 517124 642907
rect 516773 642789 516782 642807
rect 516628 642780 516782 642789
rect 512508 642432 512822 642441
rect 516347 642486 516603 642492
rect 516347 642434 516353 642486
rect 516405 642434 516417 642486
rect 516469 642434 516481 642486
rect 516533 642434 516545 642486
rect 516597 642434 516603 642486
rect 516347 642428 516603 642434
rect 509186 642391 509340 642400
rect 515757 642243 515821 642249
rect 515757 642191 515763 642243
rect 515815 642191 515821 642243
rect 515757 642179 515821 642191
rect 511254 642161 511328 642170
rect 507865 642143 507929 642149
rect 507865 642091 507871 642143
rect 507923 642133 507929 642143
rect 508053 642143 508117 642149
rect 508053 642133 508059 642143
rect 507923 642091 508059 642133
rect 508111 642133 508117 642143
rect 508511 642143 508575 642149
rect 508511 642133 508517 642143
rect 508111 642091 508517 642133
rect 508569 642133 508575 642143
rect 509427 642143 509491 642149
rect 509427 642133 509433 642143
rect 508569 642091 509433 642133
rect 509485 642091 509491 642143
rect 507865 642079 509491 642091
rect 507865 642027 507871 642079
rect 507923 642027 508059 642079
rect 508111 642027 508517 642079
rect 508569 642027 509433 642079
rect 509485 642027 509491 642079
rect 507865 642015 509491 642027
rect 507865 641963 507871 642015
rect 507923 641973 508059 642015
rect 507923 641963 507929 641973
rect 507865 641957 507929 641963
rect 508053 641963 508059 641973
rect 508111 641973 508517 642015
rect 508111 641963 508117 641973
rect 508053 641957 508117 641963
rect 508511 641963 508517 641973
rect 508569 641973 509433 642015
rect 508569 641963 508575 641973
rect 508511 641957 508575 641963
rect 509427 641963 509433 641973
rect 509485 641963 509491 642015
rect 509427 641957 509491 641963
rect 510343 642143 510407 642149
rect 510343 642091 510349 642143
rect 510401 642133 510407 642143
rect 511254 642133 511263 642161
rect 510401 642105 511263 642133
rect 511319 642105 511328 642161
rect 510401 642091 511265 642105
rect 511317 642091 511328 642105
rect 510343 642081 511328 642091
rect 510343 642079 511263 642081
rect 510343 642027 510349 642079
rect 510401 642027 511263 642079
rect 510343 642025 511263 642027
rect 511319 642025 511328 642081
rect 510343 642015 511328 642025
rect 510343 641963 510349 642015
rect 510401 642001 511265 642015
rect 511317 642001 511328 642015
rect 510401 641973 511263 642001
rect 510401 641963 510407 641973
rect 510343 641957 510407 641963
rect 511254 641945 511263 641973
rect 511319 641945 511328 642001
rect 511254 641936 511328 641945
rect 512170 642161 512244 642170
rect 512170 642105 512179 642161
rect 512235 642133 512244 642161
rect 513091 642143 513155 642149
rect 513091 642133 513097 642143
rect 512235 642105 513097 642133
rect 512170 642091 512181 642105
rect 512233 642091 513097 642105
rect 513149 642091 513155 642143
rect 512170 642081 513155 642091
rect 512170 642025 512179 642081
rect 512235 642079 513155 642081
rect 512235 642027 513097 642079
rect 513149 642027 513155 642079
rect 512235 642025 513155 642027
rect 512170 642015 513155 642025
rect 512170 642001 512181 642015
rect 512233 642001 513097 642015
rect 512170 641945 512179 642001
rect 512235 641973 513097 642001
rect 512235 641945 512244 641973
rect 513091 641963 513097 641973
rect 513149 641963 513155 642015
rect 513091 641957 513155 641963
rect 514007 642143 514071 642149
rect 514007 642091 514013 642143
rect 514065 642133 514071 642143
rect 514465 642143 514529 642149
rect 514465 642133 514471 642143
rect 514065 642121 514471 642133
rect 514523 642133 514529 642143
rect 514923 642143 514987 642149
rect 514923 642133 514929 642143
rect 514523 642121 514929 642133
rect 514981 642133 514987 642143
rect 515381 642143 515445 642149
rect 515381 642133 515387 642143
rect 514981 642121 515387 642133
rect 514065 642091 514335 642121
rect 515351 642091 515387 642121
rect 515439 642133 515445 642143
rect 515569 642143 515633 642149
rect 515569 642133 515575 642143
rect 515439 642091 515575 642133
rect 515627 642091 515633 642143
rect 514007 642079 514335 642091
rect 515351 642079 515633 642091
rect 514007 642027 514013 642079
rect 514065 642027 514335 642079
rect 515351 642027 515387 642079
rect 515439 642027 515575 642079
rect 515627 642027 515633 642079
rect 514007 642015 514335 642027
rect 515351 642015 515633 642027
rect 514007 641963 514013 642015
rect 514065 641985 514335 642015
rect 515351 641985 515387 642015
rect 514065 641973 514471 641985
rect 514065 641963 514071 641973
rect 514007 641957 514071 641963
rect 514465 641963 514471 641973
rect 514523 641973 514929 641985
rect 514523 641963 514529 641973
rect 514465 641957 514529 641963
rect 514923 641963 514929 641973
rect 514981 641973 515387 641985
rect 514981 641963 514987 641973
rect 514923 641957 514987 641963
rect 515381 641963 515387 641973
rect 515439 641973 515575 642015
rect 515439 641963 515445 641973
rect 515381 641957 515445 641963
rect 515569 641963 515575 641973
rect 515627 641963 515633 642015
rect 515569 641957 515633 641963
rect 515757 642127 515763 642179
rect 515815 642127 515821 642179
rect 515757 642115 515821 642127
rect 515757 642063 515763 642115
rect 515815 642107 515821 642115
rect 516426 642107 516526 642428
rect 515815 642063 516526 642107
rect 515757 642051 516526 642063
rect 515757 641999 515763 642051
rect 515815 642007 516526 642051
rect 516668 642285 516742 642294
rect 516668 642229 516677 642285
rect 516733 642229 516742 642285
rect 516668 642205 516679 642229
rect 516731 642205 516742 642229
rect 516668 642149 516677 642205
rect 516733 642149 516742 642205
rect 516668 642127 516679 642149
rect 516731 642127 516742 642149
rect 516668 642125 516742 642127
rect 516668 642069 516677 642125
rect 516733 642069 516742 642125
rect 516668 642063 516679 642069
rect 516731 642063 516742 642069
rect 516668 642051 516742 642063
rect 516668 642045 516679 642051
rect 516731 642045 516742 642051
rect 515815 641999 515821 642007
rect 515757 641987 515821 641999
rect 512170 641936 512244 641945
rect 515757 641935 515763 641987
rect 515815 641935 515821 641987
rect 515757 641923 515821 641935
rect 515757 641871 515763 641923
rect 515815 641871 515821 641923
rect 515757 641865 515821 641871
rect 516668 641989 516677 642045
rect 516733 641989 516742 642045
rect 516668 641987 516742 641989
rect 516668 641965 516679 641987
rect 516731 641965 516742 641987
rect 516668 641909 516677 641965
rect 516733 641909 516742 641965
rect 516668 641885 516679 641909
rect 516731 641885 516742 641909
rect 516668 641829 516677 641885
rect 516733 641829 516742 641885
rect 516668 641820 516742 641829
rect 516197 641791 516297 641797
rect 516197 641739 516221 641791
rect 516273 641739 516297 641791
rect 516197 641727 516297 641739
rect 508969 641678 509033 641684
rect 508969 641626 508975 641678
rect 509027 641668 509033 641678
rect 509885 641678 509949 641684
rect 509885 641668 509891 641678
rect 509027 641626 509891 641668
rect 509943 641668 509949 641678
rect 510801 641678 510865 641684
rect 510801 641668 510807 641678
rect 509943 641626 510807 641668
rect 510859 641668 510865 641678
rect 511717 641678 511781 641684
rect 511717 641668 511723 641678
rect 510859 641626 511723 641668
rect 511775 641668 511781 641678
rect 512633 641678 512697 641684
rect 512633 641668 512639 641678
rect 511775 641626 512639 641668
rect 512691 641668 512697 641678
rect 513549 641678 513613 641684
rect 513549 641668 513555 641678
rect 512691 641626 513555 641668
rect 513607 641626 513613 641678
rect 508969 641614 513613 641626
rect 508969 641562 508975 641614
rect 509027 641562 509891 641614
rect 509943 641562 510807 641614
rect 510859 641562 511723 641614
rect 511775 641562 512639 641614
rect 512691 641562 513555 641614
rect 513607 641562 513613 641614
rect 508969 641550 513613 641562
rect 508969 641498 508975 641550
rect 509027 641508 509891 641550
rect 509027 641498 509033 641508
rect 508969 641492 509033 641498
rect 509885 641498 509891 641508
rect 509943 641508 510807 641550
rect 509943 641498 509949 641508
rect 509885 641492 509949 641498
rect 510801 641498 510807 641508
rect 510859 641508 511723 641550
rect 510859 641498 510865 641508
rect 510801 641492 510865 641498
rect 511717 641498 511723 641508
rect 511775 641508 512639 641550
rect 511775 641498 511781 641508
rect 511717 641492 511781 641498
rect 512633 641498 512639 641508
rect 512691 641508 513555 641550
rect 512691 641498 512697 641508
rect 512633 641492 512697 641498
rect 513549 641498 513555 641508
rect 513607 641498 513613 641550
rect 513549 641492 513613 641498
rect 516197 641675 516221 641727
rect 516273 641675 516297 641727
rect 516197 641663 516297 641675
rect 516197 641611 516221 641663
rect 516273 641611 516297 641663
rect 516197 641599 516297 641611
rect 516197 641547 516221 641599
rect 516273 641547 516297 641599
rect 516197 641535 516297 641547
rect 516197 641483 516221 641535
rect 516273 641483 516297 641535
rect 509422 641206 509496 641215
rect 509422 641150 509431 641206
rect 509487 641150 509496 641206
rect 509422 641136 509433 641150
rect 509485 641136 509496 641150
rect 509422 641126 509496 641136
rect 509422 641070 509431 641126
rect 509487 641070 509496 641126
rect 509422 641060 509496 641070
rect 509422 641046 509433 641060
rect 509485 641046 509496 641060
rect 509422 640990 509431 641046
rect 509487 640990 509496 641046
rect 509422 640981 509496 640990
rect 510338 641206 510412 641215
rect 510338 641150 510347 641206
rect 510403 641150 510412 641206
rect 510338 641136 510349 641150
rect 510401 641136 510412 641150
rect 510338 641126 510412 641136
rect 510338 641070 510347 641126
rect 510403 641070 510412 641126
rect 510338 641060 510412 641070
rect 510338 641046 510349 641060
rect 510401 641046 510412 641060
rect 510338 640990 510347 641046
rect 510403 640990 510412 641046
rect 510338 640981 510412 640990
rect 513086 641206 513160 641215
rect 513086 641150 513095 641206
rect 513151 641150 513160 641206
rect 513086 641136 513097 641150
rect 513149 641136 513160 641150
rect 513086 641126 513160 641136
rect 513086 641070 513095 641126
rect 513151 641070 513160 641126
rect 513086 641060 513160 641070
rect 513086 641046 513097 641060
rect 513149 641046 513160 641060
rect 513086 640990 513095 641046
rect 513151 640990 513160 641046
rect 513086 640981 513160 640990
rect 514002 641206 514076 641215
rect 514002 641150 514011 641206
rect 514067 641150 514076 641206
rect 514002 641136 514013 641150
rect 514065 641136 514076 641150
rect 514002 641126 514076 641136
rect 514002 641070 514011 641126
rect 514067 641070 514076 641126
rect 514002 641060 514076 641070
rect 514002 641046 514013 641060
rect 514065 641046 514076 641060
rect 514002 640990 514011 641046
rect 514067 640990 514076 641046
rect 514002 640981 514076 640990
rect 509880 640852 509954 640861
rect 509880 640796 509889 640852
rect 509945 640796 509954 640852
rect 513544 640852 513618 640861
rect 509880 640794 509954 640796
rect 511259 640834 511323 640840
rect 511259 640794 511265 640834
rect 509880 640782 511265 640794
rect 511317 640782 511323 640834
rect 509880 640772 511323 640782
rect 509880 640716 509889 640772
rect 509945 640770 511323 640772
rect 509945 640718 511265 640770
rect 511317 640718 511323 640770
rect 509945 640716 511323 640718
rect 509880 640706 511323 640716
rect 509880 640694 511265 640706
rect 509880 640692 509954 640694
rect 509880 640636 509889 640692
rect 509945 640636 509954 640692
rect 511259 640654 511265 640694
rect 511317 640654 511323 640706
rect 511259 640648 511323 640654
rect 512175 640834 512239 640840
rect 512175 640782 512181 640834
rect 512233 640794 512239 640834
rect 513544 640796 513553 640852
rect 513609 640796 513618 640852
rect 513544 640794 513618 640796
rect 512233 640782 513618 640794
rect 512175 640772 513618 640782
rect 512175 640770 513553 640772
rect 512175 640718 512181 640770
rect 512233 640718 513553 640770
rect 512175 640716 513553 640718
rect 513609 640716 513618 640772
rect 512175 640706 513618 640716
rect 512175 640654 512181 640706
rect 512233 640694 513618 640706
rect 512233 640654 512239 640694
rect 512175 640648 512239 640654
rect 513544 640692 513618 640694
rect 509880 640627 509954 640636
rect 513544 640636 513553 640692
rect 513609 640636 513618 640692
rect 513544 640627 513618 640636
rect 507864 640503 507928 640509
rect 507864 640451 507870 640503
rect 507922 640493 507928 640503
rect 508053 640503 508117 640509
rect 508053 640493 508059 640503
rect 507922 640451 508059 640493
rect 508111 640493 508117 640503
rect 508511 640503 508575 640509
rect 508511 640493 508517 640503
rect 508111 640451 508517 640493
rect 508569 640493 508575 640503
rect 508969 640503 509033 640509
rect 508969 640493 508975 640503
rect 508569 640451 508975 640493
rect 509027 640493 509033 640503
rect 509885 640503 509949 640509
rect 509885 640493 509891 640503
rect 509027 640451 509891 640493
rect 509943 640493 509949 640503
rect 510801 640503 510865 640509
rect 510801 640493 510807 640503
rect 509943 640451 510807 640493
rect 510859 640493 510865 640503
rect 511717 640503 511781 640509
rect 511717 640493 511723 640503
rect 510859 640451 511723 640493
rect 511775 640493 511781 640503
rect 512633 640503 512697 640509
rect 512633 640493 512639 640503
rect 511775 640451 512639 640493
rect 512691 640493 512697 640503
rect 513549 640503 513613 640509
rect 513549 640493 513555 640503
rect 512691 640481 513555 640493
rect 513607 640493 513613 640503
rect 514465 640503 514529 640509
rect 514465 640493 514471 640503
rect 513607 640481 514471 640493
rect 512691 640451 512724 640481
rect 514300 640451 514471 640481
rect 514523 640493 514529 640503
rect 514923 640503 514987 640509
rect 514923 640493 514929 640503
rect 514523 640451 514929 640493
rect 514981 640493 514987 640503
rect 515381 640503 515445 640509
rect 515381 640493 515387 640503
rect 514981 640451 515387 640493
rect 515439 640493 515445 640503
rect 515655 640503 516039 640509
rect 515655 640493 515661 640503
rect 515439 640451 515661 640493
rect 507864 640439 512724 640451
rect 514300 640439 515661 640451
rect 507864 640387 507870 640439
rect 507922 640387 508059 640439
rect 508111 640387 508517 640439
rect 508569 640387 508975 640439
rect 509027 640387 509891 640439
rect 509943 640387 510807 640439
rect 510859 640387 511723 640439
rect 511775 640387 512639 640439
rect 512691 640387 512724 640439
rect 514300 640387 514471 640439
rect 514523 640387 514929 640439
rect 514981 640387 515387 640439
rect 515439 640387 515661 640439
rect 507864 640375 512724 640387
rect 514300 640375 515661 640387
rect 507864 640323 507870 640375
rect 507922 640333 508059 640375
rect 507922 640323 507928 640333
rect 507864 640317 507928 640323
rect 508053 640323 508059 640333
rect 508111 640333 508517 640375
rect 508111 640323 508117 640333
rect 508053 640317 508117 640323
rect 508511 640323 508517 640333
rect 508569 640333 508975 640375
rect 508569 640323 508575 640333
rect 508511 640317 508575 640323
rect 508969 640323 508975 640333
rect 509027 640333 509891 640375
rect 509027 640323 509033 640333
rect 508969 640317 509033 640323
rect 509885 640323 509891 640333
rect 509943 640333 510807 640375
rect 509943 640323 509949 640333
rect 509885 640317 509949 640323
rect 510801 640323 510807 640333
rect 510859 640333 511723 640375
rect 510859 640323 510865 640333
rect 510801 640317 510865 640323
rect 511717 640323 511723 640333
rect 511775 640333 512639 640375
rect 511775 640323 511781 640333
rect 511717 640317 511781 640323
rect 512633 640323 512639 640333
rect 512691 640345 512724 640375
rect 514300 640345 514471 640375
rect 512691 640333 513555 640345
rect 512691 640323 512697 640333
rect 512633 640317 512697 640323
rect 513549 640323 513555 640333
rect 513607 640333 514471 640345
rect 513607 640323 513613 640333
rect 513549 640317 513613 640323
rect 514465 640323 514471 640333
rect 514523 640333 514929 640375
rect 514523 640323 514529 640333
rect 514465 640317 514529 640323
rect 514923 640323 514929 640333
rect 514981 640333 515387 640375
rect 514981 640323 514987 640333
rect 514923 640317 514987 640323
rect 515381 640323 515387 640333
rect 515439 640333 515661 640375
rect 515439 640323 515445 640333
rect 515381 640317 515445 640323
rect 515655 640323 515661 640333
rect 516033 640463 516039 640503
rect 516197 640463 516297 641483
rect 516033 640363 516297 640463
rect 516033 640323 516039 640363
rect 515655 640317 516039 640323
<< via2 >>
rect 509001 645359 509027 645389
rect 509027 645359 509891 645389
rect 509891 645359 509943 645389
rect 509943 645359 510577 645389
rect 515572 645411 515628 645438
rect 515572 645382 515576 645411
rect 515576 645382 515628 645411
rect 509001 645347 510577 645359
rect 515572 645347 515628 645358
rect 509001 645295 509027 645347
rect 509027 645295 509891 645347
rect 509891 645295 509943 645347
rect 509943 645295 510577 645347
rect 515572 645302 515576 645347
rect 515576 645302 515628 645347
rect 509001 645283 510577 645295
rect 509001 645253 509027 645283
rect 509027 645253 509891 645283
rect 509891 645253 509943 645283
rect 509943 645253 510577 645283
rect 515572 645231 515576 645278
rect 515576 645231 515628 645278
rect 515572 645222 515628 645231
rect 509431 645050 509487 645106
rect 509431 644970 509487 645026
rect 509431 644890 509487 644946
rect 514011 645050 514067 645106
rect 514011 644970 514067 645026
rect 514011 644890 514067 644946
rect 509889 644738 509945 644794
rect 509889 644658 509945 644714
rect 509889 644578 509945 644634
rect 511263 644738 511319 644794
rect 511263 644658 511319 644714
rect 511263 644578 511319 644634
rect 512179 644738 512235 644794
rect 512179 644658 512235 644714
rect 512179 644578 512235 644634
rect 513553 644738 513609 644794
rect 513553 644658 513609 644714
rect 513553 644578 513609 644634
rect 516677 644559 516733 644601
rect 516677 644545 516679 644559
rect 516679 644545 516731 644559
rect 516731 644545 516733 644559
rect 516677 644507 516679 644521
rect 516679 644507 516731 644521
rect 516731 644507 516733 644521
rect 516677 644495 516733 644507
rect 516677 644465 516679 644495
rect 516679 644465 516731 644495
rect 516731 644465 516733 644495
rect 508012 643727 508059 643757
rect 508059 643727 508111 643757
rect 508111 643727 508517 643757
rect 508517 643727 508569 643757
rect 508569 643727 509108 643757
rect 508012 643715 509108 643727
rect 508012 643663 508059 643715
rect 508059 643663 508111 643715
rect 508111 643663 508517 643715
rect 508517 643663 508569 643715
rect 508569 643663 509108 643715
rect 508012 643651 509108 643663
rect 508012 643621 508059 643651
rect 508059 643621 508111 643651
rect 508111 643621 508517 643651
rect 508517 643621 508569 643651
rect 508569 643621 509108 643651
rect 510347 643779 510403 643797
rect 510347 643741 510349 643779
rect 510349 643741 510401 643779
rect 510401 643741 510403 643779
rect 510347 643715 510403 643717
rect 510347 643663 510349 643715
rect 510349 643663 510401 643715
rect 510401 643663 510403 643715
rect 510347 643661 510403 643663
rect 510347 643599 510349 643637
rect 510349 643599 510401 643637
rect 510401 643599 510403 643637
rect 510347 643581 510403 643599
rect 513095 643779 513151 643797
rect 513095 643741 513097 643779
rect 513097 643741 513149 643779
rect 513149 643741 513151 643779
rect 513095 643715 513151 643717
rect 513095 643663 513097 643715
rect 513097 643663 513149 643715
rect 513149 643663 513151 643715
rect 513095 643661 513151 643663
rect 513095 643599 513097 643637
rect 513097 643599 513149 643637
rect 513149 643599 513151 643637
rect 513095 643581 513151 643599
rect 515572 643779 515628 643805
rect 515572 643749 515575 643779
rect 515575 643749 515627 643779
rect 515627 643749 515628 643779
rect 515572 643715 515628 643725
rect 515572 643669 515575 643715
rect 515575 643669 515627 643715
rect 515627 643669 515628 643715
rect 515572 643599 515575 643645
rect 515575 643599 515627 643645
rect 515627 643599 515628 643645
rect 515572 643589 515628 643599
rect 507742 643195 507878 643331
rect 516677 644431 516733 644441
rect 516677 644385 516679 644431
rect 516679 644385 516731 644431
rect 516731 644385 516733 644431
rect 516677 644315 516679 644361
rect 516679 644315 516731 644361
rect 516731 644315 516733 644361
rect 516677 644305 516733 644315
rect 516677 644251 516679 644281
rect 516679 644251 516731 644281
rect 516731 644251 516733 644281
rect 516677 644239 516733 644251
rect 516677 644225 516679 644239
rect 516679 644225 516731 644239
rect 516731 644225 516733 644239
rect 516677 644187 516679 644201
rect 516679 644187 516731 644201
rect 516731 644187 516733 644201
rect 516677 644145 516733 644187
rect 510685 643290 510741 643292
rect 510765 643290 510821 643292
rect 510845 643290 510901 643292
rect 510925 643290 510981 643292
rect 510685 643238 510711 643290
rect 510711 643238 510741 643290
rect 510765 643238 510775 643290
rect 510775 643238 510821 643290
rect 510845 643238 510891 643290
rect 510891 643238 510901 643290
rect 510925 643238 510955 643290
rect 510955 643238 510981 643290
rect 510685 643236 510741 643238
rect 510765 643236 510821 643238
rect 510845 643236 510901 643238
rect 510925 643236 510981 643238
rect 512517 643290 512573 643292
rect 512597 643290 512653 643292
rect 512677 643290 512733 643292
rect 512757 643290 512813 643292
rect 512517 643238 512543 643290
rect 512543 643238 512573 643290
rect 512597 643238 512607 643290
rect 512607 643238 512653 643290
rect 512677 643238 512723 643290
rect 512723 643238 512733 643290
rect 512757 643238 512787 643290
rect 512787 643238 512813 643290
rect 512517 643236 512573 643238
rect 512597 643236 512653 643238
rect 512677 643236 512733 643238
rect 512757 643236 512813 643238
rect 512598 642922 512734 643058
rect 510765 642687 510901 642823
rect 513514 642782 513650 642918
rect 513971 642782 514107 642918
rect 509195 642400 509331 642536
rect 510685 642495 510741 642497
rect 510765 642495 510821 642497
rect 510845 642495 510901 642497
rect 510925 642495 510981 642497
rect 510685 642443 510711 642495
rect 510711 642443 510741 642495
rect 510765 642443 510775 642495
rect 510775 642443 510821 642495
rect 510845 642443 510891 642495
rect 510891 642443 510901 642495
rect 510925 642443 510955 642495
rect 510955 642443 510981 642495
rect 510685 642441 510741 642443
rect 510765 642441 510821 642443
rect 510845 642441 510901 642443
rect 510925 642441 510981 642443
rect 512517 642495 512573 642497
rect 512597 642495 512653 642497
rect 512677 642495 512733 642497
rect 512757 642495 512813 642497
rect 512517 642443 512543 642495
rect 512543 642443 512573 642495
rect 512597 642443 512607 642495
rect 512607 642443 512653 642495
rect 512677 642443 512723 642495
rect 512723 642443 512733 642495
rect 512757 642443 512787 642495
rect 512787 642443 512813 642495
rect 512517 642441 512573 642443
rect 512597 642441 512653 642443
rect 512677 642441 512733 642443
rect 512757 642441 512813 642443
rect 516637 642789 516773 642925
rect 511263 642143 511319 642161
rect 511263 642105 511265 642143
rect 511265 642105 511317 642143
rect 511317 642105 511319 642143
rect 511263 642079 511319 642081
rect 511263 642027 511265 642079
rect 511265 642027 511317 642079
rect 511317 642027 511319 642079
rect 511263 642025 511319 642027
rect 511263 641963 511265 642001
rect 511265 641963 511317 642001
rect 511317 641963 511319 642001
rect 511263 641945 511319 641963
rect 512179 642143 512235 642161
rect 512179 642105 512181 642143
rect 512181 642105 512233 642143
rect 512233 642105 512235 642143
rect 512179 642079 512235 642081
rect 512179 642027 512181 642079
rect 512181 642027 512233 642079
rect 512233 642027 512235 642079
rect 512179 642025 512235 642027
rect 512179 641963 512181 642001
rect 512181 641963 512233 642001
rect 512233 641963 512235 642001
rect 512179 641945 512235 641963
rect 514335 642091 514471 642121
rect 514471 642091 514523 642121
rect 514523 642091 514929 642121
rect 514929 642091 514981 642121
rect 514981 642091 515351 642121
rect 514335 642079 515351 642091
rect 514335 642027 514471 642079
rect 514471 642027 514523 642079
rect 514523 642027 514929 642079
rect 514929 642027 514981 642079
rect 514981 642027 515351 642079
rect 514335 642015 515351 642027
rect 514335 641985 514471 642015
rect 514471 641985 514523 642015
rect 514523 641985 514929 642015
rect 514929 641985 514981 642015
rect 514981 641985 515351 642015
rect 516677 642243 516733 642285
rect 516677 642229 516679 642243
rect 516679 642229 516731 642243
rect 516731 642229 516733 642243
rect 516677 642191 516679 642205
rect 516679 642191 516731 642205
rect 516731 642191 516733 642205
rect 516677 642179 516733 642191
rect 516677 642149 516679 642179
rect 516679 642149 516731 642179
rect 516731 642149 516733 642179
rect 516677 642115 516733 642125
rect 516677 642069 516679 642115
rect 516679 642069 516731 642115
rect 516731 642069 516733 642115
rect 516677 641999 516679 642045
rect 516679 641999 516731 642045
rect 516731 641999 516733 642045
rect 516677 641989 516733 641999
rect 516677 641935 516679 641965
rect 516679 641935 516731 641965
rect 516731 641935 516733 641965
rect 516677 641923 516733 641935
rect 516677 641909 516679 641923
rect 516679 641909 516731 641923
rect 516731 641909 516733 641923
rect 516677 641871 516679 641885
rect 516679 641871 516731 641885
rect 516731 641871 516733 641885
rect 516677 641829 516733 641871
rect 509431 641188 509487 641206
rect 509431 641150 509433 641188
rect 509433 641150 509485 641188
rect 509485 641150 509487 641188
rect 509431 641124 509487 641126
rect 509431 641072 509433 641124
rect 509433 641072 509485 641124
rect 509485 641072 509487 641124
rect 509431 641070 509487 641072
rect 509431 641008 509433 641046
rect 509433 641008 509485 641046
rect 509485 641008 509487 641046
rect 509431 640990 509487 641008
rect 510347 641188 510403 641206
rect 510347 641150 510349 641188
rect 510349 641150 510401 641188
rect 510401 641150 510403 641188
rect 510347 641124 510403 641126
rect 510347 641072 510349 641124
rect 510349 641072 510401 641124
rect 510401 641072 510403 641124
rect 510347 641070 510403 641072
rect 510347 641008 510349 641046
rect 510349 641008 510401 641046
rect 510401 641008 510403 641046
rect 510347 640990 510403 641008
rect 513095 641188 513151 641206
rect 513095 641150 513097 641188
rect 513097 641150 513149 641188
rect 513149 641150 513151 641188
rect 513095 641124 513151 641126
rect 513095 641072 513097 641124
rect 513097 641072 513149 641124
rect 513149 641072 513151 641124
rect 513095 641070 513151 641072
rect 513095 641008 513097 641046
rect 513097 641008 513149 641046
rect 513149 641008 513151 641046
rect 513095 640990 513151 641008
rect 514011 641188 514067 641206
rect 514011 641150 514013 641188
rect 514013 641150 514065 641188
rect 514065 641150 514067 641188
rect 514011 641124 514067 641126
rect 514011 641072 514013 641124
rect 514013 641072 514065 641124
rect 514065 641072 514067 641124
rect 514011 641070 514067 641072
rect 514011 641008 514013 641046
rect 514013 641008 514065 641046
rect 514065 641008 514067 641046
rect 514011 640990 514067 641008
rect 509889 640796 509945 640852
rect 509889 640716 509945 640772
rect 509889 640636 509945 640692
rect 513553 640796 513609 640852
rect 513553 640716 513609 640772
rect 513553 640636 513609 640692
rect 512724 640451 513555 640481
rect 513555 640451 513607 640481
rect 513607 640451 514300 640481
rect 512724 640439 514300 640451
rect 512724 640387 513555 640439
rect 513555 640387 513607 640439
rect 513607 640387 514300 640439
rect 512724 640375 514300 640387
rect 512724 640345 513555 640375
rect 513555 640345 513607 640375
rect 513607 640345 514300 640375
<< metal3 >>
rect 508533 644156 508593 645743
rect 507781 644096 508593 644156
rect 508830 644157 508890 645743
rect 515532 645438 515670 645461
rect 508981 645408 510597 645414
rect 508981 645344 508987 645408
rect 509051 645389 509097 645408
rect 509161 645389 509207 645408
rect 509271 645389 509317 645408
rect 509381 645389 509427 645408
rect 509491 645389 509537 645408
rect 509601 645389 509647 645408
rect 509711 645389 509757 645408
rect 509821 645389 509867 645408
rect 509931 645389 509977 645408
rect 510041 645389 510087 645408
rect 510151 645389 510197 645408
rect 510261 645389 510307 645408
rect 510371 645389 510417 645408
rect 510481 645389 510527 645408
rect 510591 645344 510597 645408
rect 508981 645298 509001 645344
rect 510577 645298 510597 645344
rect 508981 645234 508987 645298
rect 509051 645234 509097 645253
rect 509161 645234 509207 645253
rect 509271 645234 509317 645253
rect 509381 645234 509427 645253
rect 509491 645234 509537 645253
rect 509601 645234 509647 645253
rect 509711 645234 509757 645253
rect 509821 645234 509867 645253
rect 509931 645234 509977 645253
rect 510041 645234 510087 645253
rect 510151 645234 510197 645253
rect 510261 645234 510307 645253
rect 510371 645234 510417 645253
rect 510481 645234 510527 645253
rect 510591 645234 510597 645298
rect 508981 645228 510597 645234
rect 515532 645382 515572 645438
rect 515628 645382 515670 645438
rect 515532 645358 515670 645382
rect 515532 645302 515572 645358
rect 515628 645302 515670 645358
rect 515532 645278 515670 645302
rect 515532 645222 515572 645278
rect 515628 645222 515670 645278
rect 509409 645106 509509 645115
rect 509409 645050 509431 645106
rect 509487 645050 509509 645106
rect 509409 645026 509509 645050
rect 509409 644970 509431 645026
rect 509487 644970 509509 645026
rect 509409 644946 509509 644970
rect 509409 644890 509431 644946
rect 509487 644890 509509 644946
rect 508830 644097 509292 644157
rect 507781 643340 507841 644096
rect 507972 643776 509148 643782
rect 507972 643712 507978 643776
rect 508042 643757 508088 643776
rect 508152 643757 508198 643776
rect 508262 643757 508308 643776
rect 508372 643757 508418 643776
rect 508482 643757 508528 643776
rect 508592 643757 508638 643776
rect 508702 643757 508748 643776
rect 508812 643757 508858 643776
rect 508922 643757 508968 643776
rect 509032 643757 509078 643776
rect 509142 643712 509148 643776
rect 507972 643666 508012 643712
rect 509108 643666 509148 643712
rect 507972 643602 507978 643666
rect 508042 643602 508088 643621
rect 508152 643602 508198 643621
rect 508262 643602 508308 643621
rect 508372 643602 508418 643621
rect 508482 643602 508528 643621
rect 508592 643602 508638 643621
rect 508702 643602 508748 643621
rect 508812 643602 508858 643621
rect 508922 643602 508968 643621
rect 509032 643602 509078 643621
rect 509142 643602 509148 643666
rect 507972 643596 509148 643602
rect 507733 643331 507887 643340
rect 507733 643195 507742 643331
rect 507878 643195 507887 643331
rect 507733 643186 507887 643195
rect 509232 642545 509292 644097
rect 509186 642536 509340 642545
rect 509186 642400 509195 642536
rect 509331 642400 509340 642536
rect 509186 642391 509340 642400
rect 509409 641206 509509 644890
rect 513989 645106 514089 645115
rect 513989 645050 514011 645106
rect 514067 645050 514089 645106
rect 513989 645026 514089 645050
rect 513989 644970 514011 645026
rect 514067 644970 514089 645026
rect 513989 644946 514089 644970
rect 513989 644890 514011 644946
rect 514067 644890 514089 644946
rect 509409 641150 509431 641206
rect 509487 641150 509509 641206
rect 509409 641126 509509 641150
rect 509409 641070 509431 641126
rect 509487 641070 509509 641126
rect 509409 641046 509509 641070
rect 509409 640990 509431 641046
rect 509487 640990 509509 641046
rect 509409 640981 509509 640990
rect 509868 644794 509968 644803
rect 509868 644738 509889 644794
rect 509945 644738 509968 644794
rect 509868 644714 509968 644738
rect 509868 644658 509889 644714
rect 509945 644658 509968 644714
rect 509868 644634 509968 644658
rect 509868 644578 509889 644634
rect 509945 644578 509968 644634
rect 509868 640852 509968 644578
rect 511241 644794 511341 644803
rect 511241 644738 511263 644794
rect 511319 644738 511341 644794
rect 511241 644714 511341 644738
rect 511241 644658 511263 644714
rect 511319 644658 511341 644714
rect 511241 644634 511341 644658
rect 511241 644578 511263 644634
rect 511319 644578 511341 644634
rect 510325 643797 510425 643806
rect 510325 643741 510347 643797
rect 510403 643741 510425 643797
rect 510325 643717 510425 643741
rect 510325 643661 510347 643717
rect 510403 643661 510425 643717
rect 510325 643637 510425 643661
rect 510325 643581 510347 643637
rect 510403 643581 510425 643637
rect 510325 641206 510425 643581
rect 510676 643292 510990 643301
rect 510676 643236 510685 643292
rect 510741 643236 510765 643292
rect 510821 643236 510845 643292
rect 510901 643236 510925 643292
rect 510981 643236 510990 643292
rect 510676 643227 510990 643236
rect 510783 642832 510883 643227
rect 510756 642823 510910 642832
rect 510756 642687 510765 642823
rect 510901 642687 510910 642823
rect 510756 642678 510910 642687
rect 510783 642506 510883 642678
rect 510676 642497 510990 642506
rect 510676 642441 510685 642497
rect 510741 642441 510765 642497
rect 510821 642441 510845 642497
rect 510901 642441 510925 642497
rect 510981 642441 510990 642497
rect 510676 642432 510990 642441
rect 511241 642161 511341 644578
rect 511241 642105 511263 642161
rect 511319 642105 511341 642161
rect 511241 642081 511341 642105
rect 511241 642025 511263 642081
rect 511319 642025 511341 642081
rect 511241 642001 511341 642025
rect 511241 641945 511263 642001
rect 511319 641945 511341 642001
rect 511241 641936 511341 641945
rect 512157 644794 512257 644803
rect 512157 644738 512179 644794
rect 512235 644738 512257 644794
rect 512157 644714 512257 644738
rect 512157 644658 512179 644714
rect 512235 644658 512257 644714
rect 512157 644634 512257 644658
rect 512157 644578 512179 644634
rect 512235 644578 512257 644634
rect 512157 642161 512257 644578
rect 513531 644794 513631 644803
rect 513531 644738 513553 644794
rect 513609 644738 513631 644794
rect 513531 644714 513631 644738
rect 513531 644658 513553 644714
rect 513609 644658 513631 644714
rect 513531 644634 513631 644658
rect 513531 644578 513553 644634
rect 513609 644578 513631 644634
rect 513073 643797 513173 643806
rect 513073 643741 513095 643797
rect 513151 643741 513173 643797
rect 513073 643717 513173 643741
rect 513073 643661 513095 643717
rect 513151 643661 513173 643717
rect 513073 643637 513173 643661
rect 513073 643581 513095 643637
rect 513151 643581 513173 643637
rect 512508 643292 512822 643301
rect 512508 643236 512517 643292
rect 512573 643236 512597 643292
rect 512653 643236 512677 643292
rect 512733 643236 512757 643292
rect 512813 643236 512822 643292
rect 512508 643227 512822 643236
rect 512616 643067 512716 643227
rect 512589 643058 512743 643067
rect 512589 642922 512598 643058
rect 512734 642922 512743 643058
rect 512589 642913 512743 642922
rect 512616 642506 512716 642913
rect 512508 642497 512822 642506
rect 512508 642441 512517 642497
rect 512573 642441 512597 642497
rect 512653 642441 512677 642497
rect 512733 642441 512757 642497
rect 512813 642441 512822 642497
rect 512508 642432 512822 642441
rect 512157 642105 512179 642161
rect 512235 642105 512257 642161
rect 512157 642081 512257 642105
rect 512157 642025 512179 642081
rect 512235 642025 512257 642081
rect 512157 642001 512257 642025
rect 512157 641945 512179 642001
rect 512235 641945 512257 642001
rect 512157 641936 512257 641945
rect 510325 641150 510347 641206
rect 510403 641150 510425 641206
rect 510325 641126 510425 641150
rect 510325 641070 510347 641126
rect 510403 641070 510425 641126
rect 510325 641046 510425 641070
rect 510325 640990 510347 641046
rect 510403 640990 510425 641046
rect 510325 640981 510425 640990
rect 513073 641206 513173 643581
rect 513531 642927 513631 644578
rect 513989 642927 514089 644890
rect 515532 643805 515670 645222
rect 515532 643749 515572 643805
rect 515628 643749 515670 643805
rect 515532 643725 515670 643749
rect 515532 643669 515572 643725
rect 515628 643669 515670 643725
rect 515532 643645 515670 643669
rect 515532 643589 515572 643645
rect 515628 643589 515670 643645
rect 515532 643574 515670 643589
rect 516655 644601 516755 644610
rect 516655 644545 516677 644601
rect 516733 644545 516755 644601
rect 516655 644521 516755 644545
rect 516655 644465 516677 644521
rect 516733 644465 516755 644521
rect 516655 644441 516755 644465
rect 516655 644385 516677 644441
rect 516733 644385 516755 644441
rect 516655 644361 516755 644385
rect 516655 644305 516677 644361
rect 516733 644305 516755 644361
rect 516655 644281 516755 644305
rect 516655 644225 516677 644281
rect 516733 644225 516755 644281
rect 516655 644201 516755 644225
rect 516655 644145 516677 644201
rect 516733 644145 516755 644201
rect 516655 642934 516755 644145
rect 513505 642918 513659 642927
rect 513505 642782 513514 642918
rect 513650 642782 513659 642918
rect 513505 642773 513659 642782
rect 513962 642918 514116 642927
rect 513962 642782 513971 642918
rect 514107 642782 514116 642918
rect 513962 642773 514116 642782
rect 516628 642925 516782 642934
rect 516628 642789 516637 642925
rect 516773 642789 516782 642925
rect 516628 642780 516782 642789
rect 513073 641150 513095 641206
rect 513151 641150 513173 641206
rect 513073 641126 513173 641150
rect 513073 641070 513095 641126
rect 513151 641070 513173 641126
rect 513073 641046 513173 641070
rect 513073 640990 513095 641046
rect 513151 640990 513173 641046
rect 513073 640981 513173 640990
rect 509868 640796 509889 640852
rect 509945 640796 509968 640852
rect 509868 640772 509968 640796
rect 509868 640716 509889 640772
rect 509945 640716 509968 640772
rect 509868 640692 509968 640716
rect 509868 640636 509889 640692
rect 509945 640636 509968 640692
rect 509868 640627 509968 640636
rect 513531 640852 513631 642773
rect 513989 641206 514089 642773
rect 516655 642285 516755 642780
rect 516655 642229 516677 642285
rect 516733 642229 516755 642285
rect 516655 642205 516755 642229
rect 516655 642149 516677 642205
rect 516733 642149 516755 642205
rect 514313 642140 515379 642146
rect 514313 642076 514319 642140
rect 514383 642121 514429 642140
rect 514493 642121 514539 642140
rect 514603 642121 514649 642140
rect 514713 642121 514759 642140
rect 514823 642121 514869 642140
rect 514933 642121 514979 642140
rect 515043 642121 515089 642140
rect 515153 642121 515199 642140
rect 515263 642121 515309 642140
rect 515373 642076 515379 642140
rect 514313 642030 514335 642076
rect 515351 642030 515379 642076
rect 514313 641966 514319 642030
rect 514383 641966 514429 641985
rect 514493 641966 514539 641985
rect 514603 641966 514649 641985
rect 514713 641966 514759 641985
rect 514823 641966 514869 641985
rect 514933 641966 514979 641985
rect 515043 641966 515089 641985
rect 515153 641966 515199 641985
rect 515263 641966 515309 641985
rect 515373 641966 515379 642030
rect 514313 641960 515379 641966
rect 516655 642125 516755 642149
rect 516655 642069 516677 642125
rect 516733 642069 516755 642125
rect 516655 642045 516755 642069
rect 516655 641989 516677 642045
rect 516733 641989 516755 642045
rect 516655 641965 516755 641989
rect 516655 641909 516677 641965
rect 516733 641909 516755 641965
rect 516655 641885 516755 641909
rect 516655 641829 516677 641885
rect 516733 641829 516755 641885
rect 516655 641820 516755 641829
rect 513989 641150 514011 641206
rect 514067 641150 514089 641206
rect 513989 641126 514089 641150
rect 513989 641070 514011 641126
rect 514067 641070 514089 641126
rect 513989 641046 514089 641070
rect 513989 640990 514011 641046
rect 514067 640990 514089 641046
rect 513989 640981 514089 640990
rect 513531 640796 513553 640852
rect 513609 640796 513631 640852
rect 513531 640772 513631 640796
rect 513531 640716 513553 640772
rect 513609 640716 513631 640772
rect 513531 640692 513631 640716
rect 513531 640636 513553 640692
rect 513609 640636 513631 640692
rect 513531 640627 513631 640636
rect 512704 640500 514320 640506
rect 512704 640436 512710 640500
rect 512774 640481 512820 640500
rect 512884 640481 512930 640500
rect 512994 640481 513040 640500
rect 513104 640481 513150 640500
rect 513214 640481 513260 640500
rect 513324 640481 513370 640500
rect 513434 640481 513480 640500
rect 513544 640481 513590 640500
rect 513654 640481 513700 640500
rect 513764 640481 513810 640500
rect 513874 640481 513920 640500
rect 513984 640481 514030 640500
rect 514094 640481 514140 640500
rect 514204 640481 514250 640500
rect 514314 640436 514320 640500
rect 512704 640390 512724 640436
rect 514300 640390 514320 640436
rect 512704 640326 512710 640390
rect 512774 640326 512820 640345
rect 512884 640326 512930 640345
rect 512994 640326 513040 640345
rect 513104 640326 513150 640345
rect 513214 640326 513260 640345
rect 513324 640326 513370 640345
rect 513434 640326 513480 640345
rect 513544 640326 513590 640345
rect 513654 640326 513700 640345
rect 513764 640326 513810 640345
rect 513874 640326 513920 640345
rect 513984 640326 514030 640345
rect 514094 640326 514140 640345
rect 514204 640326 514250 640345
rect 514314 640326 514320 640390
rect 512704 640320 514320 640326
<< via3 >>
rect 508987 645389 509051 645408
rect 509097 645389 509161 645408
rect 509207 645389 509271 645408
rect 509317 645389 509381 645408
rect 509427 645389 509491 645408
rect 509537 645389 509601 645408
rect 509647 645389 509711 645408
rect 509757 645389 509821 645408
rect 509867 645389 509931 645408
rect 509977 645389 510041 645408
rect 510087 645389 510151 645408
rect 510197 645389 510261 645408
rect 510307 645389 510371 645408
rect 510417 645389 510481 645408
rect 510527 645389 510591 645408
rect 508987 645344 509001 645389
rect 509001 645344 509051 645389
rect 509097 645344 509161 645389
rect 509207 645344 509271 645389
rect 509317 645344 509381 645389
rect 509427 645344 509491 645389
rect 509537 645344 509601 645389
rect 509647 645344 509711 645389
rect 509757 645344 509821 645389
rect 509867 645344 509931 645389
rect 509977 645344 510041 645389
rect 510087 645344 510151 645389
rect 510197 645344 510261 645389
rect 510307 645344 510371 645389
rect 510417 645344 510481 645389
rect 510527 645344 510577 645389
rect 510577 645344 510591 645389
rect 508987 645253 509001 645298
rect 509001 645253 509051 645298
rect 509097 645253 509161 645298
rect 509207 645253 509271 645298
rect 509317 645253 509381 645298
rect 509427 645253 509491 645298
rect 509537 645253 509601 645298
rect 509647 645253 509711 645298
rect 509757 645253 509821 645298
rect 509867 645253 509931 645298
rect 509977 645253 510041 645298
rect 510087 645253 510151 645298
rect 510197 645253 510261 645298
rect 510307 645253 510371 645298
rect 510417 645253 510481 645298
rect 510527 645253 510577 645298
rect 510577 645253 510591 645298
rect 508987 645234 509051 645253
rect 509097 645234 509161 645253
rect 509207 645234 509271 645253
rect 509317 645234 509381 645253
rect 509427 645234 509491 645253
rect 509537 645234 509601 645253
rect 509647 645234 509711 645253
rect 509757 645234 509821 645253
rect 509867 645234 509931 645253
rect 509977 645234 510041 645253
rect 510087 645234 510151 645253
rect 510197 645234 510261 645253
rect 510307 645234 510371 645253
rect 510417 645234 510481 645253
rect 510527 645234 510591 645253
rect 507978 643757 508042 643776
rect 508088 643757 508152 643776
rect 508198 643757 508262 643776
rect 508308 643757 508372 643776
rect 508418 643757 508482 643776
rect 508528 643757 508592 643776
rect 508638 643757 508702 643776
rect 508748 643757 508812 643776
rect 508858 643757 508922 643776
rect 508968 643757 509032 643776
rect 509078 643757 509142 643776
rect 507978 643712 508012 643757
rect 508012 643712 508042 643757
rect 508088 643712 508152 643757
rect 508198 643712 508262 643757
rect 508308 643712 508372 643757
rect 508418 643712 508482 643757
rect 508528 643712 508592 643757
rect 508638 643712 508702 643757
rect 508748 643712 508812 643757
rect 508858 643712 508922 643757
rect 508968 643712 509032 643757
rect 509078 643712 509108 643757
rect 509108 643712 509142 643757
rect 507978 643621 508012 643666
rect 508012 643621 508042 643666
rect 508088 643621 508152 643666
rect 508198 643621 508262 643666
rect 508308 643621 508372 643666
rect 508418 643621 508482 643666
rect 508528 643621 508592 643666
rect 508638 643621 508702 643666
rect 508748 643621 508812 643666
rect 508858 643621 508922 643666
rect 508968 643621 509032 643666
rect 509078 643621 509108 643666
rect 509108 643621 509142 643666
rect 507978 643602 508042 643621
rect 508088 643602 508152 643621
rect 508198 643602 508262 643621
rect 508308 643602 508372 643621
rect 508418 643602 508482 643621
rect 508528 643602 508592 643621
rect 508638 643602 508702 643621
rect 508748 643602 508812 643621
rect 508858 643602 508922 643621
rect 508968 643602 509032 643621
rect 509078 643602 509142 643621
rect 514319 642121 514383 642140
rect 514429 642121 514493 642140
rect 514539 642121 514603 642140
rect 514649 642121 514713 642140
rect 514759 642121 514823 642140
rect 514869 642121 514933 642140
rect 514979 642121 515043 642140
rect 515089 642121 515153 642140
rect 515199 642121 515263 642140
rect 515309 642121 515373 642140
rect 514319 642076 514335 642121
rect 514335 642076 514383 642121
rect 514429 642076 514493 642121
rect 514539 642076 514603 642121
rect 514649 642076 514713 642121
rect 514759 642076 514823 642121
rect 514869 642076 514933 642121
rect 514979 642076 515043 642121
rect 515089 642076 515153 642121
rect 515199 642076 515263 642121
rect 515309 642076 515351 642121
rect 515351 642076 515373 642121
rect 514319 641985 514335 642030
rect 514335 641985 514383 642030
rect 514429 641985 514493 642030
rect 514539 641985 514603 642030
rect 514649 641985 514713 642030
rect 514759 641985 514823 642030
rect 514869 641985 514933 642030
rect 514979 641985 515043 642030
rect 515089 641985 515153 642030
rect 515199 641985 515263 642030
rect 515309 641985 515351 642030
rect 515351 641985 515373 642030
rect 514319 641966 514383 641985
rect 514429 641966 514493 641985
rect 514539 641966 514603 641985
rect 514649 641966 514713 641985
rect 514759 641966 514823 641985
rect 514869 641966 514933 641985
rect 514979 641966 515043 641985
rect 515089 641966 515153 641985
rect 515199 641966 515263 641985
rect 515309 641966 515373 641985
rect 512710 640481 512774 640500
rect 512820 640481 512884 640500
rect 512930 640481 512994 640500
rect 513040 640481 513104 640500
rect 513150 640481 513214 640500
rect 513260 640481 513324 640500
rect 513370 640481 513434 640500
rect 513480 640481 513544 640500
rect 513590 640481 513654 640500
rect 513700 640481 513764 640500
rect 513810 640481 513874 640500
rect 513920 640481 513984 640500
rect 514030 640481 514094 640500
rect 514140 640481 514204 640500
rect 514250 640481 514314 640500
rect 512710 640436 512724 640481
rect 512724 640436 512774 640481
rect 512820 640436 512884 640481
rect 512930 640436 512994 640481
rect 513040 640436 513104 640481
rect 513150 640436 513214 640481
rect 513260 640436 513324 640481
rect 513370 640436 513434 640481
rect 513480 640436 513544 640481
rect 513590 640436 513654 640481
rect 513700 640436 513764 640481
rect 513810 640436 513874 640481
rect 513920 640436 513984 640481
rect 514030 640436 514094 640481
rect 514140 640436 514204 640481
rect 514250 640436 514300 640481
rect 514300 640436 514314 640481
rect 512710 640345 512724 640390
rect 512724 640345 512774 640390
rect 512820 640345 512884 640390
rect 512930 640345 512994 640390
rect 513040 640345 513104 640390
rect 513150 640345 513214 640390
rect 513260 640345 513324 640390
rect 513370 640345 513434 640390
rect 513480 640345 513544 640390
rect 513590 640345 513654 640390
rect 513700 640345 513764 640390
rect 513810 640345 513874 640390
rect 513920 640345 513984 640390
rect 514030 640345 514094 640390
rect 514140 640345 514204 640390
rect 514250 640345 514300 640390
rect 514300 640345 514314 640390
rect 512710 640326 512774 640345
rect 512820 640326 512884 640345
rect 512930 640326 512994 640345
rect 513040 640326 513104 640345
rect 513150 640326 513214 640345
rect 513260 640326 513324 640345
rect 513370 640326 513434 640345
rect 513480 640326 513544 640345
rect 513590 640326 513654 640345
rect 513700 640326 513764 640345
rect 513810 640326 513874 640345
rect 513920 640326 513984 640345
rect 514030 640326 514094 640345
rect 514140 640326 514204 640345
rect 514250 640326 514314 640345
<< metal4 >>
rect 507879 645408 510679 645496
rect 507879 645344 508987 645408
rect 509051 645344 509097 645408
rect 509161 645344 509207 645408
rect 509271 645344 509317 645408
rect 509381 645344 509427 645408
rect 509491 645344 509537 645408
rect 509601 645344 509647 645408
rect 509711 645344 509757 645408
rect 509821 645344 509867 645408
rect 509931 645344 509977 645408
rect 510041 645344 510087 645408
rect 510151 645344 510197 645408
rect 510261 645344 510307 645408
rect 510371 645344 510417 645408
rect 510481 645344 510527 645408
rect 510591 645344 510679 645408
rect 507879 645298 510679 645344
rect 507879 645234 508987 645298
rect 509051 645234 509097 645298
rect 509161 645234 509207 645298
rect 509271 645234 509317 645298
rect 509381 645234 509427 645298
rect 509491 645234 509537 645298
rect 509601 645234 509647 645298
rect 509711 645234 509757 645298
rect 509821 645234 509867 645298
rect 509931 645234 509977 645298
rect 510041 645234 510087 645298
rect 510151 645234 510197 645298
rect 510261 645234 510307 645298
rect 510371 645234 510417 645298
rect 510481 645234 510527 645298
rect 510591 645234 510679 645298
rect 507879 643776 510679 645234
rect 507879 643712 507978 643776
rect 508042 643712 508088 643776
rect 508152 643712 508198 643776
rect 508262 643712 508308 643776
rect 508372 643712 508418 643776
rect 508482 643712 508528 643776
rect 508592 643712 508638 643776
rect 508702 643712 508748 643776
rect 508812 643712 508858 643776
rect 508922 643712 508968 643776
rect 509032 643712 509078 643776
rect 509142 643712 510679 643776
rect 507879 643666 510679 643712
rect 507879 643602 507978 643666
rect 508042 643602 508088 643666
rect 508152 643602 508198 643666
rect 508262 643602 508308 643666
rect 508372 643602 508418 643666
rect 508482 643602 508528 643666
rect 508592 643602 508638 643666
rect 508702 643602 508748 643666
rect 508812 643602 508858 643666
rect 508922 643602 508968 643666
rect 509032 643602 509078 643666
rect 509142 643602 510679 643666
rect 507879 640193 510679 643602
rect 512194 642140 515394 645496
rect 512194 642076 514319 642140
rect 514383 642076 514429 642140
rect 514493 642076 514539 642140
rect 514603 642076 514649 642140
rect 514713 642076 514759 642140
rect 514823 642076 514869 642140
rect 514933 642076 514979 642140
rect 515043 642076 515089 642140
rect 515153 642076 515199 642140
rect 515263 642076 515309 642140
rect 515373 642076 515394 642140
rect 512194 642030 515394 642076
rect 512194 641966 514319 642030
rect 514383 641966 514429 642030
rect 514493 641966 514539 642030
rect 514603 641966 514649 642030
rect 514713 641966 514759 642030
rect 514823 641966 514869 642030
rect 514933 641966 514979 642030
rect 515043 641966 515089 642030
rect 515153 641966 515199 642030
rect 515263 641966 515309 642030
rect 515373 641966 515394 642030
rect 512194 640500 515394 641966
rect 512194 640436 512710 640500
rect 512774 640436 512820 640500
rect 512884 640436 512930 640500
rect 512994 640436 513040 640500
rect 513104 640436 513150 640500
rect 513214 640436 513260 640500
rect 513324 640436 513370 640500
rect 513434 640436 513480 640500
rect 513544 640436 513590 640500
rect 513654 640436 513700 640500
rect 513764 640436 513810 640500
rect 513874 640436 513920 640500
rect 513984 640436 514030 640500
rect 514094 640436 514140 640500
rect 514204 640436 514250 640500
rect 514314 640436 515394 640500
rect 512194 640390 515394 640436
rect 512194 640326 512710 640390
rect 512774 640326 512820 640390
rect 512884 640326 512930 640390
rect 512994 640326 513040 640390
rect 513104 640326 513150 640390
rect 513214 640326 513260 640390
rect 513324 640326 513370 640390
rect 513434 640326 513480 640390
rect 513544 640326 513590 640390
rect 513654 640326 513700 640390
rect 513764 640326 513810 640390
rect 513874 640326 513920 640390
rect 513984 640326 514030 640390
rect 514094 640326 514140 640390
rect 514204 640326 514250 640390
rect 514314 640326 515394 640390
rect 512194 640192 515394 640326
<< labels >>
flabel metal2 s 516982 642857 516982 642857 0 FreeSans 364 0 0 0 VOUT
flabel metal2 s 507830 642468 507830 642468 0 FreeSans 364 0 0 0 VBN
flabel metal2 s 508001 640415 508001 640415 0 FreeSans 364 0 0 0 VSS
flabel metal2 s 508011 645316 508011 645316 0 FreeSans 364 0 0 0 VDD
flabel metal2 s 507825 642754 507825 642754 0 FreeSans 364 0 0 0 VINM
flabel metal2 s 507823 642989 507823 642989 0 FreeSans 364 0 0 0 VINP
flabel metal3 s 507839 643262 507839 643262 0 FreeSans 364 0 0 0 VBP
<< end >>
