* NGSPICE file created from EF_R2RVC02mf.ext - technology: sky130A

.subckt EF_R2RVC02mf a1 a2 b1 b2 vo sela selb vdd1p8 vss dvss vdd3p3
X0 a_1821_8526.t1 comparator_top_0.comparator_0.VBN.t3 comparator_top_0.comparator_0.VBN.t4 vdd3p3.t92 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=1.5e+07u
X1 vss vss.t52 vss vss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=3.335e+13p pd=2.4334e+08u as=0p ps=0u w=5e+06u l=2e+06u
X2 vss.t51 vss.t49 vss.t50 vss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X3 a_2551_4880.t5 a_2151_4783.t8 vdd3p3.t5 vdd3p3.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X4 comparator_top_0.comparator_0.VOUT a_8881_1782.t2 vdd3p3.t154 vdd3p3.t153 sky130_fd_pr__pfet_g5v0d10v5 ad=2.9e+12p pd=2.058e+07u as=0p ps=0u w=1e+07u l=2e+06u
X5 a_570_n5724.t5 a_470_n5812# dvss.t94 dvss.t93 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 b1.t1 dvss.t24 sky130_fd_pr__nfet_g5v0d10v5 ad=4.64e+12p pd=3.664e+07u as=0p ps=0u w=2e+06u l=500000u
X7 dvss.t158 a_570_n5724.t6 a_1777_n6060# dvss.t157 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X8 vdd3p3.t107 a_1821_8526.t6 a_2221_8623.t5 vdd3p3.t106 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X9 a_2093_3714.t7 comparator_top_0.comparator_0.VBP.t4 vdd3p3.t150 vdd3p3.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X10 vdd3p3.t129 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 vdd3p3.t128 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
D0 dvss EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X11 a_6351_6657# a_10811_7187# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X12 vss.t80 a_2151_594.t8 a_2551_620.t1 vss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X13 a_5299_3714.t7 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_3714.t11 vdd3p3.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X14 dvss.t164 a_3916_n5703.t6 a_5123_n6039# dvss.t163 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X15 vss.t67 comparator_top_0.comparator_0.VBN.t9 a_2093_1782.t7 vss.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X16 a_10542_n5707.t4 a_10442_n5795# dvss.t70 dvss.t69 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X17 a_2093_3714.t5 vdd3p3.t71 vdd3p3.t72 vdd3p3.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X18 dvss.t181 a_10965_3602# a_10975_4108# dvss.t180 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=6.075e+11p ps=6.12e+06u w=750000u l=500000u
X19 a_7889_n6842# a_7464_n6798# dvss.t17 dvss.t16 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X20 vdd3p3 vdd3p3.t67 vdd3p3 vdd3p3.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=4.40314e+13p pd=3.334e+08u as=0p ps=0u w=5e+06u l=2e+06u
X21 dvss.t28 a_10975_4108# vo.t1 dvss.t27 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=740000u l=150000u
X22 dvss.t124 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 dvss.t123 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X23 vdd3p3.t32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 vdd3p3.t31 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 vdd3p3.t17 vdd3p3.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A sela.t0 vdd1p8.t22 vdd1p8.t21 sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X26 dvss.t15 a_7464_n6798# a_7889_n6842# dvss.t14 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X27 vdd1p8.t24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A a_10442_n5795# vdd1p8.t23 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X28 a_7464_n6798# a_7096_n5816# vdd1p8.t28 vdd1p8.t27 sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_5123_n6039# dvss.t33 dvss.t32 sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X30 a_4184_n6773# a_3816_n5791# vdd1p8.t14 vdd1p8.t13 sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X31 vss.t48 vss.t46 comparator_top_0.comparator_0.VBN.t8 vss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X33 a_2093_3714.t10 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_5299_3714.t6 vdd3p3.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X34 vss.t58 a_5299_620.t8 a_8881_1782.t0 vss.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
D1 dvss EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X35 dvss.t22 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 dvss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X36 a_4609_n6817# a_4184_n6773# dvss.t50 dvss.t49 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X37 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_1777_n6060# vdd3p3.t127 vdd3p3.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X38 a1.t7 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=2.32e+12p ps=2.064e+07u w=1e+06u l=500000u
X39 a_838_n6794# a_470_n5812# vdd1p8.t12 vdd1p8.t11 sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X40 dvss.t120 comparator_top_0.comparator_0.VOUT a_11031_3400# dvss.t119 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.197e+11p ps=1.41e+06u w=420000u l=500000u
X41 vss vss.t42 vss vss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X42 vdd3p3.t109 a_11235_n6821# a_10542_n5707.t5 vdd3p3.t108 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X43 vdd3p3 vdd3p3.t62 vdd3p3 vdd3p3.t63 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X44 a_2151_594.t3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_3714.t0 vdd3p3.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
D2 dvss EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X45 comparator_top_0.comparator_0.VBN.t5 a_2221_8623.t6 a_1821_8526.t2 vdd3p3.t95 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X46 a_7464_n6798# a_7096_n5816# dvss.t195 dvss.t194 sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss.t168 dvss.t167 sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_11749_n6043# vdd3p3.t116 vdd3p3.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X49 vdd3p3.t146 a_570_n5724.t7 a_1777_n6060# vdd3p3.t126 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X50 a_5299_1782.t3 a_5299_1782.t2 vdd3p3.t149 vdd3p3.t145 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X51 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 a1.t6 vdd3p3.t162 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X52 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t169 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X53 a_7889_n6842# a_7464_n6798# dvss.t13 dvss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X54 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A vdd3p3.t14 vdd3p3.t13 sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X55 comparator_top_0.comparator_0.VOUT a_8881_1782.t3 vss.t82 vss.t81 sky130_fd_pr__nfet_g5v0d10v5 ad=1.45e+12p pd=1.058e+07u as=0p ps=0u w=5e+06u l=2e+06u
X56 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A sela.t1 dvss.t26 dvss.t25 sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X57 dvss.t142 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 dvss.t141 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X58 vdd1p8.t10 a_11271_4224# a_10975_4108# vdd1p8.t9 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.968e+11p ps=2.77e+06u w=1.12e+06u l=150000u
X59 a_11271_4224# a_11031_3400# dvss.t152 dvss.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=6.075e+11p pd=6.12e+06u as=0p ps=0u w=750000u l=500000u
X60 b1.t3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 b1.t2 vdd3p3.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X61 vdd3p3.t139 a_10542_n5707.t6 a_11749_n6043# vdd3p3.t115 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X62 vdd3p3.t7 a_2151_4783.t9 a_2551_4880.t4 vdd3p3.t6 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X63 a_2093_1782.t6 comparator_top_0.comparator_0.VBN.t10 vss.t65 vss.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X64 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 b2.t5 vdd3p3.t159 sky130_fd_pr__pfet_g5v0d10v5 ad=2.32e+12p pd=2.064e+07u as=0p ps=0u w=1e+06u l=500000u
X65 a_838_n6794# a_470_n5812# dvss.t92 dvss.t91 sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X66 a_2093_3714.t3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2151_594.t2 vdd3p3.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X67 a_11271_4224# a_10975_4108# vdd1p8.t2 vdd1p8.t0 sky130_fd_pr__pfet_01v8_hvt ad=2.968e+11p pd=2.77e+06u as=0p ps=0u w=1.12e+06u l=150000u
X68 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A selb.t0 vdd1p8.t16 vdd1p8.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X69 vdd3p3.t152 a_3916_n5703.t7 a_5123_n6039# vdd3p3.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X70 a_3916_n5703.t4 a_3816_n5791# dvss.t106 dvss.t105 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X71 a_5299_1782.t7 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_1782.t9 vss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X72 vss.t76 a_5299_3714.t8 a_5299_620.t4 vss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X73 dvss.t104 a_3816_n5791# a_3916_n5703.t3 dvss.t103 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X74 vdd3p3.t61 vdd3p3.t59 vdd3p3.t60 vdd3p3.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X75 vdd3p3.t171 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 vdd3p3.t170 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X76 vdd3p3.t148 a_5299_1782.t0 a_5299_1782.t1 vdd3p3.t144 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X77 comparator_top_0.comparator_0.VBN.t2 comparator_top_0.comparator_0.VBN.t1 vss.t64 vss.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X78 dvss.t179 a_10965_3602# a_10975_4108# dvss.t178 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X79 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_5123_n6039# vdd3p3.t29 vdd3p3.t28 sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X80 dvss.t108 a_7196_n5728.t6 a_8403_n6064# dvss.t107 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X81 a_2093_1782.t5 vss.t39 vss.t41 vss.t40 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X82 a_570_n5724.t4 a_470_n5812# dvss.t90 dvss.t89 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X83 a_10810_n6777# a_10442_n5795# dvss.t68 dvss.t67 sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X84 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss.t7 dvss.t6 sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X85 a_6349_9307# a_10809_9307# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X86 a2.t3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X87 a_2151_4783.t7 a_2151_4783.t6 vdd3p3.t91 vdd3p3.t27 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X88 vdd1p8.t6 selb.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A vdd1p8.t5 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X89 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A vdd3p3.t158 vdd3p3.t157 sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X90 a_6351_7717# a_10811_7187# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X91 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 vdd3p3.t114 vdd3p3.t15 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X92 dvss.t134 a_10810_n6777# a_11235_n6821# dvss.t133 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.2375e+12p ps=1.065e+07u w=1.5e+06u l=500000u
X93 dvss.t11 a_7464_n6798# a_7889_n6842# dvss.t10 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X94 a_1821_8526.t3 a_2221_8623.t7 comparator_top_0.comparator_0.VBN.t6 vdd3p3.t96 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X95 a_7889_n6842# a_7464_n6798# dvss.t9 dvss.t8 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X96 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_8403_n6064# dvss.t160 dvss.t159 sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X97 b2.t3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 b2.t2 vdd3p3.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X98 a_2093_1782.t8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_5299_1782.t6 vss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X99 dvss.t111 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 dvss.t110 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X100 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A selb.t2 dvss.t40 dvss.t39 sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X101 vss vss.t34 vss vss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X102 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 b2.t1 dvss.t23 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X103 vdd1p8.t1 a_10975_4108# vo.t0 vdd1p8.t0 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=0p ps=0u w=1.12e+06u l=150000u
X104 a_2151_4783.t0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_1782.t3 vss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X105 a2.t1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 a2.t0 dvss.t109 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X106 vdd3p3.t168 a_2551_620.t4 a_2551_620.t5 vdd3p3.t26 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X107 dvss.t151 a_11031_3400# a_10965_3602# dvss.t150 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.197e+11p ps=1.41e+06u w=420000u l=500000u
X108 vss.t1 a_5299_3714.t2 a_5299_3714.t3 vss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X109 a_2151_594.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_3714.t2 vdd3p3.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X110 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 vdd3p3.t131 vdd3p3.t130 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X111 a_1263_n6838# a_838_n6794# dvss.t80 dvss.t79 sky130_fd_pr__nfet_g5v0d10v5 ad=1.2375e+12p pd=1.065e+07u as=0p ps=0u w=1.5e+06u l=500000u
X112 vdd3p3.t58 vdd3p3.t55 vdd3p3.t57 vdd3p3.t56 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X113 dvss.t149 a_11031_3400# a_11271_4224# dvss.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X114 a_570_n5724.t3 a_470_n5812# dvss.t88 dvss.t87 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X115 dvss.t170 selb.t3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A dvss.t169 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X116 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A vdd3p3.t123 vdd3p3.t122 sky130_fd_pr__pfet_g5v0d10v5 ad=4.2e+11p pd=3.56e+06u as=0p ps=0u w=1.5e+06u l=500000u
X117 vdd3p3.t94 a_1263_n6838# a_570_n5724.t0 vdd3p3.t93 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X118 vss vss.t29 vss vss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X119 dvss.t1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 dvss.t0 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X120 vdd3p3.t105 a_1821_8526.t7 a_2221_8623.t4 vdd3p3.t104 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X121 a_6351_6657# a_1821_8526.t5 dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X122 a_11235_n6821# a_10810_n6777# dvss.t132 dvss.t131 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X123 a_6349_9307# a_10811_8247# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X124 vdd3p3 vdd3p3.t50 vdd3p3 vdd3p3.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X125 a_2093_1782.t2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2151_4783.t3 vss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X126 comparator_top_0.comparator_0.VBP.t3 comparator_top_0.comparator_0.VBP.t2 vdd3p3.t74 vdd3p3.t73 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X127 vdd3p3.t24 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 vdd3p3.t23 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X128 a_10810_n6777# a_10442_n5795# vdd1p8.t4 vdd1p8.t3 sky130_fd_pr__pfet_01v8_hvt ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X129 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t30 vdd3p3.t22 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X130 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t30 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X131 a_7196_n5728.t5 a_7096_n5816# dvss.t193 dvss.t192 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X132 vss.t28 vss.t25 vss.t27 vss.t26 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
D3 dvss EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y sky130_fd_pr__diode_pw2nd_05v5 pj=1.8e+06 area=2.025e+11
X133 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t117 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X134 dvss.t102 a_3816_n5791# a_3916_n5703.t2 dvss.t101 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X135 a2.t7 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t19 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=4.64e+12p ps=3.664e+07u w=2e+06u l=500000u
X136 dvss.t191 a_7096_n5816# a_7196_n5728.t4 dvss.t190 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X137 comparator_top_0.comparator_0.VBN.t7 a_2221_8623.t8 a_1821_8526.t4 vdd3p3.t97 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X138 vdd3p3.t3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 vdd3p3.t2 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X139 dvss.t78 a_838_n6794# a_1263_n6838# dvss.t77 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X140 a_1263_n6838# a_838_n6794# dvss.t76 dvss.t75 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X141 dvss.t86 a_470_n5812# a_570_n5724.t2 dvss.t85 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X142 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss.t118 dvss.t117 sky130_fd_pr__nfet_g5v0d10v5 ad=2.1e+11p pd=2.06e+06u as=0p ps=0u w=750000u l=500000u
X143 vss.t62 comparator_top_0.comparator_0.VBN.t11 a_2221_8623.t1 vss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X144 vdd3p3.t136 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 vdd3p3.t135 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X145 dvss.t130 a_10810_n6777# a_11235_n6821# dvss.t129 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X146 a_2551_620.t3 a_2551_620.t2 vdd3p3.t10 vdd3p3.t9 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X147 a_2093_3714.t9 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_5299_3714.t5 vdd3p3.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X148 a_4609_n6817# a_4184_n6773# dvss.t48 dvss.t47 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X149 vdd1p8.t20 sela.t2 a_470_n5812# vdd1p8.t19 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X150 a_11235_n6821# a_10810_n6777# dvss.t128 dvss.t127 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X151 vss.t73 a_2551_4880.t6 a_5299_620.t1 vss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X152 a_5299_620.t3 a_5299_3714.t9 vss.t77 vss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X153 vdd3p3.t78 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 vdd3p3.t77 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X154 a1.t5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 a1.t4 dvss.t171 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X155 dvss.t52 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 dvss.t51 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X156 a1.t3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t135 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X157 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t134 vdd3p3.t18 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X158 vdd3p3.t89 a_5299_1782.t8 a_5299_620.t2 vdd3p3.t51 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X159 b1.t4 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X160 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t19 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X161 dvss.t82 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A a_3816_n5791# dvss.t81 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X162 dvss.t189 a_7096_n5816# a_7196_n5728.t3 dvss.t188 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X163 b1.t6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 b1.t5 dvss.t140 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X164 a_3916_n5703.t1 a_3816_n5791# dvss.t100 dvss.t99 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X165 a_2221_8623.t3 a_1821_8526.t8 vdd3p3.t103 vdd3p3.t102 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X166 vdd3p3.t49 vdd3p3.t47 a_2093_3714.t4 vdd3p3.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X167 a_2151_4783.t2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_1782.t1 vss.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X168 a_7196_n5728.t2 a_7096_n5816# dvss.t187 dvss.t186 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X169 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 a1.t2 dvss.t136 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X170 dvss.t156 sela.t3 a_470_n5812# dvss.t155 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X171 vdd3p3.t88 a_570_n5724.t8 a_1263_n6838# vdd3p3.t87 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=1e+06u
X172 a_5299_620.t0 a_2551_4880.t7 vss.t75 vss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X173 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t133 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X174 a1.t1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 a1.t0 vdd3p3.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X175 a_1263_n6838# a_838_n6794# dvss.t74 dvss.t73 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X176 dvss.t84 a_470_n5812# a_570_n5724.t1 dvss.t83 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X177 a_2093_3714.t1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2151_594.t0 vdd3p3.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X178 vdd3p3.t121 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t120 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X179 vdd3p3.t141 a_10542_n5707.t7 a_11235_n6821# vdd3p3.t140 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=1e+06u
X180 vss vss.t20 vss vss.t21 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X181 a_11271_4224# a_11031_3400# dvss.t148 dvss.t147 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X182 a_11235_n6821# a_10810_n6777# dvss.t126 dvss.t125 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X183 dvss.t46 a_4184_n6773# a_4609_n6817# dvss.t45 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X184 a_2151_594.t7 a_2151_594.t6 vss.t79 vss.t5 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X185 vss.t71 a_2551_4880.t2 a_2551_4880.t3 vss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X186 a_10975_4108# a_10965_3602# dvss.t177 dvss.t176 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X187 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 a2.t2 vdd3p3.t110 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X188 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_11749_n6043# dvss.t113 dvss.t112 sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X189 a_2221_8623.t0 vss.t17 vss.t19 vss.t18 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X190 vdd3p3.t160 a_2551_620.t6 a_5299_620.t7 vdd3p3.t143 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X191 vdd3p3.t112 a_7889_n6842# a_7196_n5728.t0 vdd3p3.t111 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X192 a_5299_3714.t4 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_3714.t8 vdd3p3.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X193 b1.t0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t114 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X194 comparator_top_0.comparator_0.VBP.t0 vss.t14 vss.t16 vss.t15 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X195 a_5299_3714.t1 a_5299_3714.t0 vss.t69 vss.t68 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X196 a_10542_n5707.t3 a_10442_n5795# dvss.t66 dvss.t65 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X197 dvss.t139 a_10542_n5707.t8 a_11749_n6043# dvss.t138 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=1.9875e+11p ps=2.03e+06u w=750000u l=500000u
X198 vdd1p8.t18 sela.t4 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A vdd1p8.t17 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X199 vdd1p8.t26 selb.t4 a_7096_n5816# vdd1p8.t25 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X200 a_1821_8526.t0 a_2221_8623.t9 comparator_top_0.comparator_0.VBN.t0 vdd3p3.t8 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X201 a_10965_3602# a_11031_3400# vdd3p3.t138 vdd3p3.t137 sky130_fd_pr__pfet_g5v0d10v5 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=500000u
X202 a_11031_3400# comparator_top_0.comparator_0.VOUT vdd3p3.t125 vdd3p3.t124 sky130_fd_pr__pfet_g5v0d10v5 ad=1.113e+11p pd=1.37e+06u as=0p ps=0u w=420000u l=500000u
X203 a_2093_1782.t11 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_5299_1782.t5 vss.t72 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X204 a_2551_4880.t1 a_2551_4880.t0 vss.t70 vss.t3 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X205 dvss.t36 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 dvss.t35 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X206 dvss.t116 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss.t115 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X207 vdd1p8.t8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A a_3816_n5791# vdd1p8.t7 sky130_fd_pr__pfet_01v8_hvt ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X208 a_5299_620.t5 a_5299_1782.t9 vdd3p3.t113 vdd3p3.t48 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X209 vdd3p3 vdd3p3.t43 vdd3p3 vdd3p3.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X210 vdd3p3.t99 a_7196_n5728.t7 a_8403_n6064# vdd3p3.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=3.975e+11p ps=3.53e+06u w=1.5e+06u l=500000u
X211 a_4609_n6817# a_4184_n6773# dvss.t44 dvss.t43 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X212 dvss.t42 a_4184_n6773# a_4609_n6817# dvss.t41 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X213 dvss.t58 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss.t57 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=2.1e+11p ps=2.06e+06u w=750000u l=500000u
X214 vdd3p3.t21 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 vdd3p3.t20 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X215 vdd3p3.t90 a_2151_4783.t4 a_2151_4783.t5 vdd3p3.t25 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X216 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss.t56 dvss.t55 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X217 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_8403_n6064# vdd3p3.t147 vdd3p3.t98 sky130_fd_pr__pfet_g5v0d10v5 ad=3.975e+11p pd=3.53e+06u as=0p ps=0u w=1.5e+06u l=500000u
X218 a_2551_620.t0 a_2151_594.t9 vss.t78 vss.t66 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X219 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t34 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X220 dvss.t166 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss.t165 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X221 vss.t13 vss.t11 a_2093_1782.t4 vss.t12 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X222 a_3916_n5703.t0 a_3816_n5791# dvss.t98 dvss.t97 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X223 dvss.t173 selb.t5 a_7096_n5816# dvss.t172 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X224 vdd3p3.t132 a_10809_9307# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X225 vdd3p3.t151 comparator_top_0.comparator_0.VBP.t5 a_2093_3714.t6 vdd3p3.t4 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X226 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 vdd3p3.t119 vdd3p3.t118 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X227 b2.t4 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out vdd3p3.t16 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X228 vdd3p3.t12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t11 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X229 a_7196_n5728.t1 a_7096_n5816# dvss.t185 dvss.t184 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X230 dvss.t154 sela.t5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A dvss.t153 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X231 dvss.t146 a_11031_3400# a_11271_4224# dvss.t145 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X232 vss.t56 a_2151_594.t4 a_2151_594.t5 vss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X233 a_5299_620.t6 a_2551_620.t7 vdd3p3.t161 vdd3p3.t142 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X234 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 b1.t7 vdd3p3.t165 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X235 a_2093_1782.t0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2151_4783.t1 vss.t2 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X236 dvss.t162 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 dvss.t161 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X237 dvss.t72 a_838_n6794# a_1263_n6838# dvss.t71 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X238 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t29 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X239 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 a2.t6 dvss.t20 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X240 vdd3p3.t84 a_3916_n5703.t8 a_4609_n6817# vdd3p3.t83 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=1e+06u
X241 dvss.t175 a_10965_3602# a_10975_4108# dvss.t174 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X242 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t1 vdd3p3.t0 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X243 vss vss.t6 vss vss.t7 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X244 a_6351_7717# a_10811_8247# dvss sky130_fd_pr__res_high_po w=1.41e+06u l=2.014e+07u
X245 vdd3p3.t86 a_5299_620.t9 a_8881_1782.t1 vdd3p3.t85 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+07u l=2e+06u
X246 vdd3p3 vdd3p3.t38 vdd3p3 vdd3p3.t39 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X247 vdd3p3.t164 a_4609_n6817# a_3916_n5703.t5 vdd3p3.t163 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=420000u l=1e+06u
X248 vdd3p3.t82 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t81 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=4.2e+11p ps=3.56e+06u w=1.5e+06u l=500000u
X249 a_2221_8623.t2 a_1821_8526.t9 vdd3p3.t101 vdd3p3.t100 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X250 vdd3p3 vdd3p3.t33 vdd3p3 vdd3p3.t34 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X251 a_5299_1782.t4 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_2093_1782.t10 vss.t74 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X252 a2.t5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 a2.t4 vdd3p3.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X253 dvss.t64 a_10442_n5795# a_10542_n5707.t2 dvss.t63 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X254 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A vdd3p3.t80 vdd3p3.t79 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X255 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t76 vdd3p3.t75 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1e+06u l=500000u
X256 dvss.t183 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A a_10442_n5795# dvss.t182 sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.478e+11p ps=2.27e+06u w=840000u l=150000u
X257 dvss.t5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss.t4 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=750000u l=500000u
X258 a_4184_n6773# a_3816_n5791# dvss.t96 dvss.t95 sky130_fd_pr__nfet_01v8 ad=2.478e+11p pd=2.27e+06u as=0p ps=0u w=840000u l=150000u
X259 a_10542_n5707.t1 a_10442_n5795# dvss.t62 dvss.t61 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X260 vss.t60 comparator_top_0.comparator_0.VBN.t12 comparator_top_0.comparator_0.VBP.t1 vss.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=5e+06u l=2e+06u
X261 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_1777_n6060# dvss.t122 dvss.t121 sky130_fd_pr__nfet_g5v0d10v5 ad=1.9875e+11p pd=2.03e+06u as=0p ps=0u w=750000u l=500000u
X262 vdd3p3.t156 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y vdd3p3.t155 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
X263 vdd3p3.t167 a_7196_n5728.t8 a_7889_n6842# vdd3p3.t166 sky130_fd_pr__pfet_g5v0d10v5 ad=0p pd=0u as=1.365e+11p ps=1.49e+06u w=420000u l=1e+06u
X264 b2.t0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss.t137 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X265 b2.t7 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 b2.t6 dvss.t31 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=2e+06u l=500000u
X266 dvss.t60 a_10442_n5795# a_10542_n5707.t0 dvss.t59 sky130_fd_pr__nfet_g5v0d10v5 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=500000u
R0 comparator_top_0.comparator_0.VBN.n263 comparator_top_0.comparator_0.VBN.t1 60.25
R1 comparator_top_0.comparator_0.VBN.n284 comparator_top_0.comparator_0.VBN.t11 60.25
R2 comparator_top_0.comparator_0.VBN.n304 comparator_top_0.comparator_0.VBN.t12 60.25
R3 comparator_top_0.comparator_0.VBN.n306 comparator_top_0.comparator_0.VBN.t10 60.25
R4 comparator_top_0.comparator_0.VBN.n318 comparator_top_0.comparator_0.VBN.t9 60.25
R5 comparator_top_0.comparator_0.VBN.n97 comparator_top_0.comparator_0.VBN.n95 41.883
R6 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.t4 35.112
R7 comparator_top_0.comparator_0.VBN.n105 comparator_top_0.comparator_0.VBN.n102 26.336
R8 comparator_top_0.comparator_0.VBN.n52 comparator_top_0.comparator_0.VBN.n51 26.336
R9 comparator_top_0.comparator_0.VBN.n38 comparator_top_0.comparator_0.VBN.n35 26.336
R10 comparator_top_0.comparator_0.VBN.n97 comparator_top_0.comparator_0.VBN.n96 15.952
R11 comparator_top_0.comparator_0.VBN.n44 comparator_top_0.comparator_0.VBN.n42 12.8
R12 comparator_top_0.comparator_0.VBN.n44 comparator_top_0.comparator_0.VBN.n43 12.8
R13 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n267 9.3
R14 comparator_top_0.comparator_0.VBN.n273 comparator_top_0.comparator_0.VBN.n272 9.3
R15 comparator_top_0.comparator_0.VBN.n282 comparator_top_0.comparator_0.VBN.n281 9.3
R16 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n276 9.3
R17 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n287 9.3
R18 comparator_top_0.comparator_0.VBN.n302 comparator_top_0.comparator_0.VBN.n301 9.3
R19 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n296 9.3
R20 comparator_top_0.comparator_0.VBN.n293 comparator_top_0.comparator_0.VBN.n292 9.3
R21 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n23 9.3
R22 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n31 9.3
R23 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n40 9.3
R24 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n46 9.3
R25 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n55 9.3
R26 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n63 9.3
R27 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n71 9.3
R28 comparator_top_0.comparator_0.VBN.n15 comparator_top_0.comparator_0.VBN.n79 9.3
R29 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n87 9.3
R30 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n86 9.3
R31 comparator_top_0.comparator_0.VBN.n15 comparator_top_0.comparator_0.VBN.n85 9.3
R32 comparator_top_0.comparator_0.VBN.n85 comparator_top_0.comparator_0.VBN.n84 9.3
R33 comparator_top_0.comparator_0.VBN.n15 comparator_top_0.comparator_0.VBN.n78 9.3
R34 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n77 9.3
R35 comparator_top_0.comparator_0.VBN.n77 comparator_top_0.comparator_0.VBN.n76 9.3
R36 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n70 9.3
R37 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n69 9.3
R38 comparator_top_0.comparator_0.VBN.n69 comparator_top_0.comparator_0.VBN.n68 9.3
R39 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n62 9.3
R40 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n61 9.3
R41 comparator_top_0.comparator_0.VBN.n61 comparator_top_0.comparator_0.VBN.n60 9.3
R42 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n54 9.3
R43 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n53 9.3
R44 comparator_top_0.comparator_0.VBN.n53 comparator_top_0.comparator_0.VBN.n52 9.3
R45 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n45 9.3
R46 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n41 9.3
R47 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n39 9.3
R48 comparator_top_0.comparator_0.VBN.n39 comparator_top_0.comparator_0.VBN.n38 9.3
R49 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n32 9.3
R50 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n30 9.3
R51 comparator_top_0.comparator_0.VBN.n30 comparator_top_0.comparator_0.VBN.n29 9.3
R52 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n24 9.3
R53 comparator_top_0.comparator_0.VBN.n10 comparator_top_0.comparator_0.VBN.n22 9.3
R54 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n155 9.3
R55 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n147 9.3
R56 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n139 9.3
R57 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n131 9.3
R58 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n123 9.3
R59 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n115 9.3
R60 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n107 9.3
R61 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n98 9.3
R62 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n106 9.3
R63 comparator_top_0.comparator_0.VBN.n106 comparator_top_0.comparator_0.VBN.n105 9.3
R64 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n99 9.3
R65 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n108 9.3
R66 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n114 9.3
R67 comparator_top_0.comparator_0.VBN.n114 comparator_top_0.comparator_0.VBN.n113 9.3
R68 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n122 9.3
R69 comparator_top_0.comparator_0.VBN.n122 comparator_top_0.comparator_0.VBN.n121 9.3
R70 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n116 9.3
R71 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n124 9.3
R72 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n130 9.3
R73 comparator_top_0.comparator_0.VBN.n130 comparator_top_0.comparator_0.VBN.n129 9.3
R74 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n138 9.3
R75 comparator_top_0.comparator_0.VBN.n138 comparator_top_0.comparator_0.VBN.n137 9.3
R76 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n132 9.3
R77 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n140 9.3
R78 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n146 9.3
R79 comparator_top_0.comparator_0.VBN.n146 comparator_top_0.comparator_0.VBN.n145 9.3
R80 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n154 9.3
R81 comparator_top_0.comparator_0.VBN.n154 comparator_top_0.comparator_0.VBN.n153 9.3
R82 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n148 9.3
R83 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n156 9.3
R84 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n162 9.3
R85 comparator_top_0.comparator_0.VBN.n162 comparator_top_0.comparator_0.VBN.n161 9.3
R86 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n170 9.3
R87 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n171 9.3
R88 comparator_top_0.comparator_0.VBN.n177 comparator_top_0.comparator_0.VBN.n176 9.3
R89 comparator_top_0.comparator_0.VBN.n92 comparator_top_0.comparator_0.VBN.n91 9.3
R90 comparator_top_0.comparator_0.VBN.n167 comparator_top_0.comparator_0.VBN.n166 9.3
R91 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n315 9.3
R92 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n313 9.3
R93 comparator_top_0.comparator_0.VBN.n313 comparator_top_0.comparator_0.VBN.n312 9.3
R94 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n314 9.3
R95 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n327 9.3
R96 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n326 9.3
R97 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n325 9.3
R98 comparator_top_0.comparator_0.VBN.n325 comparator_top_0.comparator_0.VBN.n324 9.3
R99 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n246 9.3
R100 comparator_top_0.comparator_0.VBN.n252 comparator_top_0.comparator_0.VBN.n251 9.3
R101 comparator_top_0.comparator_0.VBN.n261 comparator_top_0.comparator_0.VBN.n260 9.3
R102 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n255 9.3
R103 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n242 9.3
R104 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n241 9.3
R105 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n243 9.3
R106 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n197 9.3
R107 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n192 9.3
R108 comparator_top_0.comparator_0.VBN.n285 comparator_top_0.comparator_0.VBN.n284 8.764
R109 comparator_top_0.comparator_0.VBN.n305 comparator_top_0.comparator_0.VBN.n304 8.764
R110 comparator_top_0.comparator_0.VBN.n264 comparator_top_0.comparator_0.VBN.n263 8.764
R111 comparator_top_0.comparator_0.VBN.n271 comparator_top_0.comparator_0.VBN.n270 8.215
R112 comparator_top_0.comparator_0.VBN.n280 comparator_top_0.comparator_0.VBN.n279 8.215
R113 comparator_top_0.comparator_0.VBN.n291 comparator_top_0.comparator_0.VBN.n290 8.215
R114 comparator_top_0.comparator_0.VBN.n300 comparator_top_0.comparator_0.VBN.n299 8.215
R115 comparator_top_0.comparator_0.VBN.n311 comparator_top_0.comparator_0.VBN.n310 8.215
R116 comparator_top_0.comparator_0.VBN.n323 comparator_top_0.comparator_0.VBN.n322 8.215
R117 comparator_top_0.comparator_0.VBN.n250 comparator_top_0.comparator_0.VBN.n249 8.215
R118 comparator_top_0.comparator_0.VBN.n259 comparator_top_0.comparator_0.VBN.n258 8.215
R119 comparator_top_0.comparator_0.VBN.n160 comparator_top_0.comparator_0.VBN.n159 7.95
R120 comparator_top_0.comparator_0.VBN.n165 comparator_top_0.comparator_0.VBN.n164 7.95
R121 comparator_top_0.comparator_0.VBN.n105 comparator_top_0.comparator_0.VBN.n104 7.453
R122 comparator_top_0.comparator_0.VBN.n52 comparator_top_0.comparator_0.VBN.n50 7.453
R123 comparator_top_0.comparator_0.VBN.n38 comparator_top_0.comparator_0.VBN.n37 7.453
R124 comparator_top_0.comparator_0.VBN.n152 comparator_top_0.comparator_0.VBN.n151 6.956
R125 comparator_top_0.comparator_0.VBN.n175 comparator_top_0.comparator_0.VBN.n174 6.956
R126 comparator_top_0.comparator_0.VBN.n319 comparator_top_0.comparator_0.VBN.n318 6.922
R127 comparator_top_0.comparator_0.VBN.n307 comparator_top_0.comparator_0.VBN.n306 6.92
R128 comparator_top_0.comparator_0.VBN.n113 comparator_top_0.comparator_0.VBN.n112 6.459
R129 comparator_top_0.comparator_0.VBN.n60 comparator_top_0.comparator_0.VBN.n59 6.459
R130 comparator_top_0.comparator_0.VBN.n29 comparator_top_0.comparator_0.VBN.n28 6.459
R131 comparator_top_0.comparator_0.VBN.n158 comparator_top_0.comparator_0.VBN.n157 6.023
R132 comparator_top_0.comparator_0.VBN.n144 comparator_top_0.comparator_0.VBN.n143 5.962
R133 comparator_top_0.comparator_0.VBN.n90 comparator_top_0.comparator_0.VBN.n89 5.962
R134 comparator_top_0.comparator_0.VBN.n269 comparator_top_0.comparator_0.VBN.n268 5.647
R135 comparator_top_0.comparator_0.VBN.n278 comparator_top_0.comparator_0.VBN.n277 5.647
R136 comparator_top_0.comparator_0.VBN.n289 comparator_top_0.comparator_0.VBN.n288 5.647
R137 comparator_top_0.comparator_0.VBN.n298 comparator_top_0.comparator_0.VBN.n297 5.647
R138 comparator_top_0.comparator_0.VBN.n106 comparator_top_0.comparator_0.VBN.n101 5.647
R139 comparator_top_0.comparator_0.VBN.n53 comparator_top_0.comparator_0.VBN.n48 5.647
R140 comparator_top_0.comparator_0.VBN.n39 comparator_top_0.comparator_0.VBN.n34 5.647
R141 comparator_top_0.comparator_0.VBN.n309 comparator_top_0.comparator_0.VBN.n308 5.647
R142 comparator_top_0.comparator_0.VBN.n321 comparator_top_0.comparator_0.VBN.n320 5.647
R143 comparator_top_0.comparator_0.VBN.n248 comparator_top_0.comparator_0.VBN.n247 5.647
R144 comparator_top_0.comparator_0.VBN.n257 comparator_top_0.comparator_0.VBN.n256 5.647
R145 comparator_top_0.comparator_0.VBN.n210 comparator_top_0.comparator_0.VBN.t6 5.539
R146 comparator_top_0.comparator_0.VBN.n210 comparator_top_0.comparator_0.VBN.t7 5.539
R147 comparator_top_0.comparator_0.VBN.n227 comparator_top_0.comparator_0.VBN.t0 5.539
R148 comparator_top_0.comparator_0.VBN.n227 comparator_top_0.comparator_0.VBN.t5 5.539
R149 comparator_top_0.comparator_0.VBN.n121 comparator_top_0.comparator_0.VBN.n120 5.465
R150 comparator_top_0.comparator_0.VBN.n68 comparator_top_0.comparator_0.VBN.n67 5.465
R151 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n244 5.285
R152 comparator_top_0.comparator_0.VBN.n150 comparator_top_0.comparator_0.VBN.n149 5.27
R153 comparator_top_0.comparator_0.VBN.n136 comparator_top_0.comparator_0.VBN.n135 4.969
R154 comparator_top_0.comparator_0.VBN.n83 comparator_top_0.comparator_0.VBN.n82 4.969
R155 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n266 4.908
R156 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n286 4.908
R157 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n275 4.907
R158 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n254 4.907
R159 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n295 4.906
R160 comparator_top_0.comparator_0.VBN.n114 comparator_top_0.comparator_0.VBN.n110 4.894
R161 comparator_top_0.comparator_0.VBN.n61 comparator_top_0.comparator_0.VBN.n57 4.894
R162 comparator_top_0.comparator_0.VBN.n30 comparator_top_0.comparator_0.VBN.n26 4.894
R163 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n245 4.764
R164 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n44 4.65
R165 comparator_top_0.comparator_0.VBN.n142 comparator_top_0.comparator_0.VBN.n141 4.517
R166 comparator_top_0.comparator_0.VBN.n169 comparator_top_0.comparator_0.VBN.n163 4.517
R167 comparator_top_0.comparator_0.VBN.n195 comparator_top_0.comparator_0.VBN.n194 4.517
R168 comparator_top_0.comparator_0.VBN.n206 comparator_top_0.comparator_0.VBN.n205 4.517
R169 comparator_top_0.comparator_0.VBN.n236 comparator_top_0.comparator_0.VBN.n235 4.517
R170 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n94 4.5
R171 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n182 4.5
R172 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n179 4.5
R173 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n169 4.5
R174 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n274 4.5
R175 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n283 4.5
R176 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n303 4.5
R177 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n294 4.5
R178 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n253 4.5
R179 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n262 4.5
R180 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n195 4.5
R181 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n190 4.5
R182 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n185 4.5
R183 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n239 4.5
R184 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n200 4.5
R185 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n216 4.5
R186 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n204 4.5
R187 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n213 4.5
R188 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n209 4.5
R189 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n226 4.5
R190 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n231 4.5
R191 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n234 4.5
R192 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n220 4.5
R193 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n224 4.5
R194 comparator_top_0.comparator_0.VBN.n129 comparator_top_0.comparator_0.VBN.n128 4.472
R195 comparator_top_0.comparator_0.VBN.n76 comparator_top_0.comparator_0.VBN.n75 4.472
R196 comparator_top_0.comparator_0.VBN.n21 comparator_top_0.comparator_0.VBN.n9 4.443
R197 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n316 7.328
R198 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n329 4.244
R199 comparator_top_0.comparator_0.VBN.n122 comparator_top_0.comparator_0.VBN.n118 4.141
R200 comparator_top_0.comparator_0.VBN.n69 comparator_top_0.comparator_0.VBN.n65 4.141
R201 comparator_top_0.comparator_0.VBN.n128 comparator_top_0.comparator_0.VBN.n127 3.975
R202 comparator_top_0.comparator_0.VBN.n75 comparator_top_0.comparator_0.VBN.n74 3.975
R203 comparator_top_0.comparator_0.VBN.n134 comparator_top_0.comparator_0.VBN.n133 3.764
R204 comparator_top_0.comparator_0.VBN.n179 comparator_top_0.comparator_0.VBN.n173 3.764
R205 comparator_top_0.comparator_0.VBN.n182 comparator_top_0.comparator_0.VBN.n180 3.764
R206 comparator_top_0.comparator_0.VBN.n81 comparator_top_0.comparator_0.VBN.n80 3.764
R207 comparator_top_0.comparator_0.VBN.n239 comparator_top_0.comparator_0.VBN.n238 3.764
R208 comparator_top_0.comparator_0.VBN.n137 comparator_top_0.comparator_0.VBN.n136 3.478
R209 comparator_top_0.comparator_0.VBN.n84 comparator_top_0.comparator_0.VBN.n83 3.478
R210 comparator_top_0.comparator_0.VBN.n20 comparator_top_0.comparator_0.VBN.n307 3.477
R211 comparator_top_0.comparator_0.VBN.n17 comparator_top_0.comparator_0.VBN.n319 3.476
R212 comparator_top_0.comparator_0.VBN.n130 comparator_top_0.comparator_0.VBN.n126 3.388
R213 comparator_top_0.comparator_0.VBN.n77 comparator_top_0.comparator_0.VBN.n73 3.388
R214 comparator_top_0.comparator_0.VBN.n186 comparator_top_0.comparator_0.VBN.t8 3.306
R215 comparator_top_0.comparator_0.VBN.n186 comparator_top_0.comparator_0.VBN.t2 3.306
R216 comparator_top_0.comparator_0.VBN.n190 comparator_top_0.comparator_0.VBN.n188 3.746
R217 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n187 3.158
R218 comparator_top_0.comparator_0.VBN.n2 comparator_top_0.comparator_0.VBN.n285 3.033
R219 comparator_top_0.comparator_0.VBN.n3 comparator_top_0.comparator_0.VBN.n305 3.033
R220 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n264 3.033
R221 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n206 3.033
R222 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n236 3.033
R223 comparator_top_0.comparator_0.VBN.n126 comparator_top_0.comparator_0.VBN.n125 3.011
R224 comparator_top_0.comparator_0.VBN.n94 comparator_top_0.comparator_0.VBN.n88 3.011
R225 comparator_top_0.comparator_0.VBN.n73 comparator_top_0.comparator_0.VBN.n72 3.011
R226 comparator_top_0.comparator_0.VBN.n190 comparator_top_0.comparator_0.VBN.n189 3.011
R227 comparator_top_0.comparator_0.VBN.n120 comparator_top_0.comparator_0.VBN.n119 2.981
R228 comparator_top_0.comparator_0.VBN.n67 comparator_top_0.comparator_0.VBN.n66 2.981
R229 comparator_top_0.comparator_0.VBN.n138 comparator_top_0.comparator_0.VBN.n134 2.635
R230 comparator_top_0.comparator_0.VBN.n85 comparator_top_0.comparator_0.VBN.n81 2.635
R231 comparator_top_0.comparator_0.VBN.n239 comparator_top_0.comparator_0.VBN.n237 2.635
R232 comparator_top_0.comparator_0.VBN.n204 comparator_top_0.comparator_0.VBN.n202 2.635
R233 comparator_top_0.comparator_0.VBN.n224 comparator_top_0.comparator_0.VBN.n222 2.635
R234 comparator_top_0.comparator_0.VBN.n192 comparator_top_0.comparator_0.VBN.n191 2.616
R235 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n198 2.604
R236 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n218 2.604
R237 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n183 2.525
R238 comparator_top_0.comparator_0.VBN.n145 comparator_top_0.comparator_0.VBN.n144 2.484
R239 comparator_top_0.comparator_0.VBN.n91 comparator_top_0.comparator_0.VBN.n90 2.484
R240 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n17 2.423
R241 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n20 2.395
R242 comparator_top_0.comparator_0.VBN.n118 comparator_top_0.comparator_0.VBN.n117 2.258
R243 comparator_top_0.comparator_0.VBN.n65 comparator_top_0.comparator_0.VBN.n64 2.258
R244 comparator_top_0.comparator_0.VBN.n216 comparator_top_0.comparator_0.VBN.n214 2.258
R245 comparator_top_0.comparator_0.VBN.n208 comparator_top_0.comparator_0.VBN.n207 2.258
R246 comparator_top_0.comparator_0.VBN.n234 comparator_top_0.comparator_0.VBN.n232 2.258
R247 comparator_top_0.comparator_0.VBN.n230 comparator_top_0.comparator_0.VBN.n229 2.258
R248 comparator_top_0.comparator_0.VBN.n216 comparator_top_0.comparator_0.VBN.n215 2.252
R249 comparator_top_0.comparator_0.VBN.n234 comparator_top_0.comparator_0.VBN.n233 2.252
R250 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN.n317 2.25
R251 comparator_top_0.comparator_0.VBN.n197 comparator_top_0.comparator_0.VBN.n196 2.246
R252 comparator_top_0.comparator_0.VBN.n265 comparator_top_0.comparator_0.VBN.n18 2.069
R253 comparator_top_0.comparator_bias_0.VBN comparator_top_0.comparator_0.VBN.n19 2.068
R254 comparator_top_0.comparator_0.VBN.n112 comparator_top_0.comparator_0.VBN.n111 1.987
R255 comparator_top_0.comparator_0.VBN.n59 comparator_top_0.comparator_0.VBN.n58 1.987
R256 comparator_top_0.comparator_0.VBN.n28 comparator_top_0.comparator_0.VBN.n27 1.987
R257 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n172 1.94
R258 comparator_top_0.comparator_0.VBN.n146 comparator_top_0.comparator_0.VBN.n142 1.882
R259 comparator_top_0.comparator_0.VBN.n93 comparator_top_0.comparator_0.VBN.n92 1.882
R260 comparator_top_0.comparator_0.VBN.n195 comparator_top_0.comparator_0.VBN.n193 1.882
R261 comparator_top_0.comparator_0.VBN.n204 comparator_top_0.comparator_0.VBN.n203 1.878
R262 comparator_top_0.comparator_0.VBN.n224 comparator_top_0.comparator_0.VBN.n223 1.878
R263 comparator_top_0.comparator_0.VBN.n265 comparator_top_0.comparator_0.VBN.n2 1.841
R264 comparator_top_0.comparator_0.VBN.n217 comparator_top_0.comparator_0.VBN.n1 1.738
R265 comparator_top_0.comparator_0.VBN.n21 comparator_top_0.comparator_0.VBN.n172 1.701
R266 comparator_top_0.comparator_0.VBN.n19 comparator_top_0.comparator_0.VBN.n3 1.693
R267 comparator_top_0.comparator_0.VBN.n8 comparator_top_0.comparator_0.VBN.n186 1.615
R268 comparator_top_0.comparator_0.VBN.n95 comparator_top_0.comparator_0.VBN.t3 1.606
R269 comparator_top_0.comparator_0.VBN.n9 comparator_top_0.comparator_0.VBN 1.601
R270 comparator_top_0.comparator_0.VBN.n110 comparator_top_0.comparator_0.VBN.n109 1.505
R271 comparator_top_0.comparator_0.VBN.n169 comparator_top_0.comparator_0.VBN.n168 1.505
R272 comparator_top_0.comparator_0.VBN.n179 comparator_top_0.comparator_0.VBN.n178 1.505
R273 comparator_top_0.comparator_0.VBN.n94 comparator_top_0.comparator_0.VBN.n93 1.505
R274 comparator_top_0.comparator_0.VBN.n57 comparator_top_0.comparator_0.VBN.n56 1.505
R275 comparator_top_0.comparator_0.VBN.n26 comparator_top_0.comparator_0.VBN.n25 1.505
R276 comparator_top_0.comparator_0.VBN.n213 comparator_top_0.comparator_0.VBN.n212 1.505
R277 comparator_top_0.comparator_0.VBN.n226 comparator_top_0.comparator_0.VBN.n225 1.505
R278 comparator_top_0.comparator_0.VBN.n228 comparator_top_0.comparator_0.VBN.n227 1.5
R279 comparator_top_0.comparator_0.VBN.n211 comparator_top_0.comparator_0.VBN.n210 1.5
R280 comparator_top_0.comparator_0.VBN.n153 comparator_top_0.comparator_0.VBN.n152 1.49
R281 comparator_top_0.comparator_0.VBN.n176 comparator_top_0.comparator_0.VBN.n175 1.49
R282 comparator_top_0.comparator_0.VBN.n19 comparator_top_0.comparator_0.VBN.n265 1.259
R283 comparator_top_0.comparator_0.VBN.n217 comparator_top_0.comparator_0.VBN.n0 1.196
R284 comparator_top_0.comparator_0.VBN.n19 comparator_top_0.comparator_0.VBN.n21 1.153
R285 comparator_top_0.comparator_0.VBN.n154 comparator_top_0.comparator_0.VBN.n150 1.129
R286 comparator_top_0.comparator_0.VBN.n178 comparator_top_0.comparator_0.VBN.n177 1.129
R287 comparator_top_0.comparator_0.VBN.n185 comparator_top_0.comparator_0.VBN.n184 1.129
R288 comparator_top_0.comparator_0.VBN.n272 comparator_top_0.comparator_0.VBN.n271 1.095
R289 comparator_top_0.comparator_0.VBN.n281 comparator_top_0.comparator_0.VBN.n280 1.095
R290 comparator_top_0.comparator_0.VBN.n292 comparator_top_0.comparator_0.VBN.n291 1.095
R291 comparator_top_0.comparator_0.VBN.n301 comparator_top_0.comparator_0.VBN.n300 1.095
R292 comparator_top_0.comparator_0.VBN.n312 comparator_top_0.comparator_0.VBN.n311 1.095
R293 comparator_top_0.comparator_0.VBN.n324 comparator_top_0.comparator_0.VBN.n323 1.095
R294 comparator_top_0.comparator_0.VBN.n251 comparator_top_0.comparator_0.VBN.n250 1.095
R295 comparator_top_0.comparator_0.VBN.n260 comparator_top_0.comparator_0.VBN.n259 1.095
R296 comparator_top_0.comparator_0.VBN.n14 comparator_top_0.comparator_0.VBN.n97 1.031
R297 comparator_top_0.comparator_0.VBN.n104 comparator_top_0.comparator_0.VBN.n103 0.993
R298 comparator_top_0.comparator_0.VBN.n50 comparator_top_0.comparator_0.VBN.n49 0.993
R299 comparator_top_0.comparator_0.VBN.n37 comparator_top_0.comparator_0.VBN.n36 0.993
R300 comparator_top_0.comparator_0.VBN.n183 comparator_top_0.comparator_0.VBN.n217 0.885
R301 comparator_top_0.comparator_0.VBN.n1 comparator_top_0.comparator_0.VBN.n211 0.821
R302 comparator_top_0.comparator_0.VBN.n0 comparator_top_0.comparator_0.VBN.n228 0.821
R303 comparator_top_0.comparator_0.VBN.n274 comparator_top_0.comparator_0.VBN.n273 0.752
R304 comparator_top_0.comparator_0.VBN.n273 comparator_top_0.comparator_0.VBN.n269 0.752
R305 comparator_top_0.comparator_0.VBN.n282 comparator_top_0.comparator_0.VBN.n278 0.752
R306 comparator_top_0.comparator_0.VBN.n283 comparator_top_0.comparator_0.VBN.n282 0.752
R307 comparator_top_0.comparator_0.VBN.n294 comparator_top_0.comparator_0.VBN.n293 0.752
R308 comparator_top_0.comparator_0.VBN.n293 comparator_top_0.comparator_0.VBN.n289 0.752
R309 comparator_top_0.comparator_0.VBN.n302 comparator_top_0.comparator_0.VBN.n298 0.752
R310 comparator_top_0.comparator_0.VBN.n303 comparator_top_0.comparator_0.VBN.n302 0.752
R311 comparator_top_0.comparator_0.VBN.n101 comparator_top_0.comparator_0.VBN.n100 0.752
R312 comparator_top_0.comparator_0.VBN.n48 comparator_top_0.comparator_0.VBN.n47 0.752
R313 comparator_top_0.comparator_0.VBN.n34 comparator_top_0.comparator_0.VBN.n33 0.752
R314 comparator_top_0.comparator_0.VBN.n313 comparator_top_0.comparator_0.VBN.n309 0.752
R315 comparator_top_0.comparator_0.VBN.n325 comparator_top_0.comparator_0.VBN.n321 0.752
R316 comparator_top_0.comparator_0.VBN.n253 comparator_top_0.comparator_0.VBN.n252 0.752
R317 comparator_top_0.comparator_0.VBN.n252 comparator_top_0.comparator_0.VBN.n248 0.752
R318 comparator_top_0.comparator_0.VBN.n261 comparator_top_0.comparator_0.VBN.n257 0.752
R319 comparator_top_0.comparator_0.VBN.n262 comparator_top_0.comparator_0.VBN.n261 0.752
R320 comparator_top_0.comparator_0.VBN.n200 comparator_top_0.comparator_0.VBN.n199 0.752
R321 comparator_top_0.comparator_0.VBN.n209 comparator_top_0.comparator_0.VBN.n208 0.752
R322 comparator_top_0.comparator_0.VBN.n220 comparator_top_0.comparator_0.VBN.n219 0.752
R323 comparator_top_0.comparator_0.VBN.n231 comparator_top_0.comparator_0.VBN.n230 0.752
R324 comparator_top_0.comparator_0.VBN.n329 comparator_top_0.comparator_0.VBN.n328 0.738
R325 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n15 0.691
R326 comparator_top_0.comparator_0.VBN.n5 comparator_top_0.comparator_0.VBN.n4 0.628
R327 comparator_top_0.comparator_0.VBN.n4 comparator_top_0.comparator_0.VBN.n8 0.607
R328 comparator_top_0.comparator_0.VBN.n6 comparator_top_0.comparator_0.VBN.n12 0.568
R329 comparator_top_0.comparator_0.VBN.n161 comparator_top_0.comparator_0.VBN.n160 0.496
R330 comparator_top_0.comparator_0.VBN.n166 comparator_top_0.comparator_0.VBN.n165 0.496
R331 comparator_top_0.comparator_0.VBN.n18 comparator_top_0.comparator_0.VBN.n5 0.487
R332 comparator_top_0.comparator_0.VBN.n241 comparator_top_0.comparator_0.VBN.n240 0.461
R333 comparator_top_0.comparator_0.VBN.n11 comparator_top_0.comparator_0.VBN.n10 0.423
R334 comparator_top_0.comparator_0.VBN.n13 comparator_top_0.comparator_0.VBN.n11 0.38
R335 comparator_top_0.comparator_0.VBN.n7 comparator_top_0.comparator_0.VBN.n6 0.379
R336 comparator_top_0.comparator_0.VBN.n15 comparator_top_0.comparator_0.VBN.n16 0.378
R337 comparator_top_0.comparator_0.VBN.n12 comparator_top_0.comparator_0.VBN.n14 0.378
R338 comparator_top_0.comparator_0.VBN.n16 comparator_top_0.comparator_0.VBN.n13 0.378
R339 comparator_top_0.comparator_0.VBN.n162 comparator_top_0.comparator_0.VBN.n158 0.376
R340 comparator_top_0.comparator_0.VBN.n168 comparator_top_0.comparator_0.VBN.n167 0.376
R341 comparator_top_0.comparator_0.VBN.n182 comparator_top_0.comparator_0.VBN.n181 0.376
R342 comparator_top_0.comparator_0.VBN.n202 comparator_top_0.comparator_0.VBN.n201 0.376
R343 comparator_top_0.comparator_0.VBN.n222 comparator_top_0.comparator_0.VBN.n221 0.376
R344 a_1821_8526.n114 a_1821_8526.t2 116.84
R345 a_1821_8526.n65 a_1821_8526.t3 116.84
R346 a_1821_8526.n196 a_1821_8526.t6 60.25
R347 a_1821_8526.n175 a_1821_8526.t9 60.25
R348 a_1821_8526.n155 a_1821_8526.t7 60.25
R349 a_1821_8526.n135 a_1821_8526.t8 60.25
R350 a_1821_8526.n118 a_1821_8526.n117 52.689
R351 a_1821_8526.n69 a_1821_8526.n68 52.689
R352 a_1821_8526.n126 a_1821_8526.n125 46.103
R353 a_1821_8526.n77 a_1821_8526.n76 46.103
R354 a_1821_8526.n87 a_1821_8526.n86 39.517
R355 a_1821_8526.n38 a_1821_8526.n37 39.517
R356 a_1821_8526.n94 a_1821_8526.n93 32.931
R357 a_1821_8526.n45 a_1821_8526.n44 32.931
R358 a_1821_8526.n107 a_1821_8526.n106 29.637
R359 a_1821_8526.n56 a_1821_8526.n55 29.637
R360 a_1821_8526.n34 a_1821_8526.t1 27.695
R361 a_1821_8526.n106 a_1821_8526.n105 26.344
R362 a_1821_8526.n55 a_1821_8526.n54 26.344
R363 a_1821_8526.n95 a_1821_8526.n94 23.051
R364 a_1821_8526.n46 a_1821_8526.n45 23.051
R365 a_1821_8526.n88 a_1821_8526.n87 16.465
R366 a_1821_8526.n39 a_1821_8526.n38 16.465
R367 a_1821_8526.n32 a_1821_8526.n31 13.176
R368 a_1821_8526.n127 a_1821_8526.n126 9.879
R369 a_1821_8526.n78 a_1821_8526.n77 9.879
R370 a_1821_8526.n10 a_1821_8526.n28 9.316
R371 a_1821_8526.n11 a_1821_8526.n121 9.3
R372 a_1821_8526.n1 a_1821_8526.n129 9.3
R373 a_1821_8526.n11 a_1821_8526.n120 9.3
R374 a_1821_8526.n120 a_1821_8526.n119 9.3
R375 a_1821_8526.n11 a_1821_8526.n122 9.3
R376 a_1821_8526.n1 a_1821_8526.n128 9.3
R377 a_1821_8526.n128 a_1821_8526.n127 9.3
R378 a_1821_8526.n89 a_1821_8526.n88 9.3
R379 a_1821_8526.n1 a_1821_8526.n111 9.3
R380 a_1821_8526.n1 a_1821_8526.n108 9.3
R381 a_1821_8526.n108 a_1821_8526.n107 9.3
R382 a_1821_8526.n96 a_1821_8526.n95 9.3
R383 a_1821_8526.n12 a_1821_8526.n72 9.3
R384 a_1821_8526.n0 a_1821_8526.n80 9.3
R385 a_1821_8526.n12 a_1821_8526.n71 9.3
R386 a_1821_8526.n71 a_1821_8526.n70 9.3
R387 a_1821_8526.n12 a_1821_8526.n73 9.3
R388 a_1821_8526.n0 a_1821_8526.n79 9.3
R389 a_1821_8526.n79 a_1821_8526.n78 9.3
R390 a_1821_8526.n0 a_1821_8526.n57 9.3
R391 a_1821_8526.n57 a_1821_8526.n56 9.3
R392 a_1821_8526.n0 a_1821_8526.n60 9.3
R393 a_1821_8526.n47 a_1821_8526.n46 9.3
R394 a_1821_8526.n40 a_1821_8526.n39 9.3
R395 a_1821_8526.n10 a_1821_8526.n35 9.3
R396 a_1821_8526.n9 a_1821_8526.n143 9.3
R397 a_1821_8526.n9 a_1821_8526.n144 9.3
R398 a_1821_8526.n9 a_1821_8526.n142 9.3
R399 a_1821_8526.n142 a_1821_8526.n141 9.3
R400 a_1821_8526.n7 a_1821_8526.n148 9.3
R401 a_1821_8526.n8 a_1821_8526.n163 9.3
R402 a_1821_8526.n8 a_1821_8526.n164 9.3
R403 a_1821_8526.n8 a_1821_8526.n162 9.3
R404 a_1821_8526.n162 a_1821_8526.n161 9.3
R405 a_1821_8526.n7 a_1821_8526.n154 9.3
R406 a_1821_8526.n154 a_1821_8526.n153 9.3
R407 a_1821_8526.n7 a_1821_8526.n147 9.3
R408 a_1821_8526.n5 a_1821_8526.n168 9.3
R409 a_1821_8526.n6 a_1821_8526.n183 9.3
R410 a_1821_8526.n6 a_1821_8526.n184 9.3
R411 a_1821_8526.n6 a_1821_8526.n182 9.3
R412 a_1821_8526.n182 a_1821_8526.n181 9.3
R413 a_1821_8526.n5 a_1821_8526.n174 9.3
R414 a_1821_8526.n174 a_1821_8526.n173 9.3
R415 a_1821_8526.n5 a_1821_8526.n167 9.3
R416 a_1821_8526.n4 a_1821_8526.n188 9.3
R417 a_1821_8526.n13 a_1821_8526.n195 9.3
R418 a_1821_8526.n13 a_1821_8526.n197 9.3
R419 a_1821_8526.n4 a_1821_8526.n194 9.3
R420 a_1821_8526.n194 a_1821_8526.n193 9.3
R421 a_1821_8526.n4 a_1821_8526.n187 9.3
R422 a_1821_8526.n204 a_1821_8526.n203 9.3
R423 a_1821_8526.n210 a_1821_8526.n206 9.3
R424 a_1821_8526.n210 a_1821_8526.n209 9.3
R425 a_1821_8526.n35 a_1821_8526.n34 9.02
R426 a_1821_8526.n156 a_1821_8526.n155 8.764
R427 a_1821_8526.n176 a_1821_8526.n175 8.764
R428 a_1821_8526.n197 a_1821_8526.n196 8.764
R429 a_1821_8526.n14 a_1821_8526.t5 7.506
R430 a_1821_8526.n202 a_1821_8526.n201 7.453
R431 a_1821_8526.n192 a_1821_8526.n191 7.453
R432 a_1821_8526.n180 a_1821_8526.n179 7.453
R433 a_1821_8526.n172 a_1821_8526.n171 7.453
R434 a_1821_8526.n160 a_1821_8526.n159 7.453
R435 a_1821_8526.n152 a_1821_8526.n151 7.453
R436 a_1821_8526.n140 a_1821_8526.n139 7.453
R437 a_1821_8526.n136 a_1821_8526.n135 6.8
R438 a_1821_8526.n116 a_1821_8526.n115 6.023
R439 a_1821_8526.n67 a_1821_8526.n66 6.023
R440 a_1821_8526.n190 a_1821_8526.n189 5.647
R441 a_1821_8526.n178 a_1821_8526.n177 5.647
R442 a_1821_8526.n170 a_1821_8526.n169 5.647
R443 a_1821_8526.n158 a_1821_8526.n157 5.647
R444 a_1821_8526.n150 a_1821_8526.n149 5.647
R445 a_1821_8526.n138 a_1821_8526.n137 5.647
R446 a_1821_8526.n210 a_1821_8526.t4 5.539
R447 a_1821_8526.t0 a_1821_8526.n210 5.539
R448 a_1821_8526.n124 a_1821_8526.n123 5.27
R449 a_1821_8526.n75 a_1821_8526.n74 5.27
R450 a_1821_8526.n1 a_1821_8526.n104 5.264
R451 a_1821_8526.n0 a_1821_8526.n53 5.264
R452 a_1821_8526.n4 a_1821_8526.n186 4.735
R453 a_1821_8526.n5 a_1821_8526.n166 4.735
R454 a_1821_8526.n7 a_1821_8526.n146 4.735
R455 a_1821_8526.n6 a_1821_8526.n185 4.735
R456 a_1821_8526.n8 a_1821_8526.n165 4.735
R457 a_1821_8526.n9 a_1821_8526.n145 4.735
R458 a_1821_8526.n7 a_1821_8526.n156 4.65
R459 a_1821_8526.n5 a_1821_8526.n176 4.65
R460 a_1821_8526.n2 a_1821_8526.n17 4.63
R461 a_1821_8526.n15 a_1821_8526.n134 6.761
R462 a_1821_8526.n113 a_1821_8526.n112 4.517
R463 a_1821_8526.n64 a_1821_8526.n63 4.517
R464 a_1821_8526.n26 a_1821_8526.n25 4.517
R465 a_1821_8526.n1 a_1821_8526.n131 4.5
R466 a_1821_8526.n1 a_1821_8526.n103 4.5
R467 a_1821_8526.n0 a_1821_8526.n52 4.5
R468 a_1821_8526.n0 a_1821_8526.n82 4.5
R469 a_1821_8526.n10 a_1821_8526.n30 4.5
R470 a_1821_8526.n10 a_1821_8526.n33 4.5
R471 a_1821_8526.n13 a_1821_8526.n198 4.5
R472 a_1821_8526.n199 a_1821_8526.n205 4.5
R473 a_1821_8526.n1 a_1821_8526.n101 4.5
R474 a_1821_8526.n1 a_1821_8526.n99 4.5
R475 a_1821_8526.n1 a_1821_8526.n91 4.5
R476 a_1821_8526.n0 a_1821_8526.n62 4.5
R477 a_1821_8526.n0 a_1821_8526.n50 4.5
R478 a_1821_8526.n0 a_1821_8526.n42 4.5
R479 a_1821_8526.n2 a_1821_8526.n20 4.5
R480 a_1821_8526.n2 a_1821_8526.n24 4.5
R481 a_1821_8526.n210 a_1821_8526.n16 4.357
R482 a_1821_8526.n11 a_1821_8526.n114 4.235
R483 a_1821_8526.n12 a_1821_8526.n65 4.235
R484 a_1821_8526.n91 a_1821_8526.n85 4.141
R485 a_1821_8526.n42 a_1821_8526.n36 4.141
R486 a_1821_8526.n205 a_1821_8526.n204 4.141
R487 a_1821_8526.n134 a_1821_8526.n132 3.764
R488 a_1821_8526.n9 a_1821_8526.n136 3.427
R489 a_1821_8526.n99 a_1821_8526.n92 3.388
R490 a_1821_8526.n50 a_1821_8526.n43 3.388
R491 a_1821_8526.n24 a_1821_8526.n21 3.388
R492 a_1821_8526.n208 a_1821_8526.n207 3.384
R493 a_1821_8526.n119 a_1821_8526.n118 3.293
R494 a_1821_8526.n70 a_1821_8526.n69 3.293
R495 a_1821_8526.n1 a_1821_8526.n113 3.033
R496 a_1821_8526.n0 a_1821_8526.n64 3.033
R497 a_1821_8526.n3 a_1821_8526.n26 3.033
R498 a_1821_8526.n110 a_1821_8526.n109 3.011
R499 a_1821_8526.n59 a_1821_8526.n58 3.011
R500 a_1821_8526.n98 a_1821_8526.n97 2.258
R501 a_1821_8526.n49 a_1821_8526.n48 2.258
R502 a_1821_8526.n205 a_1821_8526.n200 2.258
R503 a_1821_8526.n23 a_1821_8526.n22 2.258
R504 a_1821_8526.n15 a_1821_8526.n13 2.257
R505 a_1821_8526.n15 a_1821_8526.n199 2.29
R506 a_1821_8526.n83 a_1821_8526.n27 1.907
R507 a_1821_8526.n90 a_1821_8526.n89 1.882
R508 a_1821_8526.n111 a_1821_8526.n110 1.882
R509 a_1821_8526.n41 a_1821_8526.n40 1.882
R510 a_1821_8526.n60 a_1821_8526.n59 1.882
R511 a_1821_8526.n134 a_1821_8526.n133 1.882
R512 a_1821_8526.n210 a_1821_8526.n3 1.717
R513 a_1821_8526.n27 a_1821_8526.n10 1.666
R514 a_1821_8526.n103 a_1821_8526.n102 1.505
R515 a_1821_8526.n52 a_1821_8526.n51 1.505
R516 a_1821_8526.n209 a_1821_8526.n208 1.505
R517 a_1821_8526.n17 a_1821_8526.n18 1.505
R518 a_1821_8526.n128 a_1821_8526.n124 1.129
R519 a_1821_8526.n79 a_1821_8526.n75 1.129
R520 a_1821_8526.n83 a_1821_8526.n0 1.078
R521 a_1821_8526.n203 a_1821_8526.n202 0.993
R522 a_1821_8526.n193 a_1821_8526.n192 0.993
R523 a_1821_8526.n181 a_1821_8526.n180 0.993
R524 a_1821_8526.n173 a_1821_8526.n172 0.993
R525 a_1821_8526.n161 a_1821_8526.n160 0.993
R526 a_1821_8526.n153 a_1821_8526.n152 0.993
R527 a_1821_8526.n141 a_1821_8526.n140 0.993
R528 a_1821_8526.n3 a_1821_8526.n14 0.895
R529 a_1821_8526.n131 a_1821_8526.n130 0.752
R530 a_1821_8526.n101 a_1821_8526.n100 0.752
R531 a_1821_8526.n82 a_1821_8526.n81 0.752
R532 a_1821_8526.n62 a_1821_8526.n61 0.752
R533 a_1821_8526.n194 a_1821_8526.n190 0.752
R534 a_1821_8526.n182 a_1821_8526.n178 0.752
R535 a_1821_8526.n174 a_1821_8526.n170 0.752
R536 a_1821_8526.n162 a_1821_8526.n158 0.752
R537 a_1821_8526.n154 a_1821_8526.n150 0.752
R538 a_1821_8526.n142 a_1821_8526.n138 0.752
R539 a_1821_8526.n20 a_1821_8526.n19 0.752
R540 a_1821_8526.n84 a_1821_8526.n1 0.737
R541 a_1821_8526.n14 a_1821_8526.n84 0.716
R542 a_1821_8526.n1 a_1821_8526.n11 0.662
R543 a_1821_8526.n0 a_1821_8526.n12 0.662
R544 a_1821_8526.n7 a_1821_8526.n9 0.66
R545 a_1821_8526.n5 a_1821_8526.n8 0.66
R546 a_1821_8526.n4 a_1821_8526.n6 0.66
R547 a_1821_8526.n8 a_1821_8526.n7 0.583
R548 a_1821_8526.n6 a_1821_8526.n5 0.583
R549 a_1821_8526.n14 a_1821_8526.n83 0.532
R550 a_1821_8526.n3 a_1821_8526.n2 0.456
R551 a_1821_8526.n13 a_1821_8526.n4 0.442
R552 a_1821_8526.n84 a_1821_8526.n15 0.388
R553 a_1821_8526.n120 a_1821_8526.n116 0.376
R554 a_1821_8526.n91 a_1821_8526.n90 0.376
R555 a_1821_8526.n99 a_1821_8526.n98 0.376
R556 a_1821_8526.n97 a_1821_8526.n96 0.376
R557 a_1821_8526.n71 a_1821_8526.n67 0.376
R558 a_1821_8526.n42 a_1821_8526.n41 0.376
R559 a_1821_8526.n50 a_1821_8526.n49 0.376
R560 a_1821_8526.n48 a_1821_8526.n47 0.376
R561 a_1821_8526.n30 a_1821_8526.n29 0.376
R562 a_1821_8526.n33 a_1821_8526.n32 0.376
R563 a_1821_8526.n24 a_1821_8526.n23 0.376
R564 vdd3p3.n3386 vdd3p3.t124 840.188
R565 vdd3p3.n3386 vdd3p3.t137 840.188
R566 vdd3p3.n3383 vdd3p3.t125 403.572
R567 vdd3p3.n3382 vdd3p3.t138 403.572
R568 vdd3p3.n2844 vdd3p3.n2628 373.448
R569 vdd3p3.n2864 vdd3p3.n2632 373.448
R570 vdd3p3.n3163 vdd3p3.n3162 373.448
R571 vdd3p3.n3179 vdd3p3.n3021 373.448
R572 vdd3p3.n1998 vdd3p3.n1782 373.448
R573 vdd3p3.n2018 vdd3p3.n1786 373.448
R574 vdd3p3.n2317 vdd3p3.n2316 373.448
R575 vdd3p3.n2333 vdd3p3.n2175 373.448
R576 vdd3p3.n1153 vdd3p3.n937 373.448
R577 vdd3p3.n1173 vdd3p3.n941 373.448
R578 vdd3p3.n1472 vdd3p3.n1471 373.448
R579 vdd3p3.n1488 vdd3p3.n1330 373.448
R580 vdd3p3.n307 vdd3p3.n91 373.448
R581 vdd3p3.n327 vdd3p3.n95 373.448
R582 vdd3p3.n626 vdd3p3.n625 373.448
R583 vdd3p3.n642 vdd3p3.n484 373.448
R584 vdd3p3.n3099 vdd3p3.n3037 351.827
R585 vdd3p3.n3120 vdd3p3.n3119 351.827
R586 vdd3p3.n3342 vdd3p3.n2668 351.827
R587 vdd3p3.n3322 vdd3p3.n2664 351.827
R588 vdd3p3.n2253 vdd3p3.n2191 351.827
R589 vdd3p3.n2274 vdd3p3.n2273 351.827
R590 vdd3p3.n2496 vdd3p3.n1822 351.827
R591 vdd3p3.n2476 vdd3p3.n1818 351.827
R592 vdd3p3.n1408 vdd3p3.n1346 351.827
R593 vdd3p3.n1429 vdd3p3.n1428 351.827
R594 vdd3p3.n1651 vdd3p3.n977 351.827
R595 vdd3p3.n1631 vdd3p3.n973 351.827
R596 vdd3p3.n562 vdd3p3.n500 351.827
R597 vdd3p3.n583 vdd3p3.n582 351.827
R598 vdd3p3.n805 vdd3p3.n131 351.827
R599 vdd3p3.n785 vdd3p3.n127 351.827
R600 vdd3p3.n52 vdd3p3.n34 321.882
R601 vdd3p3.n38 vdd3p3.n33 321.882
R602 vdd3p3.n15 vdd3p3.n7 321.882
R603 vdd3p3.n28 vdd3p3.n7 321.882
R604 vdd3p3.n28 vdd3p3.n5 321.882
R605 vdd3p3.n57 vdd3p3.n5 321.882
R606 vdd3p3.n894 vdd3p3.n887 321.882
R607 vdd3p3.n886 vdd3p3.n848 321.882
R608 vdd3p3.n866 vdd3p3.n857 321.882
R609 vdd3p3.n869 vdd3p3.n857 321.882
R610 vdd3p3.n869 vdd3p3.n850 321.882
R611 vdd3p3.n882 vdd3p3.n850 321.882
R612 vdd3p3.n1743 vdd3p3.n1725 321.882
R613 vdd3p3.n1729 vdd3p3.n1724 321.882
R614 vdd3p3.n1706 vdd3p3.n1698 321.882
R615 vdd3p3.n1719 vdd3p3.n1698 321.882
R616 vdd3p3.n1719 vdd3p3.n1696 321.882
R617 vdd3p3.n1748 vdd3p3.n1696 321.882
R618 vdd3p3.n2585 vdd3p3.n2578 321.882
R619 vdd3p3.n2577 vdd3p3.n2539 321.882
R620 vdd3p3.n2557 vdd3p3.n2548 321.882
R621 vdd3p3.n2560 vdd3p3.n2548 321.882
R622 vdd3p3.n2560 vdd3p3.n2541 321.882
R623 vdd3p3.n2573 vdd3p3.n2541 321.882
R624 vdd3p3.n56 vdd3p3.n55 266.73
R625 vdd3p3.n884 vdd3p3.n883 266.73
R626 vdd3p3.n1747 vdd3p3.n1746 266.73
R627 vdd3p3.n2575 vdd3p3.n2574 266.73
R628 vdd3p3.n903 vdd3p3.t112 240.531
R629 vdd3p3.n2594 vdd3p3.t94 240.531
R630 vdd3p3.n3075 vdd3p3.n3072 239.793
R631 vdd3p3.n3072 vdd3p3.n3071 239.793
R632 vdd3p3.n3056 vdd3p3.n3047 239.793
R633 vdd3p3.n3056 vdd3p3.n3055 239.793
R634 vdd3p3.n3079 vdd3p3.n2609 239.793
R635 vdd3p3.n2638 vdd3p3.n2620 239.793
R636 vdd3p3.n3082 vdd3p3.n2612 239.793
R637 vdd3p3.n2660 vdd3p3.n2642 239.793
R638 vdd3p3.n2229 vdd3p3.n2226 239.793
R639 vdd3p3.n2226 vdd3p3.n2225 239.793
R640 vdd3p3.n2210 vdd3p3.n2201 239.793
R641 vdd3p3.n2210 vdd3p3.n2209 239.793
R642 vdd3p3.n2233 vdd3p3.n1763 239.793
R643 vdd3p3.n1792 vdd3p3.n1774 239.793
R644 vdd3p3.n2236 vdd3p3.n1766 239.793
R645 vdd3p3.n1814 vdd3p3.n1796 239.793
R646 vdd3p3.n1384 vdd3p3.n1381 239.793
R647 vdd3p3.n1381 vdd3p3.n1380 239.793
R648 vdd3p3.n1365 vdd3p3.n1356 239.793
R649 vdd3p3.n1365 vdd3p3.n1364 239.793
R650 vdd3p3.n1388 vdd3p3.n918 239.793
R651 vdd3p3.n947 vdd3p3.n929 239.793
R652 vdd3p3.n1391 vdd3p3.n921 239.793
R653 vdd3p3.n969 vdd3p3.n951 239.793
R654 vdd3p3.n538 vdd3p3.n535 239.793
R655 vdd3p3.n535 vdd3p3.n534 239.793
R656 vdd3p3.n519 vdd3p3.n510 239.793
R657 vdd3p3.n519 vdd3p3.n518 239.793
R658 vdd3p3.n542 vdd3p3.n72 239.793
R659 vdd3p3.n101 vdd3p3.n83 239.793
R660 vdd3p3.n545 vdd3p3.n75 239.793
R661 vdd3p3.n123 vdd3p3.n105 239.793
R662 vdd3p3.n45 vdd3p3.t109 239.694
R663 vdd3p3.n1736 vdd3p3.t164 239.694
R664 vdd3p3.n3079 vdd3p3.n3078 218.172
R665 vdd3p3.n3351 vdd3p3.n2638 218.172
R666 vdd3p3.n3125 vdd3p3.n3082 218.172
R667 vdd3p3.n3349 vdd3p3.n2642 218.172
R668 vdd3p3.n2233 vdd3p3.n2232 218.172
R669 vdd3p3.n2505 vdd3p3.n1792 218.172
R670 vdd3p3.n2279 vdd3p3.n2236 218.172
R671 vdd3p3.n2503 vdd3p3.n1796 218.172
R672 vdd3p3.n1388 vdd3p3.n1387 218.172
R673 vdd3p3.n1660 vdd3p3.n947 218.172
R674 vdd3p3.n1434 vdd3p3.n1391 218.172
R675 vdd3p3.n1658 vdd3p3.n951 218.172
R676 vdd3p3.n542 vdd3p3.n541 218.172
R677 vdd3p3.n814 vdd3p3.n101 218.172
R678 vdd3p3.n588 vdd3p3.n545 218.172
R679 vdd3p3.n812 vdd3p3.n105 218.172
R680 vdd3p3.n54 vdd3p3.t108 217.947
R681 vdd3p3.n896 vdd3p3.t111 217.947
R682 vdd3p3.n1745 vdd3p3.t163 217.947
R683 vdd3p3.n2587 vdd3p3.t93 217.947
R684 vdd3p3.n2910 vdd3p3.n2827 205.079
R685 vdd3p3.n2910 vdd3p3.n2909 205.079
R686 vdd3p3.n2909 vdd3p3.n2908 205.079
R687 vdd3p3.n2908 vdd3p3.n2828 205.079
R688 vdd3p3.n2902 vdd3p3.n2828 205.079
R689 vdd3p3.n2902 vdd3p3.n2901 205.079
R690 vdd3p3.n2901 vdd3p3.n2900 205.079
R691 vdd3p3.n2900 vdd3p3.n2832 205.079
R692 vdd3p3.n2894 vdd3p3.n2832 205.079
R693 vdd3p3.n2894 vdd3p3.n2893 205.079
R694 vdd3p3.n2893 vdd3p3.n2892 205.079
R695 vdd3p3.n2892 vdd3p3.n2836 205.079
R696 vdd3p3.n2886 vdd3p3.n2836 205.079
R697 vdd3p3.n2989 vdd3p3.n2785 205.079
R698 vdd3p3.n2995 vdd3p3.n2785 205.079
R699 vdd3p3.n2996 vdd3p3.n2995 205.079
R700 vdd3p3.n2997 vdd3p3.n2996 205.079
R701 vdd3p3.n2997 vdd3p3.n2781 205.079
R702 vdd3p3.n3003 vdd3p3.n2781 205.079
R703 vdd3p3.n3004 vdd3p3.n3003 205.079
R704 vdd3p3.n3005 vdd3p3.n3004 205.079
R705 vdd3p3.n3005 vdd3p3.n2777 205.079
R706 vdd3p3.n3011 vdd3p3.n2777 205.079
R707 vdd3p3.n3012 vdd3p3.n3011 205.079
R708 vdd3p3.n3014 vdd3p3.n3012 205.079
R709 vdd3p3.n3014 vdd3p3.n3013 205.079
R710 vdd3p3.n3310 vdd3p3.n2689 205.079
R711 vdd3p3.n3310 vdd3p3.n3309 205.079
R712 vdd3p3.n3309 vdd3p3.n3308 205.079
R713 vdd3p3.n3308 vdd3p3.n2690 205.079
R714 vdd3p3.n3302 vdd3p3.n2690 205.079
R715 vdd3p3.n3302 vdd3p3.n3301 205.079
R716 vdd3p3.n3301 vdd3p3.n3300 205.079
R717 vdd3p3.n3300 vdd3p3.n2694 205.079
R718 vdd3p3.n3294 vdd3p3.n2694 205.079
R719 vdd3p3.n3294 vdd3p3.n3293 205.079
R720 vdd3p3.n3293 vdd3p3.n3292 205.079
R721 vdd3p3.n3292 vdd3p3.n2698 205.079
R722 vdd3p3.n3286 vdd3p3.n2698 205.079
R723 vdd3p3.n3195 vdd3p3.n2751 205.079
R724 vdd3p3.n3196 vdd3p3.n3195 205.079
R725 vdd3p3.n3197 vdd3p3.n3196 205.079
R726 vdd3p3.n3197 vdd3p3.n2747 205.079
R727 vdd3p3.n3203 vdd3p3.n2747 205.079
R728 vdd3p3.n3204 vdd3p3.n3203 205.079
R729 vdd3p3.n3205 vdd3p3.n3204 205.079
R730 vdd3p3.n3205 vdd3p3.n2743 205.079
R731 vdd3p3.n3211 vdd3p3.n2743 205.079
R732 vdd3p3.n3212 vdd3p3.n3211 205.079
R733 vdd3p3.n3213 vdd3p3.n3212 205.079
R734 vdd3p3.n3213 vdd3p3.n2738 205.079
R735 vdd3p3.n3220 vdd3p3.n2738 205.079
R736 vdd3p3.n2064 vdd3p3.n1981 205.079
R737 vdd3p3.n2064 vdd3p3.n2063 205.079
R738 vdd3p3.n2063 vdd3p3.n2062 205.079
R739 vdd3p3.n2062 vdd3p3.n1982 205.079
R740 vdd3p3.n2056 vdd3p3.n1982 205.079
R741 vdd3p3.n2056 vdd3p3.n2055 205.079
R742 vdd3p3.n2055 vdd3p3.n2054 205.079
R743 vdd3p3.n2054 vdd3p3.n1986 205.079
R744 vdd3p3.n2048 vdd3p3.n1986 205.079
R745 vdd3p3.n2048 vdd3p3.n2047 205.079
R746 vdd3p3.n2047 vdd3p3.n2046 205.079
R747 vdd3p3.n2046 vdd3p3.n1990 205.079
R748 vdd3p3.n2040 vdd3p3.n1990 205.079
R749 vdd3p3.n2143 vdd3p3.n1939 205.079
R750 vdd3p3.n2149 vdd3p3.n1939 205.079
R751 vdd3p3.n2150 vdd3p3.n2149 205.079
R752 vdd3p3.n2151 vdd3p3.n2150 205.079
R753 vdd3p3.n2151 vdd3p3.n1935 205.079
R754 vdd3p3.n2157 vdd3p3.n1935 205.079
R755 vdd3p3.n2158 vdd3p3.n2157 205.079
R756 vdd3p3.n2159 vdd3p3.n2158 205.079
R757 vdd3p3.n2159 vdd3p3.n1931 205.079
R758 vdd3p3.n2165 vdd3p3.n1931 205.079
R759 vdd3p3.n2166 vdd3p3.n2165 205.079
R760 vdd3p3.n2168 vdd3p3.n2166 205.079
R761 vdd3p3.n2168 vdd3p3.n2167 205.079
R762 vdd3p3.n2464 vdd3p3.n1843 205.079
R763 vdd3p3.n2464 vdd3p3.n2463 205.079
R764 vdd3p3.n2463 vdd3p3.n2462 205.079
R765 vdd3p3.n2462 vdd3p3.n1844 205.079
R766 vdd3p3.n2456 vdd3p3.n1844 205.079
R767 vdd3p3.n2456 vdd3p3.n2455 205.079
R768 vdd3p3.n2455 vdd3p3.n2454 205.079
R769 vdd3p3.n2454 vdd3p3.n1848 205.079
R770 vdd3p3.n2448 vdd3p3.n1848 205.079
R771 vdd3p3.n2448 vdd3p3.n2447 205.079
R772 vdd3p3.n2447 vdd3p3.n2446 205.079
R773 vdd3p3.n2446 vdd3p3.n1852 205.079
R774 vdd3p3.n2440 vdd3p3.n1852 205.079
R775 vdd3p3.n2349 vdd3p3.n1905 205.079
R776 vdd3p3.n2350 vdd3p3.n2349 205.079
R777 vdd3p3.n2351 vdd3p3.n2350 205.079
R778 vdd3p3.n2351 vdd3p3.n1901 205.079
R779 vdd3p3.n2357 vdd3p3.n1901 205.079
R780 vdd3p3.n2358 vdd3p3.n2357 205.079
R781 vdd3p3.n2359 vdd3p3.n2358 205.079
R782 vdd3p3.n2359 vdd3p3.n1897 205.079
R783 vdd3p3.n2365 vdd3p3.n1897 205.079
R784 vdd3p3.n2366 vdd3p3.n2365 205.079
R785 vdd3p3.n2367 vdd3p3.n2366 205.079
R786 vdd3p3.n2367 vdd3p3.n1892 205.079
R787 vdd3p3.n2374 vdd3p3.n1892 205.079
R788 vdd3p3.n1219 vdd3p3.n1136 205.079
R789 vdd3p3.n1219 vdd3p3.n1218 205.079
R790 vdd3p3.n1218 vdd3p3.n1217 205.079
R791 vdd3p3.n1217 vdd3p3.n1137 205.079
R792 vdd3p3.n1211 vdd3p3.n1137 205.079
R793 vdd3p3.n1211 vdd3p3.n1210 205.079
R794 vdd3p3.n1210 vdd3p3.n1209 205.079
R795 vdd3p3.n1209 vdd3p3.n1141 205.079
R796 vdd3p3.n1203 vdd3p3.n1141 205.079
R797 vdd3p3.n1203 vdd3p3.n1202 205.079
R798 vdd3p3.n1202 vdd3p3.n1201 205.079
R799 vdd3p3.n1201 vdd3p3.n1145 205.079
R800 vdd3p3.n1195 vdd3p3.n1145 205.079
R801 vdd3p3.n1298 vdd3p3.n1094 205.079
R802 vdd3p3.n1304 vdd3p3.n1094 205.079
R803 vdd3p3.n1305 vdd3p3.n1304 205.079
R804 vdd3p3.n1306 vdd3p3.n1305 205.079
R805 vdd3p3.n1306 vdd3p3.n1090 205.079
R806 vdd3p3.n1312 vdd3p3.n1090 205.079
R807 vdd3p3.n1313 vdd3p3.n1312 205.079
R808 vdd3p3.n1314 vdd3p3.n1313 205.079
R809 vdd3p3.n1314 vdd3p3.n1086 205.079
R810 vdd3p3.n1320 vdd3p3.n1086 205.079
R811 vdd3p3.n1321 vdd3p3.n1320 205.079
R812 vdd3p3.n1323 vdd3p3.n1321 205.079
R813 vdd3p3.n1323 vdd3p3.n1322 205.079
R814 vdd3p3.n1619 vdd3p3.n998 205.079
R815 vdd3p3.n1619 vdd3p3.n1618 205.079
R816 vdd3p3.n1618 vdd3p3.n1617 205.079
R817 vdd3p3.n1617 vdd3p3.n999 205.079
R818 vdd3p3.n1611 vdd3p3.n999 205.079
R819 vdd3p3.n1611 vdd3p3.n1610 205.079
R820 vdd3p3.n1610 vdd3p3.n1609 205.079
R821 vdd3p3.n1609 vdd3p3.n1003 205.079
R822 vdd3p3.n1603 vdd3p3.n1003 205.079
R823 vdd3p3.n1603 vdd3p3.n1602 205.079
R824 vdd3p3.n1602 vdd3p3.n1601 205.079
R825 vdd3p3.n1601 vdd3p3.n1007 205.079
R826 vdd3p3.n1595 vdd3p3.n1007 205.079
R827 vdd3p3.n1504 vdd3p3.n1060 205.079
R828 vdd3p3.n1505 vdd3p3.n1504 205.079
R829 vdd3p3.n1506 vdd3p3.n1505 205.079
R830 vdd3p3.n1506 vdd3p3.n1056 205.079
R831 vdd3p3.n1512 vdd3p3.n1056 205.079
R832 vdd3p3.n1513 vdd3p3.n1512 205.079
R833 vdd3p3.n1514 vdd3p3.n1513 205.079
R834 vdd3p3.n1514 vdd3p3.n1052 205.079
R835 vdd3p3.n1520 vdd3p3.n1052 205.079
R836 vdd3p3.n1521 vdd3p3.n1520 205.079
R837 vdd3p3.n1522 vdd3p3.n1521 205.079
R838 vdd3p3.n1522 vdd3p3.n1047 205.079
R839 vdd3p3.n1529 vdd3p3.n1047 205.079
R840 vdd3p3.n373 vdd3p3.n290 205.079
R841 vdd3p3.n373 vdd3p3.n372 205.079
R842 vdd3p3.n372 vdd3p3.n371 205.079
R843 vdd3p3.n371 vdd3p3.n291 205.079
R844 vdd3p3.n365 vdd3p3.n291 205.079
R845 vdd3p3.n365 vdd3p3.n364 205.079
R846 vdd3p3.n364 vdd3p3.n363 205.079
R847 vdd3p3.n363 vdd3p3.n295 205.079
R848 vdd3p3.n357 vdd3p3.n295 205.079
R849 vdd3p3.n357 vdd3p3.n356 205.079
R850 vdd3p3.n356 vdd3p3.n355 205.079
R851 vdd3p3.n355 vdd3p3.n299 205.079
R852 vdd3p3.n349 vdd3p3.n299 205.079
R853 vdd3p3.n452 vdd3p3.n248 205.079
R854 vdd3p3.n458 vdd3p3.n248 205.079
R855 vdd3p3.n459 vdd3p3.n458 205.079
R856 vdd3p3.n460 vdd3p3.n459 205.079
R857 vdd3p3.n460 vdd3p3.n244 205.079
R858 vdd3p3.n466 vdd3p3.n244 205.079
R859 vdd3p3.n467 vdd3p3.n466 205.079
R860 vdd3p3.n468 vdd3p3.n467 205.079
R861 vdd3p3.n468 vdd3p3.n240 205.079
R862 vdd3p3.n474 vdd3p3.n240 205.079
R863 vdd3p3.n475 vdd3p3.n474 205.079
R864 vdd3p3.n477 vdd3p3.n475 205.079
R865 vdd3p3.n477 vdd3p3.n476 205.079
R866 vdd3p3.n773 vdd3p3.n152 205.079
R867 vdd3p3.n773 vdd3p3.n772 205.079
R868 vdd3p3.n772 vdd3p3.n771 205.079
R869 vdd3p3.n771 vdd3p3.n153 205.079
R870 vdd3p3.n765 vdd3p3.n153 205.079
R871 vdd3p3.n765 vdd3p3.n764 205.079
R872 vdd3p3.n764 vdd3p3.n763 205.079
R873 vdd3p3.n763 vdd3p3.n157 205.079
R874 vdd3p3.n757 vdd3p3.n157 205.079
R875 vdd3p3.n757 vdd3p3.n756 205.079
R876 vdd3p3.n756 vdd3p3.n755 205.079
R877 vdd3p3.n755 vdd3p3.n161 205.079
R878 vdd3p3.n749 vdd3p3.n161 205.079
R879 vdd3p3.n658 vdd3p3.n214 205.079
R880 vdd3p3.n659 vdd3p3.n658 205.079
R881 vdd3p3.n660 vdd3p3.n659 205.079
R882 vdd3p3.n660 vdd3p3.n210 205.079
R883 vdd3p3.n666 vdd3p3.n210 205.079
R884 vdd3p3.n667 vdd3p3.n666 205.079
R885 vdd3p3.n668 vdd3p3.n667 205.079
R886 vdd3p3.n668 vdd3p3.n206 205.079
R887 vdd3p3.n674 vdd3p3.n206 205.079
R888 vdd3p3.n675 vdd3p3.n674 205.079
R889 vdd3p3.n676 vdd3p3.n675 205.079
R890 vdd3p3.n676 vdd3p3.n201 205.079
R891 vdd3p3.n683 vdd3p3.n201 205.079
R892 vdd3p3.n3228 vdd3p3.n2733 203.785
R893 vdd3p3.n3229 vdd3p3.n3228 203.785
R894 vdd3p3.n3230 vdd3p3.n3229 203.785
R895 vdd3p3.n3230 vdd3p3.n2729 203.785
R896 vdd3p3.n3236 vdd3p3.n2729 203.785
R897 vdd3p3.n3237 vdd3p3.n3236 203.785
R898 vdd3p3.n3238 vdd3p3.n3237 203.785
R899 vdd3p3.n3238 vdd3p3.n2725 203.785
R900 vdd3p3.n3244 vdd3p3.n2725 203.785
R901 vdd3p3.n3245 vdd3p3.n3244 203.785
R902 vdd3p3.n3246 vdd3p3.n3245 203.785
R903 vdd3p3.n3246 vdd3p3.n2721 203.785
R904 vdd3p3.n3252 vdd3p3.n2721 203.785
R905 vdd3p3.n3253 vdd3p3.n3252 203.785
R906 vdd3p3.n3254 vdd3p3.n3253 203.785
R907 vdd3p3.n3254 vdd3p3.n2717 203.785
R908 vdd3p3.n3260 vdd3p3.n2717 203.785
R909 vdd3p3.n3261 vdd3p3.n3260 203.785
R910 vdd3p3.n3262 vdd3p3.n3261 203.785
R911 vdd3p3.n3262 vdd3p3.n2713 203.785
R912 vdd3p3.n3268 vdd3p3.n2713 203.785
R913 vdd3p3.n3269 vdd3p3.n3268 203.785
R914 vdd3p3.n3270 vdd3p3.n3269 203.785
R915 vdd3p3.n3270 vdd3p3.n2709 203.785
R916 vdd3p3.n3276 vdd3p3.n2709 203.785
R917 vdd3p3.n3277 vdd3p3.n3276 203.785
R918 vdd3p3.n3278 vdd3p3.n3277 203.785
R919 vdd3p3.n3278 vdd3p3.n2702 203.785
R920 vdd3p3.n2382 vdd3p3.n1887 203.785
R921 vdd3p3.n2383 vdd3p3.n2382 203.785
R922 vdd3p3.n2384 vdd3p3.n2383 203.785
R923 vdd3p3.n2384 vdd3p3.n1883 203.785
R924 vdd3p3.n2390 vdd3p3.n1883 203.785
R925 vdd3p3.n2391 vdd3p3.n2390 203.785
R926 vdd3p3.n2392 vdd3p3.n2391 203.785
R927 vdd3p3.n2392 vdd3p3.n1879 203.785
R928 vdd3p3.n2398 vdd3p3.n1879 203.785
R929 vdd3p3.n2399 vdd3p3.n2398 203.785
R930 vdd3p3.n2400 vdd3p3.n2399 203.785
R931 vdd3p3.n2400 vdd3p3.n1875 203.785
R932 vdd3p3.n2406 vdd3p3.n1875 203.785
R933 vdd3p3.n2407 vdd3p3.n2406 203.785
R934 vdd3p3.n2408 vdd3p3.n2407 203.785
R935 vdd3p3.n2408 vdd3p3.n1871 203.785
R936 vdd3p3.n2414 vdd3p3.n1871 203.785
R937 vdd3p3.n2415 vdd3p3.n2414 203.785
R938 vdd3p3.n2416 vdd3p3.n2415 203.785
R939 vdd3p3.n2416 vdd3p3.n1867 203.785
R940 vdd3p3.n2422 vdd3p3.n1867 203.785
R941 vdd3p3.n2423 vdd3p3.n2422 203.785
R942 vdd3p3.n2424 vdd3p3.n2423 203.785
R943 vdd3p3.n2424 vdd3p3.n1863 203.785
R944 vdd3p3.n2430 vdd3p3.n1863 203.785
R945 vdd3p3.n2431 vdd3p3.n2430 203.785
R946 vdd3p3.n2432 vdd3p3.n2431 203.785
R947 vdd3p3.n2432 vdd3p3.n1856 203.785
R948 vdd3p3.n1537 vdd3p3.n1042 203.785
R949 vdd3p3.n1538 vdd3p3.n1537 203.785
R950 vdd3p3.n1539 vdd3p3.n1538 203.785
R951 vdd3p3.n1539 vdd3p3.n1038 203.785
R952 vdd3p3.n1545 vdd3p3.n1038 203.785
R953 vdd3p3.n1546 vdd3p3.n1545 203.785
R954 vdd3p3.n1547 vdd3p3.n1546 203.785
R955 vdd3p3.n1547 vdd3p3.n1034 203.785
R956 vdd3p3.n1553 vdd3p3.n1034 203.785
R957 vdd3p3.n1554 vdd3p3.n1553 203.785
R958 vdd3p3.n1555 vdd3p3.n1554 203.785
R959 vdd3p3.n1555 vdd3p3.n1030 203.785
R960 vdd3p3.n1561 vdd3p3.n1030 203.785
R961 vdd3p3.n1562 vdd3p3.n1561 203.785
R962 vdd3p3.n1563 vdd3p3.n1562 203.785
R963 vdd3p3.n1563 vdd3p3.n1026 203.785
R964 vdd3p3.n1569 vdd3p3.n1026 203.785
R965 vdd3p3.n1570 vdd3p3.n1569 203.785
R966 vdd3p3.n1571 vdd3p3.n1570 203.785
R967 vdd3p3.n1571 vdd3p3.n1022 203.785
R968 vdd3p3.n1577 vdd3p3.n1022 203.785
R969 vdd3p3.n1578 vdd3p3.n1577 203.785
R970 vdd3p3.n1579 vdd3p3.n1578 203.785
R971 vdd3p3.n1579 vdd3p3.n1018 203.785
R972 vdd3p3.n1585 vdd3p3.n1018 203.785
R973 vdd3p3.n1586 vdd3p3.n1585 203.785
R974 vdd3p3.n1587 vdd3p3.n1586 203.785
R975 vdd3p3.n1587 vdd3p3.n1011 203.785
R976 vdd3p3.n691 vdd3p3.n196 203.785
R977 vdd3p3.n692 vdd3p3.n691 203.785
R978 vdd3p3.n693 vdd3p3.n692 203.785
R979 vdd3p3.n693 vdd3p3.n192 203.785
R980 vdd3p3.n699 vdd3p3.n192 203.785
R981 vdd3p3.n700 vdd3p3.n699 203.785
R982 vdd3p3.n701 vdd3p3.n700 203.785
R983 vdd3p3.n701 vdd3p3.n188 203.785
R984 vdd3p3.n707 vdd3p3.n188 203.785
R985 vdd3p3.n708 vdd3p3.n707 203.785
R986 vdd3p3.n709 vdd3p3.n708 203.785
R987 vdd3p3.n709 vdd3p3.n184 203.785
R988 vdd3p3.n715 vdd3p3.n184 203.785
R989 vdd3p3.n716 vdd3p3.n715 203.785
R990 vdd3p3.n717 vdd3p3.n716 203.785
R991 vdd3p3.n717 vdd3p3.n180 203.785
R992 vdd3p3.n723 vdd3p3.n180 203.785
R993 vdd3p3.n724 vdd3p3.n723 203.785
R994 vdd3p3.n725 vdd3p3.n724 203.785
R995 vdd3p3.n725 vdd3p3.n176 203.785
R996 vdd3p3.n731 vdd3p3.n176 203.785
R997 vdd3p3.n732 vdd3p3.n731 203.785
R998 vdd3p3.n733 vdd3p3.n732 203.785
R999 vdd3p3.n733 vdd3p3.n172 203.785
R1000 vdd3p3.n739 vdd3p3.n172 203.785
R1001 vdd3p3.n740 vdd3p3.n739 203.785
R1002 vdd3p3.n741 vdd3p3.n740 203.785
R1003 vdd3p3.n741 vdd3p3.n165 203.785
R1004 vdd3p3.n29 vdd3p3.n6 175.384
R1005 vdd3p3.n56 vdd3p3.n30 175.384
R1006 vdd3p3.n868 vdd3p3.n867 175.384
R1007 vdd3p3.n883 vdd3p3.n849 175.384
R1008 vdd3p3.n1720 vdd3p3.n1697 175.384
R1009 vdd3p3.n1747 vdd3p3.n1721 175.384
R1010 vdd3p3.n2559 vdd3p3.n2558 175.384
R1011 vdd3p3.n2574 vdd3p3.n2540 175.384
R1012 vdd3p3.n15 vdd3p3.t120 171.451
R1013 vdd3p3.t155 vdd3p3.n866 171.451
R1014 vdd3p3.n1706 vdd3p3.t11 171.451
R1015 vdd3p3.t81 vdd3p3.n2557 171.451
R1016 vdd3p3.n2885 vdd3p3.n2689 168.888
R1017 vdd3p3.n2755 vdd3p3.n2751 168.888
R1018 vdd3p3.n2039 vdd3p3.n1843 168.888
R1019 vdd3p3.n1909 vdd3p3.n1905 168.888
R1020 vdd3p3.n1194 vdd3p3.n998 168.888
R1021 vdd3p3.n1064 vdd3p3.n1060 168.888
R1022 vdd3p3.n348 vdd3p3.n152 168.888
R1023 vdd3p3.n218 vdd3p3.n214 168.888
R1024 vdd3p3.n3222 vdd3p3.n3221 164.826
R1025 vdd3p3.n2376 vdd3p3.n2375 164.826
R1026 vdd3p3.n1531 vdd3p3.n1530 164.826
R1027 vdd3p3.n685 vdd3p3.n684 164.826
R1028 vdd3p3.n3286 vdd3p3.n3285 162.857
R1029 vdd3p3.n3221 vdd3p3.n3220 162.857
R1030 vdd3p3.n2440 vdd3p3.n2439 162.857
R1031 vdd3p3.n2375 vdd3p3.n2374 162.857
R1032 vdd3p3.n1595 vdd3p3.n1594 162.857
R1033 vdd3p3.n1530 vdd3p3.n1529 162.857
R1034 vdd3p3.n749 vdd3p3.n748 162.857
R1035 vdd3p3.n684 vdd3p3.n683 162.857
R1036 vdd3p3.n3285 vdd3p3.n3284 161.829
R1037 vdd3p3.n2439 vdd3p3.n2438 161.829
R1038 vdd3p3.n1594 vdd3p3.n1593 161.829
R1039 vdd3p3.n748 vdd3p3.n747 161.829
R1040 vdd3p3.n18 vdd3p3.t121 160.741
R1041 vdd3p3.n858 vdd3p3.t156 160.741
R1042 vdd3p3.n1709 vdd3p3.t12 160.741
R1043 vdd3p3.n2549 vdd3p3.t82 160.741
R1044 vdd3p3.n3177 vdd3p3.n2755 160.256
R1045 vdd3p3.n2331 vdd3p3.n1909 160.256
R1046 vdd3p3.n1486 vdd3p3.n1064 160.256
R1047 vdd3p3.n640 vdd3p3.n218 160.256
R1048 vdd3p3.n2987 vdd3p3.n2790 159.113
R1049 vdd3p3.n2973 vdd3p3.n2790 159.113
R1050 vdd3p3.n2973 vdd3p3.n2972 159.113
R1051 vdd3p3.n2972 vdd3p3.n2971 159.113
R1052 vdd3p3.n2971 vdd3p3.n2795 159.113
R1053 vdd3p3.n2965 vdd3p3.n2795 159.113
R1054 vdd3p3.n2965 vdd3p3.n2964 159.113
R1055 vdd3p3.n2964 vdd3p3.n2963 159.113
R1056 vdd3p3.n2963 vdd3p3.n2799 159.113
R1057 vdd3p3.n2957 vdd3p3.n2799 159.113
R1058 vdd3p3.n2957 vdd3p3.n2956 159.113
R1059 vdd3p3.n2956 vdd3p3.n2955 159.113
R1060 vdd3p3.n2955 vdd3p3.n2803 159.113
R1061 vdd3p3.n2949 vdd3p3.n2803 159.113
R1062 vdd3p3.n2949 vdd3p3.n2948 159.113
R1063 vdd3p3.n2948 vdd3p3.n2947 159.113
R1064 vdd3p3.n2947 vdd3p3.n2807 159.113
R1065 vdd3p3.n2941 vdd3p3.n2807 159.113
R1066 vdd3p3.n2941 vdd3p3.n2940 159.113
R1067 vdd3p3.n2940 vdd3p3.n2939 159.113
R1068 vdd3p3.n2939 vdd3p3.n2811 159.113
R1069 vdd3p3.n2933 vdd3p3.n2811 159.113
R1070 vdd3p3.n2933 vdd3p3.n2932 159.113
R1071 vdd3p3.n2932 vdd3p3.n2931 159.113
R1072 vdd3p3.n2931 vdd3p3.n2815 159.113
R1073 vdd3p3.n2925 vdd3p3.n2815 159.113
R1074 vdd3p3.n2925 vdd3p3.n2924 159.113
R1075 vdd3p3.n2924 vdd3p3.n2923 159.113
R1076 vdd3p3.n2141 vdd3p3.n1944 159.113
R1077 vdd3p3.n2127 vdd3p3.n1944 159.113
R1078 vdd3p3.n2127 vdd3p3.n2126 159.113
R1079 vdd3p3.n2126 vdd3p3.n2125 159.113
R1080 vdd3p3.n2125 vdd3p3.n1949 159.113
R1081 vdd3p3.n2119 vdd3p3.n1949 159.113
R1082 vdd3p3.n2119 vdd3p3.n2118 159.113
R1083 vdd3p3.n2118 vdd3p3.n2117 159.113
R1084 vdd3p3.n2117 vdd3p3.n1953 159.113
R1085 vdd3p3.n2111 vdd3p3.n1953 159.113
R1086 vdd3p3.n2111 vdd3p3.n2110 159.113
R1087 vdd3p3.n2110 vdd3p3.n2109 159.113
R1088 vdd3p3.n2109 vdd3p3.n1957 159.113
R1089 vdd3p3.n2103 vdd3p3.n1957 159.113
R1090 vdd3p3.n2103 vdd3p3.n2102 159.113
R1091 vdd3p3.n2102 vdd3p3.n2101 159.113
R1092 vdd3p3.n2101 vdd3p3.n1961 159.113
R1093 vdd3p3.n2095 vdd3p3.n1961 159.113
R1094 vdd3p3.n2095 vdd3p3.n2094 159.113
R1095 vdd3p3.n2094 vdd3p3.n2093 159.113
R1096 vdd3p3.n2093 vdd3p3.n1965 159.113
R1097 vdd3p3.n2087 vdd3p3.n1965 159.113
R1098 vdd3p3.n2087 vdd3p3.n2086 159.113
R1099 vdd3p3.n2086 vdd3p3.n2085 159.113
R1100 vdd3p3.n2085 vdd3p3.n1969 159.113
R1101 vdd3p3.n2079 vdd3p3.n1969 159.113
R1102 vdd3p3.n2079 vdd3p3.n2078 159.113
R1103 vdd3p3.n2078 vdd3p3.n2077 159.113
R1104 vdd3p3.n1296 vdd3p3.n1099 159.113
R1105 vdd3p3.n1282 vdd3p3.n1099 159.113
R1106 vdd3p3.n1282 vdd3p3.n1281 159.113
R1107 vdd3p3.n1281 vdd3p3.n1280 159.113
R1108 vdd3p3.n1280 vdd3p3.n1104 159.113
R1109 vdd3p3.n1274 vdd3p3.n1104 159.113
R1110 vdd3p3.n1274 vdd3p3.n1273 159.113
R1111 vdd3p3.n1273 vdd3p3.n1272 159.113
R1112 vdd3p3.n1272 vdd3p3.n1108 159.113
R1113 vdd3p3.n1266 vdd3p3.n1108 159.113
R1114 vdd3p3.n1266 vdd3p3.n1265 159.113
R1115 vdd3p3.n1265 vdd3p3.n1264 159.113
R1116 vdd3p3.n1264 vdd3p3.n1112 159.113
R1117 vdd3p3.n1258 vdd3p3.n1112 159.113
R1118 vdd3p3.n1258 vdd3p3.n1257 159.113
R1119 vdd3p3.n1257 vdd3p3.n1256 159.113
R1120 vdd3p3.n1256 vdd3p3.n1116 159.113
R1121 vdd3p3.n1250 vdd3p3.n1116 159.113
R1122 vdd3p3.n1250 vdd3p3.n1249 159.113
R1123 vdd3p3.n1249 vdd3p3.n1248 159.113
R1124 vdd3p3.n1248 vdd3p3.n1120 159.113
R1125 vdd3p3.n1242 vdd3p3.n1120 159.113
R1126 vdd3p3.n1242 vdd3p3.n1241 159.113
R1127 vdd3p3.n1241 vdd3p3.n1240 159.113
R1128 vdd3p3.n1240 vdd3p3.n1124 159.113
R1129 vdd3p3.n1234 vdd3p3.n1124 159.113
R1130 vdd3p3.n1234 vdd3p3.n1233 159.113
R1131 vdd3p3.n1233 vdd3p3.n1232 159.113
R1132 vdd3p3.n450 vdd3p3.n253 159.113
R1133 vdd3p3.n436 vdd3p3.n253 159.113
R1134 vdd3p3.n436 vdd3p3.n435 159.113
R1135 vdd3p3.n435 vdd3p3.n434 159.113
R1136 vdd3p3.n434 vdd3p3.n258 159.113
R1137 vdd3p3.n428 vdd3p3.n258 159.113
R1138 vdd3p3.n428 vdd3p3.n427 159.113
R1139 vdd3p3.n427 vdd3p3.n426 159.113
R1140 vdd3p3.n426 vdd3p3.n262 159.113
R1141 vdd3p3.n420 vdd3p3.n262 159.113
R1142 vdd3p3.n420 vdd3p3.n419 159.113
R1143 vdd3p3.n419 vdd3p3.n418 159.113
R1144 vdd3p3.n418 vdd3p3.n266 159.113
R1145 vdd3p3.n412 vdd3p3.n266 159.113
R1146 vdd3p3.n412 vdd3p3.n411 159.113
R1147 vdd3p3.n411 vdd3p3.n410 159.113
R1148 vdd3p3.n410 vdd3p3.n270 159.113
R1149 vdd3p3.n404 vdd3p3.n270 159.113
R1150 vdd3p3.n404 vdd3p3.n403 159.113
R1151 vdd3p3.n403 vdd3p3.n402 159.113
R1152 vdd3p3.n402 vdd3p3.n274 159.113
R1153 vdd3p3.n396 vdd3p3.n274 159.113
R1154 vdd3p3.n396 vdd3p3.n395 159.113
R1155 vdd3p3.n395 vdd3p3.n394 159.113
R1156 vdd3p3.n394 vdd3p3.n278 159.113
R1157 vdd3p3.n388 vdd3p3.n278 159.113
R1158 vdd3p3.n388 vdd3p3.n387 159.113
R1159 vdd3p3.n387 vdd3p3.n386 159.113
R1160 vdd3p3.n5022 vdd3p3.n4722 158.752
R1161 vdd3p3.n10 vdd3p3.t123 158.223
R1162 vdd3p3.n879 vdd3p3.t158 158.223
R1163 vdd3p3.n1701 vdd3p3.t14 158.223
R1164 vdd3p3.n2570 vdd3p3.t80 158.223
R1165 vdd3p3.n2885 vdd3p3.n2683 154.487
R1166 vdd3p3.n2039 vdd3p3.n1837 154.487
R1167 vdd3p3.n1194 vdd3p3.n992 154.487
R1168 vdd3p3.n348 vdd3p3.n146 154.487
R1169 vdd3p3.t145 vdd3p3.t143 151.181
R1170 vdd3p3.t26 vdd3p3.t9 151.181
R1171 vdd3p3.t9 vdd3p3.t25 151.181
R1172 vdd3p3.t25 vdd3p3.t27 151.181
R1173 vdd3p3.t4 vdd3p3.t6 151.181
R1174 vdd3p3.t63 vdd3p3.t4 151.181
R1175 vdd3p3.t56 vdd3p3.t63 151.181
R1176 vdd3p3.n2986 vdd3p3.n2791 141.729
R1177 vdd3p3.n2922 vdd3p3.n2820 141.729
R1178 vdd3p3.n2140 vdd3p3.n1945 141.729
R1179 vdd3p3.n2076 vdd3p3.n1974 141.729
R1180 vdd3p3.n1295 vdd3p3.n1100 141.729
R1181 vdd3p3.n1231 vdd3p3.n1129 141.729
R1182 vdd3p3.n449 vdd3p3.n254 141.729
R1183 vdd3p3.n385 vdd3p3.n283 141.729
R1184 vdd3p3.n3223 vdd3p3.n2734 140.188
R1185 vdd3p3.n3283 vdd3p3.n2705 140.188
R1186 vdd3p3.n2377 vdd3p3.n1888 140.188
R1187 vdd3p3.n2437 vdd3p3.n1859 140.188
R1188 vdd3p3.n1532 vdd3p3.n1043 140.188
R1189 vdd3p3.n1592 vdd3p3.n1014 140.188
R1190 vdd3p3.n686 vdd3p3.n197 140.188
R1191 vdd3p3.n746 vdd3p3.n168 140.188
R1192 vdd3p3.n3140 vdd3p3.n3079 133.655
R1193 vdd3p3.n3129 vdd3p3.n3082 133.655
R1194 vdd3p3.n3058 vdd3p3.n3056 133.655
R1195 vdd3p3.n3062 vdd3p3.n3052 133.655
R1196 vdd3p3.n3065 vdd3p3.n3064 133.655
R1197 vdd3p3.n3072 vdd3p3.n3068 133.655
R1198 vdd3p3.n2865 vdd3p3.n2864 133.655
R1199 vdd3p3.n3162 vdd3p3.n3033 133.655
R1200 vdd3p3.n3154 vdd3p3.n3033 133.655
R1201 vdd3p3.n3154 vdd3p3.n3040 133.655
R1202 vdd3p3.n3146 vdd3p3.n3040 133.655
R1203 vdd3p3.n3146 vdd3p3.n3075 133.655
R1204 vdd3p3.n3071 vdd3p3.n3070 133.655
R1205 vdd3p3.n3070 vdd3p3.n2623 133.655
R1206 vdd3p3.n2631 vdd3p3.n2623 133.655
R1207 vdd3p3.n3356 vdd3p3.n2631 133.655
R1208 vdd3p3.n3356 vdd3p3.n2632 133.655
R1209 vdd3p3.n3175 vdd3p3.n3022 133.655
R1210 vdd3p3.n3167 vdd3p3.n3028 133.655
R1211 vdd3p3.n3043 vdd3p3.n3021 133.655
R1212 vdd3p3.n3152 vdd3p3.n3043 133.655
R1213 vdd3p3.n3152 vdd3p3.n3044 133.655
R1214 vdd3p3.n3148 vdd3p3.n3044 133.655
R1215 vdd3p3.n3148 vdd3p3.n3047 133.655
R1216 vdd3p3.n3055 vdd3p3.n2624 133.655
R1217 vdd3p3.n3362 vdd3p3.n2624 133.655
R1218 vdd3p3.n3362 vdd3p3.n2625 133.655
R1219 vdd3p3.n3358 vdd3p3.n2625 133.655
R1220 vdd3p3.n3358 vdd3p3.n2628 133.655
R1221 vdd3p3.n3105 vdd3p3.n3104 133.655
R1222 vdd3p3.n3111 vdd3p3.n3110 133.655
R1223 vdd3p3.n3159 vdd3p3.n3037 133.655
R1224 vdd3p3.n3159 vdd3p3.n3038 133.655
R1225 vdd3p3.n3078 vdd3p3.n3038 133.655
R1226 vdd3p3.n3374 vdd3p3.n2609 133.655
R1227 vdd3p3.n3374 vdd3p3.n2610 133.655
R1228 vdd3p3.n3366 vdd3p3.n2610 133.655
R1229 vdd3p3.n3366 vdd3p3.n3365 133.655
R1230 vdd3p3.n3365 vdd3p3.n2620 133.655
R1231 vdd3p3.n3351 vdd3p3.n2639 133.655
R1232 vdd3p3.n3343 vdd3p3.n3342 133.655
R1233 vdd3p3.n3333 vdd3p3.n3332 133.655
R1234 vdd3p3.n3324 vdd3p3.n2682 133.655
R1235 vdd3p3.n3120 vdd3p3.n3036 133.655
R1236 vdd3p3.n3124 vdd3p3.n3036 133.655
R1237 vdd3p3.n3125 vdd3p3.n3124 133.655
R1238 vdd3p3.n3372 vdd3p3.n2612 133.655
R1239 vdd3p3.n3372 vdd3p3.n2613 133.655
R1240 vdd3p3.n3368 vdd3p3.n2613 133.655
R1241 vdd3p3.n3368 vdd3p3.n2616 133.655
R1242 vdd3p3.n2660 vdd3p3.n2616 133.655
R1243 vdd3p3.n3349 vdd3p3.n2643 133.655
R1244 vdd3p3.n3345 vdd3p3.n2643 133.655
R1245 vdd3p3.n3345 vdd3p3.n2664 133.655
R1246 vdd3p3.n2647 vdd3p3.n2638 133.655
R1247 vdd3p3.n2658 vdd3p3.n2642 133.655
R1248 vdd3p3.n2294 vdd3p3.n2233 133.655
R1249 vdd3p3.n2283 vdd3p3.n2236 133.655
R1250 vdd3p3.n2212 vdd3p3.n2210 133.655
R1251 vdd3p3.n2216 vdd3p3.n2206 133.655
R1252 vdd3p3.n2219 vdd3p3.n2218 133.655
R1253 vdd3p3.n2226 vdd3p3.n2222 133.655
R1254 vdd3p3.n2019 vdd3p3.n2018 133.655
R1255 vdd3p3.n2316 vdd3p3.n2187 133.655
R1256 vdd3p3.n2308 vdd3p3.n2187 133.655
R1257 vdd3p3.n2308 vdd3p3.n2194 133.655
R1258 vdd3p3.n2300 vdd3p3.n2194 133.655
R1259 vdd3p3.n2300 vdd3p3.n2229 133.655
R1260 vdd3p3.n2225 vdd3p3.n2224 133.655
R1261 vdd3p3.n2224 vdd3p3.n1777 133.655
R1262 vdd3p3.n1785 vdd3p3.n1777 133.655
R1263 vdd3p3.n2510 vdd3p3.n1785 133.655
R1264 vdd3p3.n2510 vdd3p3.n1786 133.655
R1265 vdd3p3.n2329 vdd3p3.n2176 133.655
R1266 vdd3p3.n2321 vdd3p3.n2182 133.655
R1267 vdd3p3.n2197 vdd3p3.n2175 133.655
R1268 vdd3p3.n2306 vdd3p3.n2197 133.655
R1269 vdd3p3.n2306 vdd3p3.n2198 133.655
R1270 vdd3p3.n2302 vdd3p3.n2198 133.655
R1271 vdd3p3.n2302 vdd3p3.n2201 133.655
R1272 vdd3p3.n2209 vdd3p3.n1778 133.655
R1273 vdd3p3.n2516 vdd3p3.n1778 133.655
R1274 vdd3p3.n2516 vdd3p3.n1779 133.655
R1275 vdd3p3.n2512 vdd3p3.n1779 133.655
R1276 vdd3p3.n2512 vdd3p3.n1782 133.655
R1277 vdd3p3.n2259 vdd3p3.n2258 133.655
R1278 vdd3p3.n2265 vdd3p3.n2264 133.655
R1279 vdd3p3.n2313 vdd3p3.n2191 133.655
R1280 vdd3p3.n2313 vdd3p3.n2192 133.655
R1281 vdd3p3.n2232 vdd3p3.n2192 133.655
R1282 vdd3p3.n2528 vdd3p3.n1763 133.655
R1283 vdd3p3.n2528 vdd3p3.n1764 133.655
R1284 vdd3p3.n2520 vdd3p3.n1764 133.655
R1285 vdd3p3.n2520 vdd3p3.n2519 133.655
R1286 vdd3p3.n2519 vdd3p3.n1774 133.655
R1287 vdd3p3.n2505 vdd3p3.n1793 133.655
R1288 vdd3p3.n2497 vdd3p3.n2496 133.655
R1289 vdd3p3.n2487 vdd3p3.n2486 133.655
R1290 vdd3p3.n2478 vdd3p3.n1836 133.655
R1291 vdd3p3.n2274 vdd3p3.n2190 133.655
R1292 vdd3p3.n2278 vdd3p3.n2190 133.655
R1293 vdd3p3.n2279 vdd3p3.n2278 133.655
R1294 vdd3p3.n2526 vdd3p3.n1766 133.655
R1295 vdd3p3.n2526 vdd3p3.n1767 133.655
R1296 vdd3p3.n2522 vdd3p3.n1767 133.655
R1297 vdd3p3.n2522 vdd3p3.n1770 133.655
R1298 vdd3p3.n1814 vdd3p3.n1770 133.655
R1299 vdd3p3.n2503 vdd3p3.n1797 133.655
R1300 vdd3p3.n2499 vdd3p3.n1797 133.655
R1301 vdd3p3.n2499 vdd3p3.n1818 133.655
R1302 vdd3p3.n1801 vdd3p3.n1792 133.655
R1303 vdd3p3.n1812 vdd3p3.n1796 133.655
R1304 vdd3p3.n1449 vdd3p3.n1388 133.655
R1305 vdd3p3.n1438 vdd3p3.n1391 133.655
R1306 vdd3p3.n1367 vdd3p3.n1365 133.655
R1307 vdd3p3.n1371 vdd3p3.n1361 133.655
R1308 vdd3p3.n1374 vdd3p3.n1373 133.655
R1309 vdd3p3.n1381 vdd3p3.n1377 133.655
R1310 vdd3p3.n1174 vdd3p3.n1173 133.655
R1311 vdd3p3.n1471 vdd3p3.n1342 133.655
R1312 vdd3p3.n1463 vdd3p3.n1342 133.655
R1313 vdd3p3.n1463 vdd3p3.n1349 133.655
R1314 vdd3p3.n1455 vdd3p3.n1349 133.655
R1315 vdd3p3.n1455 vdd3p3.n1384 133.655
R1316 vdd3p3.n1380 vdd3p3.n1379 133.655
R1317 vdd3p3.n1379 vdd3p3.n932 133.655
R1318 vdd3p3.n940 vdd3p3.n932 133.655
R1319 vdd3p3.n1665 vdd3p3.n940 133.655
R1320 vdd3p3.n1665 vdd3p3.n941 133.655
R1321 vdd3p3.n1484 vdd3p3.n1331 133.655
R1322 vdd3p3.n1476 vdd3p3.n1337 133.655
R1323 vdd3p3.n1352 vdd3p3.n1330 133.655
R1324 vdd3p3.n1461 vdd3p3.n1352 133.655
R1325 vdd3p3.n1461 vdd3p3.n1353 133.655
R1326 vdd3p3.n1457 vdd3p3.n1353 133.655
R1327 vdd3p3.n1457 vdd3p3.n1356 133.655
R1328 vdd3p3.n1364 vdd3p3.n933 133.655
R1329 vdd3p3.n1671 vdd3p3.n933 133.655
R1330 vdd3p3.n1671 vdd3p3.n934 133.655
R1331 vdd3p3.n1667 vdd3p3.n934 133.655
R1332 vdd3p3.n1667 vdd3p3.n937 133.655
R1333 vdd3p3.n1414 vdd3p3.n1413 133.655
R1334 vdd3p3.n1420 vdd3p3.n1419 133.655
R1335 vdd3p3.n1468 vdd3p3.n1346 133.655
R1336 vdd3p3.n1468 vdd3p3.n1347 133.655
R1337 vdd3p3.n1387 vdd3p3.n1347 133.655
R1338 vdd3p3.n1683 vdd3p3.n918 133.655
R1339 vdd3p3.n1683 vdd3p3.n919 133.655
R1340 vdd3p3.n1675 vdd3p3.n919 133.655
R1341 vdd3p3.n1675 vdd3p3.n1674 133.655
R1342 vdd3p3.n1674 vdd3p3.n929 133.655
R1343 vdd3p3.n1660 vdd3p3.n948 133.655
R1344 vdd3p3.n1652 vdd3p3.n1651 133.655
R1345 vdd3p3.n1642 vdd3p3.n1641 133.655
R1346 vdd3p3.n1633 vdd3p3.n991 133.655
R1347 vdd3p3.n1429 vdd3p3.n1345 133.655
R1348 vdd3p3.n1433 vdd3p3.n1345 133.655
R1349 vdd3p3.n1434 vdd3p3.n1433 133.655
R1350 vdd3p3.n1681 vdd3p3.n921 133.655
R1351 vdd3p3.n1681 vdd3p3.n922 133.655
R1352 vdd3p3.n1677 vdd3p3.n922 133.655
R1353 vdd3p3.n1677 vdd3p3.n925 133.655
R1354 vdd3p3.n969 vdd3p3.n925 133.655
R1355 vdd3p3.n1658 vdd3p3.n952 133.655
R1356 vdd3p3.n1654 vdd3p3.n952 133.655
R1357 vdd3p3.n1654 vdd3p3.n973 133.655
R1358 vdd3p3.n956 vdd3p3.n947 133.655
R1359 vdd3p3.n967 vdd3p3.n951 133.655
R1360 vdd3p3.n603 vdd3p3.n542 133.655
R1361 vdd3p3.n592 vdd3p3.n545 133.655
R1362 vdd3p3.n521 vdd3p3.n519 133.655
R1363 vdd3p3.n525 vdd3p3.n515 133.655
R1364 vdd3p3.n528 vdd3p3.n527 133.655
R1365 vdd3p3.n535 vdd3p3.n531 133.655
R1366 vdd3p3.n328 vdd3p3.n327 133.655
R1367 vdd3p3.n625 vdd3p3.n496 133.655
R1368 vdd3p3.n617 vdd3p3.n496 133.655
R1369 vdd3p3.n617 vdd3p3.n503 133.655
R1370 vdd3p3.n609 vdd3p3.n503 133.655
R1371 vdd3p3.n609 vdd3p3.n538 133.655
R1372 vdd3p3.n534 vdd3p3.n533 133.655
R1373 vdd3p3.n533 vdd3p3.n86 133.655
R1374 vdd3p3.n94 vdd3p3.n86 133.655
R1375 vdd3p3.n819 vdd3p3.n94 133.655
R1376 vdd3p3.n819 vdd3p3.n95 133.655
R1377 vdd3p3.n638 vdd3p3.n485 133.655
R1378 vdd3p3.n630 vdd3p3.n491 133.655
R1379 vdd3p3.n506 vdd3p3.n484 133.655
R1380 vdd3p3.n615 vdd3p3.n506 133.655
R1381 vdd3p3.n615 vdd3p3.n507 133.655
R1382 vdd3p3.n611 vdd3p3.n507 133.655
R1383 vdd3p3.n611 vdd3p3.n510 133.655
R1384 vdd3p3.n518 vdd3p3.n87 133.655
R1385 vdd3p3.n825 vdd3p3.n87 133.655
R1386 vdd3p3.n825 vdd3p3.n88 133.655
R1387 vdd3p3.n821 vdd3p3.n88 133.655
R1388 vdd3p3.n821 vdd3p3.n91 133.655
R1389 vdd3p3.n568 vdd3p3.n567 133.655
R1390 vdd3p3.n574 vdd3p3.n573 133.655
R1391 vdd3p3.n622 vdd3p3.n500 133.655
R1392 vdd3p3.n622 vdd3p3.n501 133.655
R1393 vdd3p3.n541 vdd3p3.n501 133.655
R1394 vdd3p3.n837 vdd3p3.n72 133.655
R1395 vdd3p3.n837 vdd3p3.n73 133.655
R1396 vdd3p3.n829 vdd3p3.n73 133.655
R1397 vdd3p3.n829 vdd3p3.n828 133.655
R1398 vdd3p3.n828 vdd3p3.n83 133.655
R1399 vdd3p3.n814 vdd3p3.n102 133.655
R1400 vdd3p3.n806 vdd3p3.n805 133.655
R1401 vdd3p3.n796 vdd3p3.n795 133.655
R1402 vdd3p3.n787 vdd3p3.n145 133.655
R1403 vdd3p3.n583 vdd3p3.n499 133.655
R1404 vdd3p3.n587 vdd3p3.n499 133.655
R1405 vdd3p3.n588 vdd3p3.n587 133.655
R1406 vdd3p3.n835 vdd3p3.n75 133.655
R1407 vdd3p3.n835 vdd3p3.n76 133.655
R1408 vdd3p3.n831 vdd3p3.n76 133.655
R1409 vdd3p3.n831 vdd3p3.n79 133.655
R1410 vdd3p3.n123 vdd3p3.n79 133.655
R1411 vdd3p3.n812 vdd3p3.n106 133.655
R1412 vdd3p3.n808 vdd3p3.n106 133.655
R1413 vdd3p3.n808 vdd3p3.n127 133.655
R1414 vdd3p3.n110 vdd3p3.n101 133.655
R1415 vdd3p3.n121 vdd3p3.n105 133.655
R1416 vdd3p3.n2988 vdd3p3.n2789 128.694
R1417 vdd3p3.n2142 vdd3p3.n1943 128.694
R1418 vdd3p3.n1297 vdd3p3.n1098 128.694
R1419 vdd3p3.n451 vdd3p3.n252 128.694
R1420 vdd3p3.n5020 vdd3p3.t56 126.424
R1421 vdd3p3.n2823 vdd3p3.n2819 126.354
R1422 vdd3p3.n1977 vdd3p3.n1973 126.354
R1423 vdd3p3.n1132 vdd3p3.n1128 126.354
R1424 vdd3p3.n286 vdd3p3.n282 126.354
R1425 vdd3p3.t140 vdd3p3.n54 117.837
R1426 vdd3p3.n896 vdd3p3.t166 117.837
R1427 vdd3p3.t83 vdd3p3.n1745 117.837
R1428 vdd3p3.n2587 vdd3p3.t87 117.837
R1429 vdd3p3.n7005 vdd3p3.n7004 117.619
R1430 vdd3p3.n4952 vdd3p3.t61 116.84
R1431 vdd3p3.n8499 vdd3p3.t107 116.84
R1432 vdd3p3.n8843 vdd3p3.t103 116.84
R1433 vdd3p3.n5045 vdd3p3.t58 116.84
R1434 vdd3p3.n8754 vdd3p3.t74 116.84
R1435 vdd3p3.n2974 vdd3p3.n2792 104.756
R1436 vdd3p3.n2974 vdd3p3.n2794 104.756
R1437 vdd3p3.n2970 vdd3p3.n2794 104.756
R1438 vdd3p3.n2970 vdd3p3.n2796 104.756
R1439 vdd3p3.n2966 vdd3p3.n2796 104.756
R1440 vdd3p3.n2966 vdd3p3.n2798 104.756
R1441 vdd3p3.n2962 vdd3p3.n2798 104.756
R1442 vdd3p3.n2962 vdd3p3.n2800 104.756
R1443 vdd3p3.n2958 vdd3p3.n2800 104.756
R1444 vdd3p3.n2958 vdd3p3.n2802 104.756
R1445 vdd3p3.n2954 vdd3p3.n2802 104.756
R1446 vdd3p3.n2954 vdd3p3.n2804 104.756
R1447 vdd3p3.n2950 vdd3p3.n2804 104.756
R1448 vdd3p3.n2950 vdd3p3.n2806 104.756
R1449 vdd3p3.n2946 vdd3p3.n2806 104.756
R1450 vdd3p3.n2946 vdd3p3.n2808 104.756
R1451 vdd3p3.n2942 vdd3p3.n2808 104.756
R1452 vdd3p3.n2942 vdd3p3.n2810 104.756
R1453 vdd3p3.n2938 vdd3p3.n2810 104.756
R1454 vdd3p3.n2938 vdd3p3.n2812 104.756
R1455 vdd3p3.n2934 vdd3p3.n2812 104.756
R1456 vdd3p3.n2934 vdd3p3.n2814 104.756
R1457 vdd3p3.n2930 vdd3p3.n2814 104.756
R1458 vdd3p3.n2930 vdd3p3.n2816 104.756
R1459 vdd3p3.n2926 vdd3p3.n2816 104.756
R1460 vdd3p3.n2926 vdd3p3.n2818 104.756
R1461 vdd3p3.n2922 vdd3p3.n2818 104.756
R1462 vdd3p3.n2990 vdd3p3.n2788 104.756
R1463 vdd3p3.n2990 vdd3p3.n2786 104.756
R1464 vdd3p3.n2994 vdd3p3.n2786 104.756
R1465 vdd3p3.n2994 vdd3p3.n2784 104.756
R1466 vdd3p3.n2998 vdd3p3.n2784 104.756
R1467 vdd3p3.n2998 vdd3p3.n2782 104.756
R1468 vdd3p3.n3002 vdd3p3.n2782 104.756
R1469 vdd3p3.n3002 vdd3p3.n2780 104.756
R1470 vdd3p3.n3006 vdd3p3.n2780 104.756
R1471 vdd3p3.n3006 vdd3p3.n2778 104.756
R1472 vdd3p3.n3010 vdd3p3.n2778 104.756
R1473 vdd3p3.n3010 vdd3p3.n2776 104.756
R1474 vdd3p3.n3015 vdd3p3.n2776 104.756
R1475 vdd3p3.n3015 vdd3p3.n2774 104.756
R1476 vdd3p3.n3186 vdd3p3.n2774 104.756
R1477 vdd3p3.n3165 vdd3p3.n2766 104.756
R1478 vdd3p3.n3089 vdd3p3.n2766 104.756
R1479 vdd3p3.n3093 vdd3p3.n3092 104.756
R1480 vdd3p3.n3190 vdd3p3.n2752 104.756
R1481 vdd3p3.n3194 vdd3p3.n2752 104.756
R1482 vdd3p3.n3194 vdd3p3.n2750 104.756
R1483 vdd3p3.n3198 vdd3p3.n2750 104.756
R1484 vdd3p3.n3198 vdd3p3.n2748 104.756
R1485 vdd3p3.n3202 vdd3p3.n2748 104.756
R1486 vdd3p3.n3202 vdd3p3.n2746 104.756
R1487 vdd3p3.n3206 vdd3p3.n2746 104.756
R1488 vdd3p3.n3206 vdd3p3.n2744 104.756
R1489 vdd3p3.n3210 vdd3p3.n2744 104.756
R1490 vdd3p3.n3210 vdd3p3.n2742 104.756
R1491 vdd3p3.n3214 vdd3p3.n2742 104.756
R1492 vdd3p3.n3214 vdd3p3.n2739 104.756
R1493 vdd3p3.n3219 vdd3p3.n2739 104.756
R1494 vdd3p3.n3219 vdd3p3.n2740 104.756
R1495 vdd3p3.n3223 vdd3p3.n2736 104.756
R1496 vdd3p3.n3227 vdd3p3.n2734 104.756
R1497 vdd3p3.n3227 vdd3p3.n2732 104.756
R1498 vdd3p3.n3231 vdd3p3.n2732 104.756
R1499 vdd3p3.n3231 vdd3p3.n2730 104.756
R1500 vdd3p3.n3235 vdd3p3.n2730 104.756
R1501 vdd3p3.n3235 vdd3p3.n2728 104.756
R1502 vdd3p3.n3239 vdd3p3.n2728 104.756
R1503 vdd3p3.n3239 vdd3p3.n2726 104.756
R1504 vdd3p3.n3243 vdd3p3.n2726 104.756
R1505 vdd3p3.n3243 vdd3p3.n2724 104.756
R1506 vdd3p3.n3247 vdd3p3.n2724 104.756
R1507 vdd3p3.n3247 vdd3p3.n2722 104.756
R1508 vdd3p3.n3251 vdd3p3.n2722 104.756
R1509 vdd3p3.n3251 vdd3p3.n2720 104.756
R1510 vdd3p3.n3255 vdd3p3.n2720 104.756
R1511 vdd3p3.n3255 vdd3p3.n2718 104.756
R1512 vdd3p3.n3259 vdd3p3.n2718 104.756
R1513 vdd3p3.n3259 vdd3p3.n2716 104.756
R1514 vdd3p3.n3263 vdd3p3.n2716 104.756
R1515 vdd3p3.n3263 vdd3p3.n2714 104.756
R1516 vdd3p3.n3267 vdd3p3.n2714 104.756
R1517 vdd3p3.n3267 vdd3p3.n2712 104.756
R1518 vdd3p3.n3271 vdd3p3.n2712 104.756
R1519 vdd3p3.n3271 vdd3p3.n2710 104.756
R1520 vdd3p3.n3275 vdd3p3.n2710 104.756
R1521 vdd3p3.n3275 vdd3p3.n2708 104.756
R1522 vdd3p3.n3279 vdd3p3.n2708 104.756
R1523 vdd3p3.n3279 vdd3p3.n2705 104.756
R1524 vdd3p3.n2918 vdd3p3.n2917 104.756
R1525 vdd3p3.n2915 vdd3p3.n2824 104.756
R1526 vdd3p3.n2911 vdd3p3.n2824 104.756
R1527 vdd3p3.n2911 vdd3p3.n2826 104.756
R1528 vdd3p3.n2907 vdd3p3.n2826 104.756
R1529 vdd3p3.n2907 vdd3p3.n2829 104.756
R1530 vdd3p3.n2903 vdd3p3.n2829 104.756
R1531 vdd3p3.n2903 vdd3p3.n2831 104.756
R1532 vdd3p3.n2899 vdd3p3.n2831 104.756
R1533 vdd3p3.n2899 vdd3p3.n2833 104.756
R1534 vdd3p3.n2895 vdd3p3.n2833 104.756
R1535 vdd3p3.n2895 vdd3p3.n2835 104.756
R1536 vdd3p3.n2891 vdd3p3.n2835 104.756
R1537 vdd3p3.n2891 vdd3p3.n2837 104.756
R1538 vdd3p3.n2887 vdd3p3.n2837 104.756
R1539 vdd3p3.n2887 vdd3p3.n2884 104.756
R1540 vdd3p3.n2879 vdd3p3.n2878 104.756
R1541 vdd3p3.n2870 vdd3p3.n2848 104.756
R1542 vdd3p3.n2868 vdd3p3.n2849 104.756
R1543 vdd3p3.n2861 vdd3p3.n2860 104.756
R1544 vdd3p3.n3337 vdd3p3.n3336 104.756
R1545 vdd3p3.n3329 vdd3p3.n2679 104.756
R1546 vdd3p3.n3327 vdd3p3.n2680 104.756
R1547 vdd3p3.n3319 vdd3p3.n3318 104.756
R1548 vdd3p3.n3316 vdd3p3.n2686 104.756
R1549 vdd3p3.n3311 vdd3p3.n2686 104.756
R1550 vdd3p3.n3311 vdd3p3.n2688 104.756
R1551 vdd3p3.n3307 vdd3p3.n2688 104.756
R1552 vdd3p3.n3307 vdd3p3.n2691 104.756
R1553 vdd3p3.n3303 vdd3p3.n2691 104.756
R1554 vdd3p3.n3303 vdd3p3.n2693 104.756
R1555 vdd3p3.n3299 vdd3p3.n2693 104.756
R1556 vdd3p3.n3299 vdd3p3.n2695 104.756
R1557 vdd3p3.n3295 vdd3p3.n2695 104.756
R1558 vdd3p3.n3295 vdd3p3.n2697 104.756
R1559 vdd3p3.n3291 vdd3p3.n2697 104.756
R1560 vdd3p3.n3291 vdd3p3.n2699 104.756
R1561 vdd3p3.n3287 vdd3p3.n2699 104.756
R1562 vdd3p3.n3287 vdd3p3.n2701 104.756
R1563 vdd3p3.n3283 vdd3p3.n2704 104.756
R1564 vdd3p3.n2128 vdd3p3.n1946 104.756
R1565 vdd3p3.n2128 vdd3p3.n1948 104.756
R1566 vdd3p3.n2124 vdd3p3.n1948 104.756
R1567 vdd3p3.n2124 vdd3p3.n1950 104.756
R1568 vdd3p3.n2120 vdd3p3.n1950 104.756
R1569 vdd3p3.n2120 vdd3p3.n1952 104.756
R1570 vdd3p3.n2116 vdd3p3.n1952 104.756
R1571 vdd3p3.n2116 vdd3p3.n1954 104.756
R1572 vdd3p3.n2112 vdd3p3.n1954 104.756
R1573 vdd3p3.n2112 vdd3p3.n1956 104.756
R1574 vdd3p3.n2108 vdd3p3.n1956 104.756
R1575 vdd3p3.n2108 vdd3p3.n1958 104.756
R1576 vdd3p3.n2104 vdd3p3.n1958 104.756
R1577 vdd3p3.n2104 vdd3p3.n1960 104.756
R1578 vdd3p3.n2100 vdd3p3.n1960 104.756
R1579 vdd3p3.n2100 vdd3p3.n1962 104.756
R1580 vdd3p3.n2096 vdd3p3.n1962 104.756
R1581 vdd3p3.n2096 vdd3p3.n1964 104.756
R1582 vdd3p3.n2092 vdd3p3.n1964 104.756
R1583 vdd3p3.n2092 vdd3p3.n1966 104.756
R1584 vdd3p3.n2088 vdd3p3.n1966 104.756
R1585 vdd3p3.n2088 vdd3p3.n1968 104.756
R1586 vdd3p3.n2084 vdd3p3.n1968 104.756
R1587 vdd3p3.n2084 vdd3p3.n1970 104.756
R1588 vdd3p3.n2080 vdd3p3.n1970 104.756
R1589 vdd3p3.n2080 vdd3p3.n1972 104.756
R1590 vdd3p3.n2076 vdd3p3.n1972 104.756
R1591 vdd3p3.n2144 vdd3p3.n1942 104.756
R1592 vdd3p3.n2144 vdd3p3.n1940 104.756
R1593 vdd3p3.n2148 vdd3p3.n1940 104.756
R1594 vdd3p3.n2148 vdd3p3.n1938 104.756
R1595 vdd3p3.n2152 vdd3p3.n1938 104.756
R1596 vdd3p3.n2152 vdd3p3.n1936 104.756
R1597 vdd3p3.n2156 vdd3p3.n1936 104.756
R1598 vdd3p3.n2156 vdd3p3.n1934 104.756
R1599 vdd3p3.n2160 vdd3p3.n1934 104.756
R1600 vdd3p3.n2160 vdd3p3.n1932 104.756
R1601 vdd3p3.n2164 vdd3p3.n1932 104.756
R1602 vdd3p3.n2164 vdd3p3.n1930 104.756
R1603 vdd3p3.n2169 vdd3p3.n1930 104.756
R1604 vdd3p3.n2169 vdd3p3.n1928 104.756
R1605 vdd3p3.n2340 vdd3p3.n1928 104.756
R1606 vdd3p3.n2319 vdd3p3.n1920 104.756
R1607 vdd3p3.n2243 vdd3p3.n1920 104.756
R1608 vdd3p3.n2247 vdd3p3.n2246 104.756
R1609 vdd3p3.n2344 vdd3p3.n1906 104.756
R1610 vdd3p3.n2348 vdd3p3.n1906 104.756
R1611 vdd3p3.n2348 vdd3p3.n1904 104.756
R1612 vdd3p3.n2352 vdd3p3.n1904 104.756
R1613 vdd3p3.n2352 vdd3p3.n1902 104.756
R1614 vdd3p3.n2356 vdd3p3.n1902 104.756
R1615 vdd3p3.n2356 vdd3p3.n1900 104.756
R1616 vdd3p3.n2360 vdd3p3.n1900 104.756
R1617 vdd3p3.n2360 vdd3p3.n1898 104.756
R1618 vdd3p3.n2364 vdd3p3.n1898 104.756
R1619 vdd3p3.n2364 vdd3p3.n1896 104.756
R1620 vdd3p3.n2368 vdd3p3.n1896 104.756
R1621 vdd3p3.n2368 vdd3p3.n1893 104.756
R1622 vdd3p3.n2373 vdd3p3.n1893 104.756
R1623 vdd3p3.n2373 vdd3p3.n1894 104.756
R1624 vdd3p3.n2377 vdd3p3.n1890 104.756
R1625 vdd3p3.n2381 vdd3p3.n1888 104.756
R1626 vdd3p3.n2381 vdd3p3.n1886 104.756
R1627 vdd3p3.n2385 vdd3p3.n1886 104.756
R1628 vdd3p3.n2385 vdd3p3.n1884 104.756
R1629 vdd3p3.n2389 vdd3p3.n1884 104.756
R1630 vdd3p3.n2389 vdd3p3.n1882 104.756
R1631 vdd3p3.n2393 vdd3p3.n1882 104.756
R1632 vdd3p3.n2393 vdd3p3.n1880 104.756
R1633 vdd3p3.n2397 vdd3p3.n1880 104.756
R1634 vdd3p3.n2397 vdd3p3.n1878 104.756
R1635 vdd3p3.n2401 vdd3p3.n1878 104.756
R1636 vdd3p3.n2401 vdd3p3.n1876 104.756
R1637 vdd3p3.n2405 vdd3p3.n1876 104.756
R1638 vdd3p3.n2405 vdd3p3.n1874 104.756
R1639 vdd3p3.n2409 vdd3p3.n1874 104.756
R1640 vdd3p3.n2409 vdd3p3.n1872 104.756
R1641 vdd3p3.n2413 vdd3p3.n1872 104.756
R1642 vdd3p3.n2413 vdd3p3.n1870 104.756
R1643 vdd3p3.n2417 vdd3p3.n1870 104.756
R1644 vdd3p3.n2417 vdd3p3.n1868 104.756
R1645 vdd3p3.n2421 vdd3p3.n1868 104.756
R1646 vdd3p3.n2421 vdd3p3.n1866 104.756
R1647 vdd3p3.n2425 vdd3p3.n1866 104.756
R1648 vdd3p3.n2425 vdd3p3.n1864 104.756
R1649 vdd3p3.n2429 vdd3p3.n1864 104.756
R1650 vdd3p3.n2429 vdd3p3.n1862 104.756
R1651 vdd3p3.n2433 vdd3p3.n1862 104.756
R1652 vdd3p3.n2433 vdd3p3.n1859 104.756
R1653 vdd3p3.n2072 vdd3p3.n2071 104.756
R1654 vdd3p3.n2069 vdd3p3.n1978 104.756
R1655 vdd3p3.n2065 vdd3p3.n1978 104.756
R1656 vdd3p3.n2065 vdd3p3.n1980 104.756
R1657 vdd3p3.n2061 vdd3p3.n1980 104.756
R1658 vdd3p3.n2061 vdd3p3.n1983 104.756
R1659 vdd3p3.n2057 vdd3p3.n1983 104.756
R1660 vdd3p3.n2057 vdd3p3.n1985 104.756
R1661 vdd3p3.n2053 vdd3p3.n1985 104.756
R1662 vdd3p3.n2053 vdd3p3.n1987 104.756
R1663 vdd3p3.n2049 vdd3p3.n1987 104.756
R1664 vdd3p3.n2049 vdd3p3.n1989 104.756
R1665 vdd3p3.n2045 vdd3p3.n1989 104.756
R1666 vdd3p3.n2045 vdd3p3.n1991 104.756
R1667 vdd3p3.n2041 vdd3p3.n1991 104.756
R1668 vdd3p3.n2041 vdd3p3.n2038 104.756
R1669 vdd3p3.n2033 vdd3p3.n2032 104.756
R1670 vdd3p3.n2024 vdd3p3.n2002 104.756
R1671 vdd3p3.n2022 vdd3p3.n2003 104.756
R1672 vdd3p3.n2015 vdd3p3.n2014 104.756
R1673 vdd3p3.n2491 vdd3p3.n2490 104.756
R1674 vdd3p3.n2483 vdd3p3.n1833 104.756
R1675 vdd3p3.n2481 vdd3p3.n1834 104.756
R1676 vdd3p3.n2473 vdd3p3.n2472 104.756
R1677 vdd3p3.n2470 vdd3p3.n1840 104.756
R1678 vdd3p3.n2465 vdd3p3.n1840 104.756
R1679 vdd3p3.n2465 vdd3p3.n1842 104.756
R1680 vdd3p3.n2461 vdd3p3.n1842 104.756
R1681 vdd3p3.n2461 vdd3p3.n1845 104.756
R1682 vdd3p3.n2457 vdd3p3.n1845 104.756
R1683 vdd3p3.n2457 vdd3p3.n1847 104.756
R1684 vdd3p3.n2453 vdd3p3.n1847 104.756
R1685 vdd3p3.n2453 vdd3p3.n1849 104.756
R1686 vdd3p3.n2449 vdd3p3.n1849 104.756
R1687 vdd3p3.n2449 vdd3p3.n1851 104.756
R1688 vdd3p3.n2445 vdd3p3.n1851 104.756
R1689 vdd3p3.n2445 vdd3p3.n1853 104.756
R1690 vdd3p3.n2441 vdd3p3.n1853 104.756
R1691 vdd3p3.n2441 vdd3p3.n1855 104.756
R1692 vdd3p3.n2437 vdd3p3.n1858 104.756
R1693 vdd3p3.n1283 vdd3p3.n1101 104.756
R1694 vdd3p3.n1283 vdd3p3.n1103 104.756
R1695 vdd3p3.n1279 vdd3p3.n1103 104.756
R1696 vdd3p3.n1279 vdd3p3.n1105 104.756
R1697 vdd3p3.n1275 vdd3p3.n1105 104.756
R1698 vdd3p3.n1275 vdd3p3.n1107 104.756
R1699 vdd3p3.n1271 vdd3p3.n1107 104.756
R1700 vdd3p3.n1271 vdd3p3.n1109 104.756
R1701 vdd3p3.n1267 vdd3p3.n1109 104.756
R1702 vdd3p3.n1267 vdd3p3.n1111 104.756
R1703 vdd3p3.n1263 vdd3p3.n1111 104.756
R1704 vdd3p3.n1263 vdd3p3.n1113 104.756
R1705 vdd3p3.n1259 vdd3p3.n1113 104.756
R1706 vdd3p3.n1259 vdd3p3.n1115 104.756
R1707 vdd3p3.n1255 vdd3p3.n1115 104.756
R1708 vdd3p3.n1255 vdd3p3.n1117 104.756
R1709 vdd3p3.n1251 vdd3p3.n1117 104.756
R1710 vdd3p3.n1251 vdd3p3.n1119 104.756
R1711 vdd3p3.n1247 vdd3p3.n1119 104.756
R1712 vdd3p3.n1247 vdd3p3.n1121 104.756
R1713 vdd3p3.n1243 vdd3p3.n1121 104.756
R1714 vdd3p3.n1243 vdd3p3.n1123 104.756
R1715 vdd3p3.n1239 vdd3p3.n1123 104.756
R1716 vdd3p3.n1239 vdd3p3.n1125 104.756
R1717 vdd3p3.n1235 vdd3p3.n1125 104.756
R1718 vdd3p3.n1235 vdd3p3.n1127 104.756
R1719 vdd3p3.n1231 vdd3p3.n1127 104.756
R1720 vdd3p3.n1299 vdd3p3.n1097 104.756
R1721 vdd3p3.n1299 vdd3p3.n1095 104.756
R1722 vdd3p3.n1303 vdd3p3.n1095 104.756
R1723 vdd3p3.n1303 vdd3p3.n1093 104.756
R1724 vdd3p3.n1307 vdd3p3.n1093 104.756
R1725 vdd3p3.n1307 vdd3p3.n1091 104.756
R1726 vdd3p3.n1311 vdd3p3.n1091 104.756
R1727 vdd3p3.n1311 vdd3p3.n1089 104.756
R1728 vdd3p3.n1315 vdd3p3.n1089 104.756
R1729 vdd3p3.n1315 vdd3p3.n1087 104.756
R1730 vdd3p3.n1319 vdd3p3.n1087 104.756
R1731 vdd3p3.n1319 vdd3p3.n1085 104.756
R1732 vdd3p3.n1324 vdd3p3.n1085 104.756
R1733 vdd3p3.n1324 vdd3p3.n1083 104.756
R1734 vdd3p3.n1495 vdd3p3.n1083 104.756
R1735 vdd3p3.n1474 vdd3p3.n1075 104.756
R1736 vdd3p3.n1398 vdd3p3.n1075 104.756
R1737 vdd3p3.n1402 vdd3p3.n1401 104.756
R1738 vdd3p3.n1499 vdd3p3.n1061 104.756
R1739 vdd3p3.n1503 vdd3p3.n1061 104.756
R1740 vdd3p3.n1503 vdd3p3.n1059 104.756
R1741 vdd3p3.n1507 vdd3p3.n1059 104.756
R1742 vdd3p3.n1507 vdd3p3.n1057 104.756
R1743 vdd3p3.n1511 vdd3p3.n1057 104.756
R1744 vdd3p3.n1511 vdd3p3.n1055 104.756
R1745 vdd3p3.n1515 vdd3p3.n1055 104.756
R1746 vdd3p3.n1515 vdd3p3.n1053 104.756
R1747 vdd3p3.n1519 vdd3p3.n1053 104.756
R1748 vdd3p3.n1519 vdd3p3.n1051 104.756
R1749 vdd3p3.n1523 vdd3p3.n1051 104.756
R1750 vdd3p3.n1523 vdd3p3.n1048 104.756
R1751 vdd3p3.n1528 vdd3p3.n1048 104.756
R1752 vdd3p3.n1528 vdd3p3.n1049 104.756
R1753 vdd3p3.n1532 vdd3p3.n1045 104.756
R1754 vdd3p3.n1536 vdd3p3.n1043 104.756
R1755 vdd3p3.n1536 vdd3p3.n1041 104.756
R1756 vdd3p3.n1540 vdd3p3.n1041 104.756
R1757 vdd3p3.n1540 vdd3p3.n1039 104.756
R1758 vdd3p3.n1544 vdd3p3.n1039 104.756
R1759 vdd3p3.n1544 vdd3p3.n1037 104.756
R1760 vdd3p3.n1548 vdd3p3.n1037 104.756
R1761 vdd3p3.n1548 vdd3p3.n1035 104.756
R1762 vdd3p3.n1552 vdd3p3.n1035 104.756
R1763 vdd3p3.n1552 vdd3p3.n1033 104.756
R1764 vdd3p3.n1556 vdd3p3.n1033 104.756
R1765 vdd3p3.n1556 vdd3p3.n1031 104.756
R1766 vdd3p3.n1560 vdd3p3.n1031 104.756
R1767 vdd3p3.n1560 vdd3p3.n1029 104.756
R1768 vdd3p3.n1564 vdd3p3.n1029 104.756
R1769 vdd3p3.n1564 vdd3p3.n1027 104.756
R1770 vdd3p3.n1568 vdd3p3.n1027 104.756
R1771 vdd3p3.n1568 vdd3p3.n1025 104.756
R1772 vdd3p3.n1572 vdd3p3.n1025 104.756
R1773 vdd3p3.n1572 vdd3p3.n1023 104.756
R1774 vdd3p3.n1576 vdd3p3.n1023 104.756
R1775 vdd3p3.n1576 vdd3p3.n1021 104.756
R1776 vdd3p3.n1580 vdd3p3.n1021 104.756
R1777 vdd3p3.n1580 vdd3p3.n1019 104.756
R1778 vdd3p3.n1584 vdd3p3.n1019 104.756
R1779 vdd3p3.n1584 vdd3p3.n1017 104.756
R1780 vdd3p3.n1588 vdd3p3.n1017 104.756
R1781 vdd3p3.n1588 vdd3p3.n1014 104.756
R1782 vdd3p3.n1227 vdd3p3.n1226 104.756
R1783 vdd3p3.n1224 vdd3p3.n1133 104.756
R1784 vdd3p3.n1220 vdd3p3.n1133 104.756
R1785 vdd3p3.n1220 vdd3p3.n1135 104.756
R1786 vdd3p3.n1216 vdd3p3.n1135 104.756
R1787 vdd3p3.n1216 vdd3p3.n1138 104.756
R1788 vdd3p3.n1212 vdd3p3.n1138 104.756
R1789 vdd3p3.n1212 vdd3p3.n1140 104.756
R1790 vdd3p3.n1208 vdd3p3.n1140 104.756
R1791 vdd3p3.n1208 vdd3p3.n1142 104.756
R1792 vdd3p3.n1204 vdd3p3.n1142 104.756
R1793 vdd3p3.n1204 vdd3p3.n1144 104.756
R1794 vdd3p3.n1200 vdd3p3.n1144 104.756
R1795 vdd3p3.n1200 vdd3p3.n1146 104.756
R1796 vdd3p3.n1196 vdd3p3.n1146 104.756
R1797 vdd3p3.n1196 vdd3p3.n1193 104.756
R1798 vdd3p3.n1188 vdd3p3.n1187 104.756
R1799 vdd3p3.n1179 vdd3p3.n1157 104.756
R1800 vdd3p3.n1177 vdd3p3.n1158 104.756
R1801 vdd3p3.n1170 vdd3p3.n1169 104.756
R1802 vdd3p3.n1646 vdd3p3.n1645 104.756
R1803 vdd3p3.n1638 vdd3p3.n988 104.756
R1804 vdd3p3.n1636 vdd3p3.n989 104.756
R1805 vdd3p3.n1628 vdd3p3.n1627 104.756
R1806 vdd3p3.n1625 vdd3p3.n995 104.756
R1807 vdd3p3.n1620 vdd3p3.n995 104.756
R1808 vdd3p3.n1620 vdd3p3.n997 104.756
R1809 vdd3p3.n1616 vdd3p3.n997 104.756
R1810 vdd3p3.n1616 vdd3p3.n1000 104.756
R1811 vdd3p3.n1612 vdd3p3.n1000 104.756
R1812 vdd3p3.n1612 vdd3p3.n1002 104.756
R1813 vdd3p3.n1608 vdd3p3.n1002 104.756
R1814 vdd3p3.n1608 vdd3p3.n1004 104.756
R1815 vdd3p3.n1604 vdd3p3.n1004 104.756
R1816 vdd3p3.n1604 vdd3p3.n1006 104.756
R1817 vdd3p3.n1600 vdd3p3.n1006 104.756
R1818 vdd3p3.n1600 vdd3p3.n1008 104.756
R1819 vdd3p3.n1596 vdd3p3.n1008 104.756
R1820 vdd3p3.n1596 vdd3p3.n1010 104.756
R1821 vdd3p3.n1592 vdd3p3.n1013 104.756
R1822 vdd3p3.n437 vdd3p3.n255 104.756
R1823 vdd3p3.n437 vdd3p3.n257 104.756
R1824 vdd3p3.n433 vdd3p3.n257 104.756
R1825 vdd3p3.n433 vdd3p3.n259 104.756
R1826 vdd3p3.n429 vdd3p3.n259 104.756
R1827 vdd3p3.n429 vdd3p3.n261 104.756
R1828 vdd3p3.n425 vdd3p3.n261 104.756
R1829 vdd3p3.n425 vdd3p3.n263 104.756
R1830 vdd3p3.n421 vdd3p3.n263 104.756
R1831 vdd3p3.n421 vdd3p3.n265 104.756
R1832 vdd3p3.n417 vdd3p3.n265 104.756
R1833 vdd3p3.n417 vdd3p3.n267 104.756
R1834 vdd3p3.n413 vdd3p3.n267 104.756
R1835 vdd3p3.n413 vdd3p3.n269 104.756
R1836 vdd3p3.n409 vdd3p3.n269 104.756
R1837 vdd3p3.n409 vdd3p3.n271 104.756
R1838 vdd3p3.n405 vdd3p3.n271 104.756
R1839 vdd3p3.n405 vdd3p3.n273 104.756
R1840 vdd3p3.n401 vdd3p3.n273 104.756
R1841 vdd3p3.n401 vdd3p3.n275 104.756
R1842 vdd3p3.n397 vdd3p3.n275 104.756
R1843 vdd3p3.n397 vdd3p3.n277 104.756
R1844 vdd3p3.n393 vdd3p3.n277 104.756
R1845 vdd3p3.n393 vdd3p3.n279 104.756
R1846 vdd3p3.n389 vdd3p3.n279 104.756
R1847 vdd3p3.n389 vdd3p3.n281 104.756
R1848 vdd3p3.n385 vdd3p3.n281 104.756
R1849 vdd3p3.n453 vdd3p3.n251 104.756
R1850 vdd3p3.n453 vdd3p3.n249 104.756
R1851 vdd3p3.n457 vdd3p3.n249 104.756
R1852 vdd3p3.n457 vdd3p3.n247 104.756
R1853 vdd3p3.n461 vdd3p3.n247 104.756
R1854 vdd3p3.n461 vdd3p3.n245 104.756
R1855 vdd3p3.n465 vdd3p3.n245 104.756
R1856 vdd3p3.n465 vdd3p3.n243 104.756
R1857 vdd3p3.n469 vdd3p3.n243 104.756
R1858 vdd3p3.n469 vdd3p3.n241 104.756
R1859 vdd3p3.n473 vdd3p3.n241 104.756
R1860 vdd3p3.n473 vdd3p3.n239 104.756
R1861 vdd3p3.n478 vdd3p3.n239 104.756
R1862 vdd3p3.n478 vdd3p3.n237 104.756
R1863 vdd3p3.n649 vdd3p3.n237 104.756
R1864 vdd3p3.n628 vdd3p3.n229 104.756
R1865 vdd3p3.n552 vdd3p3.n229 104.756
R1866 vdd3p3.n556 vdd3p3.n555 104.756
R1867 vdd3p3.n653 vdd3p3.n215 104.756
R1868 vdd3p3.n657 vdd3p3.n215 104.756
R1869 vdd3p3.n657 vdd3p3.n213 104.756
R1870 vdd3p3.n661 vdd3p3.n213 104.756
R1871 vdd3p3.n661 vdd3p3.n211 104.756
R1872 vdd3p3.n665 vdd3p3.n211 104.756
R1873 vdd3p3.n665 vdd3p3.n209 104.756
R1874 vdd3p3.n669 vdd3p3.n209 104.756
R1875 vdd3p3.n669 vdd3p3.n207 104.756
R1876 vdd3p3.n673 vdd3p3.n207 104.756
R1877 vdd3p3.n673 vdd3p3.n205 104.756
R1878 vdd3p3.n677 vdd3p3.n205 104.756
R1879 vdd3p3.n677 vdd3p3.n202 104.756
R1880 vdd3p3.n682 vdd3p3.n202 104.756
R1881 vdd3p3.n682 vdd3p3.n203 104.756
R1882 vdd3p3.n686 vdd3p3.n199 104.756
R1883 vdd3p3.n690 vdd3p3.n197 104.756
R1884 vdd3p3.n690 vdd3p3.n195 104.756
R1885 vdd3p3.n694 vdd3p3.n195 104.756
R1886 vdd3p3.n694 vdd3p3.n193 104.756
R1887 vdd3p3.n698 vdd3p3.n193 104.756
R1888 vdd3p3.n698 vdd3p3.n191 104.756
R1889 vdd3p3.n702 vdd3p3.n191 104.756
R1890 vdd3p3.n702 vdd3p3.n189 104.756
R1891 vdd3p3.n706 vdd3p3.n189 104.756
R1892 vdd3p3.n706 vdd3p3.n187 104.756
R1893 vdd3p3.n710 vdd3p3.n187 104.756
R1894 vdd3p3.n710 vdd3p3.n185 104.756
R1895 vdd3p3.n714 vdd3p3.n185 104.756
R1896 vdd3p3.n714 vdd3p3.n183 104.756
R1897 vdd3p3.n718 vdd3p3.n183 104.756
R1898 vdd3p3.n718 vdd3p3.n181 104.756
R1899 vdd3p3.n722 vdd3p3.n181 104.756
R1900 vdd3p3.n722 vdd3p3.n179 104.756
R1901 vdd3p3.n726 vdd3p3.n179 104.756
R1902 vdd3p3.n726 vdd3p3.n177 104.756
R1903 vdd3p3.n730 vdd3p3.n177 104.756
R1904 vdd3p3.n730 vdd3p3.n175 104.756
R1905 vdd3p3.n734 vdd3p3.n175 104.756
R1906 vdd3p3.n734 vdd3p3.n173 104.756
R1907 vdd3p3.n738 vdd3p3.n173 104.756
R1908 vdd3p3.n738 vdd3p3.n171 104.756
R1909 vdd3p3.n742 vdd3p3.n171 104.756
R1910 vdd3p3.n742 vdd3p3.n168 104.756
R1911 vdd3p3.n381 vdd3p3.n380 104.756
R1912 vdd3p3.n378 vdd3p3.n287 104.756
R1913 vdd3p3.n374 vdd3p3.n287 104.756
R1914 vdd3p3.n374 vdd3p3.n289 104.756
R1915 vdd3p3.n370 vdd3p3.n289 104.756
R1916 vdd3p3.n370 vdd3p3.n292 104.756
R1917 vdd3p3.n366 vdd3p3.n292 104.756
R1918 vdd3p3.n366 vdd3p3.n294 104.756
R1919 vdd3p3.n362 vdd3p3.n294 104.756
R1920 vdd3p3.n362 vdd3p3.n296 104.756
R1921 vdd3p3.n358 vdd3p3.n296 104.756
R1922 vdd3p3.n358 vdd3p3.n298 104.756
R1923 vdd3p3.n354 vdd3p3.n298 104.756
R1924 vdd3p3.n354 vdd3p3.n300 104.756
R1925 vdd3p3.n350 vdd3p3.n300 104.756
R1926 vdd3p3.n350 vdd3p3.n347 104.756
R1927 vdd3p3.n342 vdd3p3.n341 104.756
R1928 vdd3p3.n333 vdd3p3.n311 104.756
R1929 vdd3p3.n331 vdd3p3.n312 104.756
R1930 vdd3p3.n324 vdd3p3.n323 104.756
R1931 vdd3p3.n800 vdd3p3.n799 104.756
R1932 vdd3p3.n792 vdd3p3.n142 104.756
R1933 vdd3p3.n790 vdd3p3.n143 104.756
R1934 vdd3p3.n782 vdd3p3.n781 104.756
R1935 vdd3p3.n779 vdd3p3.n149 104.756
R1936 vdd3p3.n774 vdd3p3.n149 104.756
R1937 vdd3p3.n774 vdd3p3.n151 104.756
R1938 vdd3p3.n770 vdd3p3.n151 104.756
R1939 vdd3p3.n770 vdd3p3.n154 104.756
R1940 vdd3p3.n766 vdd3p3.n154 104.756
R1941 vdd3p3.n766 vdd3p3.n156 104.756
R1942 vdd3p3.n762 vdd3p3.n156 104.756
R1943 vdd3p3.n762 vdd3p3.n158 104.756
R1944 vdd3p3.n758 vdd3p3.n158 104.756
R1945 vdd3p3.n758 vdd3p3.n160 104.756
R1946 vdd3p3.n754 vdd3p3.n160 104.756
R1947 vdd3p3.n754 vdd3p3.n162 104.756
R1948 vdd3p3.n750 vdd3p3.n162 104.756
R1949 vdd3p3.n750 vdd3p3.n164 104.756
R1950 vdd3p3.n746 vdd3p3.n167 104.756
R1951 vdd3p3.n2922 vdd3p3.n2921 96.863
R1952 vdd3p3.n2076 vdd3p3.n2075 96.863
R1953 vdd3p3.n1231 vdd3p3.n1230 96.863
R1954 vdd3p3.n385 vdd3p3.n384 96.863
R1955 vdd3p3.t122 vdd3p3.n29 96.826
R1956 vdd3p3.n868 vdd3p3.t157 96.826
R1957 vdd3p3.t13 vdd3p3.n1720 96.826
R1958 vdd3p3.n2559 vdd3p3.t79 96.826
R1959 vdd3p3.n2827 vdd3p3.n2819 96.507
R1960 vdd3p3.n2989 vdd3p3.n2988 96.507
R1961 vdd3p3.n1981 vdd3p3.n1973 96.507
R1962 vdd3p3.n2143 vdd3p3.n2142 96.507
R1963 vdd3p3.n1136 vdd3p3.n1128 96.507
R1964 vdd3p3.n1298 vdd3p3.n1297 96.507
R1965 vdd3p3.n290 vdd3p3.n282 96.507
R1966 vdd3p3.n452 vdd3p3.n451 96.507
R1967 vdd3p3.n3021 vdd3p3.n3018 92.5
R1968 vdd3p3.n3161 vdd3p3.n3021 92.5
R1969 vdd3p3.n2628 vdd3p3.n2627 92.5
R1970 vdd3p3.n2640 vdd3p3.n2628 92.5
R1971 vdd3p3.n3359 vdd3p3.n3358 92.5
R1972 vdd3p3.n3358 vdd3p3.n3357 92.5
R1973 vdd3p3.n3360 vdd3p3.n2625 92.5
R1974 vdd3p3.n2630 vdd3p3.n2625 92.5
R1975 vdd3p3.n3362 vdd3p3.n3361 92.5
R1976 vdd3p3.n3363 vdd3p3.n3362 92.5
R1977 vdd3p3.n2626 vdd3p3.n2624 92.5
R1978 vdd3p3.n2624 vdd3p3.n2619 92.5
R1979 vdd3p3.n3055 vdd3p3.n3054 92.5
R1980 vdd3p3.n3055 vdd3p3.n2618 92.5
R1981 vdd3p3.n3060 vdd3p3.n3052 92.5
R1982 vdd3p3.n3062 vdd3p3.n3061 92.5
R1983 vdd3p3.n3064 vdd3p3.n3051 92.5
R1984 vdd3p3.n3066 vdd3p3.n3065 92.5
R1985 vdd3p3.n3068 vdd3p3.n3067 92.5
R1986 vdd3p3.n3059 vdd3p3.n3058 92.5
R1987 vdd3p3.n3047 vdd3p3.n3046 92.5
R1988 vdd3p3.n3074 vdd3p3.n3047 92.5
R1989 vdd3p3.n3149 vdd3p3.n3148 92.5
R1990 vdd3p3.n3148 vdd3p3.n3147 92.5
R1991 vdd3p3.n3150 vdd3p3.n3044 92.5
R1992 vdd3p3.n3048 vdd3p3.n3044 92.5
R1993 vdd3p3.n3152 vdd3p3.n3151 92.5
R1994 vdd3p3.n3153 vdd3p3.n3152 92.5
R1995 vdd3p3.n3045 vdd3p3.n3043 92.5
R1996 vdd3p3.n3043 vdd3p3.n3035 92.5
R1997 vdd3p3.n3192 vdd3p3.n2752 92.5
R1998 vdd3p3.n2752 vdd3p3.n2751 92.5
R1999 vdd3p3.n3215 vdd3p3.n3214 92.5
R2000 vdd3p3.n3214 vdd3p3.n3213 92.5
R2001 vdd3p3.n2742 vdd3p3.n2741 92.5
R2002 vdd3p3.n3212 vdd3p3.n2742 92.5
R2003 vdd3p3.n3210 vdd3p3.n3209 92.5
R2004 vdd3p3.n3211 vdd3p3.n3210 92.5
R2005 vdd3p3.n3208 vdd3p3.n2744 92.5
R2006 vdd3p3.n2744 vdd3p3.n2743 92.5
R2007 vdd3p3.n3207 vdd3p3.n3206 92.5
R2008 vdd3p3.n3206 vdd3p3.n3205 92.5
R2009 vdd3p3.n2746 vdd3p3.n2745 92.5
R2010 vdd3p3.n3204 vdd3p3.n2746 92.5
R2011 vdd3p3.n3202 vdd3p3.n3201 92.5
R2012 vdd3p3.n3203 vdd3p3.n3202 92.5
R2013 vdd3p3.n3200 vdd3p3.n2748 92.5
R2014 vdd3p3.n2748 vdd3p3.n2747 92.5
R2015 vdd3p3.n3199 vdd3p3.n3198 92.5
R2016 vdd3p3.n3198 vdd3p3.n3197 92.5
R2017 vdd3p3.n2750 vdd3p3.n2749 92.5
R2018 vdd3p3.n3196 vdd3p3.n2750 92.5
R2019 vdd3p3.n3194 vdd3p3.n3193 92.5
R2020 vdd3p3.n3195 vdd3p3.n3194 92.5
R2021 vdd3p3.n3216 vdd3p3.n2739 92.5
R2022 vdd3p3.n2739 vdd3p3.n2738 92.5
R2023 vdd3p3.n3219 vdd3p3.n3218 92.5
R2024 vdd3p3.n3220 vdd3p3.n3219 92.5
R2025 vdd3p3.n3217 vdd3p3.n2740 92.5
R2026 vdd3p3.n2736 vdd3p3.n2735 92.5
R2027 vdd3p3.n3224 vdd3p3.n3223 92.5
R2028 vdd3p3.n3223 vdd3p3.n3222 92.5
R2029 vdd3p3.n3227 vdd3p3.n3226 92.5
R2030 vdd3p3.n3228 vdd3p3.n3227 92.5
R2031 vdd3p3.n2732 vdd3p3.n2731 92.5
R2032 vdd3p3.n3229 vdd3p3.n2732 92.5
R2033 vdd3p3.n3232 vdd3p3.n3231 92.5
R2034 vdd3p3.n3231 vdd3p3.n3230 92.5
R2035 vdd3p3.n3233 vdd3p3.n2730 92.5
R2036 vdd3p3.n2730 vdd3p3.n2729 92.5
R2037 vdd3p3.n3235 vdd3p3.n3234 92.5
R2038 vdd3p3.n3236 vdd3p3.n3235 92.5
R2039 vdd3p3.n2728 vdd3p3.n2727 92.5
R2040 vdd3p3.n3237 vdd3p3.n2728 92.5
R2041 vdd3p3.n3240 vdd3p3.n3239 92.5
R2042 vdd3p3.n3239 vdd3p3.n3238 92.5
R2043 vdd3p3.n3241 vdd3p3.n2726 92.5
R2044 vdd3p3.n2726 vdd3p3.n2725 92.5
R2045 vdd3p3.n3243 vdd3p3.n3242 92.5
R2046 vdd3p3.n3244 vdd3p3.n3243 92.5
R2047 vdd3p3.n2724 vdd3p3.n2723 92.5
R2048 vdd3p3.n3245 vdd3p3.n2724 92.5
R2049 vdd3p3.n3248 vdd3p3.n3247 92.5
R2050 vdd3p3.n3247 vdd3p3.n3246 92.5
R2051 vdd3p3.n3249 vdd3p3.n2722 92.5
R2052 vdd3p3.n2722 vdd3p3.n2721 92.5
R2053 vdd3p3.n3251 vdd3p3.n3250 92.5
R2054 vdd3p3.n3252 vdd3p3.n3251 92.5
R2055 vdd3p3.n2720 vdd3p3.n2719 92.5
R2056 vdd3p3.n3253 vdd3p3.n2720 92.5
R2057 vdd3p3.n3256 vdd3p3.n3255 92.5
R2058 vdd3p3.n3255 vdd3p3.n3254 92.5
R2059 vdd3p3.n3257 vdd3p3.n2718 92.5
R2060 vdd3p3.n2718 vdd3p3.n2717 92.5
R2061 vdd3p3.n3259 vdd3p3.n3258 92.5
R2062 vdd3p3.n3260 vdd3p3.n3259 92.5
R2063 vdd3p3.n2716 vdd3p3.n2715 92.5
R2064 vdd3p3.n3261 vdd3p3.n2716 92.5
R2065 vdd3p3.n3264 vdd3p3.n3263 92.5
R2066 vdd3p3.n3263 vdd3p3.n3262 92.5
R2067 vdd3p3.n3265 vdd3p3.n2714 92.5
R2068 vdd3p3.n2714 vdd3p3.n2713 92.5
R2069 vdd3p3.n3267 vdd3p3.n3266 92.5
R2070 vdd3p3.n3268 vdd3p3.n3267 92.5
R2071 vdd3p3.n2712 vdd3p3.n2711 92.5
R2072 vdd3p3.n3269 vdd3p3.n2712 92.5
R2073 vdd3p3.n3272 vdd3p3.n3271 92.5
R2074 vdd3p3.n3271 vdd3p3.n3270 92.5
R2075 vdd3p3.n3273 vdd3p3.n2710 92.5
R2076 vdd3p3.n2710 vdd3p3.n2709 92.5
R2077 vdd3p3.n3275 vdd3p3.n3274 92.5
R2078 vdd3p3.n3276 vdd3p3.n3275 92.5
R2079 vdd3p3.n2708 vdd3p3.n2707 92.5
R2080 vdd3p3.n3277 vdd3p3.n2708 92.5
R2081 vdd3p3.n3280 vdd3p3.n3279 92.5
R2082 vdd3p3.n3279 vdd3p3.n3278 92.5
R2083 vdd3p3.n3281 vdd3p3.n2705 92.5
R2084 vdd3p3.n2705 vdd3p3.n2702 92.5
R2085 vdd3p3.n3225 vdd3p3.n2734 92.5
R2086 vdd3p3.n2734 vdd3p3.n2733 92.5
R2087 vdd3p3.n2697 vdd3p3.n2696 92.5
R2088 vdd3p3.n3293 vdd3p3.n2697 92.5
R2089 vdd3p3.n3296 vdd3p3.n3295 92.5
R2090 vdd3p3.n3295 vdd3p3.n3294 92.5
R2091 vdd3p3.n3297 vdd3p3.n2695 92.5
R2092 vdd3p3.n2695 vdd3p3.n2694 92.5
R2093 vdd3p3.n3299 vdd3p3.n3298 92.5
R2094 vdd3p3.n3300 vdd3p3.n3299 92.5
R2095 vdd3p3.n2693 vdd3p3.n2692 92.5
R2096 vdd3p3.n3301 vdd3p3.n2693 92.5
R2097 vdd3p3.n3304 vdd3p3.n3303 92.5
R2098 vdd3p3.n3303 vdd3p3.n3302 92.5
R2099 vdd3p3.n3305 vdd3p3.n2691 92.5
R2100 vdd3p3.n2691 vdd3p3.n2690 92.5
R2101 vdd3p3.n3307 vdd3p3.n3306 92.5
R2102 vdd3p3.n3308 vdd3p3.n3307 92.5
R2103 vdd3p3.n2688 vdd3p3.n2687 92.5
R2104 vdd3p3.n3309 vdd3p3.n2688 92.5
R2105 vdd3p3.n3312 vdd3p3.n3311 92.5
R2106 vdd3p3.n3311 vdd3p3.n3310 92.5
R2107 vdd3p3.n3313 vdd3p3.n2686 92.5
R2108 vdd3p3.n2689 vdd3p3.n2686 92.5
R2109 vdd3p3.n3289 vdd3p3.n2699 92.5
R2110 vdd3p3.n2699 vdd3p3.n2698 92.5
R2111 vdd3p3.n3288 vdd3p3.n3287 92.5
R2112 vdd3p3.n3287 vdd3p3.n3286 92.5
R2113 vdd3p3.n2701 vdd3p3.n2700 92.5
R2114 vdd3p3.n2706 vdd3p3.n2704 92.5
R2115 vdd3p3.n3283 vdd3p3.n3282 92.5
R2116 vdd3p3.n3284 vdd3p3.n3283 92.5
R2117 vdd3p3.n3291 vdd3p3.n3290 92.5
R2118 vdd3p3.n3292 vdd3p3.n3291 92.5
R2119 vdd3p3.n3316 vdd3p3.n3315 92.5
R2120 vdd3p3.n3337 vdd3p3.n2670 92.5
R2121 vdd3p3.n3336 vdd3p3.n3335 92.5
R2122 vdd3p3.n2679 vdd3p3.n2675 92.5
R2123 vdd3p3.n3330 vdd3p3.n3329 92.5
R2124 vdd3p3.n3327 vdd3p3.n3326 92.5
R2125 vdd3p3.n2681 vdd3p3.n2680 92.5
R2126 vdd3p3.n3320 vdd3p3.n3319 92.5
R2127 vdd3p3.n3318 vdd3p3.n2684 92.5
R2128 vdd3p3.n3340 vdd3p3.n3339 92.5
R2129 vdd3p3.n2855 vdd3p3.n2669 92.5
R2130 vdd3p3.n2858 vdd3p3.n2857 92.5
R2131 vdd3p3.n2880 vdd3p3.n2879 92.5
R2132 vdd3p3.n2878 vdd3p3.n2877 92.5
R2133 vdd3p3.n2848 vdd3p3.n2843 92.5
R2134 vdd3p3.n2871 vdd3p3.n2870 92.5
R2135 vdd3p3.n2868 vdd3p3.n2867 92.5
R2136 vdd3p3.n2850 vdd3p3.n2849 92.5
R2137 vdd3p3.n2866 vdd3p3.n2865 92.5
R2138 vdd3p3.n2851 vdd3p3.n2847 92.5
R2139 vdd3p3.n2873 vdd3p3.n2872 92.5
R2140 vdd3p3.n2876 vdd3p3.n2875 92.5
R2141 vdd3p3.n2844 vdd3p3.n2841 92.5
R2142 vdd3p3.n2884 vdd3p3.n2838 92.5
R2143 vdd3p3.n2882 vdd3p3.n2881 92.5
R2144 vdd3p3.n2864 vdd3p3.n2863 92.5
R2145 vdd3p3.n2864 vdd3p3.n2641 92.5
R2146 vdd3p3.n2862 vdd3p3.n2861 92.5
R2147 vdd3p3.n2860 vdd3p3.n2853 92.5
R2148 vdd3p3.n2923 vdd3p3.n2922 92.5
R2149 vdd3p3.n2920 vdd3p3.n2820 92.5
R2150 vdd3p3.n2919 vdd3p3.n2918 92.5
R2151 vdd3p3.n2917 vdd3p3.n2821 92.5
R2152 vdd3p3.n2915 vdd3p3.n2914 92.5
R2153 vdd3p3.n2913 vdd3p3.n2824 92.5
R2154 vdd3p3.n2827 vdd3p3.n2824 92.5
R2155 vdd3p3.n2912 vdd3p3.n2911 92.5
R2156 vdd3p3.n2911 vdd3p3.n2910 92.5
R2157 vdd3p3.n2826 vdd3p3.n2825 92.5
R2158 vdd3p3.n2909 vdd3p3.n2826 92.5
R2159 vdd3p3.n2907 vdd3p3.n2906 92.5
R2160 vdd3p3.n2908 vdd3p3.n2907 92.5
R2161 vdd3p3.n2905 vdd3p3.n2829 92.5
R2162 vdd3p3.n2829 vdd3p3.n2828 92.5
R2163 vdd3p3.n2904 vdd3p3.n2903 92.5
R2164 vdd3p3.n2903 vdd3p3.n2902 92.5
R2165 vdd3p3.n2831 vdd3p3.n2830 92.5
R2166 vdd3p3.n2901 vdd3p3.n2831 92.5
R2167 vdd3p3.n2899 vdd3p3.n2898 92.5
R2168 vdd3p3.n2900 vdd3p3.n2899 92.5
R2169 vdd3p3.n2897 vdd3p3.n2833 92.5
R2170 vdd3p3.n2833 vdd3p3.n2832 92.5
R2171 vdd3p3.n2896 vdd3p3.n2895 92.5
R2172 vdd3p3.n2895 vdd3p3.n2894 92.5
R2173 vdd3p3.n2835 vdd3p3.n2834 92.5
R2174 vdd3p3.n2893 vdd3p3.n2835 92.5
R2175 vdd3p3.n2891 vdd3p3.n2890 92.5
R2176 vdd3p3.n2892 vdd3p3.n2891 92.5
R2177 vdd3p3.n2889 vdd3p3.n2837 92.5
R2178 vdd3p3.n2837 vdd3p3.n2836 92.5
R2179 vdd3p3.n2888 vdd3p3.n2887 92.5
R2180 vdd3p3.n2887 vdd3p3.n2886 92.5
R2181 vdd3p3.n2975 vdd3p3.n2974 92.5
R2182 vdd3p3.n2974 vdd3p3.n2973 92.5
R2183 vdd3p3.n2794 vdd3p3.n2793 92.5
R2184 vdd3p3.n2972 vdd3p3.n2794 92.5
R2185 vdd3p3.n2970 vdd3p3.n2969 92.5
R2186 vdd3p3.n2971 vdd3p3.n2970 92.5
R2187 vdd3p3.n2968 vdd3p3.n2796 92.5
R2188 vdd3p3.n2796 vdd3p3.n2795 92.5
R2189 vdd3p3.n2967 vdd3p3.n2966 92.5
R2190 vdd3p3.n2966 vdd3p3.n2965 92.5
R2191 vdd3p3.n2798 vdd3p3.n2797 92.5
R2192 vdd3p3.n2964 vdd3p3.n2798 92.5
R2193 vdd3p3.n2962 vdd3p3.n2961 92.5
R2194 vdd3p3.n2963 vdd3p3.n2962 92.5
R2195 vdd3p3.n2960 vdd3p3.n2800 92.5
R2196 vdd3p3.n2800 vdd3p3.n2799 92.5
R2197 vdd3p3.n2959 vdd3p3.n2958 92.5
R2198 vdd3p3.n2958 vdd3p3.n2957 92.5
R2199 vdd3p3.n2802 vdd3p3.n2801 92.5
R2200 vdd3p3.n2956 vdd3p3.n2802 92.5
R2201 vdd3p3.n2954 vdd3p3.n2953 92.5
R2202 vdd3p3.n2955 vdd3p3.n2954 92.5
R2203 vdd3p3.n2952 vdd3p3.n2804 92.5
R2204 vdd3p3.n2804 vdd3p3.n2803 92.5
R2205 vdd3p3.n2951 vdd3p3.n2950 92.5
R2206 vdd3p3.n2950 vdd3p3.n2949 92.5
R2207 vdd3p3.n2806 vdd3p3.n2805 92.5
R2208 vdd3p3.n2948 vdd3p3.n2806 92.5
R2209 vdd3p3.n2946 vdd3p3.n2945 92.5
R2210 vdd3p3.n2947 vdd3p3.n2946 92.5
R2211 vdd3p3.n2944 vdd3p3.n2808 92.5
R2212 vdd3p3.n2808 vdd3p3.n2807 92.5
R2213 vdd3p3.n2943 vdd3p3.n2942 92.5
R2214 vdd3p3.n2942 vdd3p3.n2941 92.5
R2215 vdd3p3.n2810 vdd3p3.n2809 92.5
R2216 vdd3p3.n2940 vdd3p3.n2810 92.5
R2217 vdd3p3.n2938 vdd3p3.n2937 92.5
R2218 vdd3p3.n2939 vdd3p3.n2938 92.5
R2219 vdd3p3.n2936 vdd3p3.n2812 92.5
R2220 vdd3p3.n2812 vdd3p3.n2811 92.5
R2221 vdd3p3.n2935 vdd3p3.n2934 92.5
R2222 vdd3p3.n2934 vdd3p3.n2933 92.5
R2223 vdd3p3.n2814 vdd3p3.n2813 92.5
R2224 vdd3p3.n2932 vdd3p3.n2814 92.5
R2225 vdd3p3.n2930 vdd3p3.n2929 92.5
R2226 vdd3p3.n2931 vdd3p3.n2930 92.5
R2227 vdd3p3.n2928 vdd3p3.n2816 92.5
R2228 vdd3p3.n2816 vdd3p3.n2815 92.5
R2229 vdd3p3.n2927 vdd3p3.n2926 92.5
R2230 vdd3p3.n2926 vdd3p3.n2925 92.5
R2231 vdd3p3.n2818 vdd3p3.n2817 92.5
R2232 vdd3p3.n2924 vdd3p3.n2818 92.5
R2233 vdd3p3.n2983 vdd3p3.n2791 92.5
R2234 vdd3p3.n2987 vdd3p3.n2986 92.5
R2235 vdd3p3.n2792 vdd3p3.n2790 92.5
R2236 vdd3p3.n3017 vdd3p3.n2774 92.5
R2237 vdd3p3.n3013 vdd3p3.n2774 92.5
R2238 vdd3p3.n3016 vdd3p3.n3015 92.5
R2239 vdd3p3.n3015 vdd3p3.n3014 92.5
R2240 vdd3p3.n2776 vdd3p3.n2775 92.5
R2241 vdd3p3.n3012 vdd3p3.n2776 92.5
R2242 vdd3p3.n3010 vdd3p3.n3009 92.5
R2243 vdd3p3.n3011 vdd3p3.n3010 92.5
R2244 vdd3p3.n3008 vdd3p3.n2778 92.5
R2245 vdd3p3.n2778 vdd3p3.n2777 92.5
R2246 vdd3p3.n3007 vdd3p3.n3006 92.5
R2247 vdd3p3.n3006 vdd3p3.n3005 92.5
R2248 vdd3p3.n2780 vdd3p3.n2779 92.5
R2249 vdd3p3.n3004 vdd3p3.n2780 92.5
R2250 vdd3p3.n3002 vdd3p3.n3001 92.5
R2251 vdd3p3.n3003 vdd3p3.n3002 92.5
R2252 vdd3p3.n3000 vdd3p3.n2782 92.5
R2253 vdd3p3.n2782 vdd3p3.n2781 92.5
R2254 vdd3p3.n2999 vdd3p3.n2998 92.5
R2255 vdd3p3.n2998 vdd3p3.n2997 92.5
R2256 vdd3p3.n2784 vdd3p3.n2783 92.5
R2257 vdd3p3.n2996 vdd3p3.n2784 92.5
R2258 vdd3p3.n2994 vdd3p3.n2993 92.5
R2259 vdd3p3.n2995 vdd3p3.n2994 92.5
R2260 vdd3p3.n2992 vdd3p3.n2786 92.5
R2261 vdd3p3.n2786 vdd3p3.n2785 92.5
R2262 vdd3p3.n2991 vdd3p3.n2990 92.5
R2263 vdd3p3.n2990 vdd3p3.n2989 92.5
R2264 vdd3p3.n2788 vdd3p3.n2787 92.5
R2265 vdd3p3.n2979 vdd3p3.n2976 92.5
R2266 vdd3p3.n2982 vdd3p3.n2981 92.5
R2267 vdd3p3.n3191 vdd3p3.n3190 92.5
R2268 vdd3p3.n3115 vdd3p3.n2754 92.5
R2269 vdd3p3.n3117 vdd3p3.n3116 92.5
R2270 vdd3p3.n3114 vdd3p3.n3113 92.5
R2271 vdd3p3.n3084 vdd3p3.n3083 92.5
R2272 vdd3p3.n3108 vdd3p3.n3107 92.5
R2273 vdd3p3.n3086 vdd3p3.n3085 92.5
R2274 vdd3p3.n3102 vdd3p3.n3101 92.5
R2275 vdd3p3.n3098 vdd3p3.n3097 92.5
R2276 vdd3p3.n3096 vdd3p3.n3095 92.5
R2277 vdd3p3.n3166 vdd3p3.n3165 92.5
R2278 vdd3p3.n3170 vdd3p3.n3169 92.5
R2279 vdd3p3.n3173 vdd3p3.n3172 92.5
R2280 vdd3p3.n3031 vdd3p3.n3030 92.5
R2281 vdd3p3.n3020 vdd3p3.n3019 92.5
R2282 vdd3p3.n3182 vdd3p3.n3181 92.5
R2283 vdd3p3.n3183 vdd3p3.n2773 92.5
R2284 vdd3p3.n3186 vdd3p3.n3185 92.5
R2285 vdd3p3.n3180 vdd3p3.n3179 92.5
R2286 vdd3p3.n3029 vdd3p3.n3022 92.5
R2287 vdd3p3.n3175 vdd3p3.n3174 92.5
R2288 vdd3p3.n3171 vdd3p3.n3028 92.5
R2289 vdd3p3.n3168 vdd3p3.n3167 92.5
R2290 vdd3p3.n3032 vdd3p3.n2766 92.5
R2291 vdd3p3.n3188 vdd3p3.n2766 92.5
R2292 vdd3p3.n3164 vdd3p3.n3163 92.5
R2293 vdd3p3.n3090 vdd3p3.n3089 92.5
R2294 vdd3p3.n3092 vdd3p3.n3091 92.5
R2295 vdd3p3.n3094 vdd3p3.n3093 92.5
R2296 vdd3p3.n3100 vdd3p3.n3099 92.5
R2297 vdd3p3.n3119 vdd3p3.n3118 92.5
R2298 vdd3p3.n3112 vdd3p3.n3111 92.5
R2299 vdd3p3.n3110 vdd3p3.n3109 92.5
R2300 vdd3p3.n3106 vdd3p3.n3105 92.5
R2301 vdd3p3.n3104 vdd3p3.n3103 92.5
R2302 vdd3p3.n2665 vdd3p3.n2639 92.5
R2303 vdd3p3.n3344 vdd3p3.n3343 92.5
R2304 vdd3p3.n3342 vdd3p3.n3341 92.5
R2305 vdd3p3.n3342 vdd3p3.n2666 92.5
R2306 vdd3p3.n3334 vdd3p3.n3333 92.5
R2307 vdd3p3.n3332 vdd3p3.n3331 92.5
R2308 vdd3p3.n2682 vdd3p3.n2678 92.5
R2309 vdd3p3.n3325 vdd3p3.n3324 92.5
R2310 vdd3p3.n3322 vdd3p3.n3321 92.5
R2311 vdd3p3.n2674 vdd3p3.n2668 92.5
R2312 vdd3p3.n2659 vdd3p3.n2658 92.5
R2313 vdd3p3.n2656 vdd3p3.n2644 92.5
R2314 vdd3p3.n2654 vdd3p3.n2653 92.5
R2315 vdd3p3.n2652 vdd3p3.n2651 92.5
R2316 vdd3p3.n2649 vdd3p3.n2646 92.5
R2317 vdd3p3.n2647 vdd3p3.n2636 92.5
R2318 vdd3p3.n2664 vdd3p3.n2663 92.5
R2319 vdd3p3.n2666 vdd3p3.n2664 92.5
R2320 vdd3p3.n3346 vdd3p3.n3345 92.5
R2321 vdd3p3.n3345 vdd3p3.n3344 92.5
R2322 vdd3p3.n3347 vdd3p3.n2643 92.5
R2323 vdd3p3.n2665 vdd3p3.n2643 92.5
R2324 vdd3p3.n3349 vdd3p3.n3348 92.5
R2325 vdd3p3.n3350 vdd3p3.n3349 92.5
R2326 vdd3p3.n2661 vdd3p3.n2660 92.5
R2327 vdd3p3.n2660 vdd3p3.n2622 92.5
R2328 vdd3p3.n2616 vdd3p3.n2615 92.5
R2329 vdd3p3.n3364 vdd3p3.n2616 92.5
R2330 vdd3p3.n3369 vdd3p3.n3368 92.5
R2331 vdd3p3.n3368 vdd3p3.n3367 92.5
R2332 vdd3p3.n3370 vdd3p3.n2613 92.5
R2333 vdd3p3.n2617 vdd3p3.n2613 92.5
R2334 vdd3p3.n3372 vdd3p3.n3371 92.5
R2335 vdd3p3.n3373 vdd3p3.n3372 92.5
R2336 vdd3p3.n2614 vdd3p3.n2612 92.5
R2337 vdd3p3.n3073 vdd3p3.n2612 92.5
R2338 vdd3p3.n3126 vdd3p3.n3125 92.5
R2339 vdd3p3.n3125 vdd3p3.n3042 92.5
R2340 vdd3p3.n3124 vdd3p3.n3123 92.5
R2341 vdd3p3.n3124 vdd3p3.n3041 92.5
R2342 vdd3p3.n3122 vdd3p3.n3036 92.5
R2343 vdd3p3.n3160 vdd3p3.n3036 92.5
R2344 vdd3p3.n3121 vdd3p3.n3120 92.5
R2345 vdd3p3.n3120 vdd3p3.n3023 92.5
R2346 vdd3p3.n3129 vdd3p3.n3128 92.5
R2347 vdd3p3.n3131 vdd3p3.n3081 92.5
R2348 vdd3p3.n3134 vdd3p3.n3133 92.5
R2349 vdd3p3.n3136 vdd3p3.n3135 92.5
R2350 vdd3p3.n3138 vdd3p3.n3077 92.5
R2351 vdd3p3.n3141 vdd3p3.n3140 92.5
R2352 vdd3p3.n3087 vdd3p3.n3037 92.5
R2353 vdd3p3.n3037 vdd3p3.n3023 92.5
R2354 vdd3p3.n3159 vdd3p3.n3158 92.5
R2355 vdd3p3.n3160 vdd3p3.n3159 92.5
R2356 vdd3p3.n3156 vdd3p3.n3038 92.5
R2357 vdd3p3.n3041 vdd3p3.n3038 92.5
R2358 vdd3p3.n3078 vdd3p3.n3039 92.5
R2359 vdd3p3.n3078 vdd3p3.n3042 92.5
R2360 vdd3p3.n3142 vdd3p3.n2609 92.5
R2361 vdd3p3.n3073 vdd3p3.n2609 92.5
R2362 vdd3p3.n3375 vdd3p3.n3374 92.5
R2363 vdd3p3.n3374 vdd3p3.n3373 92.5
R2364 vdd3p3.n2610 vdd3p3.n2608 92.5
R2365 vdd3p3.n2617 vdd3p3.n2610 92.5
R2366 vdd3p3.n3366 vdd3p3.n2603 92.5
R2367 vdd3p3.n3367 vdd3p3.n3366 92.5
R2368 vdd3p3.n3365 vdd3p3.n2621 92.5
R2369 vdd3p3.n3365 vdd3p3.n3364 92.5
R2370 vdd3p3.n2634 vdd3p3.n2620 92.5
R2371 vdd3p3.n2622 vdd3p3.n2620 92.5
R2372 vdd3p3.n3352 vdd3p3.n3351 92.5
R2373 vdd3p3.n3351 vdd3p3.n3350 92.5
R2374 vdd3p3.n3157 vdd3p3.n3033 92.5
R2375 vdd3p3.n3035 vdd3p3.n3033 92.5
R2376 vdd3p3.n3155 vdd3p3.n3154 92.5
R2377 vdd3p3.n3154 vdd3p3.n3153 92.5
R2378 vdd3p3.n3076 vdd3p3.n3040 92.5
R2379 vdd3p3.n3048 vdd3p3.n3040 92.5
R2380 vdd3p3.n3146 vdd3p3.n3145 92.5
R2381 vdd3p3.n3147 vdd3p3.n3146 92.5
R2382 vdd3p3.n3143 vdd3p3.n3075 92.5
R2383 vdd3p3.n3075 vdd3p3.n3074 92.5
R2384 vdd3p3.n3071 vdd3p3.n2604 92.5
R2385 vdd3p3.n3071 vdd3p3.n2618 92.5
R2386 vdd3p3.n3070 vdd3p3.n3069 92.5
R2387 vdd3p3.n3070 vdd3p3.n2619 92.5
R2388 vdd3p3.n2633 vdd3p3.n2623 92.5
R2389 vdd3p3.n3363 vdd3p3.n2623 92.5
R2390 vdd3p3.n2635 vdd3p3.n2631 92.5
R2391 vdd3p3.n2631 vdd3p3.n2630 92.5
R2392 vdd3p3.n3356 vdd3p3.n3355 92.5
R2393 vdd3p3.n3357 vdd3p3.n3356 92.5
R2394 vdd3p3.n3353 vdd3p3.n2632 92.5
R2395 vdd3p3.n2640 vdd3p3.n2632 92.5
R2396 vdd3p3.n3162 vdd3p3.n3034 92.5
R2397 vdd3p3.n3162 vdd3p3.n3161 92.5
R2398 vdd3p3.n2175 vdd3p3.n2172 92.5
R2399 vdd3p3.n2315 vdd3p3.n2175 92.5
R2400 vdd3p3.n1782 vdd3p3.n1781 92.5
R2401 vdd3p3.n1794 vdd3p3.n1782 92.5
R2402 vdd3p3.n2513 vdd3p3.n2512 92.5
R2403 vdd3p3.n2512 vdd3p3.n2511 92.5
R2404 vdd3p3.n2514 vdd3p3.n1779 92.5
R2405 vdd3p3.n1784 vdd3p3.n1779 92.5
R2406 vdd3p3.n2516 vdd3p3.n2515 92.5
R2407 vdd3p3.n2517 vdd3p3.n2516 92.5
R2408 vdd3p3.n1780 vdd3p3.n1778 92.5
R2409 vdd3p3.n1778 vdd3p3.n1773 92.5
R2410 vdd3p3.n2209 vdd3p3.n2208 92.5
R2411 vdd3p3.n2209 vdd3p3.n1772 92.5
R2412 vdd3p3.n2214 vdd3p3.n2206 92.5
R2413 vdd3p3.n2216 vdd3p3.n2215 92.5
R2414 vdd3p3.n2218 vdd3p3.n2205 92.5
R2415 vdd3p3.n2220 vdd3p3.n2219 92.5
R2416 vdd3p3.n2222 vdd3p3.n2221 92.5
R2417 vdd3p3.n2213 vdd3p3.n2212 92.5
R2418 vdd3p3.n2201 vdd3p3.n2200 92.5
R2419 vdd3p3.n2228 vdd3p3.n2201 92.5
R2420 vdd3p3.n2303 vdd3p3.n2302 92.5
R2421 vdd3p3.n2302 vdd3p3.n2301 92.5
R2422 vdd3p3.n2304 vdd3p3.n2198 92.5
R2423 vdd3p3.n2202 vdd3p3.n2198 92.5
R2424 vdd3p3.n2306 vdd3p3.n2305 92.5
R2425 vdd3p3.n2307 vdd3p3.n2306 92.5
R2426 vdd3p3.n2199 vdd3p3.n2197 92.5
R2427 vdd3p3.n2197 vdd3p3.n2189 92.5
R2428 vdd3p3.n2346 vdd3p3.n1906 92.5
R2429 vdd3p3.n1906 vdd3p3.n1905 92.5
R2430 vdd3p3.n2369 vdd3p3.n2368 92.5
R2431 vdd3p3.n2368 vdd3p3.n2367 92.5
R2432 vdd3p3.n1896 vdd3p3.n1895 92.5
R2433 vdd3p3.n2366 vdd3p3.n1896 92.5
R2434 vdd3p3.n2364 vdd3p3.n2363 92.5
R2435 vdd3p3.n2365 vdd3p3.n2364 92.5
R2436 vdd3p3.n2362 vdd3p3.n1898 92.5
R2437 vdd3p3.n1898 vdd3p3.n1897 92.5
R2438 vdd3p3.n2361 vdd3p3.n2360 92.5
R2439 vdd3p3.n2360 vdd3p3.n2359 92.5
R2440 vdd3p3.n1900 vdd3p3.n1899 92.5
R2441 vdd3p3.n2358 vdd3p3.n1900 92.5
R2442 vdd3p3.n2356 vdd3p3.n2355 92.5
R2443 vdd3p3.n2357 vdd3p3.n2356 92.5
R2444 vdd3p3.n2354 vdd3p3.n1902 92.5
R2445 vdd3p3.n1902 vdd3p3.n1901 92.5
R2446 vdd3p3.n2353 vdd3p3.n2352 92.5
R2447 vdd3p3.n2352 vdd3p3.n2351 92.5
R2448 vdd3p3.n1904 vdd3p3.n1903 92.5
R2449 vdd3p3.n2350 vdd3p3.n1904 92.5
R2450 vdd3p3.n2348 vdd3p3.n2347 92.5
R2451 vdd3p3.n2349 vdd3p3.n2348 92.5
R2452 vdd3p3.n2370 vdd3p3.n1893 92.5
R2453 vdd3p3.n1893 vdd3p3.n1892 92.5
R2454 vdd3p3.n2373 vdd3p3.n2372 92.5
R2455 vdd3p3.n2374 vdd3p3.n2373 92.5
R2456 vdd3p3.n2371 vdd3p3.n1894 92.5
R2457 vdd3p3.n1890 vdd3p3.n1889 92.5
R2458 vdd3p3.n2378 vdd3p3.n2377 92.5
R2459 vdd3p3.n2377 vdd3p3.n2376 92.5
R2460 vdd3p3.n2381 vdd3p3.n2380 92.5
R2461 vdd3p3.n2382 vdd3p3.n2381 92.5
R2462 vdd3p3.n1886 vdd3p3.n1885 92.5
R2463 vdd3p3.n2383 vdd3p3.n1886 92.5
R2464 vdd3p3.n2386 vdd3p3.n2385 92.5
R2465 vdd3p3.n2385 vdd3p3.n2384 92.5
R2466 vdd3p3.n2387 vdd3p3.n1884 92.5
R2467 vdd3p3.n1884 vdd3p3.n1883 92.5
R2468 vdd3p3.n2389 vdd3p3.n2388 92.5
R2469 vdd3p3.n2390 vdd3p3.n2389 92.5
R2470 vdd3p3.n1882 vdd3p3.n1881 92.5
R2471 vdd3p3.n2391 vdd3p3.n1882 92.5
R2472 vdd3p3.n2394 vdd3p3.n2393 92.5
R2473 vdd3p3.n2393 vdd3p3.n2392 92.5
R2474 vdd3p3.n2395 vdd3p3.n1880 92.5
R2475 vdd3p3.n1880 vdd3p3.n1879 92.5
R2476 vdd3p3.n2397 vdd3p3.n2396 92.5
R2477 vdd3p3.n2398 vdd3p3.n2397 92.5
R2478 vdd3p3.n1878 vdd3p3.n1877 92.5
R2479 vdd3p3.n2399 vdd3p3.n1878 92.5
R2480 vdd3p3.n2402 vdd3p3.n2401 92.5
R2481 vdd3p3.n2401 vdd3p3.n2400 92.5
R2482 vdd3p3.n2403 vdd3p3.n1876 92.5
R2483 vdd3p3.n1876 vdd3p3.n1875 92.5
R2484 vdd3p3.n2405 vdd3p3.n2404 92.5
R2485 vdd3p3.n2406 vdd3p3.n2405 92.5
R2486 vdd3p3.n1874 vdd3p3.n1873 92.5
R2487 vdd3p3.n2407 vdd3p3.n1874 92.5
R2488 vdd3p3.n2410 vdd3p3.n2409 92.5
R2489 vdd3p3.n2409 vdd3p3.n2408 92.5
R2490 vdd3p3.n2411 vdd3p3.n1872 92.5
R2491 vdd3p3.n1872 vdd3p3.n1871 92.5
R2492 vdd3p3.n2413 vdd3p3.n2412 92.5
R2493 vdd3p3.n2414 vdd3p3.n2413 92.5
R2494 vdd3p3.n1870 vdd3p3.n1869 92.5
R2495 vdd3p3.n2415 vdd3p3.n1870 92.5
R2496 vdd3p3.n2418 vdd3p3.n2417 92.5
R2497 vdd3p3.n2417 vdd3p3.n2416 92.5
R2498 vdd3p3.n2419 vdd3p3.n1868 92.5
R2499 vdd3p3.n1868 vdd3p3.n1867 92.5
R2500 vdd3p3.n2421 vdd3p3.n2420 92.5
R2501 vdd3p3.n2422 vdd3p3.n2421 92.5
R2502 vdd3p3.n1866 vdd3p3.n1865 92.5
R2503 vdd3p3.n2423 vdd3p3.n1866 92.5
R2504 vdd3p3.n2426 vdd3p3.n2425 92.5
R2505 vdd3p3.n2425 vdd3p3.n2424 92.5
R2506 vdd3p3.n2427 vdd3p3.n1864 92.5
R2507 vdd3p3.n1864 vdd3p3.n1863 92.5
R2508 vdd3p3.n2429 vdd3p3.n2428 92.5
R2509 vdd3p3.n2430 vdd3p3.n2429 92.5
R2510 vdd3p3.n1862 vdd3p3.n1861 92.5
R2511 vdd3p3.n2431 vdd3p3.n1862 92.5
R2512 vdd3p3.n2434 vdd3p3.n2433 92.5
R2513 vdd3p3.n2433 vdd3p3.n2432 92.5
R2514 vdd3p3.n2435 vdd3p3.n1859 92.5
R2515 vdd3p3.n1859 vdd3p3.n1856 92.5
R2516 vdd3p3.n2379 vdd3p3.n1888 92.5
R2517 vdd3p3.n1888 vdd3p3.n1887 92.5
R2518 vdd3p3.n1851 vdd3p3.n1850 92.5
R2519 vdd3p3.n2447 vdd3p3.n1851 92.5
R2520 vdd3p3.n2450 vdd3p3.n2449 92.5
R2521 vdd3p3.n2449 vdd3p3.n2448 92.5
R2522 vdd3p3.n2451 vdd3p3.n1849 92.5
R2523 vdd3p3.n1849 vdd3p3.n1848 92.5
R2524 vdd3p3.n2453 vdd3p3.n2452 92.5
R2525 vdd3p3.n2454 vdd3p3.n2453 92.5
R2526 vdd3p3.n1847 vdd3p3.n1846 92.5
R2527 vdd3p3.n2455 vdd3p3.n1847 92.5
R2528 vdd3p3.n2458 vdd3p3.n2457 92.5
R2529 vdd3p3.n2457 vdd3p3.n2456 92.5
R2530 vdd3p3.n2459 vdd3p3.n1845 92.5
R2531 vdd3p3.n1845 vdd3p3.n1844 92.5
R2532 vdd3p3.n2461 vdd3p3.n2460 92.5
R2533 vdd3p3.n2462 vdd3p3.n2461 92.5
R2534 vdd3p3.n1842 vdd3p3.n1841 92.5
R2535 vdd3p3.n2463 vdd3p3.n1842 92.5
R2536 vdd3p3.n2466 vdd3p3.n2465 92.5
R2537 vdd3p3.n2465 vdd3p3.n2464 92.5
R2538 vdd3p3.n2467 vdd3p3.n1840 92.5
R2539 vdd3p3.n1843 vdd3p3.n1840 92.5
R2540 vdd3p3.n2443 vdd3p3.n1853 92.5
R2541 vdd3p3.n1853 vdd3p3.n1852 92.5
R2542 vdd3p3.n2442 vdd3p3.n2441 92.5
R2543 vdd3p3.n2441 vdd3p3.n2440 92.5
R2544 vdd3p3.n1855 vdd3p3.n1854 92.5
R2545 vdd3p3.n1860 vdd3p3.n1858 92.5
R2546 vdd3p3.n2437 vdd3p3.n2436 92.5
R2547 vdd3p3.n2438 vdd3p3.n2437 92.5
R2548 vdd3p3.n2445 vdd3p3.n2444 92.5
R2549 vdd3p3.n2446 vdd3p3.n2445 92.5
R2550 vdd3p3.n2470 vdd3p3.n2469 92.5
R2551 vdd3p3.n2491 vdd3p3.n1824 92.5
R2552 vdd3p3.n2490 vdd3p3.n2489 92.5
R2553 vdd3p3.n1833 vdd3p3.n1829 92.5
R2554 vdd3p3.n2484 vdd3p3.n2483 92.5
R2555 vdd3p3.n2481 vdd3p3.n2480 92.5
R2556 vdd3p3.n1835 vdd3p3.n1834 92.5
R2557 vdd3p3.n2474 vdd3p3.n2473 92.5
R2558 vdd3p3.n2472 vdd3p3.n1838 92.5
R2559 vdd3p3.n2494 vdd3p3.n2493 92.5
R2560 vdd3p3.n2009 vdd3p3.n1823 92.5
R2561 vdd3p3.n2012 vdd3p3.n2011 92.5
R2562 vdd3p3.n2034 vdd3p3.n2033 92.5
R2563 vdd3p3.n2032 vdd3p3.n2031 92.5
R2564 vdd3p3.n2002 vdd3p3.n1997 92.5
R2565 vdd3p3.n2025 vdd3p3.n2024 92.5
R2566 vdd3p3.n2022 vdd3p3.n2021 92.5
R2567 vdd3p3.n2004 vdd3p3.n2003 92.5
R2568 vdd3p3.n2020 vdd3p3.n2019 92.5
R2569 vdd3p3.n2005 vdd3p3.n2001 92.5
R2570 vdd3p3.n2027 vdd3p3.n2026 92.5
R2571 vdd3p3.n2030 vdd3p3.n2029 92.5
R2572 vdd3p3.n1998 vdd3p3.n1995 92.5
R2573 vdd3p3.n2038 vdd3p3.n1992 92.5
R2574 vdd3p3.n2036 vdd3p3.n2035 92.5
R2575 vdd3p3.n2018 vdd3p3.n2017 92.5
R2576 vdd3p3.n2018 vdd3p3.n1795 92.5
R2577 vdd3p3.n2016 vdd3p3.n2015 92.5
R2578 vdd3p3.n2014 vdd3p3.n2007 92.5
R2579 vdd3p3.n2077 vdd3p3.n2076 92.5
R2580 vdd3p3.n2074 vdd3p3.n1974 92.5
R2581 vdd3p3.n2073 vdd3p3.n2072 92.5
R2582 vdd3p3.n2071 vdd3p3.n1975 92.5
R2583 vdd3p3.n2069 vdd3p3.n2068 92.5
R2584 vdd3p3.n2067 vdd3p3.n1978 92.5
R2585 vdd3p3.n1981 vdd3p3.n1978 92.5
R2586 vdd3p3.n2066 vdd3p3.n2065 92.5
R2587 vdd3p3.n2065 vdd3p3.n2064 92.5
R2588 vdd3p3.n1980 vdd3p3.n1979 92.5
R2589 vdd3p3.n2063 vdd3p3.n1980 92.5
R2590 vdd3p3.n2061 vdd3p3.n2060 92.5
R2591 vdd3p3.n2062 vdd3p3.n2061 92.5
R2592 vdd3p3.n2059 vdd3p3.n1983 92.5
R2593 vdd3p3.n1983 vdd3p3.n1982 92.5
R2594 vdd3p3.n2058 vdd3p3.n2057 92.5
R2595 vdd3p3.n2057 vdd3p3.n2056 92.5
R2596 vdd3p3.n1985 vdd3p3.n1984 92.5
R2597 vdd3p3.n2055 vdd3p3.n1985 92.5
R2598 vdd3p3.n2053 vdd3p3.n2052 92.5
R2599 vdd3p3.n2054 vdd3p3.n2053 92.5
R2600 vdd3p3.n2051 vdd3p3.n1987 92.5
R2601 vdd3p3.n1987 vdd3p3.n1986 92.5
R2602 vdd3p3.n2050 vdd3p3.n2049 92.5
R2603 vdd3p3.n2049 vdd3p3.n2048 92.5
R2604 vdd3p3.n1989 vdd3p3.n1988 92.5
R2605 vdd3p3.n2047 vdd3p3.n1989 92.5
R2606 vdd3p3.n2045 vdd3p3.n2044 92.5
R2607 vdd3p3.n2046 vdd3p3.n2045 92.5
R2608 vdd3p3.n2043 vdd3p3.n1991 92.5
R2609 vdd3p3.n1991 vdd3p3.n1990 92.5
R2610 vdd3p3.n2042 vdd3p3.n2041 92.5
R2611 vdd3p3.n2041 vdd3p3.n2040 92.5
R2612 vdd3p3.n2129 vdd3p3.n2128 92.5
R2613 vdd3p3.n2128 vdd3p3.n2127 92.5
R2614 vdd3p3.n1948 vdd3p3.n1947 92.5
R2615 vdd3p3.n2126 vdd3p3.n1948 92.5
R2616 vdd3p3.n2124 vdd3p3.n2123 92.5
R2617 vdd3p3.n2125 vdd3p3.n2124 92.5
R2618 vdd3p3.n2122 vdd3p3.n1950 92.5
R2619 vdd3p3.n1950 vdd3p3.n1949 92.5
R2620 vdd3p3.n2121 vdd3p3.n2120 92.5
R2621 vdd3p3.n2120 vdd3p3.n2119 92.5
R2622 vdd3p3.n1952 vdd3p3.n1951 92.5
R2623 vdd3p3.n2118 vdd3p3.n1952 92.5
R2624 vdd3p3.n2116 vdd3p3.n2115 92.5
R2625 vdd3p3.n2117 vdd3p3.n2116 92.5
R2626 vdd3p3.n2114 vdd3p3.n1954 92.5
R2627 vdd3p3.n1954 vdd3p3.n1953 92.5
R2628 vdd3p3.n2113 vdd3p3.n2112 92.5
R2629 vdd3p3.n2112 vdd3p3.n2111 92.5
R2630 vdd3p3.n1956 vdd3p3.n1955 92.5
R2631 vdd3p3.n2110 vdd3p3.n1956 92.5
R2632 vdd3p3.n2108 vdd3p3.n2107 92.5
R2633 vdd3p3.n2109 vdd3p3.n2108 92.5
R2634 vdd3p3.n2106 vdd3p3.n1958 92.5
R2635 vdd3p3.n1958 vdd3p3.n1957 92.5
R2636 vdd3p3.n2105 vdd3p3.n2104 92.5
R2637 vdd3p3.n2104 vdd3p3.n2103 92.5
R2638 vdd3p3.n1960 vdd3p3.n1959 92.5
R2639 vdd3p3.n2102 vdd3p3.n1960 92.5
R2640 vdd3p3.n2100 vdd3p3.n2099 92.5
R2641 vdd3p3.n2101 vdd3p3.n2100 92.5
R2642 vdd3p3.n2098 vdd3p3.n1962 92.5
R2643 vdd3p3.n1962 vdd3p3.n1961 92.5
R2644 vdd3p3.n2097 vdd3p3.n2096 92.5
R2645 vdd3p3.n2096 vdd3p3.n2095 92.5
R2646 vdd3p3.n1964 vdd3p3.n1963 92.5
R2647 vdd3p3.n2094 vdd3p3.n1964 92.5
R2648 vdd3p3.n2092 vdd3p3.n2091 92.5
R2649 vdd3p3.n2093 vdd3p3.n2092 92.5
R2650 vdd3p3.n2090 vdd3p3.n1966 92.5
R2651 vdd3p3.n1966 vdd3p3.n1965 92.5
R2652 vdd3p3.n2089 vdd3p3.n2088 92.5
R2653 vdd3p3.n2088 vdd3p3.n2087 92.5
R2654 vdd3p3.n1968 vdd3p3.n1967 92.5
R2655 vdd3p3.n2086 vdd3p3.n1968 92.5
R2656 vdd3p3.n2084 vdd3p3.n2083 92.5
R2657 vdd3p3.n2085 vdd3p3.n2084 92.5
R2658 vdd3p3.n2082 vdd3p3.n1970 92.5
R2659 vdd3p3.n1970 vdd3p3.n1969 92.5
R2660 vdd3p3.n2081 vdd3p3.n2080 92.5
R2661 vdd3p3.n2080 vdd3p3.n2079 92.5
R2662 vdd3p3.n1972 vdd3p3.n1971 92.5
R2663 vdd3p3.n2078 vdd3p3.n1972 92.5
R2664 vdd3p3.n2137 vdd3p3.n1945 92.5
R2665 vdd3p3.n2141 vdd3p3.n2140 92.5
R2666 vdd3p3.n1946 vdd3p3.n1944 92.5
R2667 vdd3p3.n2171 vdd3p3.n1928 92.5
R2668 vdd3p3.n2167 vdd3p3.n1928 92.5
R2669 vdd3p3.n2170 vdd3p3.n2169 92.5
R2670 vdd3p3.n2169 vdd3p3.n2168 92.5
R2671 vdd3p3.n1930 vdd3p3.n1929 92.5
R2672 vdd3p3.n2166 vdd3p3.n1930 92.5
R2673 vdd3p3.n2164 vdd3p3.n2163 92.5
R2674 vdd3p3.n2165 vdd3p3.n2164 92.5
R2675 vdd3p3.n2162 vdd3p3.n1932 92.5
R2676 vdd3p3.n1932 vdd3p3.n1931 92.5
R2677 vdd3p3.n2161 vdd3p3.n2160 92.5
R2678 vdd3p3.n2160 vdd3p3.n2159 92.5
R2679 vdd3p3.n1934 vdd3p3.n1933 92.5
R2680 vdd3p3.n2158 vdd3p3.n1934 92.5
R2681 vdd3p3.n2156 vdd3p3.n2155 92.5
R2682 vdd3p3.n2157 vdd3p3.n2156 92.5
R2683 vdd3p3.n2154 vdd3p3.n1936 92.5
R2684 vdd3p3.n1936 vdd3p3.n1935 92.5
R2685 vdd3p3.n2153 vdd3p3.n2152 92.5
R2686 vdd3p3.n2152 vdd3p3.n2151 92.5
R2687 vdd3p3.n1938 vdd3p3.n1937 92.5
R2688 vdd3p3.n2150 vdd3p3.n1938 92.5
R2689 vdd3p3.n2148 vdd3p3.n2147 92.5
R2690 vdd3p3.n2149 vdd3p3.n2148 92.5
R2691 vdd3p3.n2146 vdd3p3.n1940 92.5
R2692 vdd3p3.n1940 vdd3p3.n1939 92.5
R2693 vdd3p3.n2145 vdd3p3.n2144 92.5
R2694 vdd3p3.n2144 vdd3p3.n2143 92.5
R2695 vdd3p3.n1942 vdd3p3.n1941 92.5
R2696 vdd3p3.n2133 vdd3p3.n2130 92.5
R2697 vdd3p3.n2136 vdd3p3.n2135 92.5
R2698 vdd3p3.n2345 vdd3p3.n2344 92.5
R2699 vdd3p3.n2269 vdd3p3.n1908 92.5
R2700 vdd3p3.n2271 vdd3p3.n2270 92.5
R2701 vdd3p3.n2268 vdd3p3.n2267 92.5
R2702 vdd3p3.n2238 vdd3p3.n2237 92.5
R2703 vdd3p3.n2262 vdd3p3.n2261 92.5
R2704 vdd3p3.n2240 vdd3p3.n2239 92.5
R2705 vdd3p3.n2256 vdd3p3.n2255 92.5
R2706 vdd3p3.n2252 vdd3p3.n2251 92.5
R2707 vdd3p3.n2250 vdd3p3.n2249 92.5
R2708 vdd3p3.n2320 vdd3p3.n2319 92.5
R2709 vdd3p3.n2324 vdd3p3.n2323 92.5
R2710 vdd3p3.n2327 vdd3p3.n2326 92.5
R2711 vdd3p3.n2185 vdd3p3.n2184 92.5
R2712 vdd3p3.n2174 vdd3p3.n2173 92.5
R2713 vdd3p3.n2336 vdd3p3.n2335 92.5
R2714 vdd3p3.n2337 vdd3p3.n1927 92.5
R2715 vdd3p3.n2340 vdd3p3.n2339 92.5
R2716 vdd3p3.n2334 vdd3p3.n2333 92.5
R2717 vdd3p3.n2183 vdd3p3.n2176 92.5
R2718 vdd3p3.n2329 vdd3p3.n2328 92.5
R2719 vdd3p3.n2325 vdd3p3.n2182 92.5
R2720 vdd3p3.n2322 vdd3p3.n2321 92.5
R2721 vdd3p3.n2186 vdd3p3.n1920 92.5
R2722 vdd3p3.n2342 vdd3p3.n1920 92.5
R2723 vdd3p3.n2318 vdd3p3.n2317 92.5
R2724 vdd3p3.n2244 vdd3p3.n2243 92.5
R2725 vdd3p3.n2246 vdd3p3.n2245 92.5
R2726 vdd3p3.n2248 vdd3p3.n2247 92.5
R2727 vdd3p3.n2254 vdd3p3.n2253 92.5
R2728 vdd3p3.n2273 vdd3p3.n2272 92.5
R2729 vdd3p3.n2266 vdd3p3.n2265 92.5
R2730 vdd3p3.n2264 vdd3p3.n2263 92.5
R2731 vdd3p3.n2260 vdd3p3.n2259 92.5
R2732 vdd3p3.n2258 vdd3p3.n2257 92.5
R2733 vdd3p3.n1819 vdd3p3.n1793 92.5
R2734 vdd3p3.n2498 vdd3p3.n2497 92.5
R2735 vdd3p3.n2496 vdd3p3.n2495 92.5
R2736 vdd3p3.n2496 vdd3p3.n1820 92.5
R2737 vdd3p3.n2488 vdd3p3.n2487 92.5
R2738 vdd3p3.n2486 vdd3p3.n2485 92.5
R2739 vdd3p3.n1836 vdd3p3.n1832 92.5
R2740 vdd3p3.n2479 vdd3p3.n2478 92.5
R2741 vdd3p3.n2476 vdd3p3.n2475 92.5
R2742 vdd3p3.n1828 vdd3p3.n1822 92.5
R2743 vdd3p3.n1813 vdd3p3.n1812 92.5
R2744 vdd3p3.n1810 vdd3p3.n1798 92.5
R2745 vdd3p3.n1808 vdd3p3.n1807 92.5
R2746 vdd3p3.n1806 vdd3p3.n1805 92.5
R2747 vdd3p3.n1803 vdd3p3.n1800 92.5
R2748 vdd3p3.n1801 vdd3p3.n1790 92.5
R2749 vdd3p3.n1818 vdd3p3.n1817 92.5
R2750 vdd3p3.n1820 vdd3p3.n1818 92.5
R2751 vdd3p3.n2500 vdd3p3.n2499 92.5
R2752 vdd3p3.n2499 vdd3p3.n2498 92.5
R2753 vdd3p3.n2501 vdd3p3.n1797 92.5
R2754 vdd3p3.n1819 vdd3p3.n1797 92.5
R2755 vdd3p3.n2503 vdd3p3.n2502 92.5
R2756 vdd3p3.n2504 vdd3p3.n2503 92.5
R2757 vdd3p3.n1815 vdd3p3.n1814 92.5
R2758 vdd3p3.n1814 vdd3p3.n1776 92.5
R2759 vdd3p3.n1770 vdd3p3.n1769 92.5
R2760 vdd3p3.n2518 vdd3p3.n1770 92.5
R2761 vdd3p3.n2523 vdd3p3.n2522 92.5
R2762 vdd3p3.n2522 vdd3p3.n2521 92.5
R2763 vdd3p3.n2524 vdd3p3.n1767 92.5
R2764 vdd3p3.n1771 vdd3p3.n1767 92.5
R2765 vdd3p3.n2526 vdd3p3.n2525 92.5
R2766 vdd3p3.n2527 vdd3p3.n2526 92.5
R2767 vdd3p3.n1768 vdd3p3.n1766 92.5
R2768 vdd3p3.n2227 vdd3p3.n1766 92.5
R2769 vdd3p3.n2280 vdd3p3.n2279 92.5
R2770 vdd3p3.n2279 vdd3p3.n2196 92.5
R2771 vdd3p3.n2278 vdd3p3.n2277 92.5
R2772 vdd3p3.n2278 vdd3p3.n2195 92.5
R2773 vdd3p3.n2276 vdd3p3.n2190 92.5
R2774 vdd3p3.n2314 vdd3p3.n2190 92.5
R2775 vdd3p3.n2275 vdd3p3.n2274 92.5
R2776 vdd3p3.n2274 vdd3p3.n2177 92.5
R2777 vdd3p3.n2283 vdd3p3.n2282 92.5
R2778 vdd3p3.n2285 vdd3p3.n2235 92.5
R2779 vdd3p3.n2288 vdd3p3.n2287 92.5
R2780 vdd3p3.n2290 vdd3p3.n2289 92.5
R2781 vdd3p3.n2292 vdd3p3.n2231 92.5
R2782 vdd3p3.n2295 vdd3p3.n2294 92.5
R2783 vdd3p3.n2241 vdd3p3.n2191 92.5
R2784 vdd3p3.n2191 vdd3p3.n2177 92.5
R2785 vdd3p3.n2313 vdd3p3.n2312 92.5
R2786 vdd3p3.n2314 vdd3p3.n2313 92.5
R2787 vdd3p3.n2310 vdd3p3.n2192 92.5
R2788 vdd3p3.n2195 vdd3p3.n2192 92.5
R2789 vdd3p3.n2232 vdd3p3.n2193 92.5
R2790 vdd3p3.n2232 vdd3p3.n2196 92.5
R2791 vdd3p3.n2296 vdd3p3.n1763 92.5
R2792 vdd3p3.n2227 vdd3p3.n1763 92.5
R2793 vdd3p3.n2529 vdd3p3.n2528 92.5
R2794 vdd3p3.n2528 vdd3p3.n2527 92.5
R2795 vdd3p3.n1764 vdd3p3.n1762 92.5
R2796 vdd3p3.n1771 vdd3p3.n1764 92.5
R2797 vdd3p3.n2520 vdd3p3.n1757 92.5
R2798 vdd3p3.n2521 vdd3p3.n2520 92.5
R2799 vdd3p3.n2519 vdd3p3.n1775 92.5
R2800 vdd3p3.n2519 vdd3p3.n2518 92.5
R2801 vdd3p3.n1788 vdd3p3.n1774 92.5
R2802 vdd3p3.n1776 vdd3p3.n1774 92.5
R2803 vdd3p3.n2506 vdd3p3.n2505 92.5
R2804 vdd3p3.n2505 vdd3p3.n2504 92.5
R2805 vdd3p3.n2311 vdd3p3.n2187 92.5
R2806 vdd3p3.n2189 vdd3p3.n2187 92.5
R2807 vdd3p3.n2309 vdd3p3.n2308 92.5
R2808 vdd3p3.n2308 vdd3p3.n2307 92.5
R2809 vdd3p3.n2230 vdd3p3.n2194 92.5
R2810 vdd3p3.n2202 vdd3p3.n2194 92.5
R2811 vdd3p3.n2300 vdd3p3.n2299 92.5
R2812 vdd3p3.n2301 vdd3p3.n2300 92.5
R2813 vdd3p3.n2297 vdd3p3.n2229 92.5
R2814 vdd3p3.n2229 vdd3p3.n2228 92.5
R2815 vdd3p3.n2225 vdd3p3.n1758 92.5
R2816 vdd3p3.n2225 vdd3p3.n1772 92.5
R2817 vdd3p3.n2224 vdd3p3.n2223 92.5
R2818 vdd3p3.n2224 vdd3p3.n1773 92.5
R2819 vdd3p3.n1787 vdd3p3.n1777 92.5
R2820 vdd3p3.n2517 vdd3p3.n1777 92.5
R2821 vdd3p3.n1789 vdd3p3.n1785 92.5
R2822 vdd3p3.n1785 vdd3p3.n1784 92.5
R2823 vdd3p3.n2510 vdd3p3.n2509 92.5
R2824 vdd3p3.n2511 vdd3p3.n2510 92.5
R2825 vdd3p3.n2507 vdd3p3.n1786 92.5
R2826 vdd3p3.n1794 vdd3p3.n1786 92.5
R2827 vdd3p3.n2316 vdd3p3.n2188 92.5
R2828 vdd3p3.n2316 vdd3p3.n2315 92.5
R2829 vdd3p3.n1330 vdd3p3.n1327 92.5
R2830 vdd3p3.n1470 vdd3p3.n1330 92.5
R2831 vdd3p3.n937 vdd3p3.n936 92.5
R2832 vdd3p3.n949 vdd3p3.n937 92.5
R2833 vdd3p3.n1668 vdd3p3.n1667 92.5
R2834 vdd3p3.n1667 vdd3p3.n1666 92.5
R2835 vdd3p3.n1669 vdd3p3.n934 92.5
R2836 vdd3p3.n939 vdd3p3.n934 92.5
R2837 vdd3p3.n1671 vdd3p3.n1670 92.5
R2838 vdd3p3.n1672 vdd3p3.n1671 92.5
R2839 vdd3p3.n935 vdd3p3.n933 92.5
R2840 vdd3p3.n933 vdd3p3.n928 92.5
R2841 vdd3p3.n1364 vdd3p3.n1363 92.5
R2842 vdd3p3.n1364 vdd3p3.n927 92.5
R2843 vdd3p3.n1369 vdd3p3.n1361 92.5
R2844 vdd3p3.n1371 vdd3p3.n1370 92.5
R2845 vdd3p3.n1373 vdd3p3.n1360 92.5
R2846 vdd3p3.n1375 vdd3p3.n1374 92.5
R2847 vdd3p3.n1377 vdd3p3.n1376 92.5
R2848 vdd3p3.n1368 vdd3p3.n1367 92.5
R2849 vdd3p3.n1356 vdd3p3.n1355 92.5
R2850 vdd3p3.n1383 vdd3p3.n1356 92.5
R2851 vdd3p3.n1458 vdd3p3.n1457 92.5
R2852 vdd3p3.n1457 vdd3p3.n1456 92.5
R2853 vdd3p3.n1459 vdd3p3.n1353 92.5
R2854 vdd3p3.n1357 vdd3p3.n1353 92.5
R2855 vdd3p3.n1461 vdd3p3.n1460 92.5
R2856 vdd3p3.n1462 vdd3p3.n1461 92.5
R2857 vdd3p3.n1354 vdd3p3.n1352 92.5
R2858 vdd3p3.n1352 vdd3p3.n1344 92.5
R2859 vdd3p3.n1501 vdd3p3.n1061 92.5
R2860 vdd3p3.n1061 vdd3p3.n1060 92.5
R2861 vdd3p3.n1524 vdd3p3.n1523 92.5
R2862 vdd3p3.n1523 vdd3p3.n1522 92.5
R2863 vdd3p3.n1051 vdd3p3.n1050 92.5
R2864 vdd3p3.n1521 vdd3p3.n1051 92.5
R2865 vdd3p3.n1519 vdd3p3.n1518 92.5
R2866 vdd3p3.n1520 vdd3p3.n1519 92.5
R2867 vdd3p3.n1517 vdd3p3.n1053 92.5
R2868 vdd3p3.n1053 vdd3p3.n1052 92.5
R2869 vdd3p3.n1516 vdd3p3.n1515 92.5
R2870 vdd3p3.n1515 vdd3p3.n1514 92.5
R2871 vdd3p3.n1055 vdd3p3.n1054 92.5
R2872 vdd3p3.n1513 vdd3p3.n1055 92.5
R2873 vdd3p3.n1511 vdd3p3.n1510 92.5
R2874 vdd3p3.n1512 vdd3p3.n1511 92.5
R2875 vdd3p3.n1509 vdd3p3.n1057 92.5
R2876 vdd3p3.n1057 vdd3p3.n1056 92.5
R2877 vdd3p3.n1508 vdd3p3.n1507 92.5
R2878 vdd3p3.n1507 vdd3p3.n1506 92.5
R2879 vdd3p3.n1059 vdd3p3.n1058 92.5
R2880 vdd3p3.n1505 vdd3p3.n1059 92.5
R2881 vdd3p3.n1503 vdd3p3.n1502 92.5
R2882 vdd3p3.n1504 vdd3p3.n1503 92.5
R2883 vdd3p3.n1525 vdd3p3.n1048 92.5
R2884 vdd3p3.n1048 vdd3p3.n1047 92.5
R2885 vdd3p3.n1528 vdd3p3.n1527 92.5
R2886 vdd3p3.n1529 vdd3p3.n1528 92.5
R2887 vdd3p3.n1526 vdd3p3.n1049 92.5
R2888 vdd3p3.n1045 vdd3p3.n1044 92.5
R2889 vdd3p3.n1533 vdd3p3.n1532 92.5
R2890 vdd3p3.n1532 vdd3p3.n1531 92.5
R2891 vdd3p3.n1536 vdd3p3.n1535 92.5
R2892 vdd3p3.n1537 vdd3p3.n1536 92.5
R2893 vdd3p3.n1041 vdd3p3.n1040 92.5
R2894 vdd3p3.n1538 vdd3p3.n1041 92.5
R2895 vdd3p3.n1541 vdd3p3.n1540 92.5
R2896 vdd3p3.n1540 vdd3p3.n1539 92.5
R2897 vdd3p3.n1542 vdd3p3.n1039 92.5
R2898 vdd3p3.n1039 vdd3p3.n1038 92.5
R2899 vdd3p3.n1544 vdd3p3.n1543 92.5
R2900 vdd3p3.n1545 vdd3p3.n1544 92.5
R2901 vdd3p3.n1037 vdd3p3.n1036 92.5
R2902 vdd3p3.n1546 vdd3p3.n1037 92.5
R2903 vdd3p3.n1549 vdd3p3.n1548 92.5
R2904 vdd3p3.n1548 vdd3p3.n1547 92.5
R2905 vdd3p3.n1550 vdd3p3.n1035 92.5
R2906 vdd3p3.n1035 vdd3p3.n1034 92.5
R2907 vdd3p3.n1552 vdd3p3.n1551 92.5
R2908 vdd3p3.n1553 vdd3p3.n1552 92.5
R2909 vdd3p3.n1033 vdd3p3.n1032 92.5
R2910 vdd3p3.n1554 vdd3p3.n1033 92.5
R2911 vdd3p3.n1557 vdd3p3.n1556 92.5
R2912 vdd3p3.n1556 vdd3p3.n1555 92.5
R2913 vdd3p3.n1558 vdd3p3.n1031 92.5
R2914 vdd3p3.n1031 vdd3p3.n1030 92.5
R2915 vdd3p3.n1560 vdd3p3.n1559 92.5
R2916 vdd3p3.n1561 vdd3p3.n1560 92.5
R2917 vdd3p3.n1029 vdd3p3.n1028 92.5
R2918 vdd3p3.n1562 vdd3p3.n1029 92.5
R2919 vdd3p3.n1565 vdd3p3.n1564 92.5
R2920 vdd3p3.n1564 vdd3p3.n1563 92.5
R2921 vdd3p3.n1566 vdd3p3.n1027 92.5
R2922 vdd3p3.n1027 vdd3p3.n1026 92.5
R2923 vdd3p3.n1568 vdd3p3.n1567 92.5
R2924 vdd3p3.n1569 vdd3p3.n1568 92.5
R2925 vdd3p3.n1025 vdd3p3.n1024 92.5
R2926 vdd3p3.n1570 vdd3p3.n1025 92.5
R2927 vdd3p3.n1573 vdd3p3.n1572 92.5
R2928 vdd3p3.n1572 vdd3p3.n1571 92.5
R2929 vdd3p3.n1574 vdd3p3.n1023 92.5
R2930 vdd3p3.n1023 vdd3p3.n1022 92.5
R2931 vdd3p3.n1576 vdd3p3.n1575 92.5
R2932 vdd3p3.n1577 vdd3p3.n1576 92.5
R2933 vdd3p3.n1021 vdd3p3.n1020 92.5
R2934 vdd3p3.n1578 vdd3p3.n1021 92.5
R2935 vdd3p3.n1581 vdd3p3.n1580 92.5
R2936 vdd3p3.n1580 vdd3p3.n1579 92.5
R2937 vdd3p3.n1582 vdd3p3.n1019 92.5
R2938 vdd3p3.n1019 vdd3p3.n1018 92.5
R2939 vdd3p3.n1584 vdd3p3.n1583 92.5
R2940 vdd3p3.n1585 vdd3p3.n1584 92.5
R2941 vdd3p3.n1017 vdd3p3.n1016 92.5
R2942 vdd3p3.n1586 vdd3p3.n1017 92.5
R2943 vdd3p3.n1589 vdd3p3.n1588 92.5
R2944 vdd3p3.n1588 vdd3p3.n1587 92.5
R2945 vdd3p3.n1590 vdd3p3.n1014 92.5
R2946 vdd3p3.n1014 vdd3p3.n1011 92.5
R2947 vdd3p3.n1534 vdd3p3.n1043 92.5
R2948 vdd3p3.n1043 vdd3p3.n1042 92.5
R2949 vdd3p3.n1006 vdd3p3.n1005 92.5
R2950 vdd3p3.n1602 vdd3p3.n1006 92.5
R2951 vdd3p3.n1605 vdd3p3.n1604 92.5
R2952 vdd3p3.n1604 vdd3p3.n1603 92.5
R2953 vdd3p3.n1606 vdd3p3.n1004 92.5
R2954 vdd3p3.n1004 vdd3p3.n1003 92.5
R2955 vdd3p3.n1608 vdd3p3.n1607 92.5
R2956 vdd3p3.n1609 vdd3p3.n1608 92.5
R2957 vdd3p3.n1002 vdd3p3.n1001 92.5
R2958 vdd3p3.n1610 vdd3p3.n1002 92.5
R2959 vdd3p3.n1613 vdd3p3.n1612 92.5
R2960 vdd3p3.n1612 vdd3p3.n1611 92.5
R2961 vdd3p3.n1614 vdd3p3.n1000 92.5
R2962 vdd3p3.n1000 vdd3p3.n999 92.5
R2963 vdd3p3.n1616 vdd3p3.n1615 92.5
R2964 vdd3p3.n1617 vdd3p3.n1616 92.5
R2965 vdd3p3.n997 vdd3p3.n996 92.5
R2966 vdd3p3.n1618 vdd3p3.n997 92.5
R2967 vdd3p3.n1621 vdd3p3.n1620 92.5
R2968 vdd3p3.n1620 vdd3p3.n1619 92.5
R2969 vdd3p3.n1622 vdd3p3.n995 92.5
R2970 vdd3p3.n998 vdd3p3.n995 92.5
R2971 vdd3p3.n1598 vdd3p3.n1008 92.5
R2972 vdd3p3.n1008 vdd3p3.n1007 92.5
R2973 vdd3p3.n1597 vdd3p3.n1596 92.5
R2974 vdd3p3.n1596 vdd3p3.n1595 92.5
R2975 vdd3p3.n1010 vdd3p3.n1009 92.5
R2976 vdd3p3.n1015 vdd3p3.n1013 92.5
R2977 vdd3p3.n1592 vdd3p3.n1591 92.5
R2978 vdd3p3.n1593 vdd3p3.n1592 92.5
R2979 vdd3p3.n1600 vdd3p3.n1599 92.5
R2980 vdd3p3.n1601 vdd3p3.n1600 92.5
R2981 vdd3p3.n1625 vdd3p3.n1624 92.5
R2982 vdd3p3.n1646 vdd3p3.n979 92.5
R2983 vdd3p3.n1645 vdd3p3.n1644 92.5
R2984 vdd3p3.n988 vdd3p3.n984 92.5
R2985 vdd3p3.n1639 vdd3p3.n1638 92.5
R2986 vdd3p3.n1636 vdd3p3.n1635 92.5
R2987 vdd3p3.n990 vdd3p3.n989 92.5
R2988 vdd3p3.n1629 vdd3p3.n1628 92.5
R2989 vdd3p3.n1627 vdd3p3.n993 92.5
R2990 vdd3p3.n1649 vdd3p3.n1648 92.5
R2991 vdd3p3.n1164 vdd3p3.n978 92.5
R2992 vdd3p3.n1167 vdd3p3.n1166 92.5
R2993 vdd3p3.n1189 vdd3p3.n1188 92.5
R2994 vdd3p3.n1187 vdd3p3.n1186 92.5
R2995 vdd3p3.n1157 vdd3p3.n1152 92.5
R2996 vdd3p3.n1180 vdd3p3.n1179 92.5
R2997 vdd3p3.n1177 vdd3p3.n1176 92.5
R2998 vdd3p3.n1159 vdd3p3.n1158 92.5
R2999 vdd3p3.n1175 vdd3p3.n1174 92.5
R3000 vdd3p3.n1160 vdd3p3.n1156 92.5
R3001 vdd3p3.n1182 vdd3p3.n1181 92.5
R3002 vdd3p3.n1185 vdd3p3.n1184 92.5
R3003 vdd3p3.n1153 vdd3p3.n1150 92.5
R3004 vdd3p3.n1193 vdd3p3.n1147 92.5
R3005 vdd3p3.n1191 vdd3p3.n1190 92.5
R3006 vdd3p3.n1173 vdd3p3.n1172 92.5
R3007 vdd3p3.n1173 vdd3p3.n950 92.5
R3008 vdd3p3.n1171 vdd3p3.n1170 92.5
R3009 vdd3p3.n1169 vdd3p3.n1162 92.5
R3010 vdd3p3.n1232 vdd3p3.n1231 92.5
R3011 vdd3p3.n1229 vdd3p3.n1129 92.5
R3012 vdd3p3.n1228 vdd3p3.n1227 92.5
R3013 vdd3p3.n1226 vdd3p3.n1130 92.5
R3014 vdd3p3.n1224 vdd3p3.n1223 92.5
R3015 vdd3p3.n1222 vdd3p3.n1133 92.5
R3016 vdd3p3.n1136 vdd3p3.n1133 92.5
R3017 vdd3p3.n1221 vdd3p3.n1220 92.5
R3018 vdd3p3.n1220 vdd3p3.n1219 92.5
R3019 vdd3p3.n1135 vdd3p3.n1134 92.5
R3020 vdd3p3.n1218 vdd3p3.n1135 92.5
R3021 vdd3p3.n1216 vdd3p3.n1215 92.5
R3022 vdd3p3.n1217 vdd3p3.n1216 92.5
R3023 vdd3p3.n1214 vdd3p3.n1138 92.5
R3024 vdd3p3.n1138 vdd3p3.n1137 92.5
R3025 vdd3p3.n1213 vdd3p3.n1212 92.5
R3026 vdd3p3.n1212 vdd3p3.n1211 92.5
R3027 vdd3p3.n1140 vdd3p3.n1139 92.5
R3028 vdd3p3.n1210 vdd3p3.n1140 92.5
R3029 vdd3p3.n1208 vdd3p3.n1207 92.5
R3030 vdd3p3.n1209 vdd3p3.n1208 92.5
R3031 vdd3p3.n1206 vdd3p3.n1142 92.5
R3032 vdd3p3.n1142 vdd3p3.n1141 92.5
R3033 vdd3p3.n1205 vdd3p3.n1204 92.5
R3034 vdd3p3.n1204 vdd3p3.n1203 92.5
R3035 vdd3p3.n1144 vdd3p3.n1143 92.5
R3036 vdd3p3.n1202 vdd3p3.n1144 92.5
R3037 vdd3p3.n1200 vdd3p3.n1199 92.5
R3038 vdd3p3.n1201 vdd3p3.n1200 92.5
R3039 vdd3p3.n1198 vdd3p3.n1146 92.5
R3040 vdd3p3.n1146 vdd3p3.n1145 92.5
R3041 vdd3p3.n1197 vdd3p3.n1196 92.5
R3042 vdd3p3.n1196 vdd3p3.n1195 92.5
R3043 vdd3p3.n1284 vdd3p3.n1283 92.5
R3044 vdd3p3.n1283 vdd3p3.n1282 92.5
R3045 vdd3p3.n1103 vdd3p3.n1102 92.5
R3046 vdd3p3.n1281 vdd3p3.n1103 92.5
R3047 vdd3p3.n1279 vdd3p3.n1278 92.5
R3048 vdd3p3.n1280 vdd3p3.n1279 92.5
R3049 vdd3p3.n1277 vdd3p3.n1105 92.5
R3050 vdd3p3.n1105 vdd3p3.n1104 92.5
R3051 vdd3p3.n1276 vdd3p3.n1275 92.5
R3052 vdd3p3.n1275 vdd3p3.n1274 92.5
R3053 vdd3p3.n1107 vdd3p3.n1106 92.5
R3054 vdd3p3.n1273 vdd3p3.n1107 92.5
R3055 vdd3p3.n1271 vdd3p3.n1270 92.5
R3056 vdd3p3.n1272 vdd3p3.n1271 92.5
R3057 vdd3p3.n1269 vdd3p3.n1109 92.5
R3058 vdd3p3.n1109 vdd3p3.n1108 92.5
R3059 vdd3p3.n1268 vdd3p3.n1267 92.5
R3060 vdd3p3.n1267 vdd3p3.n1266 92.5
R3061 vdd3p3.n1111 vdd3p3.n1110 92.5
R3062 vdd3p3.n1265 vdd3p3.n1111 92.5
R3063 vdd3p3.n1263 vdd3p3.n1262 92.5
R3064 vdd3p3.n1264 vdd3p3.n1263 92.5
R3065 vdd3p3.n1261 vdd3p3.n1113 92.5
R3066 vdd3p3.n1113 vdd3p3.n1112 92.5
R3067 vdd3p3.n1260 vdd3p3.n1259 92.5
R3068 vdd3p3.n1259 vdd3p3.n1258 92.5
R3069 vdd3p3.n1115 vdd3p3.n1114 92.5
R3070 vdd3p3.n1257 vdd3p3.n1115 92.5
R3071 vdd3p3.n1255 vdd3p3.n1254 92.5
R3072 vdd3p3.n1256 vdd3p3.n1255 92.5
R3073 vdd3p3.n1253 vdd3p3.n1117 92.5
R3074 vdd3p3.n1117 vdd3p3.n1116 92.5
R3075 vdd3p3.n1252 vdd3p3.n1251 92.5
R3076 vdd3p3.n1251 vdd3p3.n1250 92.5
R3077 vdd3p3.n1119 vdd3p3.n1118 92.5
R3078 vdd3p3.n1249 vdd3p3.n1119 92.5
R3079 vdd3p3.n1247 vdd3p3.n1246 92.5
R3080 vdd3p3.n1248 vdd3p3.n1247 92.5
R3081 vdd3p3.n1245 vdd3p3.n1121 92.5
R3082 vdd3p3.n1121 vdd3p3.n1120 92.5
R3083 vdd3p3.n1244 vdd3p3.n1243 92.5
R3084 vdd3p3.n1243 vdd3p3.n1242 92.5
R3085 vdd3p3.n1123 vdd3p3.n1122 92.5
R3086 vdd3p3.n1241 vdd3p3.n1123 92.5
R3087 vdd3p3.n1239 vdd3p3.n1238 92.5
R3088 vdd3p3.n1240 vdd3p3.n1239 92.5
R3089 vdd3p3.n1237 vdd3p3.n1125 92.5
R3090 vdd3p3.n1125 vdd3p3.n1124 92.5
R3091 vdd3p3.n1236 vdd3p3.n1235 92.5
R3092 vdd3p3.n1235 vdd3p3.n1234 92.5
R3093 vdd3p3.n1127 vdd3p3.n1126 92.5
R3094 vdd3p3.n1233 vdd3p3.n1127 92.5
R3095 vdd3p3.n1292 vdd3p3.n1100 92.5
R3096 vdd3p3.n1296 vdd3p3.n1295 92.5
R3097 vdd3p3.n1101 vdd3p3.n1099 92.5
R3098 vdd3p3.n1326 vdd3p3.n1083 92.5
R3099 vdd3p3.n1322 vdd3p3.n1083 92.5
R3100 vdd3p3.n1325 vdd3p3.n1324 92.5
R3101 vdd3p3.n1324 vdd3p3.n1323 92.5
R3102 vdd3p3.n1085 vdd3p3.n1084 92.5
R3103 vdd3p3.n1321 vdd3p3.n1085 92.5
R3104 vdd3p3.n1319 vdd3p3.n1318 92.5
R3105 vdd3p3.n1320 vdd3p3.n1319 92.5
R3106 vdd3p3.n1317 vdd3p3.n1087 92.5
R3107 vdd3p3.n1087 vdd3p3.n1086 92.5
R3108 vdd3p3.n1316 vdd3p3.n1315 92.5
R3109 vdd3p3.n1315 vdd3p3.n1314 92.5
R3110 vdd3p3.n1089 vdd3p3.n1088 92.5
R3111 vdd3p3.n1313 vdd3p3.n1089 92.5
R3112 vdd3p3.n1311 vdd3p3.n1310 92.5
R3113 vdd3p3.n1312 vdd3p3.n1311 92.5
R3114 vdd3p3.n1309 vdd3p3.n1091 92.5
R3115 vdd3p3.n1091 vdd3p3.n1090 92.5
R3116 vdd3p3.n1308 vdd3p3.n1307 92.5
R3117 vdd3p3.n1307 vdd3p3.n1306 92.5
R3118 vdd3p3.n1093 vdd3p3.n1092 92.5
R3119 vdd3p3.n1305 vdd3p3.n1093 92.5
R3120 vdd3p3.n1303 vdd3p3.n1302 92.5
R3121 vdd3p3.n1304 vdd3p3.n1303 92.5
R3122 vdd3p3.n1301 vdd3p3.n1095 92.5
R3123 vdd3p3.n1095 vdd3p3.n1094 92.5
R3124 vdd3p3.n1300 vdd3p3.n1299 92.5
R3125 vdd3p3.n1299 vdd3p3.n1298 92.5
R3126 vdd3p3.n1097 vdd3p3.n1096 92.5
R3127 vdd3p3.n1288 vdd3p3.n1285 92.5
R3128 vdd3p3.n1291 vdd3p3.n1290 92.5
R3129 vdd3p3.n1500 vdd3p3.n1499 92.5
R3130 vdd3p3.n1424 vdd3p3.n1063 92.5
R3131 vdd3p3.n1426 vdd3p3.n1425 92.5
R3132 vdd3p3.n1423 vdd3p3.n1422 92.5
R3133 vdd3p3.n1393 vdd3p3.n1392 92.5
R3134 vdd3p3.n1417 vdd3p3.n1416 92.5
R3135 vdd3p3.n1395 vdd3p3.n1394 92.5
R3136 vdd3p3.n1411 vdd3p3.n1410 92.5
R3137 vdd3p3.n1407 vdd3p3.n1406 92.5
R3138 vdd3p3.n1405 vdd3p3.n1404 92.5
R3139 vdd3p3.n1475 vdd3p3.n1474 92.5
R3140 vdd3p3.n1479 vdd3p3.n1478 92.5
R3141 vdd3p3.n1482 vdd3p3.n1481 92.5
R3142 vdd3p3.n1340 vdd3p3.n1339 92.5
R3143 vdd3p3.n1329 vdd3p3.n1328 92.5
R3144 vdd3p3.n1491 vdd3p3.n1490 92.5
R3145 vdd3p3.n1492 vdd3p3.n1082 92.5
R3146 vdd3p3.n1495 vdd3p3.n1494 92.5
R3147 vdd3p3.n1489 vdd3p3.n1488 92.5
R3148 vdd3p3.n1338 vdd3p3.n1331 92.5
R3149 vdd3p3.n1484 vdd3p3.n1483 92.5
R3150 vdd3p3.n1480 vdd3p3.n1337 92.5
R3151 vdd3p3.n1477 vdd3p3.n1476 92.5
R3152 vdd3p3.n1341 vdd3p3.n1075 92.5
R3153 vdd3p3.n1497 vdd3p3.n1075 92.5
R3154 vdd3p3.n1473 vdd3p3.n1472 92.5
R3155 vdd3p3.n1399 vdd3p3.n1398 92.5
R3156 vdd3p3.n1401 vdd3p3.n1400 92.5
R3157 vdd3p3.n1403 vdd3p3.n1402 92.5
R3158 vdd3p3.n1409 vdd3p3.n1408 92.5
R3159 vdd3p3.n1428 vdd3p3.n1427 92.5
R3160 vdd3p3.n1421 vdd3p3.n1420 92.5
R3161 vdd3p3.n1419 vdd3p3.n1418 92.5
R3162 vdd3p3.n1415 vdd3p3.n1414 92.5
R3163 vdd3p3.n1413 vdd3p3.n1412 92.5
R3164 vdd3p3.n974 vdd3p3.n948 92.5
R3165 vdd3p3.n1653 vdd3p3.n1652 92.5
R3166 vdd3p3.n1651 vdd3p3.n1650 92.5
R3167 vdd3p3.n1651 vdd3p3.n975 92.5
R3168 vdd3p3.n1643 vdd3p3.n1642 92.5
R3169 vdd3p3.n1641 vdd3p3.n1640 92.5
R3170 vdd3p3.n991 vdd3p3.n987 92.5
R3171 vdd3p3.n1634 vdd3p3.n1633 92.5
R3172 vdd3p3.n1631 vdd3p3.n1630 92.5
R3173 vdd3p3.n983 vdd3p3.n977 92.5
R3174 vdd3p3.n968 vdd3p3.n967 92.5
R3175 vdd3p3.n965 vdd3p3.n953 92.5
R3176 vdd3p3.n963 vdd3p3.n962 92.5
R3177 vdd3p3.n961 vdd3p3.n960 92.5
R3178 vdd3p3.n958 vdd3p3.n955 92.5
R3179 vdd3p3.n956 vdd3p3.n945 92.5
R3180 vdd3p3.n973 vdd3p3.n972 92.5
R3181 vdd3p3.n975 vdd3p3.n973 92.5
R3182 vdd3p3.n1655 vdd3p3.n1654 92.5
R3183 vdd3p3.n1654 vdd3p3.n1653 92.5
R3184 vdd3p3.n1656 vdd3p3.n952 92.5
R3185 vdd3p3.n974 vdd3p3.n952 92.5
R3186 vdd3p3.n1658 vdd3p3.n1657 92.5
R3187 vdd3p3.n1659 vdd3p3.n1658 92.5
R3188 vdd3p3.n970 vdd3p3.n969 92.5
R3189 vdd3p3.n969 vdd3p3.n931 92.5
R3190 vdd3p3.n925 vdd3p3.n924 92.5
R3191 vdd3p3.n1673 vdd3p3.n925 92.5
R3192 vdd3p3.n1678 vdd3p3.n1677 92.5
R3193 vdd3p3.n1677 vdd3p3.n1676 92.5
R3194 vdd3p3.n1679 vdd3p3.n922 92.5
R3195 vdd3p3.n926 vdd3p3.n922 92.5
R3196 vdd3p3.n1681 vdd3p3.n1680 92.5
R3197 vdd3p3.n1682 vdd3p3.n1681 92.5
R3198 vdd3p3.n923 vdd3p3.n921 92.5
R3199 vdd3p3.n1382 vdd3p3.n921 92.5
R3200 vdd3p3.n1435 vdd3p3.n1434 92.5
R3201 vdd3p3.n1434 vdd3p3.n1351 92.5
R3202 vdd3p3.n1433 vdd3p3.n1432 92.5
R3203 vdd3p3.n1433 vdd3p3.n1350 92.5
R3204 vdd3p3.n1431 vdd3p3.n1345 92.5
R3205 vdd3p3.n1469 vdd3p3.n1345 92.5
R3206 vdd3p3.n1430 vdd3p3.n1429 92.5
R3207 vdd3p3.n1429 vdd3p3.n1332 92.5
R3208 vdd3p3.n1438 vdd3p3.n1437 92.5
R3209 vdd3p3.n1440 vdd3p3.n1390 92.5
R3210 vdd3p3.n1443 vdd3p3.n1442 92.5
R3211 vdd3p3.n1445 vdd3p3.n1444 92.5
R3212 vdd3p3.n1447 vdd3p3.n1386 92.5
R3213 vdd3p3.n1450 vdd3p3.n1449 92.5
R3214 vdd3p3.n1396 vdd3p3.n1346 92.5
R3215 vdd3p3.n1346 vdd3p3.n1332 92.5
R3216 vdd3p3.n1468 vdd3p3.n1467 92.5
R3217 vdd3p3.n1469 vdd3p3.n1468 92.5
R3218 vdd3p3.n1465 vdd3p3.n1347 92.5
R3219 vdd3p3.n1350 vdd3p3.n1347 92.5
R3220 vdd3p3.n1387 vdd3p3.n1348 92.5
R3221 vdd3p3.n1387 vdd3p3.n1351 92.5
R3222 vdd3p3.n1451 vdd3p3.n918 92.5
R3223 vdd3p3.n1382 vdd3p3.n918 92.5
R3224 vdd3p3.n1684 vdd3p3.n1683 92.5
R3225 vdd3p3.n1683 vdd3p3.n1682 92.5
R3226 vdd3p3.n919 vdd3p3.n917 92.5
R3227 vdd3p3.n926 vdd3p3.n919 92.5
R3228 vdd3p3.n1675 vdd3p3.n912 92.5
R3229 vdd3p3.n1676 vdd3p3.n1675 92.5
R3230 vdd3p3.n1674 vdd3p3.n930 92.5
R3231 vdd3p3.n1674 vdd3p3.n1673 92.5
R3232 vdd3p3.n943 vdd3p3.n929 92.5
R3233 vdd3p3.n931 vdd3p3.n929 92.5
R3234 vdd3p3.n1661 vdd3p3.n1660 92.5
R3235 vdd3p3.n1660 vdd3p3.n1659 92.5
R3236 vdd3p3.n1466 vdd3p3.n1342 92.5
R3237 vdd3p3.n1344 vdd3p3.n1342 92.5
R3238 vdd3p3.n1464 vdd3p3.n1463 92.5
R3239 vdd3p3.n1463 vdd3p3.n1462 92.5
R3240 vdd3p3.n1385 vdd3p3.n1349 92.5
R3241 vdd3p3.n1357 vdd3p3.n1349 92.5
R3242 vdd3p3.n1455 vdd3p3.n1454 92.5
R3243 vdd3p3.n1456 vdd3p3.n1455 92.5
R3244 vdd3p3.n1452 vdd3p3.n1384 92.5
R3245 vdd3p3.n1384 vdd3p3.n1383 92.5
R3246 vdd3p3.n1380 vdd3p3.n913 92.5
R3247 vdd3p3.n1380 vdd3p3.n927 92.5
R3248 vdd3p3.n1379 vdd3p3.n1378 92.5
R3249 vdd3p3.n1379 vdd3p3.n928 92.5
R3250 vdd3p3.n942 vdd3p3.n932 92.5
R3251 vdd3p3.n1672 vdd3p3.n932 92.5
R3252 vdd3p3.n944 vdd3p3.n940 92.5
R3253 vdd3p3.n940 vdd3p3.n939 92.5
R3254 vdd3p3.n1665 vdd3p3.n1664 92.5
R3255 vdd3p3.n1666 vdd3p3.n1665 92.5
R3256 vdd3p3.n1662 vdd3p3.n941 92.5
R3257 vdd3p3.n949 vdd3p3.n941 92.5
R3258 vdd3p3.n1471 vdd3p3.n1343 92.5
R3259 vdd3p3.n1471 vdd3p3.n1470 92.5
R3260 vdd3p3.n484 vdd3p3.n481 92.5
R3261 vdd3p3.n624 vdd3p3.n484 92.5
R3262 vdd3p3.n91 vdd3p3.n90 92.5
R3263 vdd3p3.n103 vdd3p3.n91 92.5
R3264 vdd3p3.n822 vdd3p3.n821 92.5
R3265 vdd3p3.n821 vdd3p3.n820 92.5
R3266 vdd3p3.n823 vdd3p3.n88 92.5
R3267 vdd3p3.n93 vdd3p3.n88 92.5
R3268 vdd3p3.n825 vdd3p3.n824 92.5
R3269 vdd3p3.n826 vdd3p3.n825 92.5
R3270 vdd3p3.n89 vdd3p3.n87 92.5
R3271 vdd3p3.n87 vdd3p3.n82 92.5
R3272 vdd3p3.n518 vdd3p3.n517 92.5
R3273 vdd3p3.n518 vdd3p3.n81 92.5
R3274 vdd3p3.n523 vdd3p3.n515 92.5
R3275 vdd3p3.n525 vdd3p3.n524 92.5
R3276 vdd3p3.n527 vdd3p3.n514 92.5
R3277 vdd3p3.n529 vdd3p3.n528 92.5
R3278 vdd3p3.n531 vdd3p3.n530 92.5
R3279 vdd3p3.n522 vdd3p3.n521 92.5
R3280 vdd3p3.n510 vdd3p3.n509 92.5
R3281 vdd3p3.n537 vdd3p3.n510 92.5
R3282 vdd3p3.n612 vdd3p3.n611 92.5
R3283 vdd3p3.n611 vdd3p3.n610 92.5
R3284 vdd3p3.n613 vdd3p3.n507 92.5
R3285 vdd3p3.n511 vdd3p3.n507 92.5
R3286 vdd3p3.n615 vdd3p3.n614 92.5
R3287 vdd3p3.n616 vdd3p3.n615 92.5
R3288 vdd3p3.n508 vdd3p3.n506 92.5
R3289 vdd3p3.n506 vdd3p3.n498 92.5
R3290 vdd3p3.n655 vdd3p3.n215 92.5
R3291 vdd3p3.n215 vdd3p3.n214 92.5
R3292 vdd3p3.n678 vdd3p3.n677 92.5
R3293 vdd3p3.n677 vdd3p3.n676 92.5
R3294 vdd3p3.n205 vdd3p3.n204 92.5
R3295 vdd3p3.n675 vdd3p3.n205 92.5
R3296 vdd3p3.n673 vdd3p3.n672 92.5
R3297 vdd3p3.n674 vdd3p3.n673 92.5
R3298 vdd3p3.n671 vdd3p3.n207 92.5
R3299 vdd3p3.n207 vdd3p3.n206 92.5
R3300 vdd3p3.n670 vdd3p3.n669 92.5
R3301 vdd3p3.n669 vdd3p3.n668 92.5
R3302 vdd3p3.n209 vdd3p3.n208 92.5
R3303 vdd3p3.n667 vdd3p3.n209 92.5
R3304 vdd3p3.n665 vdd3p3.n664 92.5
R3305 vdd3p3.n666 vdd3p3.n665 92.5
R3306 vdd3p3.n663 vdd3p3.n211 92.5
R3307 vdd3p3.n211 vdd3p3.n210 92.5
R3308 vdd3p3.n662 vdd3p3.n661 92.5
R3309 vdd3p3.n661 vdd3p3.n660 92.5
R3310 vdd3p3.n213 vdd3p3.n212 92.5
R3311 vdd3p3.n659 vdd3p3.n213 92.5
R3312 vdd3p3.n657 vdd3p3.n656 92.5
R3313 vdd3p3.n658 vdd3p3.n657 92.5
R3314 vdd3p3.n679 vdd3p3.n202 92.5
R3315 vdd3p3.n202 vdd3p3.n201 92.5
R3316 vdd3p3.n682 vdd3p3.n681 92.5
R3317 vdd3p3.n683 vdd3p3.n682 92.5
R3318 vdd3p3.n680 vdd3p3.n203 92.5
R3319 vdd3p3.n199 vdd3p3.n198 92.5
R3320 vdd3p3.n687 vdd3p3.n686 92.5
R3321 vdd3p3.n686 vdd3p3.n685 92.5
R3322 vdd3p3.n690 vdd3p3.n689 92.5
R3323 vdd3p3.n691 vdd3p3.n690 92.5
R3324 vdd3p3.n195 vdd3p3.n194 92.5
R3325 vdd3p3.n692 vdd3p3.n195 92.5
R3326 vdd3p3.n695 vdd3p3.n694 92.5
R3327 vdd3p3.n694 vdd3p3.n693 92.5
R3328 vdd3p3.n696 vdd3p3.n193 92.5
R3329 vdd3p3.n193 vdd3p3.n192 92.5
R3330 vdd3p3.n698 vdd3p3.n697 92.5
R3331 vdd3p3.n699 vdd3p3.n698 92.5
R3332 vdd3p3.n191 vdd3p3.n190 92.5
R3333 vdd3p3.n700 vdd3p3.n191 92.5
R3334 vdd3p3.n703 vdd3p3.n702 92.5
R3335 vdd3p3.n702 vdd3p3.n701 92.5
R3336 vdd3p3.n704 vdd3p3.n189 92.5
R3337 vdd3p3.n189 vdd3p3.n188 92.5
R3338 vdd3p3.n706 vdd3p3.n705 92.5
R3339 vdd3p3.n707 vdd3p3.n706 92.5
R3340 vdd3p3.n187 vdd3p3.n186 92.5
R3341 vdd3p3.n708 vdd3p3.n187 92.5
R3342 vdd3p3.n711 vdd3p3.n710 92.5
R3343 vdd3p3.n710 vdd3p3.n709 92.5
R3344 vdd3p3.n712 vdd3p3.n185 92.5
R3345 vdd3p3.n185 vdd3p3.n184 92.5
R3346 vdd3p3.n714 vdd3p3.n713 92.5
R3347 vdd3p3.n715 vdd3p3.n714 92.5
R3348 vdd3p3.n183 vdd3p3.n182 92.5
R3349 vdd3p3.n716 vdd3p3.n183 92.5
R3350 vdd3p3.n719 vdd3p3.n718 92.5
R3351 vdd3p3.n718 vdd3p3.n717 92.5
R3352 vdd3p3.n720 vdd3p3.n181 92.5
R3353 vdd3p3.n181 vdd3p3.n180 92.5
R3354 vdd3p3.n722 vdd3p3.n721 92.5
R3355 vdd3p3.n723 vdd3p3.n722 92.5
R3356 vdd3p3.n179 vdd3p3.n178 92.5
R3357 vdd3p3.n724 vdd3p3.n179 92.5
R3358 vdd3p3.n727 vdd3p3.n726 92.5
R3359 vdd3p3.n726 vdd3p3.n725 92.5
R3360 vdd3p3.n728 vdd3p3.n177 92.5
R3361 vdd3p3.n177 vdd3p3.n176 92.5
R3362 vdd3p3.n730 vdd3p3.n729 92.5
R3363 vdd3p3.n731 vdd3p3.n730 92.5
R3364 vdd3p3.n175 vdd3p3.n174 92.5
R3365 vdd3p3.n732 vdd3p3.n175 92.5
R3366 vdd3p3.n735 vdd3p3.n734 92.5
R3367 vdd3p3.n734 vdd3p3.n733 92.5
R3368 vdd3p3.n736 vdd3p3.n173 92.5
R3369 vdd3p3.n173 vdd3p3.n172 92.5
R3370 vdd3p3.n738 vdd3p3.n737 92.5
R3371 vdd3p3.n739 vdd3p3.n738 92.5
R3372 vdd3p3.n171 vdd3p3.n170 92.5
R3373 vdd3p3.n740 vdd3p3.n171 92.5
R3374 vdd3p3.n743 vdd3p3.n742 92.5
R3375 vdd3p3.n742 vdd3p3.n741 92.5
R3376 vdd3p3.n744 vdd3p3.n168 92.5
R3377 vdd3p3.n168 vdd3p3.n165 92.5
R3378 vdd3p3.n688 vdd3p3.n197 92.5
R3379 vdd3p3.n197 vdd3p3.n196 92.5
R3380 vdd3p3.n160 vdd3p3.n159 92.5
R3381 vdd3p3.n756 vdd3p3.n160 92.5
R3382 vdd3p3.n759 vdd3p3.n758 92.5
R3383 vdd3p3.n758 vdd3p3.n757 92.5
R3384 vdd3p3.n760 vdd3p3.n158 92.5
R3385 vdd3p3.n158 vdd3p3.n157 92.5
R3386 vdd3p3.n762 vdd3p3.n761 92.5
R3387 vdd3p3.n763 vdd3p3.n762 92.5
R3388 vdd3p3.n156 vdd3p3.n155 92.5
R3389 vdd3p3.n764 vdd3p3.n156 92.5
R3390 vdd3p3.n767 vdd3p3.n766 92.5
R3391 vdd3p3.n766 vdd3p3.n765 92.5
R3392 vdd3p3.n768 vdd3p3.n154 92.5
R3393 vdd3p3.n154 vdd3p3.n153 92.5
R3394 vdd3p3.n770 vdd3p3.n769 92.5
R3395 vdd3p3.n771 vdd3p3.n770 92.5
R3396 vdd3p3.n151 vdd3p3.n150 92.5
R3397 vdd3p3.n772 vdd3p3.n151 92.5
R3398 vdd3p3.n775 vdd3p3.n774 92.5
R3399 vdd3p3.n774 vdd3p3.n773 92.5
R3400 vdd3p3.n776 vdd3p3.n149 92.5
R3401 vdd3p3.n152 vdd3p3.n149 92.5
R3402 vdd3p3.n752 vdd3p3.n162 92.5
R3403 vdd3p3.n162 vdd3p3.n161 92.5
R3404 vdd3p3.n751 vdd3p3.n750 92.5
R3405 vdd3p3.n750 vdd3p3.n749 92.5
R3406 vdd3p3.n164 vdd3p3.n163 92.5
R3407 vdd3p3.n169 vdd3p3.n167 92.5
R3408 vdd3p3.n746 vdd3p3.n745 92.5
R3409 vdd3p3.n747 vdd3p3.n746 92.5
R3410 vdd3p3.n754 vdd3p3.n753 92.5
R3411 vdd3p3.n755 vdd3p3.n754 92.5
R3412 vdd3p3.n779 vdd3p3.n778 92.5
R3413 vdd3p3.n800 vdd3p3.n133 92.5
R3414 vdd3p3.n799 vdd3p3.n798 92.5
R3415 vdd3p3.n142 vdd3p3.n138 92.5
R3416 vdd3p3.n793 vdd3p3.n792 92.5
R3417 vdd3p3.n790 vdd3p3.n789 92.5
R3418 vdd3p3.n144 vdd3p3.n143 92.5
R3419 vdd3p3.n783 vdd3p3.n782 92.5
R3420 vdd3p3.n781 vdd3p3.n147 92.5
R3421 vdd3p3.n803 vdd3p3.n802 92.5
R3422 vdd3p3.n318 vdd3p3.n132 92.5
R3423 vdd3p3.n321 vdd3p3.n320 92.5
R3424 vdd3p3.n343 vdd3p3.n342 92.5
R3425 vdd3p3.n341 vdd3p3.n340 92.5
R3426 vdd3p3.n311 vdd3p3.n306 92.5
R3427 vdd3p3.n334 vdd3p3.n333 92.5
R3428 vdd3p3.n331 vdd3p3.n330 92.5
R3429 vdd3p3.n313 vdd3p3.n312 92.5
R3430 vdd3p3.n329 vdd3p3.n328 92.5
R3431 vdd3p3.n314 vdd3p3.n310 92.5
R3432 vdd3p3.n336 vdd3p3.n335 92.5
R3433 vdd3p3.n339 vdd3p3.n338 92.5
R3434 vdd3p3.n307 vdd3p3.n304 92.5
R3435 vdd3p3.n347 vdd3p3.n301 92.5
R3436 vdd3p3.n345 vdd3p3.n344 92.5
R3437 vdd3p3.n327 vdd3p3.n326 92.5
R3438 vdd3p3.n327 vdd3p3.n104 92.5
R3439 vdd3p3.n325 vdd3p3.n324 92.5
R3440 vdd3p3.n323 vdd3p3.n316 92.5
R3441 vdd3p3.n386 vdd3p3.n385 92.5
R3442 vdd3p3.n383 vdd3p3.n283 92.5
R3443 vdd3p3.n382 vdd3p3.n381 92.5
R3444 vdd3p3.n380 vdd3p3.n284 92.5
R3445 vdd3p3.n378 vdd3p3.n377 92.5
R3446 vdd3p3.n376 vdd3p3.n287 92.5
R3447 vdd3p3.n290 vdd3p3.n287 92.5
R3448 vdd3p3.n375 vdd3p3.n374 92.5
R3449 vdd3p3.n374 vdd3p3.n373 92.5
R3450 vdd3p3.n289 vdd3p3.n288 92.5
R3451 vdd3p3.n372 vdd3p3.n289 92.5
R3452 vdd3p3.n370 vdd3p3.n369 92.5
R3453 vdd3p3.n371 vdd3p3.n370 92.5
R3454 vdd3p3.n368 vdd3p3.n292 92.5
R3455 vdd3p3.n292 vdd3p3.n291 92.5
R3456 vdd3p3.n367 vdd3p3.n366 92.5
R3457 vdd3p3.n366 vdd3p3.n365 92.5
R3458 vdd3p3.n294 vdd3p3.n293 92.5
R3459 vdd3p3.n364 vdd3p3.n294 92.5
R3460 vdd3p3.n362 vdd3p3.n361 92.5
R3461 vdd3p3.n363 vdd3p3.n362 92.5
R3462 vdd3p3.n360 vdd3p3.n296 92.5
R3463 vdd3p3.n296 vdd3p3.n295 92.5
R3464 vdd3p3.n359 vdd3p3.n358 92.5
R3465 vdd3p3.n358 vdd3p3.n357 92.5
R3466 vdd3p3.n298 vdd3p3.n297 92.5
R3467 vdd3p3.n356 vdd3p3.n298 92.5
R3468 vdd3p3.n354 vdd3p3.n353 92.5
R3469 vdd3p3.n355 vdd3p3.n354 92.5
R3470 vdd3p3.n352 vdd3p3.n300 92.5
R3471 vdd3p3.n300 vdd3p3.n299 92.5
R3472 vdd3p3.n351 vdd3p3.n350 92.5
R3473 vdd3p3.n350 vdd3p3.n349 92.5
R3474 vdd3p3.n438 vdd3p3.n437 92.5
R3475 vdd3p3.n437 vdd3p3.n436 92.5
R3476 vdd3p3.n257 vdd3p3.n256 92.5
R3477 vdd3p3.n435 vdd3p3.n257 92.5
R3478 vdd3p3.n433 vdd3p3.n432 92.5
R3479 vdd3p3.n434 vdd3p3.n433 92.5
R3480 vdd3p3.n431 vdd3p3.n259 92.5
R3481 vdd3p3.n259 vdd3p3.n258 92.5
R3482 vdd3p3.n430 vdd3p3.n429 92.5
R3483 vdd3p3.n429 vdd3p3.n428 92.5
R3484 vdd3p3.n261 vdd3p3.n260 92.5
R3485 vdd3p3.n427 vdd3p3.n261 92.5
R3486 vdd3p3.n425 vdd3p3.n424 92.5
R3487 vdd3p3.n426 vdd3p3.n425 92.5
R3488 vdd3p3.n423 vdd3p3.n263 92.5
R3489 vdd3p3.n263 vdd3p3.n262 92.5
R3490 vdd3p3.n422 vdd3p3.n421 92.5
R3491 vdd3p3.n421 vdd3p3.n420 92.5
R3492 vdd3p3.n265 vdd3p3.n264 92.5
R3493 vdd3p3.n419 vdd3p3.n265 92.5
R3494 vdd3p3.n417 vdd3p3.n416 92.5
R3495 vdd3p3.n418 vdd3p3.n417 92.5
R3496 vdd3p3.n415 vdd3p3.n267 92.5
R3497 vdd3p3.n267 vdd3p3.n266 92.5
R3498 vdd3p3.n414 vdd3p3.n413 92.5
R3499 vdd3p3.n413 vdd3p3.n412 92.5
R3500 vdd3p3.n269 vdd3p3.n268 92.5
R3501 vdd3p3.n411 vdd3p3.n269 92.5
R3502 vdd3p3.n409 vdd3p3.n408 92.5
R3503 vdd3p3.n410 vdd3p3.n409 92.5
R3504 vdd3p3.n407 vdd3p3.n271 92.5
R3505 vdd3p3.n271 vdd3p3.n270 92.5
R3506 vdd3p3.n406 vdd3p3.n405 92.5
R3507 vdd3p3.n405 vdd3p3.n404 92.5
R3508 vdd3p3.n273 vdd3p3.n272 92.5
R3509 vdd3p3.n403 vdd3p3.n273 92.5
R3510 vdd3p3.n401 vdd3p3.n400 92.5
R3511 vdd3p3.n402 vdd3p3.n401 92.5
R3512 vdd3p3.n399 vdd3p3.n275 92.5
R3513 vdd3p3.n275 vdd3p3.n274 92.5
R3514 vdd3p3.n398 vdd3p3.n397 92.5
R3515 vdd3p3.n397 vdd3p3.n396 92.5
R3516 vdd3p3.n277 vdd3p3.n276 92.5
R3517 vdd3p3.n395 vdd3p3.n277 92.5
R3518 vdd3p3.n393 vdd3p3.n392 92.5
R3519 vdd3p3.n394 vdd3p3.n393 92.5
R3520 vdd3p3.n391 vdd3p3.n279 92.5
R3521 vdd3p3.n279 vdd3p3.n278 92.5
R3522 vdd3p3.n390 vdd3p3.n389 92.5
R3523 vdd3p3.n389 vdd3p3.n388 92.5
R3524 vdd3p3.n281 vdd3p3.n280 92.5
R3525 vdd3p3.n387 vdd3p3.n281 92.5
R3526 vdd3p3.n446 vdd3p3.n254 92.5
R3527 vdd3p3.n450 vdd3p3.n449 92.5
R3528 vdd3p3.n255 vdd3p3.n253 92.5
R3529 vdd3p3.n480 vdd3p3.n237 92.5
R3530 vdd3p3.n476 vdd3p3.n237 92.5
R3531 vdd3p3.n479 vdd3p3.n478 92.5
R3532 vdd3p3.n478 vdd3p3.n477 92.5
R3533 vdd3p3.n239 vdd3p3.n238 92.5
R3534 vdd3p3.n475 vdd3p3.n239 92.5
R3535 vdd3p3.n473 vdd3p3.n472 92.5
R3536 vdd3p3.n474 vdd3p3.n473 92.5
R3537 vdd3p3.n471 vdd3p3.n241 92.5
R3538 vdd3p3.n241 vdd3p3.n240 92.5
R3539 vdd3p3.n470 vdd3p3.n469 92.5
R3540 vdd3p3.n469 vdd3p3.n468 92.5
R3541 vdd3p3.n243 vdd3p3.n242 92.5
R3542 vdd3p3.n467 vdd3p3.n243 92.5
R3543 vdd3p3.n465 vdd3p3.n464 92.5
R3544 vdd3p3.n466 vdd3p3.n465 92.5
R3545 vdd3p3.n463 vdd3p3.n245 92.5
R3546 vdd3p3.n245 vdd3p3.n244 92.5
R3547 vdd3p3.n462 vdd3p3.n461 92.5
R3548 vdd3p3.n461 vdd3p3.n460 92.5
R3549 vdd3p3.n247 vdd3p3.n246 92.5
R3550 vdd3p3.n459 vdd3p3.n247 92.5
R3551 vdd3p3.n457 vdd3p3.n456 92.5
R3552 vdd3p3.n458 vdd3p3.n457 92.5
R3553 vdd3p3.n455 vdd3p3.n249 92.5
R3554 vdd3p3.n249 vdd3p3.n248 92.5
R3555 vdd3p3.n454 vdd3p3.n453 92.5
R3556 vdd3p3.n453 vdd3p3.n452 92.5
R3557 vdd3p3.n251 vdd3p3.n250 92.5
R3558 vdd3p3.n442 vdd3p3.n439 92.5
R3559 vdd3p3.n445 vdd3p3.n444 92.5
R3560 vdd3p3.n654 vdd3p3.n653 92.5
R3561 vdd3p3.n578 vdd3p3.n217 92.5
R3562 vdd3p3.n580 vdd3p3.n579 92.5
R3563 vdd3p3.n577 vdd3p3.n576 92.5
R3564 vdd3p3.n547 vdd3p3.n546 92.5
R3565 vdd3p3.n571 vdd3p3.n570 92.5
R3566 vdd3p3.n549 vdd3p3.n548 92.5
R3567 vdd3p3.n565 vdd3p3.n564 92.5
R3568 vdd3p3.n561 vdd3p3.n560 92.5
R3569 vdd3p3.n559 vdd3p3.n558 92.5
R3570 vdd3p3.n629 vdd3p3.n628 92.5
R3571 vdd3p3.n633 vdd3p3.n632 92.5
R3572 vdd3p3.n636 vdd3p3.n635 92.5
R3573 vdd3p3.n494 vdd3p3.n493 92.5
R3574 vdd3p3.n483 vdd3p3.n482 92.5
R3575 vdd3p3.n645 vdd3p3.n644 92.5
R3576 vdd3p3.n646 vdd3p3.n236 92.5
R3577 vdd3p3.n649 vdd3p3.n648 92.5
R3578 vdd3p3.n643 vdd3p3.n642 92.5
R3579 vdd3p3.n492 vdd3p3.n485 92.5
R3580 vdd3p3.n638 vdd3p3.n637 92.5
R3581 vdd3p3.n634 vdd3p3.n491 92.5
R3582 vdd3p3.n631 vdd3p3.n630 92.5
R3583 vdd3p3.n495 vdd3p3.n229 92.5
R3584 vdd3p3.n651 vdd3p3.n229 92.5
R3585 vdd3p3.n627 vdd3p3.n626 92.5
R3586 vdd3p3.n553 vdd3p3.n552 92.5
R3587 vdd3p3.n555 vdd3p3.n554 92.5
R3588 vdd3p3.n557 vdd3p3.n556 92.5
R3589 vdd3p3.n563 vdd3p3.n562 92.5
R3590 vdd3p3.n582 vdd3p3.n581 92.5
R3591 vdd3p3.n575 vdd3p3.n574 92.5
R3592 vdd3p3.n573 vdd3p3.n572 92.5
R3593 vdd3p3.n569 vdd3p3.n568 92.5
R3594 vdd3p3.n567 vdd3p3.n566 92.5
R3595 vdd3p3.n128 vdd3p3.n102 92.5
R3596 vdd3p3.n807 vdd3p3.n806 92.5
R3597 vdd3p3.n805 vdd3p3.n804 92.5
R3598 vdd3p3.n805 vdd3p3.n129 92.5
R3599 vdd3p3.n797 vdd3p3.n796 92.5
R3600 vdd3p3.n795 vdd3p3.n794 92.5
R3601 vdd3p3.n145 vdd3p3.n141 92.5
R3602 vdd3p3.n788 vdd3p3.n787 92.5
R3603 vdd3p3.n785 vdd3p3.n784 92.5
R3604 vdd3p3.n137 vdd3p3.n131 92.5
R3605 vdd3p3.n122 vdd3p3.n121 92.5
R3606 vdd3p3.n119 vdd3p3.n107 92.5
R3607 vdd3p3.n117 vdd3p3.n116 92.5
R3608 vdd3p3.n115 vdd3p3.n114 92.5
R3609 vdd3p3.n112 vdd3p3.n109 92.5
R3610 vdd3p3.n110 vdd3p3.n99 92.5
R3611 vdd3p3.n127 vdd3p3.n126 92.5
R3612 vdd3p3.n129 vdd3p3.n127 92.5
R3613 vdd3p3.n809 vdd3p3.n808 92.5
R3614 vdd3p3.n808 vdd3p3.n807 92.5
R3615 vdd3p3.n810 vdd3p3.n106 92.5
R3616 vdd3p3.n128 vdd3p3.n106 92.5
R3617 vdd3p3.n812 vdd3p3.n811 92.5
R3618 vdd3p3.n813 vdd3p3.n812 92.5
R3619 vdd3p3.n124 vdd3p3.n123 92.5
R3620 vdd3p3.n123 vdd3p3.n85 92.5
R3621 vdd3p3.n79 vdd3p3.n78 92.5
R3622 vdd3p3.n827 vdd3p3.n79 92.5
R3623 vdd3p3.n832 vdd3p3.n831 92.5
R3624 vdd3p3.n831 vdd3p3.n830 92.5
R3625 vdd3p3.n833 vdd3p3.n76 92.5
R3626 vdd3p3.n80 vdd3p3.n76 92.5
R3627 vdd3p3.n835 vdd3p3.n834 92.5
R3628 vdd3p3.n836 vdd3p3.n835 92.5
R3629 vdd3p3.n77 vdd3p3.n75 92.5
R3630 vdd3p3.n536 vdd3p3.n75 92.5
R3631 vdd3p3.n589 vdd3p3.n588 92.5
R3632 vdd3p3.n588 vdd3p3.n505 92.5
R3633 vdd3p3.n587 vdd3p3.n586 92.5
R3634 vdd3p3.n587 vdd3p3.n504 92.5
R3635 vdd3p3.n585 vdd3p3.n499 92.5
R3636 vdd3p3.n623 vdd3p3.n499 92.5
R3637 vdd3p3.n584 vdd3p3.n583 92.5
R3638 vdd3p3.n583 vdd3p3.n486 92.5
R3639 vdd3p3.n592 vdd3p3.n591 92.5
R3640 vdd3p3.n594 vdd3p3.n544 92.5
R3641 vdd3p3.n597 vdd3p3.n596 92.5
R3642 vdd3p3.n599 vdd3p3.n598 92.5
R3643 vdd3p3.n601 vdd3p3.n540 92.5
R3644 vdd3p3.n604 vdd3p3.n603 92.5
R3645 vdd3p3.n550 vdd3p3.n500 92.5
R3646 vdd3p3.n500 vdd3p3.n486 92.5
R3647 vdd3p3.n622 vdd3p3.n621 92.5
R3648 vdd3p3.n623 vdd3p3.n622 92.5
R3649 vdd3p3.n619 vdd3p3.n501 92.5
R3650 vdd3p3.n504 vdd3p3.n501 92.5
R3651 vdd3p3.n541 vdd3p3.n502 92.5
R3652 vdd3p3.n541 vdd3p3.n505 92.5
R3653 vdd3p3.n605 vdd3p3.n72 92.5
R3654 vdd3p3.n536 vdd3p3.n72 92.5
R3655 vdd3p3.n838 vdd3p3.n837 92.5
R3656 vdd3p3.n837 vdd3p3.n836 92.5
R3657 vdd3p3.n73 vdd3p3.n71 92.5
R3658 vdd3p3.n80 vdd3p3.n73 92.5
R3659 vdd3p3.n829 vdd3p3.n66 92.5
R3660 vdd3p3.n830 vdd3p3.n829 92.5
R3661 vdd3p3.n828 vdd3p3.n84 92.5
R3662 vdd3p3.n828 vdd3p3.n827 92.5
R3663 vdd3p3.n97 vdd3p3.n83 92.5
R3664 vdd3p3.n85 vdd3p3.n83 92.5
R3665 vdd3p3.n815 vdd3p3.n814 92.5
R3666 vdd3p3.n814 vdd3p3.n813 92.5
R3667 vdd3p3.n620 vdd3p3.n496 92.5
R3668 vdd3p3.n498 vdd3p3.n496 92.5
R3669 vdd3p3.n618 vdd3p3.n617 92.5
R3670 vdd3p3.n617 vdd3p3.n616 92.5
R3671 vdd3p3.n539 vdd3p3.n503 92.5
R3672 vdd3p3.n511 vdd3p3.n503 92.5
R3673 vdd3p3.n609 vdd3p3.n608 92.5
R3674 vdd3p3.n610 vdd3p3.n609 92.5
R3675 vdd3p3.n606 vdd3p3.n538 92.5
R3676 vdd3p3.n538 vdd3p3.n537 92.5
R3677 vdd3p3.n534 vdd3p3.n67 92.5
R3678 vdd3p3.n534 vdd3p3.n81 92.5
R3679 vdd3p3.n533 vdd3p3.n532 92.5
R3680 vdd3p3.n533 vdd3p3.n82 92.5
R3681 vdd3p3.n96 vdd3p3.n86 92.5
R3682 vdd3p3.n826 vdd3p3.n86 92.5
R3683 vdd3p3.n98 vdd3p3.n94 92.5
R3684 vdd3p3.n94 vdd3p3.n93 92.5
R3685 vdd3p3.n819 vdd3p3.n818 92.5
R3686 vdd3p3.n820 vdd3p3.n819 92.5
R3687 vdd3p3.n816 vdd3p3.n95 92.5
R3688 vdd3p3.n103 vdd3p3.n95 92.5
R3689 vdd3p3.n625 vdd3p3.n497 92.5
R3690 vdd3p3.n625 vdd3p3.n624 92.5
R3691 vdd3p3.n8704 vdd3p3.n8703 92.5
R3692 vdd3p3.n8702 vdd3p3.n8701 92.5
R3693 vdd3p3.n6390 vdd3p3.n6389 92.5
R3694 vdd3p3.n5340 vdd3p3.n5339 92.5
R3695 vdd3p3.n6713 vdd3p3.n6712 92.5
R3696 vdd3p3.n6709 vdd3p3.n6708 92.5
R3697 vdd3p3.n6705 vdd3p3.n6704 92.5
R3698 vdd3p3.n6701 vdd3p3.n6700 92.5
R3699 vdd3p3.n6697 vdd3p3.n6696 92.5
R3700 vdd3p3.n6693 vdd3p3.n6692 92.5
R3701 vdd3p3.n6692 vdd3p3.n6691 92.5
R3702 vdd3p3.n6688 vdd3p3.n6687 92.5
R3703 vdd3p3.n6687 vdd3p3.n6686 92.5
R3704 vdd3p3.n6680 vdd3p3.n6679 92.5
R3705 vdd3p3.n6679 vdd3p3.n6678 92.5
R3706 vdd3p3.n6683 vdd3p3.n6682 92.5
R3707 vdd3p3.n6682 vdd3p3.n6681 92.5
R3708 vdd3p3.n6675 vdd3p3.n6674 92.5
R3709 vdd3p3.n6674 vdd3p3.n6673 92.5
R3710 vdd3p3.n6670 vdd3p3.n6669 92.5
R3711 vdd3p3.n6669 vdd3p3.n6668 92.5
R3712 vdd3p3.n6665 vdd3p3.n6664 92.5
R3713 vdd3p3.n6664 vdd3p3.n6663 92.5
R3714 vdd3p3.n6660 vdd3p3.n6659 92.5
R3715 vdd3p3.n6659 vdd3p3.n6658 92.5
R3716 vdd3p3.n6655 vdd3p3.n6654 92.5
R3717 vdd3p3.n6654 vdd3p3.n6653 92.5
R3718 vdd3p3.n6650 vdd3p3.n6649 92.5
R3719 vdd3p3.n6649 vdd3p3.n6648 92.5
R3720 vdd3p3.n6645 vdd3p3.n6644 92.5
R3721 vdd3p3.n6644 vdd3p3.n6643 92.5
R3722 vdd3p3.n6640 vdd3p3.n6639 92.5
R3723 vdd3p3.n6639 vdd3p3.n6638 92.5
R3724 vdd3p3.n6635 vdd3p3.n6634 92.5
R3725 vdd3p3.n6634 vdd3p3.n6633 92.5
R3726 vdd3p3.n6630 vdd3p3.n6629 92.5
R3727 vdd3p3.n6629 vdd3p3.n6628 92.5
R3728 vdd3p3.n6625 vdd3p3.n6624 92.5
R3729 vdd3p3.n6624 vdd3p3.n6623 92.5
R3730 vdd3p3.n6620 vdd3p3.n6619 92.5
R3731 vdd3p3.n6619 vdd3p3.n6618 92.5
R3732 vdd3p3.n6615 vdd3p3.n6614 92.5
R3733 vdd3p3.n6614 vdd3p3.n6613 92.5
R3734 vdd3p3.n6610 vdd3p3.n6609 92.5
R3735 vdd3p3.n6609 vdd3p3.n6608 92.5
R3736 vdd3p3.n6605 vdd3p3.n6604 92.5
R3737 vdd3p3.n6604 vdd3p3.n6603 92.5
R3738 vdd3p3.n6600 vdd3p3.n6599 92.5
R3739 vdd3p3.n6599 vdd3p3.n6598 92.5
R3740 vdd3p3.n6592 vdd3p3.n6591 92.5
R3741 vdd3p3.n6591 vdd3p3.n6590 92.5
R3742 vdd3p3.n6595 vdd3p3.n6594 92.5
R3743 vdd3p3.n6594 vdd3p3.n6593 92.5
R3744 vdd3p3.n6587 vdd3p3.n6586 92.5
R3745 vdd3p3.n6583 vdd3p3.n6582 92.5
R3746 vdd3p3.n6579 vdd3p3.n6578 92.5
R3747 vdd3p3.n6575 vdd3p3.n6574 92.5
R3748 vdd3p3.n6571 vdd3p3.n6570 92.5
R3749 vdd3p3.n6567 vdd3p3.n6566 92.5
R3750 vdd3p3.n6563 vdd3p3.n6562 92.5
R3751 vdd3p3.n6546 vdd3p3.n6545 92.5
R3752 vdd3p3.n6542 vdd3p3.n6541 92.5
R3753 vdd3p3.n6538 vdd3p3.n6537 92.5
R3754 vdd3p3.n6534 vdd3p3.n6533 92.5
R3755 vdd3p3.n6530 vdd3p3.n6529 92.5
R3756 vdd3p3.n6526 vdd3p3.n6525 92.5
R3757 vdd3p3.n6522 vdd3p3.n6521 92.5
R3758 vdd3p3.n6521 vdd3p3.n6520 92.5
R3759 vdd3p3.n6517 vdd3p3.n6516 92.5
R3760 vdd3p3.n6516 vdd3p3.n6515 92.5
R3761 vdd3p3.n6512 vdd3p3.n6511 92.5
R3762 vdd3p3.n6511 vdd3p3.n6510 92.5
R3763 vdd3p3.n6504 vdd3p3.n6503 92.5
R3764 vdd3p3.n6503 vdd3p3.n6502 92.5
R3765 vdd3p3.n6507 vdd3p3.n6506 92.5
R3766 vdd3p3.n6506 vdd3p3.n6505 92.5
R3767 vdd3p3.n6499 vdd3p3.n6498 92.5
R3768 vdd3p3.n6498 vdd3p3.n6497 92.5
R3769 vdd3p3.n6494 vdd3p3.n6493 92.5
R3770 vdd3p3.n6493 vdd3p3.n6492 92.5
R3771 vdd3p3.n6489 vdd3p3.n6488 92.5
R3772 vdd3p3.n6488 vdd3p3.n6487 92.5
R3773 vdd3p3.n6484 vdd3p3.n6483 92.5
R3774 vdd3p3.n6483 vdd3p3.n6482 92.5
R3775 vdd3p3.n6479 vdd3p3.n6478 92.5
R3776 vdd3p3.n6478 vdd3p3.n6477 92.5
R3777 vdd3p3.n6474 vdd3p3.n6473 92.5
R3778 vdd3p3.n6473 vdd3p3.n6472 92.5
R3779 vdd3p3.n6469 vdd3p3.n6468 92.5
R3780 vdd3p3.n6468 vdd3p3.n6467 92.5
R3781 vdd3p3.n6464 vdd3p3.n6463 92.5
R3782 vdd3p3.n6463 vdd3p3.n6462 92.5
R3783 vdd3p3.n6459 vdd3p3.n6458 92.5
R3784 vdd3p3.n6458 vdd3p3.n6457 92.5
R3785 vdd3p3.n6454 vdd3p3.n6453 92.5
R3786 vdd3p3.n6453 vdd3p3.n6452 92.5
R3787 vdd3p3.n6449 vdd3p3.n6448 92.5
R3788 vdd3p3.n6448 vdd3p3.n6447 92.5
R3789 vdd3p3.n6444 vdd3p3.n6443 92.5
R3790 vdd3p3.n6443 vdd3p3.n6442 92.5
R3791 vdd3p3.n6439 vdd3p3.n6438 92.5
R3792 vdd3p3.n6438 vdd3p3.n6437 92.5
R3793 vdd3p3.n6434 vdd3p3.n6433 92.5
R3794 vdd3p3.n6433 vdd3p3.n6432 92.5
R3795 vdd3p3.n6429 vdd3p3.n6428 92.5
R3796 vdd3p3.n6428 vdd3p3.n6427 92.5
R3797 vdd3p3.n6424 vdd3p3.n6423 92.5
R3798 vdd3p3.n6423 vdd3p3.n6422 92.5
R3799 vdd3p3.n6417 vdd3p3.n6416 92.5
R3800 vdd3p3.n6419 vdd3p3.n6418 92.5
R3801 vdd3p3.n6413 vdd3p3.n6412 92.5
R3802 vdd3p3.n6409 vdd3p3.n6408 92.5
R3803 vdd3p3.n6405 vdd3p3.n6404 92.5
R3804 vdd3p3.n8710 vdd3p3.n8709 92.5
R3805 vdd3p3.n8713 vdd3p3.n8712 92.5
R3806 vdd3p3.n8707 vdd3p3.n8706 92.5
R3807 vdd3p3.n7498 vdd3p3.n7497 92.5
R3808 vdd3p3.n7500 vdd3p3.n7499 92.5
R3809 vdd3p3.n7502 vdd3p3.n7501 92.5
R3810 vdd3p3.n7504 vdd3p3.n7503 92.5
R3811 vdd3p3.n7506 vdd3p3.n7505 92.5
R3812 vdd3p3.n7509 vdd3p3.n7508 92.5
R3813 vdd3p3.n8459 vdd3p3.n8446 92.5
R3814 vdd3p3.n7955 vdd3p3.n7954 92.5
R3815 vdd3p3.n7961 vdd3p3.n7960 92.5
R3816 vdd3p3.n7968 vdd3p3.n7967 92.5
R3817 vdd3p3.n7975 vdd3p3.n7974 92.5
R3818 vdd3p3.n7977 vdd3p3.n7976 92.5
R3819 vdd3p3.n7984 vdd3p3.n7983 92.5
R3820 vdd3p3.n7991 vdd3p3.n7990 92.5
R3821 vdd3p3.n7998 vdd3p3.n7997 92.5
R3822 vdd3p3.n8005 vdd3p3.n8004 92.5
R3823 vdd3p3.n8012 vdd3p3.n8011 92.5
R3824 vdd3p3.n8019 vdd3p3.n8018 92.5
R3825 vdd3p3.n8031 vdd3p3.n8030 92.5
R3826 vdd3p3.n7947 vdd3p3.n7946 92.5
R3827 vdd3p3.n7952 vdd3p3.n7951 92.5
R3828 vdd3p3.n7959 vdd3p3.n7958 92.5
R3829 vdd3p3.n7963 vdd3p3.n7962 92.5
R3830 vdd3p3.n7971 vdd3p3.n7970 92.5
R3831 vdd3p3.n7979 vdd3p3.n7978 92.5
R3832 vdd3p3.n7987 vdd3p3.n7986 92.5
R3833 vdd3p3.n7993 vdd3p3.n7992 92.5
R3834 vdd3p3.n8001 vdd3p3.n8000 92.5
R3835 vdd3p3.n8007 vdd3p3.n8006 92.5
R3836 vdd3p3.n8015 vdd3p3.n8014 92.5
R3837 vdd3p3.n8022 vdd3p3.n8021 92.5
R3838 vdd3p3.n8026 vdd3p3.n8025 92.5
R3839 vdd3p3.n8035 vdd3p3.n8034 92.5
R3840 vdd3p3.n7944 vdd3p3.n7943 92.5
R3841 vdd3p3.n7927 vdd3p3.n7926 92.5
R3842 vdd3p3.n7926 vdd3p3.n7925 92.5
R3843 vdd3p3.n7919 vdd3p3.n7918 92.5
R3844 vdd3p3.n7918 vdd3p3.n7917 92.5
R3845 vdd3p3.n7911 vdd3p3.n7910 92.5
R3846 vdd3p3.n7910 vdd3p3.n7909 92.5
R3847 vdd3p3.n7903 vdd3p3.n7902 92.5
R3848 vdd3p3.n7902 vdd3p3.n7901 92.5
R3849 vdd3p3.n7895 vdd3p3.n7894 92.5
R3850 vdd3p3.n7894 vdd3p3.n7893 92.5
R3851 vdd3p3.n7887 vdd3p3.n7886 92.5
R3852 vdd3p3.n7886 vdd3p3.n7885 92.5
R3853 vdd3p3.n7879 vdd3p3.n7878 92.5
R3854 vdd3p3.n7878 vdd3p3.n7877 92.5
R3855 vdd3p3.n7871 vdd3p3.n7870 92.5
R3856 vdd3p3.n7870 vdd3p3.n7869 92.5
R3857 vdd3p3.n7860 vdd3p3.n7859 92.5
R3858 vdd3p3.n7859 vdd3p3.n7858 92.5
R3859 vdd3p3.n7866 vdd3p3.n7865 92.5
R3860 vdd3p3.n7865 vdd3p3.n7864 92.5
R3861 vdd3p3.n7855 vdd3p3.n7854 92.5
R3862 vdd3p3.n7854 vdd3p3.n7853 92.5
R3863 vdd3p3.n7847 vdd3p3.n7846 92.5
R3864 vdd3p3.n7846 vdd3p3.n7845 92.5
R3865 vdd3p3.n7836 vdd3p3.n7835 92.5
R3866 vdd3p3.n7835 vdd3p3.n7834 92.5
R3867 vdd3p3.n7828 vdd3p3.n7827 92.5
R3868 vdd3p3.n7827 vdd3p3.n7826 92.5
R3869 vdd3p3.n7820 vdd3p3.n7819 92.5
R3870 vdd3p3.n7819 vdd3p3.n7818 92.5
R3871 vdd3p3.n7812 vdd3p3.n7811 92.5
R3872 vdd3p3.n7811 vdd3p3.n7810 92.5
R3873 vdd3p3.n7804 vdd3p3.n7803 92.5
R3874 vdd3p3.n7803 vdd3p3.n7802 92.5
R3875 vdd3p3.n7796 vdd3p3.n7795 92.5
R3876 vdd3p3.n7795 vdd3p3.n7794 92.5
R3877 vdd3p3.n7785 vdd3p3.n7784 92.5
R3878 vdd3p3.n7784 vdd3p3.n7783 92.5
R3879 vdd3p3.n7777 vdd3p3.n7776 92.5
R3880 vdd3p3.n7776 vdd3p3.n7775 92.5
R3881 vdd3p3.n7769 vdd3p3.n7768 92.5
R3882 vdd3p3.n7768 vdd3p3.n7767 92.5
R3883 vdd3p3.n7761 vdd3p3.n7760 92.5
R3884 vdd3p3.n7760 vdd3p3.n7759 92.5
R3885 vdd3p3.n7753 vdd3p3.n7752 92.5
R3886 vdd3p3.n7752 vdd3p3.n7751 92.5
R3887 vdd3p3.n7745 vdd3p3.n7744 92.5
R3888 vdd3p3.n7744 vdd3p3.n7743 92.5
R3889 vdd3p3.n7737 vdd3p3.n7736 92.5
R3890 vdd3p3.n7736 vdd3p3.n7735 92.5
R3891 vdd3p3.n7729 vdd3p3.n7728 92.5
R3892 vdd3p3.n7728 vdd3p3.n7727 92.5
R3893 vdd3p3.n7719 vdd3p3.n7718 92.5
R3894 vdd3p3.n7718 vdd3p3.n7717 92.5
R3895 vdd3p3.n7724 vdd3p3.n7723 92.5
R3896 vdd3p3.n7714 vdd3p3.n7713 92.5
R3897 vdd3p3.n7708 vdd3p3.n7707 92.5
R3898 vdd3p3.n7700 vdd3p3.n7699 92.5
R3899 vdd3p3.n7694 vdd3p3.n7693 92.5
R3900 vdd3p3.n7688 vdd3p3.n7687 92.5
R3901 vdd3p3.n7687 vdd3p3.n7686 92.5
R3902 vdd3p3.n7680 vdd3p3.n7679 92.5
R3903 vdd3p3.n7679 vdd3p3.n7678 92.5
R3904 vdd3p3.n7672 vdd3p3.n7671 92.5
R3905 vdd3p3.n7671 vdd3p3.n7670 92.5
R3906 vdd3p3.n7664 vdd3p3.n7663 92.5
R3907 vdd3p3.n7663 vdd3p3.n7662 92.5
R3908 vdd3p3.n7653 vdd3p3.n7652 92.5
R3909 vdd3p3.n7652 vdd3p3.n7651 92.5
R3910 vdd3p3.n7645 vdd3p3.n7644 92.5
R3911 vdd3p3.n7644 vdd3p3.n7643 92.5
R3912 vdd3p3.n7637 vdd3p3.n7636 92.5
R3913 vdd3p3.n7636 vdd3p3.n7635 92.5
R3914 vdd3p3.n7629 vdd3p3.n7628 92.5
R3915 vdd3p3.n7628 vdd3p3.n7627 92.5
R3916 vdd3p3.n7621 vdd3p3.n7620 92.5
R3917 vdd3p3.n7620 vdd3p3.n7619 92.5
R3918 vdd3p3.n7613 vdd3p3.n7612 92.5
R3919 vdd3p3.n7612 vdd3p3.n7611 92.5
R3920 vdd3p3.n7605 vdd3p3.n7604 92.5
R3921 vdd3p3.n7604 vdd3p3.n7603 92.5
R3922 vdd3p3.n7597 vdd3p3.n7596 92.5
R3923 vdd3p3.n7596 vdd3p3.n7595 92.5
R3924 vdd3p3.n7586 vdd3p3.n7585 92.5
R3925 vdd3p3.n7585 vdd3p3.n7584 92.5
R3926 vdd3p3.n7592 vdd3p3.n7591 92.5
R3927 vdd3p3.n7591 vdd3p3.n7590 92.5
R3928 vdd3p3.n7581 vdd3p3.n7580 92.5
R3929 vdd3p3.n7580 vdd3p3.n7579 92.5
R3930 vdd3p3.n7573 vdd3p3.n7572 92.5
R3931 vdd3p3.n7572 vdd3p3.n7571 92.5
R3932 vdd3p3.n7562 vdd3p3.n7561 92.5
R3933 vdd3p3.n7561 vdd3p3.n7560 92.5
R3934 vdd3p3.n7554 vdd3p3.n7553 92.5
R3935 vdd3p3.n7553 vdd3p3.n7552 92.5
R3936 vdd3p3.n7546 vdd3p3.n7545 92.5
R3937 vdd3p3.n7545 vdd3p3.n7544 92.5
R3938 vdd3p3.n7538 vdd3p3.n7537 92.5
R3939 vdd3p3.n7537 vdd3p3.n7536 92.5
R3940 vdd3p3.n7525 vdd3p3.n7524 92.5
R3941 vdd3p3.n7524 vdd3p3.n7523 92.5
R3942 vdd3p3.n7530 vdd3p3.n7529 92.5
R3943 vdd3p3.n7529 vdd3p3.n7528 92.5
R3944 vdd3p3.n7535 vdd3p3.n7534 92.5
R3945 vdd3p3.n7534 vdd3p3.n7533 92.5
R3946 vdd3p3.n7543 vdd3p3.n7542 92.5
R3947 vdd3p3.n7542 vdd3p3.n7541 92.5
R3948 vdd3p3.n7551 vdd3p3.n7550 92.5
R3949 vdd3p3.n7550 vdd3p3.n7549 92.5
R3950 vdd3p3.n7559 vdd3p3.n7558 92.5
R3951 vdd3p3.n7558 vdd3p3.n7557 92.5
R3952 vdd3p3.n7570 vdd3p3.n7569 92.5
R3953 vdd3p3.n7569 vdd3p3.n7568 92.5
R3954 vdd3p3.n7567 vdd3p3.n7566 92.5
R3955 vdd3p3.n7566 vdd3p3.n7565 92.5
R3956 vdd3p3.n7578 vdd3p3.n7577 92.5
R3957 vdd3p3.n7577 vdd3p3.n7576 92.5
R3958 vdd3p3.n7589 vdd3p3.n7588 92.5
R3959 vdd3p3.n7588 vdd3p3.n7587 92.5
R3960 vdd3p3.n7600 vdd3p3.n7599 92.5
R3961 vdd3p3.n7599 vdd3p3.n7598 92.5
R3962 vdd3p3.n7608 vdd3p3.n7607 92.5
R3963 vdd3p3.n7607 vdd3p3.n7606 92.5
R3964 vdd3p3.n7616 vdd3p3.n7615 92.5
R3965 vdd3p3.n7615 vdd3p3.n7614 92.5
R3966 vdd3p3.n7624 vdd3p3.n7623 92.5
R3967 vdd3p3.n7623 vdd3p3.n7622 92.5
R3968 vdd3p3.n7632 vdd3p3.n7631 92.5
R3969 vdd3p3.n7631 vdd3p3.n7630 92.5
R3970 vdd3p3.n7640 vdd3p3.n7639 92.5
R3971 vdd3p3.n7639 vdd3p3.n7638 92.5
R3972 vdd3p3.n7648 vdd3p3.n7647 92.5
R3973 vdd3p3.n7647 vdd3p3.n7646 92.5
R3974 vdd3p3.n7656 vdd3p3.n7655 92.5
R3975 vdd3p3.n7655 vdd3p3.n7654 92.5
R3976 vdd3p3.n7661 vdd3p3.n7660 92.5
R3977 vdd3p3.n7660 vdd3p3.n7659 92.5
R3978 vdd3p3.n7669 vdd3p3.n7668 92.5
R3979 vdd3p3.n7668 vdd3p3.n7667 92.5
R3980 vdd3p3.n7677 vdd3p3.n7676 92.5
R3981 vdd3p3.n7676 vdd3p3.n7675 92.5
R3982 vdd3p3.n7685 vdd3p3.n7684 92.5
R3983 vdd3p3.n7684 vdd3p3.n7683 92.5
R3984 vdd3p3.n7692 vdd3p3.n7691 92.5
R3985 vdd3p3.n7698 vdd3p3.n7697 92.5
R3986 vdd3p3.n7706 vdd3p3.n7705 92.5
R3987 vdd3p3.n7704 vdd3p3.n7703 92.5
R3988 vdd3p3.n7712 vdd3p3.n7711 92.5
R3989 vdd3p3.n7722 vdd3p3.n7721 92.5
R3990 vdd3p3.n7721 vdd3p3.n7720 92.5
R3991 vdd3p3.n7732 vdd3p3.n7731 92.5
R3992 vdd3p3.n7731 vdd3p3.n7730 92.5
R3993 vdd3p3.n7740 vdd3p3.n7739 92.5
R3994 vdd3p3.n7739 vdd3p3.n7738 92.5
R3995 vdd3p3.n7748 vdd3p3.n7747 92.5
R3996 vdd3p3.n7747 vdd3p3.n7746 92.5
R3997 vdd3p3.n7756 vdd3p3.n7755 92.5
R3998 vdd3p3.n7755 vdd3p3.n7754 92.5
R3999 vdd3p3.n7764 vdd3p3.n7763 92.5
R4000 vdd3p3.n7763 vdd3p3.n7762 92.5
R4001 vdd3p3.n7772 vdd3p3.n7771 92.5
R4002 vdd3p3.n7771 vdd3p3.n7770 92.5
R4003 vdd3p3.n7780 vdd3p3.n7779 92.5
R4004 vdd3p3.n7779 vdd3p3.n7778 92.5
R4005 vdd3p3.n7788 vdd3p3.n7787 92.5
R4006 vdd3p3.n7787 vdd3p3.n7786 92.5
R4007 vdd3p3.n7793 vdd3p3.n7792 92.5
R4008 vdd3p3.n7792 vdd3p3.n7791 92.5
R4009 vdd3p3.n7801 vdd3p3.n7800 92.5
R4010 vdd3p3.n7800 vdd3p3.n7799 92.5
R4011 vdd3p3.n7809 vdd3p3.n7808 92.5
R4012 vdd3p3.n7808 vdd3p3.n7807 92.5
R4013 vdd3p3.n7817 vdd3p3.n7816 92.5
R4014 vdd3p3.n7816 vdd3p3.n7815 92.5
R4015 vdd3p3.n7825 vdd3p3.n7824 92.5
R4016 vdd3p3.n7824 vdd3p3.n7823 92.5
R4017 vdd3p3.n7833 vdd3p3.n7832 92.5
R4018 vdd3p3.n7832 vdd3p3.n7831 92.5
R4019 vdd3p3.n7844 vdd3p3.n7843 92.5
R4020 vdd3p3.n7843 vdd3p3.n7842 92.5
R4021 vdd3p3.n7841 vdd3p3.n7840 92.5
R4022 vdd3p3.n7840 vdd3p3.n7839 92.5
R4023 vdd3p3.n7852 vdd3p3.n7851 92.5
R4024 vdd3p3.n7851 vdd3p3.n7850 92.5
R4025 vdd3p3.n7863 vdd3p3.n7862 92.5
R4026 vdd3p3.n7862 vdd3p3.n7861 92.5
R4027 vdd3p3.n7874 vdd3p3.n7873 92.5
R4028 vdd3p3.n7873 vdd3p3.n7872 92.5
R4029 vdd3p3.n7882 vdd3p3.n7881 92.5
R4030 vdd3p3.n7881 vdd3p3.n7880 92.5
R4031 vdd3p3.n7890 vdd3p3.n7889 92.5
R4032 vdd3p3.n7889 vdd3p3.n7888 92.5
R4033 vdd3p3.n7898 vdd3p3.n7897 92.5
R4034 vdd3p3.n7897 vdd3p3.n7896 92.5
R4035 vdd3p3.n7906 vdd3p3.n7905 92.5
R4036 vdd3p3.n7905 vdd3p3.n7904 92.5
R4037 vdd3p3.n7914 vdd3p3.n7913 92.5
R4038 vdd3p3.n7913 vdd3p3.n7912 92.5
R4039 vdd3p3.n7922 vdd3p3.n7921 92.5
R4040 vdd3p3.n7921 vdd3p3.n7920 92.5
R4041 vdd3p3.n7933 vdd3p3.n7932 92.5
R4042 vdd3p3.n7932 vdd3p3.n7931 92.5
R4043 vdd3p3.n7930 vdd3p3.n7929 92.5
R4044 vdd3p3.n7929 vdd3p3.n7928 92.5
R4045 vdd3p3.n7942 vdd3p3.n7941 92.5
R4046 vdd3p3.n7470 vdd3p3.n7469 92.5
R4047 vdd3p3.n7469 vdd3p3.n7468 92.5
R4048 vdd3p3.n7458 vdd3p3.n7457 92.5
R4049 vdd3p3.n7457 vdd3p3.n7456 92.5
R4050 vdd3p3.n7475 vdd3p3.n7474 92.5
R4051 vdd3p3.n7474 vdd3p3.n7473 92.5
R4052 vdd3p3.n7480 vdd3p3.n7479 92.5
R4053 vdd3p3.n7479 vdd3p3.n7478 92.5
R4054 vdd3p3.n7485 vdd3p3.n7484 92.5
R4055 vdd3p3.n7484 vdd3p3.n7483 92.5
R4056 vdd3p3.n7490 vdd3p3.n7489 92.5
R4057 vdd3p3.n7489 vdd3p3.n7488 92.5
R4058 vdd3p3.n7391 vdd3p3.n7390 92.5
R4059 vdd3p3.n7395 vdd3p3.n7394 92.5
R4060 vdd3p3.n7400 vdd3p3.n7399 92.5
R4061 vdd3p3.n7405 vdd3p3.n7404 92.5
R4062 vdd3p3.n7410 vdd3p3.n7409 92.5
R4063 vdd3p3.n7415 vdd3p3.n7414 92.5
R4064 vdd3p3.n7420 vdd3p3.n7419 92.5
R4065 vdd3p3.n7426 vdd3p3.n7425 92.5
R4066 vdd3p3.n7431 vdd3p3.n7430 92.5
R4067 vdd3p3.n7436 vdd3p3.n7435 92.5
R4068 vdd3p3.n7441 vdd3p3.n7440 92.5
R4069 vdd3p3.n7446 vdd3p3.n7445 92.5
R4070 vdd3p3.n7453 vdd3p3.n7452 92.5
R4071 vdd3p3.n7450 vdd3p3.n7449 92.5
R4072 vdd3p3.n7466 vdd3p3.n7465 92.5
R4073 vdd3p3.n7460 vdd3p3.n7459 92.5
R4074 vdd3p3.n7462 vdd3p3.n7461 92.5
R4075 vdd3p3.n6396 vdd3p3.n6395 92.5
R4076 vdd3p3.n6386 vdd3p3.n6385 92.5
R4077 vdd3p3.n6381 vdd3p3.n6380 92.5
R4078 vdd3p3.n6377 vdd3p3.n6376 92.5
R4079 vdd3p3.n6372 vdd3p3.n6371 92.5
R4080 vdd3p3.n6368 vdd3p3.n6367 92.5
R4081 vdd3p3.n6363 vdd3p3.n6362 92.5
R4082 vdd3p3.n6356 vdd3p3.n6355 92.5
R4083 vdd3p3.n6359 vdd3p3.n6358 92.5
R4084 vdd3p3.n6352 vdd3p3.n6351 92.5
R4085 vdd3p3.n6348 vdd3p3.n6347 92.5
R4086 vdd3p3.n6343 vdd3p3.n6342 92.5
R4087 vdd3p3.n6339 vdd3p3.n6338 92.5
R4088 vdd3p3.n6334 vdd3p3.n6333 92.5
R4089 vdd3p3.n6330 vdd3p3.n6329 92.5
R4090 vdd3p3.n6325 vdd3p3.n6324 92.5
R4091 vdd3p3.n6321 vdd3p3.n6320 92.5
R4092 vdd3p3.n6316 vdd3p3.n6315 92.5
R4093 vdd3p3.n6311 vdd3p3.n6310 92.5
R4094 vdd3p3.n6307 vdd3p3.n6306 92.5
R4095 vdd3p3.n6302 vdd3p3.n6301 92.5
R4096 vdd3p3.n6298 vdd3p3.n6297 92.5
R4097 vdd3p3.n6293 vdd3p3.n6292 92.5
R4098 vdd3p3.n6289 vdd3p3.n6288 92.5
R4099 vdd3p3.n6284 vdd3p3.n6283 92.5
R4100 vdd3p3.n6277 vdd3p3.n6276 92.5
R4101 vdd3p3.n6280 vdd3p3.n6279 92.5
R4102 vdd3p3.n6273 vdd3p3.n6272 92.5
R4103 vdd3p3.n6269 vdd3p3.n6268 92.5
R4104 vdd3p3.n6264 vdd3p3.n6263 92.5
R4105 vdd3p3.n6263 vdd3p3.n6262 92.5
R4106 vdd3p3.n6259 vdd3p3.n6258 92.5
R4107 vdd3p3.n6258 vdd3p3.n6257 92.5
R4108 vdd3p3.n6254 vdd3p3.n6253 92.5
R4109 vdd3p3.n6253 vdd3p3.n6252 92.5
R4110 vdd3p3.n6249 vdd3p3.n6248 92.5
R4111 vdd3p3.n6248 vdd3p3.n6247 92.5
R4112 vdd3p3.n6244 vdd3p3.n6243 92.5
R4113 vdd3p3.n6243 vdd3p3.n6242 92.5
R4114 vdd3p3.n6239 vdd3p3.n6238 92.5
R4115 vdd3p3.n6238 vdd3p3.n6237 92.5
R4116 vdd3p3.n6234 vdd3p3.n6233 92.5
R4117 vdd3p3.n6233 vdd3p3.n6232 92.5
R4118 vdd3p3.n6229 vdd3p3.n6228 92.5
R4119 vdd3p3.n6228 vdd3p3.n6227 92.5
R4120 vdd3p3.n6224 vdd3p3.n6223 92.5
R4121 vdd3p3.n6223 vdd3p3.n6222 92.5
R4122 vdd3p3.n6219 vdd3p3.n6218 92.5
R4123 vdd3p3.n6218 vdd3p3.n6217 92.5
R4124 vdd3p3.n6214 vdd3p3.n6213 92.5
R4125 vdd3p3.n6213 vdd3p3.n6212 92.5
R4126 vdd3p3.n6209 vdd3p3.n6208 92.5
R4127 vdd3p3.n6208 vdd3p3.n6207 92.5
R4128 vdd3p3.n6204 vdd3p3.n6203 92.5
R4129 vdd3p3.n6203 vdd3p3.n6202 92.5
R4130 vdd3p3.n6199 vdd3p3.n6198 92.5
R4131 vdd3p3.n6198 vdd3p3.n6197 92.5
R4132 vdd3p3.n6191 vdd3p3.n6190 92.5
R4133 vdd3p3.n6190 vdd3p3.n6189 92.5
R4134 vdd3p3.n6194 vdd3p3.n6193 92.5
R4135 vdd3p3.n6193 vdd3p3.n6192 92.5
R4136 vdd3p3.n6186 vdd3p3.n6185 92.5
R4137 vdd3p3.n6185 vdd3p3.n6184 92.5
R4138 vdd3p3.n6181 vdd3p3.n6180 92.5
R4139 vdd3p3.n6180 vdd3p3.n6179 92.5
R4140 vdd3p3.n6176 vdd3p3.n6175 92.5
R4141 vdd3p3.n6175 vdd3p3.n6174 92.5
R4142 vdd3p3.n6171 vdd3p3.n6170 92.5
R4143 vdd3p3.n6170 vdd3p3.n6169 92.5
R4144 vdd3p3.n6166 vdd3p3.n6165 92.5
R4145 vdd3p3.n6165 vdd3p3.n6164 92.5
R4146 vdd3p3.n6161 vdd3p3.n6160 92.5
R4147 vdd3p3.n6160 vdd3p3.n6159 92.5
R4148 vdd3p3.n6156 vdd3p3.n6155 92.5
R4149 vdd3p3.n6155 vdd3p3.n6154 92.5
R4150 vdd3p3.n6151 vdd3p3.n6150 92.5
R4151 vdd3p3.n6150 vdd3p3.n6149 92.5
R4152 vdd3p3.n6146 vdd3p3.n6145 92.5
R4153 vdd3p3.n6145 vdd3p3.n6144 92.5
R4154 vdd3p3.n6141 vdd3p3.n6140 92.5
R4155 vdd3p3.n6140 vdd3p3.n6139 92.5
R4156 vdd3p3.n6136 vdd3p3.n6135 92.5
R4157 vdd3p3.n6135 vdd3p3.n6134 92.5
R4158 vdd3p3.n6131 vdd3p3.n6130 92.5
R4159 vdd3p3.n6130 vdd3p3.n6129 92.5
R4160 vdd3p3.n6126 vdd3p3.n6125 92.5
R4161 vdd3p3.n6125 vdd3p3.n6124 92.5
R4162 vdd3p3.n6121 vdd3p3.n6120 92.5
R4163 vdd3p3.n6120 vdd3p3.n6119 92.5
R4164 vdd3p3.n5958 vdd3p3.n5957 92.5
R4165 vdd3p3.n6116 vdd3p3.n6115 92.5
R4166 vdd3p3.n6112 vdd3p3.n6111 92.5
R4167 vdd3p3.n6106 vdd3p3.n6105 92.5
R4168 vdd3p3.n6108 vdd3p3.n6107 92.5
R4169 vdd3p3.n6102 vdd3p3.n6101 92.5
R4170 vdd3p3.n6098 vdd3p3.n6097 92.5
R4171 vdd3p3.n6094 vdd3p3.n6093 92.5
R4172 vdd3p3.n6090 vdd3p3.n6089 92.5
R4173 vdd3p3.n6086 vdd3p3.n6085 92.5
R4174 vdd3p3.n6082 vdd3p3.n6081 92.5
R4175 vdd3p3.n6078 vdd3p3.n6077 92.5
R4176 vdd3p3.n6074 vdd3p3.n6073 92.5
R4177 vdd3p3.n6070 vdd3p3.n6069 92.5
R4178 vdd3p3.n6066 vdd3p3.n6065 92.5
R4179 vdd3p3.n6062 vdd3p3.n6061 92.5
R4180 vdd3p3.n6058 vdd3p3.n6057 92.5
R4181 vdd3p3.n6054 vdd3p3.n6053 92.5
R4182 vdd3p3.n6050 vdd3p3.n6049 92.5
R4183 vdd3p3.n6046 vdd3p3.n6045 92.5
R4184 vdd3p3.n6042 vdd3p3.n6041 92.5
R4185 vdd3p3.n6036 vdd3p3.n6035 92.5
R4186 vdd3p3.n6038 vdd3p3.n6037 92.5
R4187 vdd3p3.n6032 vdd3p3.n6031 92.5
R4188 vdd3p3.n6028 vdd3p3.n6027 92.5
R4189 vdd3p3.n6024 vdd3p3.n6023 92.5
R4190 vdd3p3.n6020 vdd3p3.n6019 92.5
R4191 vdd3p3.n6016 vdd3p3.n6015 92.5
R4192 vdd3p3.n6012 vdd3p3.n6011 92.5
R4193 vdd3p3.n6008 vdd3p3.n6007 92.5
R4194 vdd3p3.n6004 vdd3p3.n6003 92.5
R4195 vdd3p3.n6000 vdd3p3.n5999 92.5
R4196 vdd3p3.n5996 vdd3p3.n5995 92.5
R4197 vdd3p3.n5992 vdd3p3.n5991 92.5
R4198 vdd3p3.n5988 vdd3p3.n5987 92.5
R4199 vdd3p3.n5984 vdd3p3.n5983 92.5
R4200 vdd3p3.n5980 vdd3p3.n5979 92.5
R4201 vdd3p3.n5976 vdd3p3.n5975 92.5
R4202 vdd3p3.n5972 vdd3p3.n5971 92.5
R4203 vdd3p3.n5966 vdd3p3.n5965 92.5
R4204 vdd3p3.n5968 vdd3p3.n5967 92.5
R4205 vdd3p3.n5962 vdd3p3.n5961 92.5
R4206 vdd3p3.n5954 vdd3p3.n5953 92.5
R4207 vdd3p3.n5950 vdd3p3.n5949 92.5
R4208 vdd3p3.n5949 vdd3p3.n5948 92.5
R4209 vdd3p3.n5945 vdd3p3.n5944 92.5
R4210 vdd3p3.n5944 vdd3p3.n5943 92.5
R4211 vdd3p3.n5940 vdd3p3.n5939 92.5
R4212 vdd3p3.n5939 vdd3p3.n5938 92.5
R4213 vdd3p3.n5935 vdd3p3.n5934 92.5
R4214 vdd3p3.n5934 vdd3p3.n5933 92.5
R4215 vdd3p3.n5930 vdd3p3.n5929 92.5
R4216 vdd3p3.n5929 vdd3p3.n5928 92.5
R4217 vdd3p3.n5925 vdd3p3.n5924 92.5
R4218 vdd3p3.n5924 vdd3p3.n5923 92.5
R4219 vdd3p3.n5920 vdd3p3.n5919 92.5
R4220 vdd3p3.n5919 vdd3p3.n5918 92.5
R4221 vdd3p3.n5915 vdd3p3.n5914 92.5
R4222 vdd3p3.n5914 vdd3p3.n5913 92.5
R4223 vdd3p3.n5910 vdd3p3.n5909 92.5
R4224 vdd3p3.n5909 vdd3p3.n5908 92.5
R4225 vdd3p3.n5905 vdd3p3.n5904 92.5
R4226 vdd3p3.n5904 vdd3p3.n5903 92.5
R4227 vdd3p3.n5900 vdd3p3.n5899 92.5
R4228 vdd3p3.n5899 vdd3p3.n5898 92.5
R4229 vdd3p3.n5895 vdd3p3.n5894 92.5
R4230 vdd3p3.n5894 vdd3p3.n5893 92.5
R4231 vdd3p3.n5890 vdd3p3.n5889 92.5
R4232 vdd3p3.n5889 vdd3p3.n5888 92.5
R4233 vdd3p3.n5882 vdd3p3.n5881 92.5
R4234 vdd3p3.n5881 vdd3p3.n5880 92.5
R4235 vdd3p3.n5885 vdd3p3.n5884 92.5
R4236 vdd3p3.n5884 vdd3p3.n5883 92.5
R4237 vdd3p3.n5877 vdd3p3.n5876 92.5
R4238 vdd3p3.n5876 vdd3p3.n5875 92.5
R4239 vdd3p3.n5872 vdd3p3.n5871 92.5
R4240 vdd3p3.n5871 vdd3p3.n5870 92.5
R4241 vdd3p3.n5867 vdd3p3.n5866 92.5
R4242 vdd3p3.n5866 vdd3p3.n5865 92.5
R4243 vdd3p3.n5862 vdd3p3.n5861 92.5
R4244 vdd3p3.n5861 vdd3p3.n5860 92.5
R4245 vdd3p3.n5857 vdd3p3.n5856 92.5
R4246 vdd3p3.n5856 vdd3p3.n5855 92.5
R4247 vdd3p3.n5852 vdd3p3.n5851 92.5
R4248 vdd3p3.n5851 vdd3p3.n5850 92.5
R4249 vdd3p3.n5847 vdd3p3.n5846 92.5
R4250 vdd3p3.n5846 vdd3p3.n5845 92.5
R4251 vdd3p3.n5842 vdd3p3.n5841 92.5
R4252 vdd3p3.n5841 vdd3p3.n5840 92.5
R4253 vdd3p3.n5837 vdd3p3.n5836 92.5
R4254 vdd3p3.n5836 vdd3p3.n5835 92.5
R4255 vdd3p3.n5832 vdd3p3.n5831 92.5
R4256 vdd3p3.n5831 vdd3p3.n5830 92.5
R4257 vdd3p3.n5827 vdd3p3.n5826 92.5
R4258 vdd3p3.n5826 vdd3p3.n5825 92.5
R4259 vdd3p3.n5822 vdd3p3.n5821 92.5
R4260 vdd3p3.n5821 vdd3p3.n5820 92.5
R4261 vdd3p3.n5817 vdd3p3.n5816 92.5
R4262 vdd3p3.n5816 vdd3p3.n5815 92.5
R4263 vdd3p3.n5812 vdd3p3.n5811 92.5
R4264 vdd3p3.n5811 vdd3p3.n5810 92.5
R4265 vdd3p3.n5807 vdd3p3.n5806 92.5
R4266 vdd3p3.n5806 vdd3p3.n5805 92.5
R4267 vdd3p3.n5802 vdd3p3.n5801 92.5
R4268 vdd3p3.n5801 vdd3p3.n5800 92.5
R4269 vdd3p3.n5794 vdd3p3.n5793 92.5
R4270 vdd3p3.n5793 vdd3p3.n5792 92.5
R4271 vdd3p3.n5797 vdd3p3.n5796 92.5
R4272 vdd3p3.n5796 vdd3p3.n5795 92.5
R4273 vdd3p3.n5789 vdd3p3.n5788 92.5
R4274 vdd3p3.n5788 vdd3p3.n5787 92.5
R4275 vdd3p3.n5784 vdd3p3.n5783 92.5
R4276 vdd3p3.n5783 vdd3p3.n5782 92.5
R4277 vdd3p3.n5779 vdd3p3.n5778 92.5
R4278 vdd3p3.n5778 vdd3p3.n5777 92.5
R4279 vdd3p3.n5774 vdd3p3.n5773 92.5
R4280 vdd3p3.n5773 vdd3p3.n5772 92.5
R4281 vdd3p3.n5769 vdd3p3.n5768 92.5
R4282 vdd3p3.n5768 vdd3p3.n5767 92.5
R4283 vdd3p3.n5764 vdd3p3.n5763 92.5
R4284 vdd3p3.n5763 vdd3p3.n5762 92.5
R4285 vdd3p3.n5759 vdd3p3.n5758 92.5
R4286 vdd3p3.n5758 vdd3p3.n5757 92.5
R4287 vdd3p3.n5754 vdd3p3.n5753 92.5
R4288 vdd3p3.n5753 vdd3p3.n5752 92.5
R4289 vdd3p3.n5749 vdd3p3.n5748 92.5
R4290 vdd3p3.n5748 vdd3p3.n5747 92.5
R4291 vdd3p3.n5744 vdd3p3.n5743 92.5
R4292 vdd3p3.n5743 vdd3p3.n5742 92.5
R4293 vdd3p3.n5731 vdd3p3.n5730 92.5
R4294 vdd3p3.n5730 vdd3p3.n5729 92.5
R4295 vdd3p3.n7010 vdd3p3.n7009 92.5
R4296 vdd3p3.n7018 vdd3p3.n7017 92.5
R4297 vdd3p3.n7022 vdd3p3.n7021 92.5
R4298 vdd3p3.n5736 vdd3p3.n5735 92.5
R4299 vdd3p3.n5734 vdd3p3.n5733 92.5
R4300 vdd3p3.n5733 vdd3p3.n5732 92.5
R4301 vdd3p3.n5725 vdd3p3.n5724 92.5
R4302 vdd3p3.n5724 vdd3p3.n5723 92.5
R4303 vdd3p3.n5720 vdd3p3.n5719 92.5
R4304 vdd3p3.n5719 vdd3p3.n5718 92.5
R4305 vdd3p3.n5715 vdd3p3.n5714 92.5
R4306 vdd3p3.n5714 vdd3p3.n5713 92.5
R4307 vdd3p3.n5710 vdd3p3.n5709 92.5
R4308 vdd3p3.n5709 vdd3p3.n5708 92.5
R4309 vdd3p3.n5705 vdd3p3.n5704 92.5
R4310 vdd3p3.n5704 vdd3p3.n5703 92.5
R4311 vdd3p3.n5700 vdd3p3.n5699 92.5
R4312 vdd3p3.n5699 vdd3p3.n5698 92.5
R4313 vdd3p3.n5695 vdd3p3.n5694 92.5
R4314 vdd3p3.n5694 vdd3p3.n5693 92.5
R4315 vdd3p3.n5690 vdd3p3.n5689 92.5
R4316 vdd3p3.n5689 vdd3p3.n5688 92.5
R4317 vdd3p3.n5685 vdd3p3.n5684 92.5
R4318 vdd3p3.n5684 vdd3p3.n5683 92.5
R4319 vdd3p3.n5680 vdd3p3.n5679 92.5
R4320 vdd3p3.n5679 vdd3p3.n5678 92.5
R4321 vdd3p3.n5675 vdd3p3.n5674 92.5
R4322 vdd3p3.n5674 vdd3p3.n5673 92.5
R4323 vdd3p3.n5672 vdd3p3.n5671 92.5
R4324 vdd3p3.n5671 vdd3p3.n5670 92.5
R4325 vdd3p3.n5667 vdd3p3.n5666 92.5
R4326 vdd3p3.n5666 vdd3p3.n5665 92.5
R4327 vdd3p3.n5662 vdd3p3.n5661 92.5
R4328 vdd3p3.n5661 vdd3p3.n5660 92.5
R4329 vdd3p3.n5657 vdd3p3.n5656 92.5
R4330 vdd3p3.n5656 vdd3p3.n5655 92.5
R4331 vdd3p3.n5652 vdd3p3.n5651 92.5
R4332 vdd3p3.n5651 vdd3p3.n5650 92.5
R4333 vdd3p3.n5647 vdd3p3.n5646 92.5
R4334 vdd3p3.n5646 vdd3p3.n5645 92.5
R4335 vdd3p3.n5642 vdd3p3.n5641 92.5
R4336 vdd3p3.n5641 vdd3p3.n5640 92.5
R4337 vdd3p3.n5637 vdd3p3.n5636 92.5
R4338 vdd3p3.n5636 vdd3p3.n5635 92.5
R4339 vdd3p3.n5632 vdd3p3.n5631 92.5
R4340 vdd3p3.n5631 vdd3p3.n5630 92.5
R4341 vdd3p3.n5627 vdd3p3.n5626 92.5
R4342 vdd3p3.n5626 vdd3p3.n5625 92.5
R4343 vdd3p3.n5622 vdd3p3.n5621 92.5
R4344 vdd3p3.n5621 vdd3p3.n5620 92.5
R4345 vdd3p3.n5617 vdd3p3.n5616 92.5
R4346 vdd3p3.n5616 vdd3p3.n5615 92.5
R4347 vdd3p3.n5612 vdd3p3.n5611 92.5
R4348 vdd3p3.n5611 vdd3p3.n5610 92.5
R4349 vdd3p3.n5607 vdd3p3.n5606 92.5
R4350 vdd3p3.n5606 vdd3p3.n5605 92.5
R4351 vdd3p3.n5602 vdd3p3.n5601 92.5
R4352 vdd3p3.n5601 vdd3p3.n5600 92.5
R4353 vdd3p3.n5597 vdd3p3.n5596 92.5
R4354 vdd3p3.n5596 vdd3p3.n5595 92.5
R4355 vdd3p3.n5592 vdd3p3.n5591 92.5
R4356 vdd3p3.n5591 vdd3p3.n5590 92.5
R4357 vdd3p3.n5587 vdd3p3.n5586 92.5
R4358 vdd3p3.n5586 vdd3p3.n5585 92.5
R4359 vdd3p3.n5584 vdd3p3.n5583 92.5
R4360 vdd3p3.n5583 vdd3p3.n5582 92.5
R4361 vdd3p3.n5579 vdd3p3.n5578 92.5
R4362 vdd3p3.n5578 vdd3p3.n5577 92.5
R4363 vdd3p3.n5574 vdd3p3.n5573 92.5
R4364 vdd3p3.n5573 vdd3p3.n5572 92.5
R4365 vdd3p3.n5569 vdd3p3.n5568 92.5
R4366 vdd3p3.n5568 vdd3p3.n5567 92.5
R4367 vdd3p3.n5564 vdd3p3.n5563 92.5
R4368 vdd3p3.n5563 vdd3p3.n5562 92.5
R4369 vdd3p3.n5559 vdd3p3.n5558 92.5
R4370 vdd3p3.n5558 vdd3p3.n5557 92.5
R4371 vdd3p3.n5554 vdd3p3.n5553 92.5
R4372 vdd3p3.n5553 vdd3p3.n5552 92.5
R4373 vdd3p3.n5549 vdd3p3.n5548 92.5
R4374 vdd3p3.n5548 vdd3p3.n5547 92.5
R4375 vdd3p3.n5544 vdd3p3.n5543 92.5
R4376 vdd3p3.n5543 vdd3p3.n5542 92.5
R4377 vdd3p3.n5539 vdd3p3.n5538 92.5
R4378 vdd3p3.n5538 vdd3p3.n5537 92.5
R4379 vdd3p3.n5534 vdd3p3.n5533 92.5
R4380 vdd3p3.n5533 vdd3p3.n5532 92.5
R4381 vdd3p3.n5529 vdd3p3.n5528 92.5
R4382 vdd3p3.n5528 vdd3p3.n5527 92.5
R4383 vdd3p3.n5524 vdd3p3.n5523 92.5
R4384 vdd3p3.n5523 vdd3p3.n5522 92.5
R4385 vdd3p3.n5519 vdd3p3.n5518 92.5
R4386 vdd3p3.n5518 vdd3p3.n5517 92.5
R4387 vdd3p3.n5514 vdd3p3.n5513 92.5
R4388 vdd3p3.n5513 vdd3p3.n5512 92.5
R4389 vdd3p3.n5509 vdd3p3.n5508 92.5
R4390 vdd3p3.n5508 vdd3p3.n5507 92.5
R4391 vdd3p3.n5504 vdd3p3.n5503 92.5
R4392 vdd3p3.n5503 vdd3p3.n5502 92.5
R4393 vdd3p3.n5499 vdd3p3.n5498 92.5
R4394 vdd3p3.n5498 vdd3p3.n5497 92.5
R4395 vdd3p3.n5496 vdd3p3.n5495 92.5
R4396 vdd3p3.n5495 vdd3p3.n5494 92.5
R4397 vdd3p3.n5491 vdd3p3.n5490 92.5
R4398 vdd3p3.n5490 vdd3p3.n5489 92.5
R4399 vdd3p3.n5486 vdd3p3.n5485 92.5
R4400 vdd3p3.n5485 vdd3p3.n5484 92.5
R4401 vdd3p3.n5481 vdd3p3.n5480 92.5
R4402 vdd3p3.n5480 vdd3p3.n5479 92.5
R4403 vdd3p3.n5476 vdd3p3.n5475 92.5
R4404 vdd3p3.n5475 vdd3p3.n5474 92.5
R4405 vdd3p3.n5471 vdd3p3.n5470 92.5
R4406 vdd3p3.n5470 vdd3p3.n5469 92.5
R4407 vdd3p3.n5466 vdd3p3.n5465 92.5
R4408 vdd3p3.n5465 vdd3p3.n5464 92.5
R4409 vdd3p3.n5461 vdd3p3.n5460 92.5
R4410 vdd3p3.n5460 vdd3p3.n5459 92.5
R4411 vdd3p3.n5456 vdd3p3.n5455 92.5
R4412 vdd3p3.n5455 vdd3p3.n5454 92.5
R4413 vdd3p3.n5451 vdd3p3.n5450 92.5
R4414 vdd3p3.n5450 vdd3p3.n5449 92.5
R4415 vdd3p3.n5446 vdd3p3.n5445 92.5
R4416 vdd3p3.n5445 vdd3p3.n5444 92.5
R4417 vdd3p3.n5441 vdd3p3.n5440 92.5
R4418 vdd3p3.n5440 vdd3p3.n5439 92.5
R4419 vdd3p3.n5436 vdd3p3.n5435 92.5
R4420 vdd3p3.n5435 vdd3p3.n5434 92.5
R4421 vdd3p3.n5431 vdd3p3.n5430 92.5
R4422 vdd3p3.n5430 vdd3p3.n5429 92.5
R4423 vdd3p3.n5426 vdd3p3.n5425 92.5
R4424 vdd3p3.n5425 vdd3p3.n5424 92.5
R4425 vdd3p3.n5421 vdd3p3.n5420 92.5
R4426 vdd3p3.n5420 vdd3p3.n5419 92.5
R4427 vdd3p3.n5416 vdd3p3.n5415 92.5
R4428 vdd3p3.n5415 vdd3p3.n5414 92.5
R4429 vdd3p3.n5411 vdd3p3.n5410 92.5
R4430 vdd3p3.n5410 vdd3p3.n5409 92.5
R4431 vdd3p3.n5408 vdd3p3.n5407 92.5
R4432 vdd3p3.n5407 vdd3p3.n5406 92.5
R4433 vdd3p3.n5403 vdd3p3.n5402 92.5
R4434 vdd3p3.n5402 vdd3p3.n5401 92.5
R4435 vdd3p3.n5398 vdd3p3.n5397 92.5
R4436 vdd3p3.n5397 vdd3p3.n5396 92.5
R4437 vdd3p3.n5393 vdd3p3.n5392 92.5
R4438 vdd3p3.n5392 vdd3p3.n5391 92.5
R4439 vdd3p3.n5388 vdd3p3.n5387 92.5
R4440 vdd3p3.n5387 vdd3p3.n5386 92.5
R4441 vdd3p3.n5383 vdd3p3.n5382 92.5
R4442 vdd3p3.n5382 vdd3p3.n5381 92.5
R4443 vdd3p3.n5378 vdd3p3.n5377 92.5
R4444 vdd3p3.n5377 vdd3p3.n5376 92.5
R4445 vdd3p3.n5373 vdd3p3.n5372 92.5
R4446 vdd3p3.n5372 vdd3p3.n5371 92.5
R4447 vdd3p3.n5368 vdd3p3.n5367 92.5
R4448 vdd3p3.n5367 vdd3p3.n5366 92.5
R4449 vdd3p3.n5363 vdd3p3.n5362 92.5
R4450 vdd3p3.n5362 vdd3p3.n5361 92.5
R4451 vdd3p3.n5358 vdd3p3.n5357 92.5
R4452 vdd3p3.n5357 vdd3p3.n5356 92.5
R4453 vdd3p3.n5353 vdd3p3.n5352 92.5
R4454 vdd3p3.n5352 vdd3p3.n5351 92.5
R4455 vdd3p3.n5348 vdd3p3.n5347 92.5
R4456 vdd3p3.n5347 vdd3p3.n5346 92.5
R4457 vdd3p3.n6720 vdd3p3.n6719 92.5
R4458 vdd3p3.n6719 vdd3p3.n6718 92.5
R4459 vdd3p3.n6725 vdd3p3.n6724 92.5
R4460 vdd3p3.n6724 vdd3p3.n6723 92.5
R4461 vdd3p3.n6730 vdd3p3.n6729 92.5
R4462 vdd3p3.n6729 vdd3p3.n6728 92.5
R4463 vdd3p3.n6735 vdd3p3.n6734 92.5
R4464 vdd3p3.n6734 vdd3p3.n6733 92.5
R4465 vdd3p3.n6743 vdd3p3.n6742 92.5
R4466 vdd3p3.n6742 vdd3p3.n6741 92.5
R4467 vdd3p3.n6740 vdd3p3.n6739 92.5
R4468 vdd3p3.n6739 vdd3p3.n6738 92.5
R4469 vdd3p3.n6748 vdd3p3.n6747 92.5
R4470 vdd3p3.n6747 vdd3p3.n6746 92.5
R4471 vdd3p3.n6753 vdd3p3.n6752 92.5
R4472 vdd3p3.n6752 vdd3p3.n6751 92.5
R4473 vdd3p3.n6758 vdd3p3.n6757 92.5
R4474 vdd3p3.n6757 vdd3p3.n6756 92.5
R4475 vdd3p3.n6763 vdd3p3.n6762 92.5
R4476 vdd3p3.n6762 vdd3p3.n6761 92.5
R4477 vdd3p3.n6768 vdd3p3.n6767 92.5
R4478 vdd3p3.n6767 vdd3p3.n6766 92.5
R4479 vdd3p3.n6773 vdd3p3.n6772 92.5
R4480 vdd3p3.n6772 vdd3p3.n6771 92.5
R4481 vdd3p3.n6778 vdd3p3.n6777 92.5
R4482 vdd3p3.n6777 vdd3p3.n6776 92.5
R4483 vdd3p3.n6783 vdd3p3.n6782 92.5
R4484 vdd3p3.n6782 vdd3p3.n6781 92.5
R4485 vdd3p3.n6788 vdd3p3.n6787 92.5
R4486 vdd3p3.n6787 vdd3p3.n6786 92.5
R4487 vdd3p3.n6793 vdd3p3.n6792 92.5
R4488 vdd3p3.n6792 vdd3p3.n6791 92.5
R4489 vdd3p3.n6798 vdd3p3.n6797 92.5
R4490 vdd3p3.n6797 vdd3p3.n6796 92.5
R4491 vdd3p3.n6803 vdd3p3.n6802 92.5
R4492 vdd3p3.n6802 vdd3p3.n6801 92.5
R4493 vdd3p3.n6808 vdd3p3.n6807 92.5
R4494 vdd3p3.n6807 vdd3p3.n6806 92.5
R4495 vdd3p3.n6813 vdd3p3.n6812 92.5
R4496 vdd3p3.n6812 vdd3p3.n6811 92.5
R4497 vdd3p3.n6818 vdd3p3.n6817 92.5
R4498 vdd3p3.n6817 vdd3p3.n6816 92.5
R4499 vdd3p3.n6823 vdd3p3.n6822 92.5
R4500 vdd3p3.n6822 vdd3p3.n6821 92.5
R4501 vdd3p3.n6831 vdd3p3.n6830 92.5
R4502 vdd3p3.n6830 vdd3p3.n6829 92.5
R4503 vdd3p3.n6828 vdd3p3.n6827 92.5
R4504 vdd3p3.n6827 vdd3p3.n6826 92.5
R4505 vdd3p3.n6836 vdd3p3.n6835 92.5
R4506 vdd3p3.n6835 vdd3p3.n6834 92.5
R4507 vdd3p3.n6841 vdd3p3.n6840 92.5
R4508 vdd3p3.n6840 vdd3p3.n6839 92.5
R4509 vdd3p3.n6846 vdd3p3.n6845 92.5
R4510 vdd3p3.n6845 vdd3p3.n6844 92.5
R4511 vdd3p3.n6851 vdd3p3.n6850 92.5
R4512 vdd3p3.n6850 vdd3p3.n6849 92.5
R4513 vdd3p3.n6856 vdd3p3.n6855 92.5
R4514 vdd3p3.n6855 vdd3p3.n6854 92.5
R4515 vdd3p3.n6861 vdd3p3.n6860 92.5
R4516 vdd3p3.n6860 vdd3p3.n6859 92.5
R4517 vdd3p3.n6866 vdd3p3.n6865 92.5
R4518 vdd3p3.n6865 vdd3p3.n6864 92.5
R4519 vdd3p3.n6871 vdd3p3.n6870 92.5
R4520 vdd3p3.n6870 vdd3p3.n6869 92.5
R4521 vdd3p3.n6876 vdd3p3.n6875 92.5
R4522 vdd3p3.n6875 vdd3p3.n6874 92.5
R4523 vdd3p3.n6881 vdd3p3.n6880 92.5
R4524 vdd3p3.n6880 vdd3p3.n6879 92.5
R4525 vdd3p3.n6886 vdd3p3.n6885 92.5
R4526 vdd3p3.n6885 vdd3p3.n6884 92.5
R4527 vdd3p3.n6891 vdd3p3.n6890 92.5
R4528 vdd3p3.n6890 vdd3p3.n6889 92.5
R4529 vdd3p3.n6896 vdd3p3.n6895 92.5
R4530 vdd3p3.n6895 vdd3p3.n6894 92.5
R4531 vdd3p3.n6901 vdd3p3.n6900 92.5
R4532 vdd3p3.n6900 vdd3p3.n6899 92.5
R4533 vdd3p3.n6906 vdd3p3.n6905 92.5
R4534 vdd3p3.n6905 vdd3p3.n6904 92.5
R4535 vdd3p3.n6911 vdd3p3.n6910 92.5
R4536 vdd3p3.n6910 vdd3p3.n6909 92.5
R4537 vdd3p3.n6919 vdd3p3.n6918 92.5
R4538 vdd3p3.n6918 vdd3p3.n6917 92.5
R4539 vdd3p3.n6916 vdd3p3.n6915 92.5
R4540 vdd3p3.n6915 vdd3p3.n6914 92.5
R4541 vdd3p3.n6924 vdd3p3.n6923 92.5
R4542 vdd3p3.n6923 vdd3p3.n6922 92.5
R4543 vdd3p3.n6929 vdd3p3.n6928 92.5
R4544 vdd3p3.n6928 vdd3p3.n6927 92.5
R4545 vdd3p3.n6934 vdd3p3.n6933 92.5
R4546 vdd3p3.n6933 vdd3p3.n6932 92.5
R4547 vdd3p3.n6939 vdd3p3.n6938 92.5
R4548 vdd3p3.n6938 vdd3p3.n6937 92.5
R4549 vdd3p3.n6944 vdd3p3.n6943 92.5
R4550 vdd3p3.n6943 vdd3p3.n6942 92.5
R4551 vdd3p3.n6949 vdd3p3.n6948 92.5
R4552 vdd3p3.n6948 vdd3p3.n6947 92.5
R4553 vdd3p3.n6954 vdd3p3.n6953 92.5
R4554 vdd3p3.n6953 vdd3p3.n6952 92.5
R4555 vdd3p3.n6959 vdd3p3.n6958 92.5
R4556 vdd3p3.n6958 vdd3p3.n6957 92.5
R4557 vdd3p3.n6964 vdd3p3.n6963 92.5
R4558 vdd3p3.n6963 vdd3p3.n6962 92.5
R4559 vdd3p3.n6969 vdd3p3.n6968 92.5
R4560 vdd3p3.n6968 vdd3p3.n6967 92.5
R4561 vdd3p3.n6974 vdd3p3.n6973 92.5
R4562 vdd3p3.n6973 vdd3p3.n6972 92.5
R4563 vdd3p3.n6979 vdd3p3.n6978 92.5
R4564 vdd3p3.n6978 vdd3p3.n6977 92.5
R4565 vdd3p3.n6984 vdd3p3.n6983 92.5
R4566 vdd3p3.n6983 vdd3p3.n6982 92.5
R4567 vdd3p3.n6989 vdd3p3.n6988 92.5
R4568 vdd3p3.n6988 vdd3p3.n6987 92.5
R4569 vdd3p3.n6994 vdd3p3.n6993 92.5
R4570 vdd3p3.n6993 vdd3p3.n6992 92.5
R4571 vdd3p3.n6999 vdd3p3.n6998 92.5
R4572 vdd3p3.n6998 vdd3p3.n6997 92.5
R4573 vdd3p3.n7014 vdd3p3.n7013 92.5
R4574 vdd3p3.n7013 vdd3p3.n7012 92.5
R4575 vdd3p3.n7003 vdd3p3.n7002 92.5
R4576 vdd3p3.n7006 vdd3p3.n7005 92.5
R4577 vdd3p3.n7027 vdd3p3.n7026 92.5
R4578 vdd3p3.n7026 vdd3p3.n7025 92.5
R4579 vdd3p3.n7032 vdd3p3.n7031 92.5
R4580 vdd3p3.n7031 vdd3p3.n7030 92.5
R4581 vdd3p3.n7037 vdd3p3.n7036 92.5
R4582 vdd3p3.n7036 vdd3p3.n7035 92.5
R4583 vdd3p3.n7042 vdd3p3.n7041 92.5
R4584 vdd3p3.n7041 vdd3p3.n7040 92.5
R4585 vdd3p3.n7047 vdd3p3.n7046 92.5
R4586 vdd3p3.n7046 vdd3p3.n7045 92.5
R4587 vdd3p3.n7052 vdd3p3.n7051 92.5
R4588 vdd3p3.n7051 vdd3p3.n7050 92.5
R4589 vdd3p3.n7057 vdd3p3.n7056 92.5
R4590 vdd3p3.n7056 vdd3p3.n7055 92.5
R4591 vdd3p3.n7065 vdd3p3.n7064 92.5
R4592 vdd3p3.n7064 vdd3p3.n7063 92.5
R4593 vdd3p3.n7062 vdd3p3.n7061 92.5
R4594 vdd3p3.n7061 vdd3p3.n7060 92.5
R4595 vdd3p3.n7070 vdd3p3.n7069 92.5
R4596 vdd3p3.n7069 vdd3p3.n7068 92.5
R4597 vdd3p3.n7075 vdd3p3.n7074 92.5
R4598 vdd3p3.n7074 vdd3p3.n7073 92.5
R4599 vdd3p3.n7080 vdd3p3.n7079 92.5
R4600 vdd3p3.n7079 vdd3p3.n7078 92.5
R4601 vdd3p3.n7085 vdd3p3.n7084 92.5
R4602 vdd3p3.n7084 vdd3p3.n7083 92.5
R4603 vdd3p3.n7090 vdd3p3.n7089 92.5
R4604 vdd3p3.n7089 vdd3p3.n7088 92.5
R4605 vdd3p3.n7095 vdd3p3.n7094 92.5
R4606 vdd3p3.n7094 vdd3p3.n7093 92.5
R4607 vdd3p3.n7100 vdd3p3.n7099 92.5
R4608 vdd3p3.n7099 vdd3p3.n7098 92.5
R4609 vdd3p3.n7105 vdd3p3.n7104 92.5
R4610 vdd3p3.n7104 vdd3p3.n7103 92.5
R4611 vdd3p3.n7109 vdd3p3.n7108 92.5
R4612 vdd3p3.n7108 vdd3p3.n7107 92.5
R4613 vdd3p3.n7114 vdd3p3.n7113 92.5
R4614 vdd3p3.n7113 vdd3p3.n7112 92.5
R4615 vdd3p3.n7119 vdd3p3.n7118 92.5
R4616 vdd3p3.n7118 vdd3p3.n7117 92.5
R4617 vdd3p3.n7124 vdd3p3.n7123 92.5
R4618 vdd3p3.n7123 vdd3p3.n7122 92.5
R4619 vdd3p3.n7129 vdd3p3.n7128 92.5
R4620 vdd3p3.n7128 vdd3p3.n7127 92.5
R4621 vdd3p3.n7134 vdd3p3.n7133 92.5
R4622 vdd3p3.n7133 vdd3p3.n7132 92.5
R4623 vdd3p3.n7139 vdd3p3.n7138 92.5
R4624 vdd3p3.n7138 vdd3p3.n7137 92.5
R4625 vdd3p3.n7144 vdd3p3.n7143 92.5
R4626 vdd3p3.n7143 vdd3p3.n7142 92.5
R4627 vdd3p3.n7152 vdd3p3.n7151 92.5
R4628 vdd3p3.n7151 vdd3p3.n7150 92.5
R4629 vdd3p3.n7149 vdd3p3.n7148 92.5
R4630 vdd3p3.n7148 vdd3p3.n7147 92.5
R4631 vdd3p3.n7157 vdd3p3.n7156 92.5
R4632 vdd3p3.n7156 vdd3p3.n7155 92.5
R4633 vdd3p3.n7162 vdd3p3.n7161 92.5
R4634 vdd3p3.n7161 vdd3p3.n7160 92.5
R4635 vdd3p3.n7167 vdd3p3.n7166 92.5
R4636 vdd3p3.n7166 vdd3p3.n7165 92.5
R4637 vdd3p3.n7172 vdd3p3.n7171 92.5
R4638 vdd3p3.n7171 vdd3p3.n7170 92.5
R4639 vdd3p3.n7177 vdd3p3.n7176 92.5
R4640 vdd3p3.n7176 vdd3p3.n7175 92.5
R4641 vdd3p3.n7182 vdd3p3.n7181 92.5
R4642 vdd3p3.n7181 vdd3p3.n7180 92.5
R4643 vdd3p3.n7187 vdd3p3.n7186 92.5
R4644 vdd3p3.n7186 vdd3p3.n7185 92.5
R4645 vdd3p3.n7192 vdd3p3.n7191 92.5
R4646 vdd3p3.n7191 vdd3p3.n7190 92.5
R4647 vdd3p3.n7196 vdd3p3.n7195 92.5
R4648 vdd3p3.n7195 vdd3p3.n7194 92.5
R4649 vdd3p3.n7201 vdd3p3.n7200 92.5
R4650 vdd3p3.n7200 vdd3p3.n7199 92.5
R4651 vdd3p3.n7206 vdd3p3.n7205 92.5
R4652 vdd3p3.n7205 vdd3p3.n7204 92.5
R4653 vdd3p3.n7211 vdd3p3.n7210 92.5
R4654 vdd3p3.n7210 vdd3p3.n7209 92.5
R4655 vdd3p3.n7216 vdd3p3.n7215 92.5
R4656 vdd3p3.n7215 vdd3p3.n7214 92.5
R4657 vdd3p3.n7221 vdd3p3.n7220 92.5
R4658 vdd3p3.n7220 vdd3p3.n7219 92.5
R4659 vdd3p3.n7226 vdd3p3.n7225 92.5
R4660 vdd3p3.n7225 vdd3p3.n7224 92.5
R4661 vdd3p3.n7231 vdd3p3.n7230 92.5
R4662 vdd3p3.n7230 vdd3p3.n7229 92.5
R4663 vdd3p3.n7237 vdd3p3.n7236 92.5
R4664 vdd3p3.n5196 vdd3p3.n5195 92.5
R4665 vdd3p3.n5198 vdd3p3.n5197 92.5
R4666 vdd3p3.n5200 vdd3p3.n5199 92.5
R4667 vdd3p3.n5202 vdd3p3.n5201 92.5
R4668 vdd3p3.n5204 vdd3p3.n5203 92.5
R4669 vdd3p3.n5207 vdd3p3.n5206 92.5
R4670 vdd3p3.n5210 vdd3p3.n5209 92.5
R4671 vdd3p3.n5213 vdd3p3.n5212 92.5
R4672 vdd3p3.n5216 vdd3p3.n5215 92.5
R4673 vdd3p3.n5219 vdd3p3.n5218 92.5
R4674 vdd3p3.n5222 vdd3p3.n5221 92.5
R4675 vdd3p3.n5225 vdd3p3.n5224 92.5
R4676 vdd3p3.n5228 vdd3p3.n5227 92.5
R4677 vdd3p3.n5231 vdd3p3.n5230 92.5
R4678 vdd3p3.n5234 vdd3p3.n5233 92.5
R4679 vdd3p3.n5237 vdd3p3.n5236 92.5
R4680 vdd3p3.n5240 vdd3p3.n5239 92.5
R4681 vdd3p3.n5243 vdd3p3.n5242 92.5
R4682 vdd3p3.n5246 vdd3p3.n5245 92.5
R4683 vdd3p3.n5249 vdd3p3.n5248 92.5
R4684 vdd3p3.n5252 vdd3p3.n5251 92.5
R4685 vdd3p3.n5255 vdd3p3.n5254 92.5
R4686 vdd3p3.n5258 vdd3p3.n5257 92.5
R4687 vdd3p3.n5261 vdd3p3.n5260 92.5
R4688 vdd3p3.n5265 vdd3p3.n5264 92.5
R4689 vdd3p3.n5179 vdd3p3.n5178 92.5
R4690 vdd3p3.n5176 vdd3p3.n5175 92.5
R4691 vdd3p3.n5173 vdd3p3.n5172 92.5
R4692 vdd3p3.n5170 vdd3p3.n5169 92.5
R4693 vdd3p3.n5167 vdd3p3.n5166 92.5
R4694 vdd3p3.n5164 vdd3p3.n5163 92.5
R4695 vdd3p3.n5302 vdd3p3.n5301 92.5
R4696 vdd3p3.n5305 vdd3p3.n5304 92.5
R4697 vdd3p3.n5308 vdd3p3.n5307 92.5
R4698 vdd3p3.n5311 vdd3p3.n5310 92.5
R4699 vdd3p3.n5314 vdd3p3.n5313 92.5
R4700 vdd3p3.n5317 vdd3p3.n5316 92.5
R4701 vdd3p3.n5320 vdd3p3.n5319 92.5
R4702 vdd3p3.n5300 vdd3p3.n5299 92.5
R4703 vdd3p3.n5296 vdd3p3.n5295 92.5
R4704 vdd3p3.n5293 vdd3p3.n5292 92.5
R4705 vdd3p3.n5290 vdd3p3.n5289 92.5
R4706 vdd3p3.n5287 vdd3p3.n5286 92.5
R4707 vdd3p3.n5284 vdd3p3.n5283 92.5
R4708 vdd3p3.n5281 vdd3p3.n5280 92.5
R4709 vdd3p3.n5323 vdd3p3.n5322 92.5
R4710 vdd3p3.n5326 vdd3p3.n5325 92.5
R4711 vdd3p3.n5329 vdd3p3.n5328 92.5
R4712 vdd3p3.n5332 vdd3p3.n5331 92.5
R4713 vdd3p3.n5335 vdd3p3.n5334 92.5
R4714 vdd3p3.n5338 vdd3p3.n5337 92.5
R4715 vdd3p3.n5194 vdd3p3.n5193 92.5
R4716 vdd3p3.n5192 vdd3p3.n5191 92.5
R4717 vdd3p3.n5190 vdd3p3.n5189 92.5
R4718 vdd3p3.n5188 vdd3p3.n5187 92.5
R4719 vdd3p3.n8408 vdd3p3.n8407 92.5
R4720 vdd3p3.n8399 vdd3p3.n8398 92.5
R4721 vdd3p3.n8390 vdd3p3.n8389 92.5
R4722 vdd3p3.n8382 vdd3p3.n8381 92.5
R4723 vdd3p3.n8373 vdd3p3.n8372 92.5
R4724 vdd3p3.n8361 vdd3p3.n8360 92.5
R4725 vdd3p3.n8352 vdd3p3.n8351 92.5
R4726 vdd3p3.n8342 vdd3p3.n8341 92.5
R4727 vdd3p3.n8343 vdd3p3.n8342 92.5
R4728 vdd3p3.n8332 vdd3p3.n8331 92.5
R4729 vdd3p3.n8333 vdd3p3.n8332 92.5
R4730 vdd3p3.n8322 vdd3p3.n8321 92.5
R4731 vdd3p3.n8323 vdd3p3.n8322 92.5
R4732 vdd3p3.n8312 vdd3p3.n8311 92.5
R4733 vdd3p3.n8313 vdd3p3.n8312 92.5
R4734 vdd3p3.n8302 vdd3p3.n8301 92.5
R4735 vdd3p3.n8303 vdd3p3.n8302 92.5
R4736 vdd3p3.n4067 vdd3p3.n4066 92.5
R4737 vdd3p3.n4068 vdd3p3.n4067 92.5
R4738 vdd3p3.n4071 vdd3p3.n4070 92.5
R4739 vdd3p3.n4072 vdd3p3.n4071 92.5
R4740 vdd3p3.n4075 vdd3p3.n4074 92.5
R4741 vdd3p3.n4076 vdd3p3.n4075 92.5
R4742 vdd3p3.n4079 vdd3p3.n4078 92.5
R4743 vdd3p3.n4080 vdd3p3.n4079 92.5
R4744 vdd3p3.n4083 vdd3p3.n4082 92.5
R4745 vdd3p3.n4084 vdd3p3.n4083 92.5
R4746 vdd3p3.n4087 vdd3p3.n4086 92.5
R4747 vdd3p3.n4088 vdd3p3.n4087 92.5
R4748 vdd3p3.n4091 vdd3p3.n4090 92.5
R4749 vdd3p3.n4092 vdd3p3.n4091 92.5
R4750 vdd3p3.n4095 vdd3p3.n4094 92.5
R4751 vdd3p3.n4096 vdd3p3.n4095 92.5
R4752 vdd3p3.n4099 vdd3p3.n4098 92.5
R4753 vdd3p3.n4100 vdd3p3.n4099 92.5
R4754 vdd3p3.n4103 vdd3p3.n4102 92.5
R4755 vdd3p3.n4104 vdd3p3.n4103 92.5
R4756 vdd3p3.n4107 vdd3p3.n4106 92.5
R4757 vdd3p3.n4108 vdd3p3.n4107 92.5
R4758 vdd3p3.n4111 vdd3p3.n4110 92.5
R4759 vdd3p3.n4112 vdd3p3.n4111 92.5
R4760 vdd3p3.n4115 vdd3p3.n4114 92.5
R4761 vdd3p3.n4116 vdd3p3.n4115 92.5
R4762 vdd3p3.n4119 vdd3p3.n4118 92.5
R4763 vdd3p3.n4120 vdd3p3.n4119 92.5
R4764 vdd3p3.n4123 vdd3p3.n4122 92.5
R4765 vdd3p3.n4124 vdd3p3.n4123 92.5
R4766 vdd3p3.n4127 vdd3p3.n4126 92.5
R4767 vdd3p3.n4128 vdd3p3.n4127 92.5
R4768 vdd3p3.n4131 vdd3p3.n4130 92.5
R4769 vdd3p3.n4132 vdd3p3.n4131 92.5
R4770 vdd3p3.n4135 vdd3p3.n4134 92.5
R4771 vdd3p3.n4136 vdd3p3.n4135 92.5
R4772 vdd3p3.n4139 vdd3p3.n4138 92.5
R4773 vdd3p3.n4140 vdd3p3.n4139 92.5
R4774 vdd3p3.n4143 vdd3p3.n4142 92.5
R4775 vdd3p3.n4144 vdd3p3.n4143 92.5
R4776 vdd3p3.n4060 vdd3p3.n4059 92.5
R4777 vdd3p3.n4061 vdd3p3.n4060 92.5
R4778 vdd3p3.n4055 vdd3p3.n4054 92.5
R4779 vdd3p3.n4056 vdd3p3.n4055 92.5
R4780 vdd3p3.n4051 vdd3p3.n4050 92.5
R4781 vdd3p3.n4052 vdd3p3.n4051 92.5
R4782 vdd3p3.n4047 vdd3p3.n4046 92.5
R4783 vdd3p3.n4048 vdd3p3.n4047 92.5
R4784 vdd3p3.n4043 vdd3p3.n4042 92.5
R4785 vdd3p3.n4044 vdd3p3.n4043 92.5
R4786 vdd3p3.n4039 vdd3p3.n4038 92.5
R4787 vdd3p3.n4040 vdd3p3.n4039 92.5
R4788 vdd3p3.n4020 vdd3p3.n4019 92.5
R4789 vdd3p3.n4021 vdd3p3.n4020 92.5
R4790 vdd3p3.n4024 vdd3p3.n4023 92.5
R4791 vdd3p3.n4025 vdd3p3.n4024 92.5
R4792 vdd3p3.n4028 vdd3p3.n4027 92.5
R4793 vdd3p3.n4029 vdd3p3.n4028 92.5
R4794 vdd3p3.n4032 vdd3p3.n4031 92.5
R4795 vdd3p3.n4033 vdd3p3.n4032 92.5
R4796 vdd3p3.n4017 vdd3p3.n4016 92.5
R4797 vdd3p3.n4018 vdd3p3.n4017 92.5
R4798 vdd3p3.n4013 vdd3p3.n4012 92.5
R4799 vdd3p3.n4014 vdd3p3.n4013 92.5
R4800 vdd3p3.n4009 vdd3p3.n4008 92.5
R4801 vdd3p3.n4010 vdd3p3.n4009 92.5
R4802 vdd3p3.n4005 vdd3p3.n4004 92.5
R4803 vdd3p3.n4006 vdd3p3.n4005 92.5
R4804 vdd3p3.n3877 vdd3p3.n3876 92.5
R4805 vdd3p3.n3878 vdd3p3.n3877 92.5
R4806 vdd3p3.n3881 vdd3p3.n3880 92.5
R4807 vdd3p3.n3882 vdd3p3.n3881 92.5
R4808 vdd3p3.n3885 vdd3p3.n3884 92.5
R4809 vdd3p3.n3886 vdd3p3.n3885 92.5
R4810 vdd3p3.n3889 vdd3p3.n3888 92.5
R4811 vdd3p3.n3890 vdd3p3.n3889 92.5
R4812 vdd3p3.n3893 vdd3p3.n3892 92.5
R4813 vdd3p3.n3894 vdd3p3.n3893 92.5
R4814 vdd3p3.n3976 vdd3p3.n3975 92.5
R4815 vdd3p3.n3977 vdd3p3.n3976 92.5
R4816 vdd3p3.n3971 vdd3p3.n3970 92.5
R4817 vdd3p3.n3972 vdd3p3.n3971 92.5
R4818 vdd3p3.n3967 vdd3p3.n3966 92.5
R4819 vdd3p3.n3968 vdd3p3.n3967 92.5
R4820 vdd3p3.n3963 vdd3p3.n3962 92.5
R4821 vdd3p3.n3964 vdd3p3.n3963 92.5
R4822 vdd3p3.n3958 vdd3p3.n3957 92.5
R4823 vdd3p3.n3959 vdd3p3.n3958 92.5
R4824 vdd3p3.n3917 vdd3p3.n3916 92.5
R4825 vdd3p3.n3918 vdd3p3.n3917 92.5
R4826 vdd3p3.n3913 vdd3p3.n3912 92.5
R4827 vdd3p3.n3914 vdd3p3.n3913 92.5
R4828 vdd3p3.n7235 vdd3p3.n7234 92.5
R4829 vdd3p3.n7241 vdd3p3.n7240 92.5
R4830 vdd3p3.n7245 vdd3p3.n7244 92.5
R4831 vdd3p3.n7249 vdd3p3.n7248 92.5
R4832 vdd3p3.n7253 vdd3p3.n7252 92.5
R4833 vdd3p3.n7257 vdd3p3.n7256 92.5
R4834 vdd3p3.n7261 vdd3p3.n7260 92.5
R4835 vdd3p3.n7265 vdd3p3.n7264 92.5
R4836 vdd3p3.n7269 vdd3p3.n7268 92.5
R4837 vdd3p3.n7272 vdd3p3.n7271 92.5
R4838 vdd3p3.n7276 vdd3p3.n7275 92.5
R4839 vdd3p3.n7280 vdd3p3.n7279 92.5
R4840 vdd3p3.n7284 vdd3p3.n7283 92.5
R4841 vdd3p3.n7288 vdd3p3.n7287 92.5
R4842 vdd3p3.n7292 vdd3p3.n7291 92.5
R4843 vdd3p3.n7296 vdd3p3.n7295 92.5
R4844 vdd3p3.n7300 vdd3p3.n7299 92.5
R4845 vdd3p3.n7306 vdd3p3.n7305 92.5
R4846 vdd3p3.n7304 vdd3p3.n7303 92.5
R4847 vdd3p3.n7310 vdd3p3.n7309 92.5
R4848 vdd3p3.n7314 vdd3p3.n7313 92.5
R4849 vdd3p3.n7318 vdd3p3.n7317 92.5
R4850 vdd3p3.n7322 vdd3p3.n7321 92.5
R4851 vdd3p3.n7326 vdd3p3.n7325 92.5
R4852 vdd3p3.n7330 vdd3p3.n7329 92.5
R4853 vdd3p3.n7334 vdd3p3.n7333 92.5
R4854 vdd3p3.n7338 vdd3p3.n7337 92.5
R4855 vdd3p3.n7341 vdd3p3.n7340 92.5
R4856 vdd3p3.n7345 vdd3p3.n7344 92.5
R4857 vdd3p3.n7349 vdd3p3.n7348 92.5
R4858 vdd3p3.n7353 vdd3p3.n7352 92.5
R4859 vdd3p3.n7357 vdd3p3.n7356 92.5
R4860 vdd3p3.n7361 vdd3p3.n7360 92.5
R4861 vdd3p3.n7365 vdd3p3.n7364 92.5
R4862 vdd3p3.n7369 vdd3p3.n7368 92.5
R4863 vdd3p3.n7375 vdd3p3.n7374 92.5
R4864 vdd3p3.n7373 vdd3p3.n7372 92.5
R4865 vdd3p3.n7385 vdd3p3.n7384 92.5
R4866 vdd3p3.n8037 vdd3p3.n8036 92.5
R4867 vdd3p3.n8042 vdd3p3.n8041 92.5
R4868 vdd3p3.n8048 vdd3p3.n8047 92.5
R4869 vdd3p3.n8054 vdd3p3.n8053 92.5
R4870 vdd3p3.n8060 vdd3p3.n8059 92.5
R4871 vdd3p3.n8066 vdd3p3.n8065 92.5
R4872 vdd3p3.n8072 vdd3p3.n8071 92.5
R4873 vdd3p3.n8078 vdd3p3.n8077 92.5
R4874 vdd3p3.n8084 vdd3p3.n8083 92.5
R4875 vdd3p3.n8090 vdd3p3.n8089 92.5
R4876 vdd3p3.n8092 vdd3p3.n8091 92.5
R4877 vdd3p3.n8098 vdd3p3.n8097 92.5
R4878 vdd3p3.n8104 vdd3p3.n8103 92.5
R4879 vdd3p3.n8110 vdd3p3.n8109 92.5
R4880 vdd3p3.n8116 vdd3p3.n8115 92.5
R4881 vdd3p3.n8122 vdd3p3.n8121 92.5
R4882 vdd3p3.n8128 vdd3p3.n8127 92.5
R4883 vdd3p3.n8136 vdd3p3.n8135 92.5
R4884 vdd3p3.n8142 vdd3p3.n8141 92.5
R4885 vdd3p3.n8147 vdd3p3.n8146 92.5
R4886 vdd3p3.n8153 vdd3p3.n8152 92.5
R4887 vdd3p3.n8159 vdd3p3.n8158 92.5
R4888 vdd3p3.n8165 vdd3p3.n8164 92.5
R4889 vdd3p3.n8171 vdd3p3.n8170 92.5
R4890 vdd3p3.n8177 vdd3p3.n8176 92.5
R4891 vdd3p3.n8183 vdd3p3.n8182 92.5
R4892 vdd3p3.n8189 vdd3p3.n8188 92.5
R4893 vdd3p3.n8195 vdd3p3.n8194 92.5
R4894 vdd3p3.n8197 vdd3p3.n8196 92.5
R4895 vdd3p3.n8203 vdd3p3.n8202 92.5
R4896 vdd3p3.n8209 vdd3p3.n8208 92.5
R4897 vdd3p3.n8215 vdd3p3.n8214 92.5
R4898 vdd3p3.n8221 vdd3p3.n8220 92.5
R4899 vdd3p3.n8227 vdd3p3.n8226 92.5
R4900 vdd3p3.n8233 vdd3p3.n8232 92.5
R4901 vdd3p3.n8241 vdd3p3.n8240 92.5
R4902 vdd3p3.n8247 vdd3p3.n8246 92.5
R4903 vdd3p3.n8252 vdd3p3.n8251 92.5
R4904 vdd3p3.n8258 vdd3p3.n8257 92.5
R4905 vdd3p3.n8264 vdd3p3.n8263 92.5
R4906 vdd3p3.n8270 vdd3p3.n8269 92.5
R4907 vdd3p3.n8276 vdd3p3.n8275 92.5
R4908 vdd3p3.n8282 vdd3p3.n8281 92.5
R4909 vdd3p3.n8288 vdd3p3.n8287 92.5
R4910 vdd3p3.n8294 vdd3p3.n8293 92.5
R4911 vdd3p3.n8300 vdd3p3.n8299 92.5
R4912 vdd3p3.n8305 vdd3p3.n8304 92.5
R4913 vdd3p3.n8304 vdd3p3.n8303 92.5
R4914 vdd3p3.n8315 vdd3p3.n8314 92.5
R4915 vdd3p3.n8314 vdd3p3.n8313 92.5
R4916 vdd3p3.n8325 vdd3p3.n8324 92.5
R4917 vdd3p3.n8324 vdd3p3.n8323 92.5
R4918 vdd3p3.n8335 vdd3p3.n8334 92.5
R4919 vdd3p3.n8334 vdd3p3.n8333 92.5
R4920 vdd3p3.n8345 vdd3p3.n8344 92.5
R4921 vdd3p3.n8344 vdd3p3.n8343 92.5
R4922 vdd3p3.n8354 vdd3p3.n8353 92.5
R4923 vdd3p3.n8353 vdd3p3.n8352 92.5
R4924 vdd3p3.n8363 vdd3p3.n8362 92.5
R4925 vdd3p3.n8362 vdd3p3.n8361 92.5
R4926 vdd3p3.n8375 vdd3p3.n8374 92.5
R4927 vdd3p3.n8374 vdd3p3.n8373 92.5
R4928 vdd3p3.n8384 vdd3p3.n8383 92.5
R4929 vdd3p3.n8383 vdd3p3.n8382 92.5
R4930 vdd3p3.n8392 vdd3p3.n8391 92.5
R4931 vdd3p3.n8391 vdd3p3.n8390 92.5
R4932 vdd3p3.n8401 vdd3p3.n8400 92.5
R4933 vdd3p3.n8400 vdd3p3.n8399 92.5
R4934 vdd3p3.n8410 vdd3p3.n8409 92.5
R4935 vdd3p3.n8409 vdd3p3.n8408 92.5
R4936 vdd3p3.n8418 vdd3p3.n8417 92.5
R4937 vdd3p3.n8417 vdd3p3.n8416 92.5
R4938 vdd3p3.n8426 vdd3p3.n8425 92.5
R4939 vdd3p3.n8425 vdd3p3.n8424 92.5
R4940 vdd3p3.n8432 vdd3p3.n8431 92.5
R4941 vdd3p3.n8040 vdd3p3.n8039 92.5
R4942 vdd3p3.n8046 vdd3p3.n8045 92.5
R4943 vdd3p3.n8052 vdd3p3.n8051 92.5
R4944 vdd3p3.n8058 vdd3p3.n8057 92.5
R4945 vdd3p3.n8064 vdd3p3.n8063 92.5
R4946 vdd3p3.n8070 vdd3p3.n8069 92.5
R4947 vdd3p3.n8076 vdd3p3.n8075 92.5
R4948 vdd3p3.n8080 vdd3p3.n8079 92.5
R4949 vdd3p3.n8086 vdd3p3.n8085 92.5
R4950 vdd3p3.n8094 vdd3p3.n8093 92.5
R4951 vdd3p3.n8100 vdd3p3.n8099 92.5
R4952 vdd3p3.n8106 vdd3p3.n8105 92.5
R4953 vdd3p3.n8112 vdd3p3.n8111 92.5
R4954 vdd3p3.n8118 vdd3p3.n8117 92.5
R4955 vdd3p3.n8124 vdd3p3.n8123 92.5
R4956 vdd3p3.n8130 vdd3p3.n8129 92.5
R4957 vdd3p3.n8134 vdd3p3.n8133 92.5
R4958 vdd3p3.n8140 vdd3p3.n8139 92.5
R4959 vdd3p3.n8145 vdd3p3.n8144 92.5
R4960 vdd3p3.n8151 vdd3p3.n8150 92.5
R4961 vdd3p3.n8157 vdd3p3.n8156 92.5
R4962 vdd3p3.n8163 vdd3p3.n8162 92.5
R4963 vdd3p3.n8169 vdd3p3.n8168 92.5
R4964 vdd3p3.n8175 vdd3p3.n8174 92.5
R4965 vdd3p3.n8181 vdd3p3.n8180 92.5
R4966 vdd3p3.n8185 vdd3p3.n8184 92.5
R4967 vdd3p3.n8191 vdd3p3.n8190 92.5
R4968 vdd3p3.n8199 vdd3p3.n8198 92.5
R4969 vdd3p3.n8205 vdd3p3.n8204 92.5
R4970 vdd3p3.n8211 vdd3p3.n8210 92.5
R4971 vdd3p3.n8217 vdd3p3.n8216 92.5
R4972 vdd3p3.n8223 vdd3p3.n8222 92.5
R4973 vdd3p3.n8229 vdd3p3.n8228 92.5
R4974 vdd3p3.n8235 vdd3p3.n8234 92.5
R4975 vdd3p3.n8239 vdd3p3.n8238 92.5
R4976 vdd3p3.n8245 vdd3p3.n8244 92.5
R4977 vdd3p3.n8250 vdd3p3.n8249 92.5
R4978 vdd3p3.n8256 vdd3p3.n8255 92.5
R4979 vdd3p3.n8262 vdd3p3.n8261 92.5
R4980 vdd3p3.n8268 vdd3p3.n8267 92.5
R4981 vdd3p3.n8274 vdd3p3.n8273 92.5
R4982 vdd3p3.n8280 vdd3p3.n8279 92.5
R4983 vdd3p3.n8286 vdd3p3.n8285 92.5
R4984 vdd3p3.n8290 vdd3p3.n8289 92.5
R4985 vdd3p3.n8296 vdd3p3.n8295 92.5
R4986 vdd3p3.n8308 vdd3p3.n8307 92.5
R4987 vdd3p3.n8307 vdd3p3.n8306 92.5
R4988 vdd3p3.n8318 vdd3p3.n8317 92.5
R4989 vdd3p3.n8317 vdd3p3.n8316 92.5
R4990 vdd3p3.n8328 vdd3p3.n8327 92.5
R4991 vdd3p3.n8327 vdd3p3.n8326 92.5
R4992 vdd3p3.n8338 vdd3p3.n8337 92.5
R4993 vdd3p3.n8337 vdd3p3.n8336 92.5
R4994 vdd3p3.n8348 vdd3p3.n8347 92.5
R4995 vdd3p3.n8347 vdd3p3.n8346 92.5
R4996 vdd3p3.n8357 vdd3p3.n8356 92.5
R4997 vdd3p3.n8356 vdd3p3.n8355 92.5
R4998 vdd3p3.n8366 vdd3p3.n8365 92.5
R4999 vdd3p3.n8365 vdd3p3.n8364 92.5
R5000 vdd3p3.n8371 vdd3p3.n8370 92.5
R5001 vdd3p3.n8370 vdd3p3.n8369 92.5
R5002 vdd3p3.n8380 vdd3p3.n8379 92.5
R5003 vdd3p3.n8379 vdd3p3.n8378 92.5
R5004 vdd3p3.n8388 vdd3p3.n8387 92.5
R5005 vdd3p3.n8387 vdd3p3.n8386 92.5
R5006 vdd3p3.n8397 vdd3p3.n8396 92.5
R5007 vdd3p3.n8396 vdd3p3.n8395 92.5
R5008 vdd3p3.n8406 vdd3p3.n8405 92.5
R5009 vdd3p3.n8405 vdd3p3.n8404 92.5
R5010 vdd3p3.n8415 vdd3p3.n8414 92.5
R5011 vdd3p3.n8414 vdd3p3.n8413 92.5
R5012 vdd3p3.n8423 vdd3p3.n8422 92.5
R5013 vdd3p3.n8422 vdd3p3.n8421 92.5
R5014 vdd3p3.n8430 vdd3p3.n8429 92.5
R5015 vdd3p3.n8461 vdd3p3.n8460 92.5
R5016 vdd3p3.n8457 vdd3p3.n8456 92.5
R5017 vdd3p3.n41 vdd3p3.t141 91.871
R5018 vdd3p3.n901 vdd3p3.t167 91.871
R5019 vdd3p3.n1732 vdd3p3.t84 91.871
R5020 vdd3p3.n2592 vdd3p3.t88 91.871
R5021 vdd3p3.n55 vdd3p3.t115 84.467
R5022 vdd3p3.n884 vdd3p3.t98 84.467
R5023 vdd3p3.n1746 vdd3p3.t28 84.467
R5024 vdd3p3.n2575 vdd3p3.t126 84.467
R5025 vdd3p3.n41 vdd3p3.n40 83.1
R5026 vdd3p3.n901 vdd3p3.n900 83.1
R5027 vdd3p3.n1732 vdd3p3.n1731 83.1
R5028 vdd3p3.n2592 vdd3p3.n2591 83.1
R5029 vdd3p3.n30 vdd3p3.t122 78.557
R5030 vdd3p3.t157 vdd3p3.n849 78.557
R5031 vdd3p3.n1721 vdd3p3.t13 78.557
R5032 vdd3p3.t79 vdd3p3.n2540 78.557
R5033 vdd3p3.n2886 vdd3p3.n2885 78.412
R5034 vdd3p3.n3013 vdd3p3.n2755 78.412
R5035 vdd3p3.n2040 vdd3p3.n2039 78.412
R5036 vdd3p3.n2167 vdd3p3.n1909 78.412
R5037 vdd3p3.n1195 vdd3p3.n1194 78.412
R5038 vdd3p3.n1322 vdd3p3.n1064 78.412
R5039 vdd3p3.n349 vdd3p3.n348 78.412
R5040 vdd3p3.n476 vdd3p3.n218 78.412
R5041 vdd3p3.n4722 vdd3p3.t142 75.59
R5042 vdd3p3.n4722 vdd3p3.t26 75.59
R5043 vdd3p3.n4719 vdd3p3.n4718 74.6
R5044 vdd3p3.n2672 vdd3p3.n2671 72.09
R5045 vdd3p3.n2856 vdd3p3.n2672 72.09
R5046 vdd3p3.n2980 vdd3p3.n2789 72.09
R5047 vdd3p3.n3188 vdd3p3.n2756 72.09
R5048 vdd3p3.n3188 vdd3p3.n2757 72.09
R5049 vdd3p3.n3188 vdd3p3.n2758 72.09
R5050 vdd3p3.n3188 vdd3p3.n2759 72.09
R5051 vdd3p3.n3188 vdd3p3.n2760 72.09
R5052 vdd3p3.n3188 vdd3p3.n2761 72.09
R5053 vdd3p3.n3188 vdd3p3.n2762 72.09
R5054 vdd3p3.n3188 vdd3p3.n2763 72.09
R5055 vdd3p3.n3188 vdd3p3.n2768 72.09
R5056 vdd3p3.n3188 vdd3p3.n2769 72.09
R5057 vdd3p3.n3188 vdd3p3.n2770 72.09
R5058 vdd3p3.n3188 vdd3p3.n2771 72.09
R5059 vdd3p3.n3188 vdd3p3.n2772 72.09
R5060 vdd3p3.n1826 vdd3p3.n1825 72.09
R5061 vdd3p3.n2010 vdd3p3.n1826 72.09
R5062 vdd3p3.n2134 vdd3p3.n1943 72.09
R5063 vdd3p3.n2342 vdd3p3.n1910 72.09
R5064 vdd3p3.n2342 vdd3p3.n1911 72.09
R5065 vdd3p3.n2342 vdd3p3.n1912 72.09
R5066 vdd3p3.n2342 vdd3p3.n1913 72.09
R5067 vdd3p3.n2342 vdd3p3.n1914 72.09
R5068 vdd3p3.n2342 vdd3p3.n1915 72.09
R5069 vdd3p3.n2342 vdd3p3.n1916 72.09
R5070 vdd3p3.n2342 vdd3p3.n1917 72.09
R5071 vdd3p3.n2342 vdd3p3.n1922 72.09
R5072 vdd3p3.n2342 vdd3p3.n1923 72.09
R5073 vdd3p3.n2342 vdd3p3.n1924 72.09
R5074 vdd3p3.n2342 vdd3p3.n1925 72.09
R5075 vdd3p3.n2342 vdd3p3.n1926 72.09
R5076 vdd3p3.n981 vdd3p3.n980 72.09
R5077 vdd3p3.n1165 vdd3p3.n981 72.09
R5078 vdd3p3.n1289 vdd3p3.n1098 72.09
R5079 vdd3p3.n1497 vdd3p3.n1065 72.09
R5080 vdd3p3.n1497 vdd3p3.n1066 72.09
R5081 vdd3p3.n1497 vdd3p3.n1067 72.09
R5082 vdd3p3.n1497 vdd3p3.n1068 72.09
R5083 vdd3p3.n1497 vdd3p3.n1069 72.09
R5084 vdd3p3.n1497 vdd3p3.n1070 72.09
R5085 vdd3p3.n1497 vdd3p3.n1071 72.09
R5086 vdd3p3.n1497 vdd3p3.n1072 72.09
R5087 vdd3p3.n1497 vdd3p3.n1077 72.09
R5088 vdd3p3.n1497 vdd3p3.n1078 72.09
R5089 vdd3p3.n1497 vdd3p3.n1079 72.09
R5090 vdd3p3.n1497 vdd3p3.n1080 72.09
R5091 vdd3p3.n1497 vdd3p3.n1081 72.09
R5092 vdd3p3.n135 vdd3p3.n134 72.09
R5093 vdd3p3.n319 vdd3p3.n135 72.09
R5094 vdd3p3.n443 vdd3p3.n252 72.09
R5095 vdd3p3.n651 vdd3p3.n219 72.09
R5096 vdd3p3.n651 vdd3p3.n220 72.09
R5097 vdd3p3.n651 vdd3p3.n221 72.09
R5098 vdd3p3.n651 vdd3p3.n222 72.09
R5099 vdd3p3.n651 vdd3p3.n223 72.09
R5100 vdd3p3.n651 vdd3p3.n224 72.09
R5101 vdd3p3.n651 vdd3p3.n225 72.09
R5102 vdd3p3.n651 vdd3p3.n226 72.09
R5103 vdd3p3.n651 vdd3p3.n231 72.09
R5104 vdd3p3.n651 vdd3p3.n232 72.09
R5105 vdd3p3.n651 vdd3p3.n233 72.09
R5106 vdd3p3.n651 vdd3p3.n234 72.09
R5107 vdd3p3.n651 vdd3p3.n235 72.09
R5108 vdd3p3.n3955 vdd3p3.n3920 72.09
R5109 vdd3p3.n3955 vdd3p3.n3921 72.09
R5110 vdd3p3.n3955 vdd3p3.n3922 72.09
R5111 vdd3p3.n3955 vdd3p3.n3923 72.09
R5112 vdd3p3.n3955 vdd3p3.n3924 72.09
R5113 vdd3p3.n3955 vdd3p3.n3925 72.09
R5114 vdd3p3.n3955 vdd3p3.n3926 72.09
R5115 vdd3p3.n3955 vdd3p3.n3927 72.09
R5116 vdd3p3.n3955 vdd3p3.n3928 72.09
R5117 vdd3p3.n3955 vdd3p3.n3929 72.09
R5118 vdd3p3.n3955 vdd3p3.n3930 72.09
R5119 vdd3p3.n3955 vdd3p3.n3931 72.09
R5120 vdd3p3.n3955 vdd3p3.n3932 72.09
R5121 vdd3p3.n3955 vdd3p3.n3933 72.09
R5122 vdd3p3.n3955 vdd3p3.n3934 72.09
R5123 vdd3p3.n3955 vdd3p3.n3935 72.09
R5124 vdd3p3.n3955 vdd3p3.n3936 72.09
R5125 vdd3p3.n3955 vdd3p3.n3937 72.09
R5126 vdd3p3.n3955 vdd3p3.n3938 72.09
R5127 vdd3p3.n3955 vdd3p3.n3939 72.09
R5128 vdd3p3.n3955 vdd3p3.n3940 72.09
R5129 vdd3p3.n3955 vdd3p3.n3941 72.09
R5130 vdd3p3.n3955 vdd3p3.n3942 72.09
R5131 vdd3p3.n3955 vdd3p3.n3943 72.09
R5132 vdd3p3.n3955 vdd3p3.n3944 72.09
R5133 vdd3p3.n3955 vdd3p3.n3945 72.09
R5134 vdd3p3.n3955 vdd3p3.n3946 72.09
R5135 vdd3p3.n3955 vdd3p3.n3947 72.09
R5136 vdd3p3.n3955 vdd3p3.n3948 72.09
R5137 vdd3p3.n3955 vdd3p3.n3949 72.09
R5138 vdd3p3.n3955 vdd3p3.n3950 72.09
R5139 vdd3p3.n3955 vdd3p3.n3951 72.09
R5140 vdd3p3.n3955 vdd3p3.n3952 72.09
R5141 vdd3p3.n3955 vdd3p3.n3953 72.09
R5142 vdd3p3.n3177 vdd3p3.n3023 71.153
R5143 vdd3p3.n2683 vdd3p3.n2666 71.153
R5144 vdd3p3.n2331 vdd3p3.n2177 71.153
R5145 vdd3p3.n1837 vdd3p3.n1820 71.153
R5146 vdd3p3.n1486 vdd3p3.n1332 71.153
R5147 vdd3p3.n992 vdd3p3.n975 71.153
R5148 vdd3p3.n640 vdd3p3.n486 71.153
R5149 vdd3p3.n146 vdd3p3.n129 71.153
R5150 vdd3p3.n5283 vdd3p3.n5282 70.536
R5151 vdd3p3.n5286 vdd3p3.n5285 70.536
R5152 vdd3p3.n5289 vdd3p3.n5288 70.536
R5153 vdd3p3.n5292 vdd3p3.n5291 70.536
R5154 vdd3p3.n5295 vdd3p3.n5294 70.536
R5155 vdd3p3.n5299 vdd3p3.n5297 70.536
R5156 vdd3p3.n5163 vdd3p3.n5162 70.536
R5157 vdd3p3.n5166 vdd3p3.n5165 70.536
R5158 vdd3p3.n5169 vdd3p3.n5168 70.536
R5159 vdd3p3.n5172 vdd3p3.n5171 70.536
R5160 vdd3p3.n5175 vdd3p3.n5174 70.536
R5161 vdd3p3.n5178 vdd3p3.n5177 70.536
R5162 vdd3p3.n5264 vdd3p3.n5262 70.536
R5163 vdd3p3.n5206 vdd3p3.n5205 70.536
R5164 vdd3p3.n5209 vdd3p3.n5208 70.536
R5165 vdd3p3.n5212 vdd3p3.n5211 70.536
R5166 vdd3p3.n5215 vdd3p3.n5214 70.536
R5167 vdd3p3.n5218 vdd3p3.n5217 70.536
R5168 vdd3p3.n5221 vdd3p3.n5220 70.536
R5169 vdd3p3.n5224 vdd3p3.n5223 70.536
R5170 vdd3p3.n5227 vdd3p3.n5226 70.536
R5171 vdd3p3.n5230 vdd3p3.n5229 70.536
R5172 vdd3p3.n5233 vdd3p3.n5232 70.536
R5173 vdd3p3.n5236 vdd3p3.n5235 70.536
R5174 vdd3p3.n5239 vdd3p3.n5238 70.536
R5175 vdd3p3.n5242 vdd3p3.n5241 70.536
R5176 vdd3p3.n5245 vdd3p3.n5244 70.536
R5177 vdd3p3.n5248 vdd3p3.n5247 70.536
R5178 vdd3p3.n5251 vdd3p3.n5250 70.536
R5179 vdd3p3.n5254 vdd3p3.n5253 70.536
R5180 vdd3p3.n5257 vdd3p3.n5256 70.536
R5181 vdd3p3.n5260 vdd3p3.n5259 70.536
R5182 vdd3p3.n5264 vdd3p3.n5263 70.536
R5183 vdd3p3.n5304 vdd3p3.n5303 70.536
R5184 vdd3p3.n5307 vdd3p3.n5306 70.536
R5185 vdd3p3.n5310 vdd3p3.n5309 70.536
R5186 vdd3p3.n5313 vdd3p3.n5312 70.536
R5187 vdd3p3.n5316 vdd3p3.n5315 70.536
R5188 vdd3p3.n5319 vdd3p3.n5318 70.536
R5189 vdd3p3.n5299 vdd3p3.n5298 70.536
R5190 vdd3p3.n5322 vdd3p3.n5321 70.536
R5191 vdd3p3.n5325 vdd3p3.n5324 70.536
R5192 vdd3p3.n5328 vdd3p3.n5327 70.536
R5193 vdd3p3.n5331 vdd3p3.n5330 70.536
R5194 vdd3p3.n5334 vdd3p3.n5333 70.536
R5195 vdd3p3.n2846 vdd3p3.n2641 67.954
R5196 vdd3p3.n2874 vdd3p3.n2641 67.954
R5197 vdd3p3.n2655 vdd3p3.n2629 67.954
R5198 vdd3p3.n2645 vdd3p3.n2629 67.954
R5199 vdd3p3.n2650 vdd3p3.n2629 67.954
R5200 vdd3p3.n3132 vdd3p3.n3049 67.954
R5201 vdd3p3.n3080 vdd3p3.n3049 67.954
R5202 vdd3p3.n3137 vdd3p3.n3049 67.954
R5203 vdd3p3.n2000 vdd3p3.n1795 67.954
R5204 vdd3p3.n2028 vdd3p3.n1795 67.954
R5205 vdd3p3.n1809 vdd3p3.n1783 67.954
R5206 vdd3p3.n1799 vdd3p3.n1783 67.954
R5207 vdd3p3.n1804 vdd3p3.n1783 67.954
R5208 vdd3p3.n2286 vdd3p3.n2203 67.954
R5209 vdd3p3.n2234 vdd3p3.n2203 67.954
R5210 vdd3p3.n2291 vdd3p3.n2203 67.954
R5211 vdd3p3.n1155 vdd3p3.n950 67.954
R5212 vdd3p3.n1183 vdd3p3.n950 67.954
R5213 vdd3p3.n964 vdd3p3.n938 67.954
R5214 vdd3p3.n954 vdd3p3.n938 67.954
R5215 vdd3p3.n959 vdd3p3.n938 67.954
R5216 vdd3p3.n1441 vdd3p3.n1358 67.954
R5217 vdd3p3.n1389 vdd3p3.n1358 67.954
R5218 vdd3p3.n1446 vdd3p3.n1358 67.954
R5219 vdd3p3.n309 vdd3p3.n104 67.954
R5220 vdd3p3.n337 vdd3p3.n104 67.954
R5221 vdd3p3.n118 vdd3p3.n92 67.954
R5222 vdd3p3.n108 vdd3p3.n92 67.954
R5223 vdd3p3.n113 vdd3p3.n92 67.954
R5224 vdd3p3.n595 vdd3p3.n512 67.954
R5225 vdd3p3.n543 vdd3p3.n512 67.954
R5226 vdd3p3.n600 vdd3p3.n512 67.954
R5227 vdd3p3.n6393 vdd3p3.n6392 66.885
R5228 vdd3p3.n7940 vdd3p3.n7939 66.885
R5229 vdd3p3.n4255 vdd3p3.t38 60.25
R5230 vdd3p3.n4271 vdd3p3.t67 60.25
R5231 vdd3p3.n4575 vdd3p3.t62 60.25
R5232 vdd3p3.n4591 vdd3p3.t55 60.25
R5233 vdd3p3.n3532 vdd3p3.t33 60.25
R5234 vdd3p3.n3517 vdd3p3.t43 60.25
R5235 vdd3p3.n3701 vdd3p3.t47 60.25
R5236 vdd3p3.n3629 vdd3p3.t50 60.25
R5237 vdd3p3.n4766 vdd3p3.t71 60.25
R5238 vdd3p3.n4907 vdd3p3.t59 60.25
R5239 vdd3p3.n2875 vdd3p3.n2845 60.14
R5240 vdd3p3.n2649 vdd3p3.n2648 60.14
R5241 vdd3p3.n3139 vdd3p3.n3138 60.14
R5242 vdd3p3.n2029 vdd3p3.n1999 60.14
R5243 vdd3p3.n1803 vdd3p3.n1802 60.14
R5244 vdd3p3.n2293 vdd3p3.n2292 60.14
R5245 vdd3p3.n1184 vdd3p3.n1154 60.14
R5246 vdd3p3.n958 vdd3p3.n957 60.14
R5247 vdd3p3.n1448 vdd3p3.n1447 60.14
R5248 vdd3p3.n338 vdd3p3.n308 60.14
R5249 vdd3p3.n112 vdd3p3.n111 60.14
R5250 vdd3p3.n602 vdd3p3.n601 60.14
R5251 vdd3p3.n2852 vdd3p3.n2851 60.139
R5252 vdd3p3.n2657 vdd3p3.n2656 60.139
R5253 vdd3p3.n3131 vdd3p3.n3130 60.139
R5254 vdd3p3.n2006 vdd3p3.n2005 60.139
R5255 vdd3p3.n1811 vdd3p3.n1810 60.139
R5256 vdd3p3.n2285 vdd3p3.n2284 60.139
R5257 vdd3p3.n1161 vdd3p3.n1160 60.139
R5258 vdd3p3.n966 vdd3p3.n965 60.139
R5259 vdd3p3.n1440 vdd3p3.n1439 60.139
R5260 vdd3p3.n315 vdd3p3.n314 60.139
R5261 vdd3p3.n120 vdd3p3.n119 60.139
R5262 vdd3p3.n594 vdd3p3.n593 60.139
R5263 vdd3p3.n3572 vdd3p3.n3571 59.275
R5264 vdd3p3.n8455 vdd3p3.n8452 57.233
R5265 vdd3p3.n8455 vdd3p3.n8453 57.233
R5266 vdd3p3.n8455 vdd3p3.n8454 57.233
R5267 vdd3p3.n3074 vdd3p3.n3073 55.128
R5268 vdd3p3.n2228 vdd3p3.n2227 55.128
R5269 vdd3p3.n1383 vdd3p3.n1382 55.128
R5270 vdd3p3.n537 vdd3p3.n536 55.128
R5271 vdd3p3.n7938 vdd3p3.n7937 54.625
R5272 vdd3p3.n4197 vdd3p3.n4196 52.689
R5273 vdd3p3.n5049 vdd3p3.n5048 52.689
R5274 vdd3p3.n4956 vdd3p3.n4955 52.689
R5275 vdd3p3.n8503 vdd3p3.n8502 52.689
R5276 vdd3p3.n8847 vdd3p3.n8846 52.689
R5277 vdd3p3.n8758 vdd3p3.n8757 52.689
R5278 vdd3p3.n7954 vdd3p3.n7953 51.067
R5279 vdd3p3.n7967 vdd3p3.n7966 51.067
R5280 vdd3p3.n7983 vdd3p3.n7982 51.066
R5281 vdd3p3.n7997 vdd3p3.n7996 51.066
R5282 vdd3p3.n8011 vdd3p3.n8010 51.066
R5283 vdd3p3.n8030 vdd3p3.n8029 51.066
R5284 vdd3p3.n7508 vdd3p3.n7507 51.066
R5285 vdd3p3.n7515 vdd3p3.n7513 51.066
R5286 vdd3p3.n7518 vdd3p3.n7516 51.066
R5287 vdd3p3.n7521 vdd3p3.n7519 51.066
R5288 vdd3p3.n7521 vdd3p3.n7520 51.066
R5289 vdd3p3.n7518 vdd3p3.n7517 51.066
R5290 vdd3p3.n7515 vdd3p3.n7514 51.066
R5291 vdd3p3.n2859 vdd3p3.n2858 50.7
R5292 vdd3p3.n3187 vdd3p3.n2773 50.7
R5293 vdd3p3.n3095 vdd3p3.n2764 50.7
R5294 vdd3p3.n2013 vdd3p3.n2012 50.7
R5295 vdd3p3.n2341 vdd3p3.n1927 50.7
R5296 vdd3p3.n2249 vdd3p3.n1918 50.7
R5297 vdd3p3.n1168 vdd3p3.n1167 50.7
R5298 vdd3p3.n1496 vdd3p3.n1082 50.7
R5299 vdd3p3.n1404 vdd3p3.n1073 50.7
R5300 vdd3p3.n322 vdd3p3.n321 50.7
R5301 vdd3p3.n650 vdd3p3.n236 50.7
R5302 vdd3p3.n558 vdd3p3.n227 50.7
R5303 vdd3p3.n3339 vdd3p3.n3338 50.699
R5304 vdd3p3.n2882 vdd3p3.n2839 50.699
R5305 vdd3p3.n2883 vdd3p3.n2882 50.699
R5306 vdd3p3.n2981 vdd3p3.n2977 50.699
R5307 vdd3p3.n2979 vdd3p3.n2978 50.699
R5308 vdd3p3.n3189 vdd3p3.n2754 50.699
R5309 vdd3p3.n3169 vdd3p3.n2767 50.699
R5310 vdd3p3.n2493 vdd3p3.n2492 50.699
R5311 vdd3p3.n2036 vdd3p3.n1993 50.699
R5312 vdd3p3.n2037 vdd3p3.n2036 50.699
R5313 vdd3p3.n2135 vdd3p3.n2131 50.699
R5314 vdd3p3.n2133 vdd3p3.n2132 50.699
R5315 vdd3p3.n2343 vdd3p3.n1908 50.699
R5316 vdd3p3.n2323 vdd3p3.n1921 50.699
R5317 vdd3p3.n1648 vdd3p3.n1647 50.699
R5318 vdd3p3.n1191 vdd3p3.n1148 50.699
R5319 vdd3p3.n1192 vdd3p3.n1191 50.699
R5320 vdd3p3.n1290 vdd3p3.n1286 50.699
R5321 vdd3p3.n1288 vdd3p3.n1287 50.699
R5322 vdd3p3.n1498 vdd3p3.n1063 50.699
R5323 vdd3p3.n1478 vdd3p3.n1076 50.699
R5324 vdd3p3.n802 vdd3p3.n801 50.699
R5325 vdd3p3.n345 vdd3p3.n302 50.699
R5326 vdd3p3.n346 vdd3p3.n345 50.699
R5327 vdd3p3.n444 vdd3p3.n440 50.699
R5328 vdd3p3.n442 vdd3p3.n441 50.699
R5329 vdd3p3.n652 vdd3p3.n217 50.699
R5330 vdd3p3.n632 vdd3p3.n230 50.699
R5331 vdd3p3.n8458 vdd3p3.n8447 50.699
R5332 vdd3p3.n3137 vdd3p3.n3136 49.094
R5333 vdd3p3.n3133 vdd3p3.n3080 49.094
R5334 vdd3p3.n3132 vdd3p3.n3131 49.094
R5335 vdd3p3.n2874 vdd3p3.n2873 49.094
R5336 vdd3p3.n2851 vdd3p3.n2846 49.094
R5337 vdd3p3.n2873 vdd3p3.n2846 49.094
R5338 vdd3p3.n2875 vdd3p3.n2874 49.094
R5339 vdd3p3.n2651 vdd3p3.n2650 49.094
R5340 vdd3p3.n2654 vdd3p3.n2645 49.094
R5341 vdd3p3.n2656 vdd3p3.n2655 49.094
R5342 vdd3p3.n2655 vdd3p3.n2654 49.094
R5343 vdd3p3.n2651 vdd3p3.n2645 49.094
R5344 vdd3p3.n2650 vdd3p3.n2649 49.094
R5345 vdd3p3.n3133 vdd3p3.n3132 49.094
R5346 vdd3p3.n3136 vdd3p3.n3080 49.094
R5347 vdd3p3.n3138 vdd3p3.n3137 49.094
R5348 vdd3p3.n2291 vdd3p3.n2290 49.094
R5349 vdd3p3.n2287 vdd3p3.n2234 49.094
R5350 vdd3p3.n2286 vdd3p3.n2285 49.094
R5351 vdd3p3.n2028 vdd3p3.n2027 49.094
R5352 vdd3p3.n2005 vdd3p3.n2000 49.094
R5353 vdd3p3.n2027 vdd3p3.n2000 49.094
R5354 vdd3p3.n2029 vdd3p3.n2028 49.094
R5355 vdd3p3.n1805 vdd3p3.n1804 49.094
R5356 vdd3p3.n1808 vdd3p3.n1799 49.094
R5357 vdd3p3.n1810 vdd3p3.n1809 49.094
R5358 vdd3p3.n1809 vdd3p3.n1808 49.094
R5359 vdd3p3.n1805 vdd3p3.n1799 49.094
R5360 vdd3p3.n1804 vdd3p3.n1803 49.094
R5361 vdd3p3.n2287 vdd3p3.n2286 49.094
R5362 vdd3p3.n2290 vdd3p3.n2234 49.094
R5363 vdd3p3.n2292 vdd3p3.n2291 49.094
R5364 vdd3p3.n1446 vdd3p3.n1445 49.094
R5365 vdd3p3.n1442 vdd3p3.n1389 49.094
R5366 vdd3p3.n1441 vdd3p3.n1440 49.094
R5367 vdd3p3.n1183 vdd3p3.n1182 49.094
R5368 vdd3p3.n1160 vdd3p3.n1155 49.094
R5369 vdd3p3.n1182 vdd3p3.n1155 49.094
R5370 vdd3p3.n1184 vdd3p3.n1183 49.094
R5371 vdd3p3.n960 vdd3p3.n959 49.094
R5372 vdd3p3.n963 vdd3p3.n954 49.094
R5373 vdd3p3.n965 vdd3p3.n964 49.094
R5374 vdd3p3.n964 vdd3p3.n963 49.094
R5375 vdd3p3.n960 vdd3p3.n954 49.094
R5376 vdd3p3.n959 vdd3p3.n958 49.094
R5377 vdd3p3.n1442 vdd3p3.n1441 49.094
R5378 vdd3p3.n1445 vdd3p3.n1389 49.094
R5379 vdd3p3.n1447 vdd3p3.n1446 49.094
R5380 vdd3p3.n600 vdd3p3.n599 49.094
R5381 vdd3p3.n596 vdd3p3.n543 49.094
R5382 vdd3p3.n595 vdd3p3.n594 49.094
R5383 vdd3p3.n337 vdd3p3.n336 49.094
R5384 vdd3p3.n314 vdd3p3.n309 49.094
R5385 vdd3p3.n336 vdd3p3.n309 49.094
R5386 vdd3p3.n338 vdd3p3.n337 49.094
R5387 vdd3p3.n114 vdd3p3.n113 49.094
R5388 vdd3p3.n117 vdd3p3.n108 49.094
R5389 vdd3p3.n119 vdd3p3.n118 49.094
R5390 vdd3p3.n118 vdd3p3.n117 49.094
R5391 vdd3p3.n114 vdd3p3.n108 49.094
R5392 vdd3p3.n113 vdd3p3.n112 49.094
R5393 vdd3p3.n596 vdd3p3.n595 49.094
R5394 vdd3p3.n599 vdd3p3.n543 49.094
R5395 vdd3p3.n601 vdd3p3.n600 49.094
R5396 vdd3p3.n3901 vdd3p3.n3900 49.083
R5397 vdd3p3.n3903 vdd3p3.n3902 49.083
R5398 vdd3p3.n3908 vdd3p3.n3907 49.083
R5399 vdd3p3.n3906 vdd3p3.n3905 49.083
R5400 vdd3p3.n3385 vdd3p3.n3384 48.36
R5401 vdd3p3.n3350 vdd3p3.n2640 48.076
R5402 vdd3p3.n2504 vdd3p3.n1794 48.076
R5403 vdd3p3.n1659 vdd3p3.n949 48.076
R5404 vdd3p3.n813 vdd3p3.n103 48.076
R5405 vdd3p3.n5194 vdd3p3.n5192 46.418
R5406 vdd3p3.n4208 vdd3p3.n4207 46.103
R5407 vdd3p3.n5060 vdd3p3.n5059 46.103
R5408 vdd3p3.n3485 vdd3p3.n3484 46.103
R5409 vdd3p3.n4967 vdd3p3.n4966 46.103
R5410 vdd3p3.n8514 vdd3p3.n8513 46.103
R5411 vdd3p3.n8858 vdd3p3.n8857 46.103
R5412 vdd3p3.n8769 vdd3p3.n8768 46.103
R5413 vdd3p3.n4242 vdd3p3.n4241 44.967
R5414 vdd3p3.n5102 vdd3p3.n5101 44.967
R5415 vdd3p3.n2859 vdd3p3.n2672 44.768
R5416 vdd3p3.n3188 vdd3p3.n2764 44.768
R5417 vdd3p3.n2013 vdd3p3.n1826 44.768
R5418 vdd3p3.n2342 vdd3p3.n1918 44.768
R5419 vdd3p3.n1168 vdd3p3.n981 44.768
R5420 vdd3p3.n1497 vdd3p3.n1073 44.768
R5421 vdd3p3.n322 vdd3p3.n135 44.768
R5422 vdd3p3.n651 vdd3p3.n227 44.768
R5423 vdd3p3.n3188 vdd3p3.n3187 44.768
R5424 vdd3p3.n2342 vdd3p3.n2341 44.768
R5425 vdd3p3.n1497 vdd3p3.n1496 44.768
R5426 vdd3p3.n651 vdd3p3.n650 44.768
R5427 vdd3p3.n7020 vdd3p3.n7019 44.768
R5428 vdd3p3.n3955 vdd3p3.n3954 44.768
R5429 vdd3p3.n3338 vdd3p3.n2672 44.768
R5430 vdd3p3.n2839 vdd3p3.n2672 44.768
R5431 vdd3p3.n2883 vdd3p3.n2672 44.768
R5432 vdd3p3.n2977 vdd3p3.n2789 44.768
R5433 vdd3p3.n2978 vdd3p3.n2789 44.768
R5434 vdd3p3.n3189 vdd3p3.n3188 44.768
R5435 vdd3p3.n3188 vdd3p3.n2767 44.768
R5436 vdd3p3.n2492 vdd3p3.n1826 44.768
R5437 vdd3p3.n1993 vdd3p3.n1826 44.768
R5438 vdd3p3.n2037 vdd3p3.n1826 44.768
R5439 vdd3p3.n2131 vdd3p3.n1943 44.768
R5440 vdd3p3.n2132 vdd3p3.n1943 44.768
R5441 vdd3p3.n2343 vdd3p3.n2342 44.768
R5442 vdd3p3.n2342 vdd3p3.n1921 44.768
R5443 vdd3p3.n1647 vdd3p3.n981 44.768
R5444 vdd3p3.n1148 vdd3p3.n981 44.768
R5445 vdd3p3.n1192 vdd3p3.n981 44.768
R5446 vdd3p3.n1286 vdd3p3.n1098 44.768
R5447 vdd3p3.n1287 vdd3p3.n1098 44.768
R5448 vdd3p3.n1498 vdd3p3.n1497 44.768
R5449 vdd3p3.n1497 vdd3p3.n1076 44.768
R5450 vdd3p3.n801 vdd3p3.n135 44.768
R5451 vdd3p3.n302 vdd3p3.n135 44.768
R5452 vdd3p3.n346 vdd3p3.n135 44.768
R5453 vdd3p3.n440 vdd3p3.n252 44.768
R5454 vdd3p3.n441 vdd3p3.n252 44.768
R5455 vdd3p3.n652 vdd3p3.n651 44.768
R5456 vdd3p3.n651 vdd3p3.n230 44.768
R5457 vdd3p3.n8459 vdd3p3.n8439 44.768
R5458 vdd3p3.n7389 vdd3p3.n7388 44.768
R5459 vdd3p3.n3955 vdd3p3.n3919 44.768
R5460 vdd3p3.n8459 vdd3p3.n8458 44.768
R5461 vdd3p3.n3344 vdd3p3.n2666 43.589
R5462 vdd3p3.n2498 vdd3p3.n1820 43.589
R5463 vdd3p3.n1653 vdd3p3.n975 43.589
R5464 vdd3p3.n807 vdd3p3.n129 43.589
R5465 vdd3p3.n3282 vdd3p3.n3281 41.788
R5466 vdd3p3.n3225 vdd3p3.n3224 41.788
R5467 vdd3p3.n2436 vdd3p3.n2435 41.788
R5468 vdd3p3.n2379 vdd3p3.n2378 41.788
R5469 vdd3p3.n1591 vdd3p3.n1590 41.788
R5470 vdd3p3.n1534 vdd3p3.n1533 41.788
R5471 vdd3p3.n745 vdd3p3.n744 41.788
R5472 vdd3p3.n688 vdd3p3.n687 41.788
R5473 vdd3p3.n5337 vdd3p3.n5336 41.722
R5474 vdd3p3.n2845 vdd3p3.n2641 41.621
R5475 vdd3p3.n2648 vdd3p3.n2629 41.621
R5476 vdd3p3.n3139 vdd3p3.n3049 41.621
R5477 vdd3p3.n1999 vdd3p3.n1795 41.621
R5478 vdd3p3.n1802 vdd3p3.n1783 41.621
R5479 vdd3p3.n2293 vdd3p3.n2203 41.621
R5480 vdd3p3.n1154 vdd3p3.n950 41.621
R5481 vdd3p3.n957 vdd3p3.n938 41.621
R5482 vdd3p3.n1448 vdd3p3.n1358 41.621
R5483 vdd3p3.n308 vdd3p3.n104 41.621
R5484 vdd3p3.n111 vdd3p3.n92 41.621
R5485 vdd3p3.n602 vdd3p3.n512 41.621
R5486 vdd3p3.n2852 vdd3p3.n2641 41.621
R5487 vdd3p3.n2657 vdd3p3.n2629 41.621
R5488 vdd3p3.n3130 vdd3p3.n3049 41.621
R5489 vdd3p3.n2006 vdd3p3.n1795 41.621
R5490 vdd3p3.n1811 vdd3p3.n1783 41.621
R5491 vdd3p3.n2284 vdd3p3.n2203 41.621
R5492 vdd3p3.n1161 vdd3p3.n950 41.621
R5493 vdd3p3.n966 vdd3p3.n938 41.621
R5494 vdd3p3.n1439 vdd3p3.n1358 41.621
R5495 vdd3p3.n315 vdd3p3.n104 41.621
R5496 vdd3p3.n120 vdd3p3.n92 41.621
R5497 vdd3p3.n593 vdd3p3.n512 41.621
R5498 vdd3p3.n2980 vdd3p3.n2979 40.821
R5499 vdd3p3.n3181 vdd3p3.n2772 40.821
R5500 vdd3p3.n3019 vdd3p3.n2771 40.821
R5501 vdd3p3.n3030 vdd3p3.n2770 40.821
R5502 vdd3p3.n3172 vdd3p3.n2769 40.821
R5503 vdd3p3.n3169 vdd3p3.n2768 40.821
R5504 vdd3p3.n3097 vdd3p3.n2763 40.821
R5505 vdd3p3.n3101 vdd3p3.n2762 40.821
R5506 vdd3p3.n3085 vdd3p3.n2761 40.821
R5507 vdd3p3.n3107 vdd3p3.n2760 40.821
R5508 vdd3p3.n3083 vdd3p3.n2759 40.821
R5509 vdd3p3.n3113 vdd3p3.n2758 40.821
R5510 vdd3p3.n3116 vdd3p3.n2757 40.821
R5511 vdd3p3.n2756 vdd3p3.n2754 40.821
R5512 vdd3p3.n2856 vdd3p3.n2855 40.821
R5513 vdd3p3.n3339 vdd3p3.n2671 40.821
R5514 vdd3p3.n2855 vdd3p3.n2671 40.821
R5515 vdd3p3.n2858 vdd3p3.n2856 40.821
R5516 vdd3p3.n2981 vdd3p3.n2980 40.821
R5517 vdd3p3.n3095 vdd3p3.n2763 40.821
R5518 vdd3p3.n3097 vdd3p3.n2762 40.821
R5519 vdd3p3.n3101 vdd3p3.n2761 40.821
R5520 vdd3p3.n3085 vdd3p3.n2760 40.821
R5521 vdd3p3.n3107 vdd3p3.n2759 40.821
R5522 vdd3p3.n3083 vdd3p3.n2758 40.821
R5523 vdd3p3.n3113 vdd3p3.n2757 40.821
R5524 vdd3p3.n3116 vdd3p3.n2756 40.821
R5525 vdd3p3.n2773 vdd3p3.n2772 40.821
R5526 vdd3p3.n3181 vdd3p3.n2771 40.821
R5527 vdd3p3.n3019 vdd3p3.n2770 40.821
R5528 vdd3p3.n3030 vdd3p3.n2769 40.821
R5529 vdd3p3.n3172 vdd3p3.n2768 40.821
R5530 vdd3p3.n2134 vdd3p3.n2133 40.821
R5531 vdd3p3.n2335 vdd3p3.n1926 40.821
R5532 vdd3p3.n2173 vdd3p3.n1925 40.821
R5533 vdd3p3.n2184 vdd3p3.n1924 40.821
R5534 vdd3p3.n2326 vdd3p3.n1923 40.821
R5535 vdd3p3.n2323 vdd3p3.n1922 40.821
R5536 vdd3p3.n2251 vdd3p3.n1917 40.821
R5537 vdd3p3.n2255 vdd3p3.n1916 40.821
R5538 vdd3p3.n2239 vdd3p3.n1915 40.821
R5539 vdd3p3.n2261 vdd3p3.n1914 40.821
R5540 vdd3p3.n2237 vdd3p3.n1913 40.821
R5541 vdd3p3.n2267 vdd3p3.n1912 40.821
R5542 vdd3p3.n2270 vdd3p3.n1911 40.821
R5543 vdd3p3.n1910 vdd3p3.n1908 40.821
R5544 vdd3p3.n2010 vdd3p3.n2009 40.821
R5545 vdd3p3.n2493 vdd3p3.n1825 40.821
R5546 vdd3p3.n2009 vdd3p3.n1825 40.821
R5547 vdd3p3.n2012 vdd3p3.n2010 40.821
R5548 vdd3p3.n2135 vdd3p3.n2134 40.821
R5549 vdd3p3.n2249 vdd3p3.n1917 40.821
R5550 vdd3p3.n2251 vdd3p3.n1916 40.821
R5551 vdd3p3.n2255 vdd3p3.n1915 40.821
R5552 vdd3p3.n2239 vdd3p3.n1914 40.821
R5553 vdd3p3.n2261 vdd3p3.n1913 40.821
R5554 vdd3p3.n2237 vdd3p3.n1912 40.821
R5555 vdd3p3.n2267 vdd3p3.n1911 40.821
R5556 vdd3p3.n2270 vdd3p3.n1910 40.821
R5557 vdd3p3.n1927 vdd3p3.n1926 40.821
R5558 vdd3p3.n2335 vdd3p3.n1925 40.821
R5559 vdd3p3.n2173 vdd3p3.n1924 40.821
R5560 vdd3p3.n2184 vdd3p3.n1923 40.821
R5561 vdd3p3.n2326 vdd3p3.n1922 40.821
R5562 vdd3p3.n1289 vdd3p3.n1288 40.821
R5563 vdd3p3.n1490 vdd3p3.n1081 40.821
R5564 vdd3p3.n1328 vdd3p3.n1080 40.821
R5565 vdd3p3.n1339 vdd3p3.n1079 40.821
R5566 vdd3p3.n1481 vdd3p3.n1078 40.821
R5567 vdd3p3.n1478 vdd3p3.n1077 40.821
R5568 vdd3p3.n1406 vdd3p3.n1072 40.821
R5569 vdd3p3.n1410 vdd3p3.n1071 40.821
R5570 vdd3p3.n1394 vdd3p3.n1070 40.821
R5571 vdd3p3.n1416 vdd3p3.n1069 40.821
R5572 vdd3p3.n1392 vdd3p3.n1068 40.821
R5573 vdd3p3.n1422 vdd3p3.n1067 40.821
R5574 vdd3p3.n1425 vdd3p3.n1066 40.821
R5575 vdd3p3.n1065 vdd3p3.n1063 40.821
R5576 vdd3p3.n1165 vdd3p3.n1164 40.821
R5577 vdd3p3.n1648 vdd3p3.n980 40.821
R5578 vdd3p3.n1164 vdd3p3.n980 40.821
R5579 vdd3p3.n1167 vdd3p3.n1165 40.821
R5580 vdd3p3.n1290 vdd3p3.n1289 40.821
R5581 vdd3p3.n1404 vdd3p3.n1072 40.821
R5582 vdd3p3.n1406 vdd3p3.n1071 40.821
R5583 vdd3p3.n1410 vdd3p3.n1070 40.821
R5584 vdd3p3.n1394 vdd3p3.n1069 40.821
R5585 vdd3p3.n1416 vdd3p3.n1068 40.821
R5586 vdd3p3.n1392 vdd3p3.n1067 40.821
R5587 vdd3p3.n1422 vdd3p3.n1066 40.821
R5588 vdd3p3.n1425 vdd3p3.n1065 40.821
R5589 vdd3p3.n1082 vdd3p3.n1081 40.821
R5590 vdd3p3.n1490 vdd3p3.n1080 40.821
R5591 vdd3p3.n1328 vdd3p3.n1079 40.821
R5592 vdd3p3.n1339 vdd3p3.n1078 40.821
R5593 vdd3p3.n1481 vdd3p3.n1077 40.821
R5594 vdd3p3.n443 vdd3p3.n442 40.821
R5595 vdd3p3.n644 vdd3p3.n235 40.821
R5596 vdd3p3.n482 vdd3p3.n234 40.821
R5597 vdd3p3.n493 vdd3p3.n233 40.821
R5598 vdd3p3.n635 vdd3p3.n232 40.821
R5599 vdd3p3.n632 vdd3p3.n231 40.821
R5600 vdd3p3.n560 vdd3p3.n226 40.821
R5601 vdd3p3.n564 vdd3p3.n225 40.821
R5602 vdd3p3.n548 vdd3p3.n224 40.821
R5603 vdd3p3.n570 vdd3p3.n223 40.821
R5604 vdd3p3.n546 vdd3p3.n222 40.821
R5605 vdd3p3.n576 vdd3p3.n221 40.821
R5606 vdd3p3.n579 vdd3p3.n220 40.821
R5607 vdd3p3.n219 vdd3p3.n217 40.821
R5608 vdd3p3.n319 vdd3p3.n318 40.821
R5609 vdd3p3.n802 vdd3p3.n134 40.821
R5610 vdd3p3.n318 vdd3p3.n134 40.821
R5611 vdd3p3.n321 vdd3p3.n319 40.821
R5612 vdd3p3.n444 vdd3p3.n443 40.821
R5613 vdd3p3.n558 vdd3p3.n226 40.821
R5614 vdd3p3.n560 vdd3p3.n225 40.821
R5615 vdd3p3.n564 vdd3p3.n224 40.821
R5616 vdd3p3.n548 vdd3p3.n223 40.821
R5617 vdd3p3.n570 vdd3p3.n222 40.821
R5618 vdd3p3.n546 vdd3p3.n221 40.821
R5619 vdd3p3.n576 vdd3p3.n220 40.821
R5620 vdd3p3.n579 vdd3p3.n219 40.821
R5621 vdd3p3.n236 vdd3p3.n235 40.821
R5622 vdd3p3.n644 vdd3p3.n234 40.821
R5623 vdd3p3.n482 vdd3p3.n233 40.821
R5624 vdd3p3.n493 vdd3p3.n232 40.821
R5625 vdd3p3.n635 vdd3p3.n231 40.821
R5626 vdd3p3.n7452 vdd3p3.n7451 40.821
R5627 vdd3p3.n7445 vdd3p3.n7444 40.821
R5628 vdd3p3.n7440 vdd3p3.n7439 40.821
R5629 vdd3p3.n7435 vdd3p3.n7434 40.821
R5630 vdd3p3.n7430 vdd3p3.n7429 40.821
R5631 vdd3p3.n7425 vdd3p3.n7423 40.821
R5632 vdd3p3.n7399 vdd3p3.n7398 40.821
R5633 vdd3p3.n7404 vdd3p3.n7403 40.821
R5634 vdd3p3.n7409 vdd3p3.n7408 40.821
R5635 vdd3p3.n7414 vdd3p3.n7413 40.821
R5636 vdd3p3.n7419 vdd3p3.n7418 40.821
R5637 vdd3p3.n7425 vdd3p3.n7424 40.821
R5638 vdd3p3.n4219 vdd3p3.n4218 39.517
R5639 vdd3p3.n5071 vdd3p3.n5070 39.517
R5640 vdd3p3.n3501 vdd3p3.n3500 39.517
R5641 vdd3p3.n4983 vdd3p3.n4982 39.517
R5642 vdd3p3.n8493 vdd3p3.n8492 39.517
R5643 vdd3p3.n8837 vdd3p3.n8836 39.517
R5644 vdd3p3.n8779 vdd3p3.n8778 39.517
R5645 vdd3p3.n3960 vdd3p3.n3898 39.206
R5646 vdd3p3.n3057 vdd3p3.n3052 38.799
R5647 vdd3p3.n3063 vdd3p3.n3062 38.799
R5648 vdd3p3.n3065 vdd3p3.n3050 38.799
R5649 vdd3p3.n3179 vdd3p3.n3178 38.799
R5650 vdd3p3.n2667 vdd3p3.n2639 38.799
R5651 vdd3p3.n3333 vdd3p3.n2676 38.799
R5652 vdd3p3.n3332 vdd3p3.n2677 38.799
R5653 vdd3p3.n3324 vdd3p3.n3323 38.799
R5654 vdd3p3.n2211 vdd3p3.n2206 38.799
R5655 vdd3p3.n2217 vdd3p3.n2216 38.799
R5656 vdd3p3.n2219 vdd3p3.n2204 38.799
R5657 vdd3p3.n2333 vdd3p3.n2332 38.799
R5658 vdd3p3.n1821 vdd3p3.n1793 38.799
R5659 vdd3p3.n2487 vdd3p3.n1830 38.799
R5660 vdd3p3.n2486 vdd3p3.n1831 38.799
R5661 vdd3p3.n2478 vdd3p3.n2477 38.799
R5662 vdd3p3.n1366 vdd3p3.n1361 38.799
R5663 vdd3p3.n1372 vdd3p3.n1371 38.799
R5664 vdd3p3.n1374 vdd3p3.n1359 38.799
R5665 vdd3p3.n1488 vdd3p3.n1487 38.799
R5666 vdd3p3.n976 vdd3p3.n948 38.799
R5667 vdd3p3.n1642 vdd3p3.n985 38.799
R5668 vdd3p3.n1641 vdd3p3.n986 38.799
R5669 vdd3p3.n1633 vdd3p3.n1632 38.799
R5670 vdd3p3.n520 vdd3p3.n515 38.799
R5671 vdd3p3.n526 vdd3p3.n525 38.799
R5672 vdd3p3.n528 vdd3p3.n513 38.799
R5673 vdd3p3.n642 vdd3p3.n641 38.799
R5674 vdd3p3.n130 vdd3p3.n102 38.799
R5675 vdd3p3.n796 vdd3p3.n139 38.799
R5676 vdd3p3.n795 vdd3p3.n140 38.799
R5677 vdd3p3.n787 vdd3p3.n786 38.799
R5678 vdd3p3.n3064 vdd3p3.n3063 38.798
R5679 vdd3p3.n3068 vdd3p3.n3050 38.798
R5680 vdd3p3.n3058 vdd3p3.n3057 38.798
R5681 vdd3p3.n3343 vdd3p3.n2667 38.798
R5682 vdd3p3.n3323 vdd3p3.n3322 38.798
R5683 vdd3p3.n2682 vdd3p3.n2677 38.798
R5684 vdd3p3.n2676 vdd3p3.n2668 38.798
R5685 vdd3p3.n2218 vdd3p3.n2217 38.798
R5686 vdd3p3.n2222 vdd3p3.n2204 38.798
R5687 vdd3p3.n2212 vdd3p3.n2211 38.798
R5688 vdd3p3.n2497 vdd3p3.n1821 38.798
R5689 vdd3p3.n2477 vdd3p3.n2476 38.798
R5690 vdd3p3.n1836 vdd3p3.n1831 38.798
R5691 vdd3p3.n1830 vdd3p3.n1822 38.798
R5692 vdd3p3.n1373 vdd3p3.n1372 38.798
R5693 vdd3p3.n1377 vdd3p3.n1359 38.798
R5694 vdd3p3.n1367 vdd3p3.n1366 38.798
R5695 vdd3p3.n1652 vdd3p3.n976 38.798
R5696 vdd3p3.n1632 vdd3p3.n1631 38.798
R5697 vdd3p3.n991 vdd3p3.n986 38.798
R5698 vdd3p3.n985 vdd3p3.n977 38.798
R5699 vdd3p3.n527 vdd3p3.n526 38.798
R5700 vdd3p3.n531 vdd3p3.n513 38.798
R5701 vdd3p3.n521 vdd3p3.n520 38.798
R5702 vdd3p3.n806 vdd3p3.n130 38.798
R5703 vdd3p3.n786 vdd3p3.n785 38.798
R5704 vdd3p3.n145 vdd3p3.n140 38.798
R5705 vdd3p3.n139 vdd3p3.n131 38.798
R5706 vdd3p3.n3178 vdd3p3.n3022 38.798
R5707 vdd3p3.n2332 vdd3p3.n2176 38.798
R5708 vdd3p3.n1487 vdd3p3.n1331 38.798
R5709 vdd3p3.n641 vdd3p3.n485 38.798
R5710 vdd3p3.n3176 vdd3p3.n3028 38.798
R5711 vdd3p3.n3163 vdd3p3.n3027 38.798
R5712 vdd3p3.n3176 vdd3p3.n3175 38.798
R5713 vdd3p3.n3167 vdd3p3.n3027 38.798
R5714 vdd3p3.n3104 vdd3p3.n3026 38.798
R5715 vdd3p3.n3110 vdd3p3.n3025 38.798
R5716 vdd3p3.n3119 vdd3p3.n3024 38.798
R5717 vdd3p3.n3111 vdd3p3.n3024 38.798
R5718 vdd3p3.n3105 vdd3p3.n3025 38.798
R5719 vdd3p3.n3099 vdd3p3.n3026 38.798
R5720 vdd3p3.n2330 vdd3p3.n2182 38.798
R5721 vdd3p3.n2317 vdd3p3.n2181 38.798
R5722 vdd3p3.n2330 vdd3p3.n2329 38.798
R5723 vdd3p3.n2321 vdd3p3.n2181 38.798
R5724 vdd3p3.n2258 vdd3p3.n2180 38.798
R5725 vdd3p3.n2264 vdd3p3.n2179 38.798
R5726 vdd3p3.n2273 vdd3p3.n2178 38.798
R5727 vdd3p3.n2265 vdd3p3.n2178 38.798
R5728 vdd3p3.n2259 vdd3p3.n2179 38.798
R5729 vdd3p3.n2253 vdd3p3.n2180 38.798
R5730 vdd3p3.n1485 vdd3p3.n1337 38.798
R5731 vdd3p3.n1472 vdd3p3.n1336 38.798
R5732 vdd3p3.n1485 vdd3p3.n1484 38.798
R5733 vdd3p3.n1476 vdd3p3.n1336 38.798
R5734 vdd3p3.n1413 vdd3p3.n1335 38.798
R5735 vdd3p3.n1419 vdd3p3.n1334 38.798
R5736 vdd3p3.n1428 vdd3p3.n1333 38.798
R5737 vdd3p3.n1420 vdd3p3.n1333 38.798
R5738 vdd3p3.n1414 vdd3p3.n1334 38.798
R5739 vdd3p3.n1408 vdd3p3.n1335 38.798
R5740 vdd3p3.n639 vdd3p3.n491 38.798
R5741 vdd3p3.n626 vdd3p3.n490 38.798
R5742 vdd3p3.n639 vdd3p3.n638 38.798
R5743 vdd3p3.n630 vdd3p3.n490 38.798
R5744 vdd3p3.n567 vdd3p3.n489 38.798
R5745 vdd3p3.n573 vdd3p3.n488 38.798
R5746 vdd3p3.n582 vdd3p3.n487 38.798
R5747 vdd3p3.n574 vdd3p3.n487 38.798
R5748 vdd3p3.n568 vdd3p3.n488 38.798
R5749 vdd3p3.n562 vdd3p3.n489 38.798
R5750 vdd3p3.n7510 vdd3p3.n7509 38.776
R5751 vdd3p3.n3161 vdd3p3.n3160 36.538
R5752 vdd3p3.n3153 vdd3p3.n3042 36.538
R5753 vdd3p3.n2315 vdd3p3.n2314 36.538
R5754 vdd3p3.n2307 vdd3p3.n2196 36.538
R5755 vdd3p3.n1470 vdd3p3.n1469 36.538
R5756 vdd3p3.n1462 vdd3p3.n1351 36.538
R5757 vdd3p3.n624 vdd3p3.n623 36.538
R5758 vdd3p3.n616 vdd3p3.n505 36.538
R5759 vdd3p3.n4932 vdd3p3.n4931 36.224
R5760 vdd3p3.n51 vdd3p3.n35 36.141
R5761 vdd3p3.n51 vdd3p3.n50 36.141
R5762 vdd3p3.n50 vdd3p3.n39 36.141
R5763 vdd3p3.n46 vdd3p3.n39 36.141
R5764 vdd3p3.n16 vdd3p3.n8 36.141
R5765 vdd3p3.n27 vdd3p3.n8 36.141
R5766 vdd3p3.n27 vdd3p3.n4 36.141
R5767 vdd3p3.n58 vdd3p3.n4 36.141
R5768 vdd3p3.n893 vdd3p3.n888 36.141
R5769 vdd3p3.n893 vdd3p3.n892 36.141
R5770 vdd3p3.n892 vdd3p3.n847 36.141
R5771 vdd3p3.n898 vdd3p3.n847 36.141
R5772 vdd3p3.n865 vdd3p3.n856 36.141
R5773 vdd3p3.n870 vdd3p3.n856 36.141
R5774 vdd3p3.n870 vdd3p3.n851 36.141
R5775 vdd3p3.n881 vdd3p3.n851 36.141
R5776 vdd3p3.n1742 vdd3p3.n1726 36.141
R5777 vdd3p3.n1742 vdd3p3.n1741 36.141
R5778 vdd3p3.n1741 vdd3p3.n1730 36.141
R5779 vdd3p3.n1737 vdd3p3.n1730 36.141
R5780 vdd3p3.n1707 vdd3p3.n1699 36.141
R5781 vdd3p3.n1718 vdd3p3.n1699 36.141
R5782 vdd3p3.n1718 vdd3p3.n1695 36.141
R5783 vdd3p3.n1749 vdd3p3.n1695 36.141
R5784 vdd3p3.n2584 vdd3p3.n2579 36.141
R5785 vdd3p3.n2584 vdd3p3.n2583 36.141
R5786 vdd3p3.n2583 vdd3p3.n2538 36.141
R5787 vdd3p3.n2589 vdd3p3.n2538 36.141
R5788 vdd3p3.n2556 vdd3p3.n2547 36.141
R5789 vdd3p3.n2561 vdd3p3.n2547 36.141
R5790 vdd3p3.n2561 vdd3p3.n2542 36.141
R5791 vdd3p3.n2572 vdd3p3.n2542 36.141
R5792 vdd3p3.n3285 vdd3p3.n2702 35.962
R5793 vdd3p3.n2439 vdd3p3.n1856 35.962
R5794 vdd3p3.n1594 vdd3p3.n1011 35.962
R5795 vdd3p3.n748 vdd3p3.n165 35.962
R5796 vdd3p3.n3188 vdd3p3.n2755 35.256
R5797 vdd3p3.n2342 vdd3p3.n1909 35.256
R5798 vdd3p3.n1497 vdd3p3.n1064 35.256
R5799 vdd3p3.n651 vdd3p3.n218 35.256
R5800 vdd3p3.n6394 vdd3p3.n6393 34.635
R5801 vdd3p3.n2885 vdd3p3.n2672 34.615
R5802 vdd3p3.n2039 vdd3p3.n1826 34.615
R5803 vdd3p3.n1194 vdd3p3.n981 34.615
R5804 vdd3p3.n348 vdd3p3.n135 34.615
R5805 vdd3p3.n7010 vdd3p3.n7007 34.38
R5806 vdd3p3.n5739 vdd3p3.n5738 34.338
R5807 vdd3p3.n7467 vdd3p3.n7463 34.298
R5808 vdd3p3.n7942 vdd3p3.n7940 33.902
R5809 vdd3p3.n8455 vdd3p3.n8451 33.853
R5810 vdd3p3.n2740 vdd3p3.n2737 33.443
R5811 vdd3p3.n2703 vdd3p3.n2701 33.443
R5812 vdd3p3.n3317 vdd3p3.n3316 33.443
R5813 vdd3p3.n3336 vdd3p3.n2673 33.443
R5814 vdd3p3.n3329 vdd3p3.n3328 33.443
R5815 vdd3p3.n2685 vdd3p3.n2680 33.443
R5816 vdd3p3.n2878 vdd3p3.n2842 33.443
R5817 vdd3p3.n2870 vdd3p3.n2869 33.443
R5818 vdd3p3.n2854 vdd3p3.n2849 33.443
R5819 vdd3p3.n2822 vdd3p3.n2820 33.443
R5820 vdd3p3.n2917 vdd3p3.n2916 33.443
R5821 vdd3p3.n2986 vdd3p3.n2985 33.443
R5822 vdd3p3.n1894 vdd3p3.n1891 33.443
R5823 vdd3p3.n1857 vdd3p3.n1855 33.443
R5824 vdd3p3.n2471 vdd3p3.n2470 33.443
R5825 vdd3p3.n2490 vdd3p3.n1827 33.443
R5826 vdd3p3.n2483 vdd3p3.n2482 33.443
R5827 vdd3p3.n1839 vdd3p3.n1834 33.443
R5828 vdd3p3.n2032 vdd3p3.n1996 33.443
R5829 vdd3p3.n2024 vdd3p3.n2023 33.443
R5830 vdd3p3.n2008 vdd3p3.n2003 33.443
R5831 vdd3p3.n1976 vdd3p3.n1974 33.443
R5832 vdd3p3.n2071 vdd3p3.n2070 33.443
R5833 vdd3p3.n2140 vdd3p3.n2139 33.443
R5834 vdd3p3.n1049 vdd3p3.n1046 33.443
R5835 vdd3p3.n1012 vdd3p3.n1010 33.443
R5836 vdd3p3.n1626 vdd3p3.n1625 33.443
R5837 vdd3p3.n1645 vdd3p3.n982 33.443
R5838 vdd3p3.n1638 vdd3p3.n1637 33.443
R5839 vdd3p3.n994 vdd3p3.n989 33.443
R5840 vdd3p3.n1187 vdd3p3.n1151 33.443
R5841 vdd3p3.n1179 vdd3p3.n1178 33.443
R5842 vdd3p3.n1163 vdd3p3.n1158 33.443
R5843 vdd3p3.n1131 vdd3p3.n1129 33.443
R5844 vdd3p3.n1226 vdd3p3.n1225 33.443
R5845 vdd3p3.n1295 vdd3p3.n1294 33.443
R5846 vdd3p3.n203 vdd3p3.n200 33.443
R5847 vdd3p3.n166 vdd3p3.n164 33.443
R5848 vdd3p3.n780 vdd3p3.n779 33.443
R5849 vdd3p3.n799 vdd3p3.n136 33.443
R5850 vdd3p3.n792 vdd3p3.n791 33.443
R5851 vdd3p3.n148 vdd3p3.n143 33.443
R5852 vdd3p3.n341 vdd3p3.n305 33.443
R5853 vdd3p3.n333 vdd3p3.n332 33.443
R5854 vdd3p3.n317 vdd3p3.n312 33.443
R5855 vdd3p3.n285 vdd3p3.n283 33.443
R5856 vdd3p3.n380 vdd3p3.n379 33.443
R5857 vdd3p3.n449 vdd3p3.n448 33.443
R5858 vdd3p3.n8442 vdd3p3.n8440 33.443
R5859 vdd3p3.n8445 vdd3p3.n8443 33.443
R5860 vdd3p3.n7951 vdd3p3.n7950 33.443
R5861 vdd3p3.n8021 vdd3p3.n8020 33.443
R5862 vdd3p3.n7940 vdd3p3.n7936 33.443
R5863 vdd3p3.n7463 vdd3p3.n7460 33.443
R5864 vdd3p3.n5738 vdd3p3.n5736 33.443
R5865 vdd3p3.n7007 vdd3p3.n7003 33.443
R5866 vdd3p3.n2737 vdd3p3.n2736 33.442
R5867 vdd3p3.n2704 vdd3p3.n2703 33.442
R5868 vdd3p3.n3318 vdd3p3.n3317 33.442
R5869 vdd3p3.n3319 vdd3p3.n2685 33.442
R5870 vdd3p3.n3328 vdd3p3.n3327 33.442
R5871 vdd3p3.n2679 vdd3p3.n2673 33.442
R5872 vdd3p3.n2861 vdd3p3.n2854 33.442
R5873 vdd3p3.n2869 vdd3p3.n2868 33.442
R5874 vdd3p3.n2848 vdd3p3.n2842 33.442
R5875 vdd3p3.n2916 vdd3p3.n2915 33.442
R5876 vdd3p3.n2918 vdd3p3.n2822 33.442
R5877 vdd3p3.n2985 vdd3p3.n2792 33.442
R5878 vdd3p3.n1891 vdd3p3.n1890 33.442
R5879 vdd3p3.n1858 vdd3p3.n1857 33.442
R5880 vdd3p3.n2472 vdd3p3.n2471 33.442
R5881 vdd3p3.n2473 vdd3p3.n1839 33.442
R5882 vdd3p3.n2482 vdd3p3.n2481 33.442
R5883 vdd3p3.n1833 vdd3p3.n1827 33.442
R5884 vdd3p3.n2015 vdd3p3.n2008 33.442
R5885 vdd3p3.n2023 vdd3p3.n2022 33.442
R5886 vdd3p3.n2002 vdd3p3.n1996 33.442
R5887 vdd3p3.n2070 vdd3p3.n2069 33.442
R5888 vdd3p3.n2072 vdd3p3.n1976 33.442
R5889 vdd3p3.n2139 vdd3p3.n1946 33.442
R5890 vdd3p3.n1046 vdd3p3.n1045 33.442
R5891 vdd3p3.n1013 vdd3p3.n1012 33.442
R5892 vdd3p3.n1627 vdd3p3.n1626 33.442
R5893 vdd3p3.n1628 vdd3p3.n994 33.442
R5894 vdd3p3.n1637 vdd3p3.n1636 33.442
R5895 vdd3p3.n988 vdd3p3.n982 33.442
R5896 vdd3p3.n1170 vdd3p3.n1163 33.442
R5897 vdd3p3.n1178 vdd3p3.n1177 33.442
R5898 vdd3p3.n1157 vdd3p3.n1151 33.442
R5899 vdd3p3.n1225 vdd3p3.n1224 33.442
R5900 vdd3p3.n1227 vdd3p3.n1131 33.442
R5901 vdd3p3.n1294 vdd3p3.n1101 33.442
R5902 vdd3p3.n200 vdd3p3.n199 33.442
R5903 vdd3p3.n167 vdd3p3.n166 33.442
R5904 vdd3p3.n781 vdd3p3.n780 33.442
R5905 vdd3p3.n782 vdd3p3.n148 33.442
R5906 vdd3p3.n791 vdd3p3.n790 33.442
R5907 vdd3p3.n142 vdd3p3.n136 33.442
R5908 vdd3p3.n324 vdd3p3.n317 33.442
R5909 vdd3p3.n332 vdd3p3.n331 33.442
R5910 vdd3p3.n311 vdd3p3.n305 33.442
R5911 vdd3p3.n379 vdd3p3.n378 33.442
R5912 vdd3p3.n381 vdd3p3.n285 33.442
R5913 vdd3p3.n448 vdd3p3.n255 33.442
R5914 vdd3p3.n6393 vdd3p3.n6391 33.442
R5915 vdd3p3.n8442 vdd3p3.n8441 33.442
R5916 vdd3p3.n8445 vdd3p3.n8444 33.442
R5917 vdd3p3.n7970 vdd3p3.n7969 33.442
R5918 vdd3p3.n7986 vdd3p3.n7985 33.442
R5919 vdd3p3.n8000 vdd3p3.n7999 33.442
R5920 vdd3p3.n8014 vdd3p3.n8013 33.442
R5921 vdd3p3.n7463 vdd3p3.n7462 33.442
R5922 vdd3p3.n5738 vdd3p3.n5737 33.442
R5923 vdd3p3.n7007 vdd3p3.n7006 33.442
R5924 vdd3p3.n3092 vdd3p3.n2765 33.442
R5925 vdd3p3.n3089 vdd3p3.n2765 33.442
R5926 vdd3p3.n2246 vdd3p3.n1919 33.442
R5927 vdd3p3.n2243 vdd3p3.n1919 33.442
R5928 vdd3p3.n1401 vdd3p3.n1074 33.442
R5929 vdd3p3.n1398 vdd3p3.n1074 33.442
R5930 vdd3p3.n555 vdd3p3.n228 33.442
R5931 vdd3p3.n552 vdd3p3.n228 33.442
R5932 vdd3p3.n6358 vdd3p3.n6357 33.442
R5933 vdd3p3.n6347 vdd3p3.n6346 33.442
R5934 vdd3p3.n6338 vdd3p3.n6337 33.442
R5935 vdd3p3.n6329 vdd3p3.n6328 33.442
R5936 vdd3p3.n6320 vdd3p3.n6319 33.442
R5937 vdd3p3.n6279 vdd3p3.n6278 33.442
R5938 vdd3p3.n6268 vdd3p3.n6267 33.442
R5939 vdd3p3.n6288 vdd3p3.n6287 33.442
R5940 vdd3p3.n6297 vdd3p3.n6296 33.442
R5941 vdd3p3.n6306 vdd3p3.n6305 33.442
R5942 vdd3p3.n6315 vdd3p3.n6314 33.442
R5943 vdd3p3.n6367 vdd3p3.n6366 33.442
R5944 vdd3p3.n6376 vdd3p3.n6375 33.442
R5945 vdd3p3.n6385 vdd3p3.n6384 33.442
R5946 vdd3p3.n3221 vdd3p3.n2733 32.965
R5947 vdd3p3.n2375 vdd3p3.n1887 32.965
R5948 vdd3p3.n1530 vdd3p3.n1042 32.965
R5949 vdd3p3.n684 vdd3p3.n196 32.965
R5950 vdd3p3.n4189 vdd3p3.n4188 32.931
R5951 vdd3p3.n5085 vdd3p3.n5084 32.931
R5952 vdd3p3.n4902 vdd3p3.n4901 32.931
R5953 vdd3p3.n8530 vdd3p3.n8529 32.931
R5954 vdd3p3.n8875 vdd3p3.n8874 32.931
R5955 vdd3p3.n8792 vdd3p3.n8791 32.931
R5956 vdd3p3.n2985 vdd3p3.n2984 32.66
R5957 vdd3p3.n2139 vdd3p3.n2138 32.66
R5958 vdd3p3.n1294 vdd3p3.n1293 32.66
R5959 vdd3p3.n448 vdd3p3.n447 32.66
R5960 vdd3p3.n3350 vdd3p3.n2641 30.128
R5961 vdd3p3.n2504 vdd3p3.n1795 30.128
R5962 vdd3p3.n1659 vdd3p3.n950 30.128
R5963 vdd3p3.n813 vdd3p3.n104 30.128
R5964 vdd3p3.n3059 vdd3p3.n3053 30.117
R5965 vdd3p3.n3354 vdd3p3.n2636 30.117
R5966 vdd3p3.n2662 vdd3p3.n2659 30.117
R5967 vdd3p3.n3144 vdd3p3.n3141 30.117
R5968 vdd3p3.n3128 vdd3p3.n3127 30.117
R5969 vdd3p3.n2213 vdd3p3.n2207 30.117
R5970 vdd3p3.n2508 vdd3p3.n1790 30.117
R5971 vdd3p3.n1816 vdd3p3.n1813 30.117
R5972 vdd3p3.n2298 vdd3p3.n2295 30.117
R5973 vdd3p3.n2282 vdd3p3.n2281 30.117
R5974 vdd3p3.n1368 vdd3p3.n1362 30.117
R5975 vdd3p3.n1663 vdd3p3.n945 30.117
R5976 vdd3p3.n971 vdd3p3.n968 30.117
R5977 vdd3p3.n1453 vdd3p3.n1450 30.117
R5978 vdd3p3.n1437 vdd3p3.n1436 30.117
R5979 vdd3p3.n522 vdd3p3.n516 30.117
R5980 vdd3p3.n817 vdd3p3.n99 30.117
R5981 vdd3p3.n125 vdd3p3.n122 30.117
R5982 vdd3p3.n607 vdd3p3.n604 30.117
R5983 vdd3p3.n591 vdd3p3.n590 30.117
R5984 vdd3p3.n2845 vdd3p3.n2844 30.07
R5985 vdd3p3.n2648 vdd3p3.n2647 30.07
R5986 vdd3p3.n3140 vdd3p3.n3139 30.07
R5987 vdd3p3.n1999 vdd3p3.n1998 30.07
R5988 vdd3p3.n1802 vdd3p3.n1801 30.07
R5989 vdd3p3.n2294 vdd3p3.n2293 30.07
R5990 vdd3p3.n1154 vdd3p3.n1153 30.07
R5991 vdd3p3.n957 vdd3p3.n956 30.07
R5992 vdd3p3.n1449 vdd3p3.n1448 30.07
R5993 vdd3p3.n308 vdd3p3.n307 30.07
R5994 vdd3p3.n111 vdd3p3.n110 30.07
R5995 vdd3p3.n603 vdd3p3.n602 30.07
R5996 vdd3p3.n3130 vdd3p3.n3129 30.07
R5997 vdd3p3.n2865 vdd3p3.n2852 30.07
R5998 vdd3p3.n2658 vdd3p3.n2657 30.07
R5999 vdd3p3.n2284 vdd3p3.n2283 30.07
R6000 vdd3p3.n2019 vdd3p3.n2006 30.07
R6001 vdd3p3.n1812 vdd3p3.n1811 30.07
R6002 vdd3p3.n1439 vdd3p3.n1438 30.07
R6003 vdd3p3.n1174 vdd3p3.n1161 30.07
R6004 vdd3p3.n967 vdd3p3.n966 30.07
R6005 vdd3p3.n593 vdd3p3.n592 30.07
R6006 vdd3p3.n328 vdd3p3.n315 30.07
R6007 vdd3p3.n121 vdd3p3.n120 30.07
R6008 vdd3p3.n4182 vdd3p3.n4181 29.637
R6009 vdd3p3.n5042 vdd3p3.n5041 29.637
R6010 vdd3p3.n4943 vdd3p3.n4942 29.637
R6011 vdd3p3.n8550 vdd3p3.n8549 29.637
R6012 vdd3p3.n8629 vdd3p3.n8628 29.637
R6013 vdd3p3.n8812 vdd3p3.n8811 29.637
R6014 vdd3p3.n3222 vdd3p3.n2737 29.53
R6015 vdd3p3.n3284 vdd3p3.n2703 29.53
R6016 vdd3p3.n2673 vdd3p3.n2672 29.53
R6017 vdd3p3.n3328 vdd3p3.n2672 29.53
R6018 vdd3p3.n2685 vdd3p3.n2672 29.53
R6019 vdd3p3.n3317 vdd3p3.n2672 29.53
R6020 vdd3p3.n2842 vdd3p3.n2672 29.53
R6021 vdd3p3.n2869 vdd3p3.n2672 29.53
R6022 vdd3p3.n2854 vdd3p3.n2672 29.53
R6023 vdd3p3.n2823 vdd3p3.n2822 29.53
R6024 vdd3p3.n2916 vdd3p3.n2823 29.53
R6025 vdd3p3.n2376 vdd3p3.n1891 29.53
R6026 vdd3p3.n2438 vdd3p3.n1857 29.53
R6027 vdd3p3.n1827 vdd3p3.n1826 29.53
R6028 vdd3p3.n2482 vdd3p3.n1826 29.53
R6029 vdd3p3.n1839 vdd3p3.n1826 29.53
R6030 vdd3p3.n2471 vdd3p3.n1826 29.53
R6031 vdd3p3.n1996 vdd3p3.n1826 29.53
R6032 vdd3p3.n2023 vdd3p3.n1826 29.53
R6033 vdd3p3.n2008 vdd3p3.n1826 29.53
R6034 vdd3p3.n1977 vdd3p3.n1976 29.53
R6035 vdd3p3.n2070 vdd3p3.n1977 29.53
R6036 vdd3p3.n1531 vdd3p3.n1046 29.53
R6037 vdd3p3.n1593 vdd3p3.n1012 29.53
R6038 vdd3p3.n982 vdd3p3.n981 29.53
R6039 vdd3p3.n1637 vdd3p3.n981 29.53
R6040 vdd3p3.n994 vdd3p3.n981 29.53
R6041 vdd3p3.n1626 vdd3p3.n981 29.53
R6042 vdd3p3.n1151 vdd3p3.n981 29.53
R6043 vdd3p3.n1178 vdd3p3.n981 29.53
R6044 vdd3p3.n1163 vdd3p3.n981 29.53
R6045 vdd3p3.n1132 vdd3p3.n1131 29.53
R6046 vdd3p3.n1225 vdd3p3.n1132 29.53
R6047 vdd3p3.n685 vdd3p3.n200 29.53
R6048 vdd3p3.n747 vdd3p3.n166 29.53
R6049 vdd3p3.n136 vdd3p3.n135 29.53
R6050 vdd3p3.n791 vdd3p3.n135 29.53
R6051 vdd3p3.n148 vdd3p3.n135 29.53
R6052 vdd3p3.n780 vdd3p3.n135 29.53
R6053 vdd3p3.n305 vdd3p3.n135 29.53
R6054 vdd3p3.n332 vdd3p3.n135 29.53
R6055 vdd3p3.n317 vdd3p3.n135 29.53
R6056 vdd3p3.n286 vdd3p3.n285 29.53
R6057 vdd3p3.n379 vdd3p3.n286 29.53
R6058 vdd3p3.n8459 vdd3p3.n8442 29.53
R6059 vdd3p3.n8459 vdd3p3.n8445 29.53
R6060 vdd3p3.n7939 vdd3p3.n7938 29.53
R6061 vdd3p3.n4716 vdd3p3.n4715 29.53
R6062 vdd3p3.n3188 vdd3p3.n2765 29.53
R6063 vdd3p3.n2342 vdd3p3.n1919 29.53
R6064 vdd3p3.n1497 vdd3p3.n1074 29.53
R6065 vdd3p3.n651 vdd3p3.n228 29.53
R6066 vdd3p3.n4716 vdd3p3.n4714 29.53
R6067 vdd3p3.n4716 vdd3p3.n4713 29.53
R6068 vdd3p3.n4716 vdd3p3.n4712 29.53
R6069 vdd3p3.n4716 vdd3p3.n4711 29.53
R6070 vdd3p3.n4716 vdd3p3.n4710 29.53
R6071 vdd3p3.n4716 vdd3p3.n4709 29.53
R6072 vdd3p3.n4716 vdd3p3.n4708 29.53
R6073 vdd3p3.n4716 vdd3p3.n4707 29.53
R6074 vdd3p3.n4716 vdd3p3.n4706 29.53
R6075 vdd3p3.n4716 vdd3p3.n4705 29.53
R6076 vdd3p3.n4716 vdd3p3.n4704 29.53
R6077 vdd3p3.n4716 vdd3p3.n4703 29.53
R6078 vdd3p3.n4716 vdd3p3.n4702 29.53
R6079 vdd3p3.n4716 vdd3p3.n4701 29.53
R6080 vdd3p3.n4716 vdd3p3.n4700 29.53
R6081 vdd3p3.n4716 vdd3p3.n4699 29.53
R6082 vdd3p3.n4716 vdd3p3.n4698 29.53
R6083 vdd3p3.n4716 vdd3p3.n4697 29.53
R6084 vdd3p3.n4716 vdd3p3.n4696 29.53
R6085 vdd3p3.n4716 vdd3p3.n4695 29.53
R6086 vdd3p3.n3367 vdd3p3.n2618 29.487
R6087 vdd3p3.n3363 vdd3p3.n2622 29.487
R6088 vdd3p3.n2521 vdd3p3.n1772 29.487
R6089 vdd3p3.n2517 vdd3p3.n1776 29.487
R6090 vdd3p3.n1676 vdd3p3.n927 29.487
R6091 vdd3p3.n1672 vdd3p3.n931 29.487
R6092 vdd3p3.n830 vdd3p3.n81 29.487
R6093 vdd3p3.n826 vdd3p3.n85 29.487
R6094 vdd3p3.t2 vdd3p3.n3048 28.846
R6095 vdd3p3.n2617 vdd3p3.t162 28.846
R6096 vdd3p3.n2630 vdd3p3.t128 28.846
R6097 vdd3p3.t77 vdd3p3.n2202 28.846
R6098 vdd3p3.n1771 vdd3p3.t110 28.846
R6099 vdd3p3.n1784 vdd3p3.t170 28.846
R6100 vdd3p3.t31 vdd3p3.n1357 28.846
R6101 vdd3p3.n926 vdd3p3.t165 28.846
R6102 vdd3p3.n939 vdd3p3.t23 28.846
R6103 vdd3p3.t135 vdd3p3.n511 28.846
R6104 vdd3p3.n80 vdd3p3.t159 28.846
R6105 vdd3p3.n93 vdd3p3.t20 28.846
R6106 vdd3p3.n5276 vdd3p3.n5275 28.596
R6107 vdd3p3.n5277 vdd3p3.n5276 28.596
R6108 vdd3p3.n5278 vdd3p3.n5277 28.596
R6109 vdd3p3.n5279 vdd3p3.n5278 28.596
R6110 vdd3p3.n5272 vdd3p3.n5271 28.596
R6111 vdd3p3.n5271 vdd3p3.n5270 28.596
R6112 vdd3p3.n5270 vdd3p3.n5269 28.596
R6113 vdd3p3.n5269 vdd3p3.n5268 28.596
R6114 vdd3p3.n5268 vdd3p3.n5267 28.596
R6115 vdd3p3.n6550 vdd3p3.n6549 28.596
R6116 vdd3p3.n6551 vdd3p3.n6550 28.596
R6117 vdd3p3.n6552 vdd3p3.n6551 28.596
R6118 vdd3p3.n6553 vdd3p3.n6552 28.596
R6119 vdd3p3.n6554 vdd3p3.n6553 28.596
R6120 vdd3p3.n6561 vdd3p3.n6560 28.596
R6121 vdd3p3.n6560 vdd3p3.n6559 28.596
R6122 vdd3p3.n6559 vdd3p3.n6558 28.596
R6123 vdd3p3.n6558 vdd3p3.n6557 28.596
R6124 vdd3p3.n6557 vdd3p3.n6556 28.596
R6125 vdd3p3.n6556 vdd3p3.n6555 28.596
R6126 vdd3p3.n8647 vdd3p3.n8646 28.596
R6127 vdd3p3.n8648 vdd3p3.n8647 28.596
R6128 vdd3p3.n8649 vdd3p3.n8648 28.596
R6129 vdd3p3.n8650 vdd3p3.n8649 28.596
R6130 vdd3p3.n8725 vdd3p3.n8724 28.596
R6131 vdd3p3.n8724 vdd3p3.n8723 28.596
R6132 vdd3p3.n8723 vdd3p3.n8722 28.596
R6133 vdd3p3.n8651 vdd3p3.n8650 28.176
R6134 vdd3p3.n55 vdd3p3.t140 28.155
R6135 vdd3p3.t166 vdd3p3.n884 28.155
R6136 vdd3p3.n1746 vdd3p3.t83 28.155
R6137 vdd3p3.t87 vdd3p3.n2575 28.155
R6138 vdd3p3.n2923 vdd3p3.n2819 28.078
R6139 vdd3p3.n2077 vdd3p3.n1973 28.078
R6140 vdd3p3.n1232 vdd3p3.n1128 28.078
R6141 vdd3p3.n386 vdd3p3.n282 28.078
R6142 vdd3p3.n2605 vdd3p3.t1 27.695
R6143 vdd3p3.n2605 vdd3p3.t3 27.695
R6144 vdd3p3.n2602 vdd3p3.t131 27.695
R6145 vdd3p3.n2602 vdd3p3.t129 27.695
R6146 vdd3p3.n1759 vdd3p3.t76 27.695
R6147 vdd3p3.n1759 vdd3p3.t78 27.695
R6148 vdd3p3.n1756 vdd3p3.t114 27.695
R6149 vdd3p3.n1756 vdd3p3.t171 27.695
R6150 vdd3p3.n914 vdd3p3.t30 27.695
R6151 vdd3p3.n914 vdd3p3.t32 27.695
R6152 vdd3p3.n911 vdd3p3.t119 27.695
R6153 vdd3p3.n911 vdd3p3.t24 27.695
R6154 vdd3p3.n68 vdd3p3.t134 27.695
R6155 vdd3p3.n68 vdd3p3.t136 27.695
R6156 vdd3p3.n65 vdd3p3.t17 27.695
R6157 vdd3p3.n65 vdd3p3.t21 27.695
R6158 vdd3p3.n3063 vdd3p3.n2611 26.852
R6159 vdd3p3.n3050 vdd3p3.n2611 26.852
R6160 vdd3p3.n3057 vdd3p3.n2611 26.852
R6161 vdd3p3.n3341 vdd3p3.n2667 26.852
R6162 vdd3p3.n2683 vdd3p3.n2677 26.852
R6163 vdd3p3.n3323 vdd3p3.n2683 26.852
R6164 vdd3p3.n2683 vdd3p3.n2676 26.852
R6165 vdd3p3.n2217 vdd3p3.n1765 26.852
R6166 vdd3p3.n2204 vdd3p3.n1765 26.852
R6167 vdd3p3.n2211 vdd3p3.n1765 26.852
R6168 vdd3p3.n2495 vdd3p3.n1821 26.852
R6169 vdd3p3.n1837 vdd3p3.n1831 26.852
R6170 vdd3p3.n2477 vdd3p3.n1837 26.852
R6171 vdd3p3.n1837 vdd3p3.n1830 26.852
R6172 vdd3p3.n1372 vdd3p3.n920 26.852
R6173 vdd3p3.n1359 vdd3p3.n920 26.852
R6174 vdd3p3.n1366 vdd3p3.n920 26.852
R6175 vdd3p3.n1650 vdd3p3.n976 26.852
R6176 vdd3p3.n992 vdd3p3.n986 26.852
R6177 vdd3p3.n1632 vdd3p3.n992 26.852
R6178 vdd3p3.n992 vdd3p3.n985 26.852
R6179 vdd3p3.n526 vdd3p3.n74 26.852
R6180 vdd3p3.n513 vdd3p3.n74 26.852
R6181 vdd3p3.n520 vdd3p3.n74 26.852
R6182 vdd3p3.n804 vdd3p3.n130 26.852
R6183 vdd3p3.n146 vdd3p3.n140 26.852
R6184 vdd3p3.n786 vdd3p3.n146 26.852
R6185 vdd3p3.n146 vdd3p3.n139 26.852
R6186 vdd3p3.n3178 vdd3p3.n3177 26.852
R6187 vdd3p3.n2332 vdd3p3.n2331 26.852
R6188 vdd3p3.n1487 vdd3p3.n1486 26.852
R6189 vdd3p3.n641 vdd3p3.n640 26.852
R6190 vdd3p3.n3177 vdd3p3.n3176 26.852
R6191 vdd3p3.n3177 vdd3p3.n3027 26.852
R6192 vdd3p3.n3177 vdd3p3.n3024 26.852
R6193 vdd3p3.n3177 vdd3p3.n3025 26.852
R6194 vdd3p3.n3177 vdd3p3.n3026 26.852
R6195 vdd3p3.n2331 vdd3p3.n2330 26.852
R6196 vdd3p3.n2331 vdd3p3.n2181 26.852
R6197 vdd3p3.n2331 vdd3p3.n2178 26.852
R6198 vdd3p3.n2331 vdd3p3.n2179 26.852
R6199 vdd3p3.n2331 vdd3p3.n2180 26.852
R6200 vdd3p3.n1486 vdd3p3.n1485 26.852
R6201 vdd3p3.n1486 vdd3p3.n1336 26.852
R6202 vdd3p3.n1486 vdd3p3.n1333 26.852
R6203 vdd3p3.n1486 vdd3p3.n1334 26.852
R6204 vdd3p3.n1486 vdd3p3.n1335 26.852
R6205 vdd3p3.n640 vdd3p3.n639 26.852
R6206 vdd3p3.n640 vdd3p3.n490 26.852
R6207 vdd3p3.n640 vdd3p3.n487 26.852
R6208 vdd3p3.n640 vdd3p3.n488 26.852
R6209 vdd3p3.n640 vdd3p3.n489 26.852
R6210 vdd3p3.n3067 vdd3p3.n2607 26.352
R6211 vdd3p3.n2221 vdd3p3.n1761 26.352
R6212 vdd3p3.n1376 vdd3p3.n916 26.352
R6213 vdd3p3.n530 vdd3p3.n70 26.352
R6214 vdd3p3.n4181 vdd3p3.n4180 26.344
R6215 vdd3p3.n5041 vdd3p3.n5040 26.344
R6216 vdd3p3.n4942 vdd3p3.n4941 26.344
R6217 vdd3p3.n8549 vdd3p3.n8548 26.344
R6218 vdd3p3.n8628 vdd3p3.n8627 26.344
R6219 vdd3p3.n8811 vdd3p3.n8810 26.344
R6220 vdd3p3.n3392 vdd3p3.n3391 25.987
R6221 vdd3p3.n2988 vdd3p3.n2987 25.738
R6222 vdd3p3.n2142 vdd3p3.n2141 25.738
R6223 vdd3p3.n1297 vdd3p3.n1296 25.738
R6224 vdd3p3.n451 vdd3p3.n450 25.738
R6225 vdd3p3.n3060 vdd3p3.n3059 25.6
R6226 vdd3p3.n3061 vdd3p3.n3060 25.6
R6227 vdd3p3.n3061 vdd3p3.n3051 25.6
R6228 vdd3p3.n3066 vdd3p3.n3051 25.6
R6229 vdd3p3.n3067 vdd3p3.n3066 25.6
R6230 vdd3p3.n3289 vdd3p3.n3288 25.6
R6231 vdd3p3.n3288 vdd3p3.n2700 25.6
R6232 vdd3p3.n2706 vdd3p3.n2700 25.6
R6233 vdd3p3.n3282 vdd3p3.n2706 25.6
R6234 vdd3p3.n3226 vdd3p3.n3225 25.6
R6235 vdd3p3.n3226 vdd3p3.n2731 25.6
R6236 vdd3p3.n3232 vdd3p3.n2731 25.6
R6237 vdd3p3.n3233 vdd3p3.n3232 25.6
R6238 vdd3p3.n3234 vdd3p3.n3233 25.6
R6239 vdd3p3.n3234 vdd3p3.n2727 25.6
R6240 vdd3p3.n3240 vdd3p3.n2727 25.6
R6241 vdd3p3.n3241 vdd3p3.n3240 25.6
R6242 vdd3p3.n3242 vdd3p3.n3241 25.6
R6243 vdd3p3.n3242 vdd3p3.n2723 25.6
R6244 vdd3p3.n3248 vdd3p3.n2723 25.6
R6245 vdd3p3.n3249 vdd3p3.n3248 25.6
R6246 vdd3p3.n3250 vdd3p3.n3249 25.6
R6247 vdd3p3.n3250 vdd3p3.n2719 25.6
R6248 vdd3p3.n3256 vdd3p3.n2719 25.6
R6249 vdd3p3.n3257 vdd3p3.n3256 25.6
R6250 vdd3p3.n3258 vdd3p3.n3257 25.6
R6251 vdd3p3.n3258 vdd3p3.n2715 25.6
R6252 vdd3p3.n3264 vdd3p3.n2715 25.6
R6253 vdd3p3.n3265 vdd3p3.n3264 25.6
R6254 vdd3p3.n3266 vdd3p3.n3265 25.6
R6255 vdd3p3.n3266 vdd3p3.n2711 25.6
R6256 vdd3p3.n3272 vdd3p3.n2711 25.6
R6257 vdd3p3.n3273 vdd3p3.n3272 25.6
R6258 vdd3p3.n3274 vdd3p3.n3273 25.6
R6259 vdd3p3.n3274 vdd3p3.n2707 25.6
R6260 vdd3p3.n3280 vdd3p3.n2707 25.6
R6261 vdd3p3.n3281 vdd3p3.n3280 25.6
R6262 vdd3p3.n3218 vdd3p3.n3216 25.6
R6263 vdd3p3.n3218 vdd3p3.n3217 25.6
R6264 vdd3p3.n3217 vdd3p3.n2735 25.6
R6265 vdd3p3.n3224 vdd3p3.n2735 25.6
R6266 vdd3p3.n2646 vdd3p3.n2636 25.6
R6267 vdd3p3.n2652 vdd3p3.n2646 25.6
R6268 vdd3p3.n2653 vdd3p3.n2652 25.6
R6269 vdd3p3.n2653 vdd3p3.n2644 25.6
R6270 vdd3p3.n2659 vdd3p3.n2644 25.6
R6271 vdd3p3.n3141 vdd3p3.n3077 25.6
R6272 vdd3p3.n3135 vdd3p3.n3077 25.6
R6273 vdd3p3.n3135 vdd3p3.n3134 25.6
R6274 vdd3p3.n3134 vdd3p3.n3081 25.6
R6275 vdd3p3.n3128 vdd3p3.n3081 25.6
R6276 vdd3p3.n2214 vdd3p3.n2213 25.6
R6277 vdd3p3.n2215 vdd3p3.n2214 25.6
R6278 vdd3p3.n2215 vdd3p3.n2205 25.6
R6279 vdd3p3.n2220 vdd3p3.n2205 25.6
R6280 vdd3p3.n2221 vdd3p3.n2220 25.6
R6281 vdd3p3.n2443 vdd3p3.n2442 25.6
R6282 vdd3p3.n2442 vdd3p3.n1854 25.6
R6283 vdd3p3.n1860 vdd3p3.n1854 25.6
R6284 vdd3p3.n2436 vdd3p3.n1860 25.6
R6285 vdd3p3.n2380 vdd3p3.n2379 25.6
R6286 vdd3p3.n2380 vdd3p3.n1885 25.6
R6287 vdd3p3.n2386 vdd3p3.n1885 25.6
R6288 vdd3p3.n2387 vdd3p3.n2386 25.6
R6289 vdd3p3.n2388 vdd3p3.n2387 25.6
R6290 vdd3p3.n2388 vdd3p3.n1881 25.6
R6291 vdd3p3.n2394 vdd3p3.n1881 25.6
R6292 vdd3p3.n2395 vdd3p3.n2394 25.6
R6293 vdd3p3.n2396 vdd3p3.n2395 25.6
R6294 vdd3p3.n2396 vdd3p3.n1877 25.6
R6295 vdd3p3.n2402 vdd3p3.n1877 25.6
R6296 vdd3p3.n2403 vdd3p3.n2402 25.6
R6297 vdd3p3.n2404 vdd3p3.n2403 25.6
R6298 vdd3p3.n2404 vdd3p3.n1873 25.6
R6299 vdd3p3.n2410 vdd3p3.n1873 25.6
R6300 vdd3p3.n2411 vdd3p3.n2410 25.6
R6301 vdd3p3.n2412 vdd3p3.n2411 25.6
R6302 vdd3p3.n2412 vdd3p3.n1869 25.6
R6303 vdd3p3.n2418 vdd3p3.n1869 25.6
R6304 vdd3p3.n2419 vdd3p3.n2418 25.6
R6305 vdd3p3.n2420 vdd3p3.n2419 25.6
R6306 vdd3p3.n2420 vdd3p3.n1865 25.6
R6307 vdd3p3.n2426 vdd3p3.n1865 25.6
R6308 vdd3p3.n2427 vdd3p3.n2426 25.6
R6309 vdd3p3.n2428 vdd3p3.n2427 25.6
R6310 vdd3p3.n2428 vdd3p3.n1861 25.6
R6311 vdd3p3.n2434 vdd3p3.n1861 25.6
R6312 vdd3p3.n2435 vdd3p3.n2434 25.6
R6313 vdd3p3.n2372 vdd3p3.n2370 25.6
R6314 vdd3p3.n2372 vdd3p3.n2371 25.6
R6315 vdd3p3.n2371 vdd3p3.n1889 25.6
R6316 vdd3p3.n2378 vdd3p3.n1889 25.6
R6317 vdd3p3.n1800 vdd3p3.n1790 25.6
R6318 vdd3p3.n1806 vdd3p3.n1800 25.6
R6319 vdd3p3.n1807 vdd3p3.n1806 25.6
R6320 vdd3p3.n1807 vdd3p3.n1798 25.6
R6321 vdd3p3.n1813 vdd3p3.n1798 25.6
R6322 vdd3p3.n2295 vdd3p3.n2231 25.6
R6323 vdd3p3.n2289 vdd3p3.n2231 25.6
R6324 vdd3p3.n2289 vdd3p3.n2288 25.6
R6325 vdd3p3.n2288 vdd3p3.n2235 25.6
R6326 vdd3p3.n2282 vdd3p3.n2235 25.6
R6327 vdd3p3.n1369 vdd3p3.n1368 25.6
R6328 vdd3p3.n1370 vdd3p3.n1369 25.6
R6329 vdd3p3.n1370 vdd3p3.n1360 25.6
R6330 vdd3p3.n1375 vdd3p3.n1360 25.6
R6331 vdd3p3.n1376 vdd3p3.n1375 25.6
R6332 vdd3p3.n1598 vdd3p3.n1597 25.6
R6333 vdd3p3.n1597 vdd3p3.n1009 25.6
R6334 vdd3p3.n1015 vdd3p3.n1009 25.6
R6335 vdd3p3.n1591 vdd3p3.n1015 25.6
R6336 vdd3p3.n1535 vdd3p3.n1534 25.6
R6337 vdd3p3.n1535 vdd3p3.n1040 25.6
R6338 vdd3p3.n1541 vdd3p3.n1040 25.6
R6339 vdd3p3.n1542 vdd3p3.n1541 25.6
R6340 vdd3p3.n1543 vdd3p3.n1542 25.6
R6341 vdd3p3.n1543 vdd3p3.n1036 25.6
R6342 vdd3p3.n1549 vdd3p3.n1036 25.6
R6343 vdd3p3.n1550 vdd3p3.n1549 25.6
R6344 vdd3p3.n1551 vdd3p3.n1550 25.6
R6345 vdd3p3.n1551 vdd3p3.n1032 25.6
R6346 vdd3p3.n1557 vdd3p3.n1032 25.6
R6347 vdd3p3.n1558 vdd3p3.n1557 25.6
R6348 vdd3p3.n1559 vdd3p3.n1558 25.6
R6349 vdd3p3.n1559 vdd3p3.n1028 25.6
R6350 vdd3p3.n1565 vdd3p3.n1028 25.6
R6351 vdd3p3.n1566 vdd3p3.n1565 25.6
R6352 vdd3p3.n1567 vdd3p3.n1566 25.6
R6353 vdd3p3.n1567 vdd3p3.n1024 25.6
R6354 vdd3p3.n1573 vdd3p3.n1024 25.6
R6355 vdd3p3.n1574 vdd3p3.n1573 25.6
R6356 vdd3p3.n1575 vdd3p3.n1574 25.6
R6357 vdd3p3.n1575 vdd3p3.n1020 25.6
R6358 vdd3p3.n1581 vdd3p3.n1020 25.6
R6359 vdd3p3.n1582 vdd3p3.n1581 25.6
R6360 vdd3p3.n1583 vdd3p3.n1582 25.6
R6361 vdd3p3.n1583 vdd3p3.n1016 25.6
R6362 vdd3p3.n1589 vdd3p3.n1016 25.6
R6363 vdd3p3.n1590 vdd3p3.n1589 25.6
R6364 vdd3p3.n1527 vdd3p3.n1525 25.6
R6365 vdd3p3.n1527 vdd3p3.n1526 25.6
R6366 vdd3p3.n1526 vdd3p3.n1044 25.6
R6367 vdd3p3.n1533 vdd3p3.n1044 25.6
R6368 vdd3p3.n955 vdd3p3.n945 25.6
R6369 vdd3p3.n961 vdd3p3.n955 25.6
R6370 vdd3p3.n962 vdd3p3.n961 25.6
R6371 vdd3p3.n962 vdd3p3.n953 25.6
R6372 vdd3p3.n968 vdd3p3.n953 25.6
R6373 vdd3p3.n1450 vdd3p3.n1386 25.6
R6374 vdd3p3.n1444 vdd3p3.n1386 25.6
R6375 vdd3p3.n1444 vdd3p3.n1443 25.6
R6376 vdd3p3.n1443 vdd3p3.n1390 25.6
R6377 vdd3p3.n1437 vdd3p3.n1390 25.6
R6378 vdd3p3.n523 vdd3p3.n522 25.6
R6379 vdd3p3.n524 vdd3p3.n523 25.6
R6380 vdd3p3.n524 vdd3p3.n514 25.6
R6381 vdd3p3.n529 vdd3p3.n514 25.6
R6382 vdd3p3.n530 vdd3p3.n529 25.6
R6383 vdd3p3.n752 vdd3p3.n751 25.6
R6384 vdd3p3.n751 vdd3p3.n163 25.6
R6385 vdd3p3.n169 vdd3p3.n163 25.6
R6386 vdd3p3.n745 vdd3p3.n169 25.6
R6387 vdd3p3.n689 vdd3p3.n688 25.6
R6388 vdd3p3.n689 vdd3p3.n194 25.6
R6389 vdd3p3.n695 vdd3p3.n194 25.6
R6390 vdd3p3.n696 vdd3p3.n695 25.6
R6391 vdd3p3.n697 vdd3p3.n696 25.6
R6392 vdd3p3.n697 vdd3p3.n190 25.6
R6393 vdd3p3.n703 vdd3p3.n190 25.6
R6394 vdd3p3.n704 vdd3p3.n703 25.6
R6395 vdd3p3.n705 vdd3p3.n704 25.6
R6396 vdd3p3.n705 vdd3p3.n186 25.6
R6397 vdd3p3.n711 vdd3p3.n186 25.6
R6398 vdd3p3.n712 vdd3p3.n711 25.6
R6399 vdd3p3.n713 vdd3p3.n712 25.6
R6400 vdd3p3.n713 vdd3p3.n182 25.6
R6401 vdd3p3.n719 vdd3p3.n182 25.6
R6402 vdd3p3.n720 vdd3p3.n719 25.6
R6403 vdd3p3.n721 vdd3p3.n720 25.6
R6404 vdd3p3.n721 vdd3p3.n178 25.6
R6405 vdd3p3.n727 vdd3p3.n178 25.6
R6406 vdd3p3.n728 vdd3p3.n727 25.6
R6407 vdd3p3.n729 vdd3p3.n728 25.6
R6408 vdd3p3.n729 vdd3p3.n174 25.6
R6409 vdd3p3.n735 vdd3p3.n174 25.6
R6410 vdd3p3.n736 vdd3p3.n735 25.6
R6411 vdd3p3.n737 vdd3p3.n736 25.6
R6412 vdd3p3.n737 vdd3p3.n170 25.6
R6413 vdd3p3.n743 vdd3p3.n170 25.6
R6414 vdd3p3.n744 vdd3p3.n743 25.6
R6415 vdd3p3.n681 vdd3p3.n679 25.6
R6416 vdd3p3.n681 vdd3p3.n680 25.6
R6417 vdd3p3.n680 vdd3p3.n198 25.6
R6418 vdd3p3.n687 vdd3p3.n198 25.6
R6419 vdd3p3.n109 vdd3p3.n99 25.6
R6420 vdd3p3.n115 vdd3p3.n109 25.6
R6421 vdd3p3.n116 vdd3p3.n115 25.6
R6422 vdd3p3.n116 vdd3p3.n107 25.6
R6423 vdd3p3.n122 vdd3p3.n107 25.6
R6424 vdd3p3.n604 vdd3p3.n540 25.6
R6425 vdd3p3.n598 vdd3p3.n540 25.6
R6426 vdd3p3.n598 vdd3p3.n597 25.6
R6427 vdd3p3.n597 vdd3p3.n544 25.6
R6428 vdd3p3.n591 vdd3p3.n544 25.6
R6429 vdd3p3.n7509 vdd3p3.n7506 25.6
R6430 vdd3p3.n7506 vdd3p3.n7504 25.6
R6431 vdd3p3.n7504 vdd3p3.n7502 25.6
R6432 vdd3p3.n7502 vdd3p3.n7500 25.6
R6433 vdd3p3.n7500 vdd3p3.n7498 25.6
R6434 vdd3p3.n7498 vdd3p3.n7496 25.6
R6435 vdd3p3.n7496 vdd3p3.n7495 25.6
R6436 vdd3p3.n7495 vdd3p3.n7494 25.6
R6437 vdd3p3.n7494 vdd3p3.n7493 25.6
R6438 vdd3p3.n3911 vdd3p3.n3910 25.6
R6439 vdd3p3.n3912 vdd3p3.n3911 25.6
R6440 vdd3p3.n5181 vdd3p3.n5180 25.6
R6441 vdd3p3.n5182 vdd3p3.n5181 25.6
R6442 vdd3p3.n5183 vdd3p3.n5182 25.6
R6443 vdd3p3.n5184 vdd3p3.n5183 25.6
R6444 vdd3p3.n5185 vdd3p3.n5184 25.6
R6445 vdd3p3.n5186 vdd3p3.n5185 25.6
R6446 vdd3p3.n5188 vdd3p3.n5186 25.6
R6447 vdd3p3.n5190 vdd3p3.n5188 25.6
R6448 vdd3p3.n5192 vdd3p3.n5190 25.6
R6449 vdd3p3.n2860 vdd3p3.n2859 25.35
R6450 vdd3p3.n3093 vdd3p3.n2764 25.35
R6451 vdd3p3.n2014 vdd3p3.n2013 25.35
R6452 vdd3p3.n2247 vdd3p3.n1918 25.35
R6453 vdd3p3.n1169 vdd3p3.n1168 25.35
R6454 vdd3p3.n1402 vdd3p3.n1073 25.35
R6455 vdd3p3.n323 vdd3p3.n322 25.35
R6456 vdd3p3.n556 vdd3p3.n227 25.35
R6457 vdd3p3.n3187 vdd3p3.n3186 25.35
R6458 vdd3p3.n2341 vdd3p3.n2340 25.35
R6459 vdd3p3.n1496 vdd3p3.n1495 25.35
R6460 vdd3p3.n650 vdd3p3.n649 25.35
R6461 vdd3p3.n7465 vdd3p3.n7464 25.35
R6462 vdd3p3.n7021 vdd3p3.n7020 25.35
R6463 vdd3p3.n2977 vdd3p3.n2791 25.35
R6464 vdd3p3.n2978 vdd3p3.n2788 25.35
R6465 vdd3p3.n3165 vdd3p3.n2767 25.35
R6466 vdd3p3.n3190 vdd3p3.n3189 25.35
R6467 vdd3p3.n2884 vdd3p3.n2883 25.35
R6468 vdd3p3.n2879 vdd3p3.n2839 25.35
R6469 vdd3p3.n3338 vdd3p3.n3337 25.35
R6470 vdd3p3.n2131 vdd3p3.n1945 25.35
R6471 vdd3p3.n2132 vdd3p3.n1942 25.35
R6472 vdd3p3.n2319 vdd3p3.n1921 25.35
R6473 vdd3p3.n2344 vdd3p3.n2343 25.35
R6474 vdd3p3.n2038 vdd3p3.n2037 25.35
R6475 vdd3p3.n2033 vdd3p3.n1993 25.35
R6476 vdd3p3.n2492 vdd3p3.n2491 25.35
R6477 vdd3p3.n1286 vdd3p3.n1100 25.35
R6478 vdd3p3.n1287 vdd3p3.n1097 25.35
R6479 vdd3p3.n1474 vdd3p3.n1076 25.35
R6480 vdd3p3.n1499 vdd3p3.n1498 25.35
R6481 vdd3p3.n1193 vdd3p3.n1192 25.35
R6482 vdd3p3.n1188 vdd3p3.n1148 25.35
R6483 vdd3p3.n1647 vdd3p3.n1646 25.35
R6484 vdd3p3.n440 vdd3p3.n254 25.35
R6485 vdd3p3.n441 vdd3p3.n251 25.35
R6486 vdd3p3.n628 vdd3p3.n230 25.35
R6487 vdd3p3.n653 vdd3p3.n652 25.35
R6488 vdd3p3.n347 vdd3p3.n346 25.35
R6489 vdd3p3.n342 vdd3p3.n302 25.35
R6490 vdd3p3.n801 vdd3p3.n800 25.35
R6491 vdd3p3.n8458 vdd3p3.n8457 25.35
R6492 vdd3p3.n8439 vdd3p3.n8438 25.35
R6493 vdd3p3.n7390 vdd3p3.n7389 25.35
R6494 vdd3p3.n7009 vdd3p3.n7008 25.35
R6495 vdd3p3.n5267 vdd3p3.t96 24.811
R6496 vdd3p3.n5275 vdd3p3.n5274 23.97
R6497 vdd3p3.n40 vdd3p3.t139 23.556
R6498 vdd3p3.n900 vdd3p3.t99 23.556
R6499 vdd3p3.n1731 vdd3p3.t152 23.556
R6500 vdd3p3.n2591 vdd3p3.t146 23.556
R6501 vdd3p3.n3391 vdd3p3.n3390 23.47
R6502 vdd3p3.n3074 vdd3p3.n3049 23.076
R6503 vdd3p3.n3073 vdd3p3.n2611 23.076
R6504 vdd3p3.n2640 vdd3p3.n2629 23.076
R6505 vdd3p3.n2228 vdd3p3.n2203 23.076
R6506 vdd3p3.n2227 vdd3p3.n1765 23.076
R6507 vdd3p3.n1794 vdd3p3.n1783 23.076
R6508 vdd3p3.n1383 vdd3p3.n1358 23.076
R6509 vdd3p3.n1382 vdd3p3.n920 23.076
R6510 vdd3p3.n949 vdd3p3.n938 23.076
R6511 vdd3p3.n537 vdd3p3.n512 23.076
R6512 vdd3p3.n536 vdd3p3.n74 23.076
R6513 vdd3p3.n103 vdd3p3.n92 23.076
R6514 vdd3p3.n4190 vdd3p3.n4189 23.051
R6515 vdd3p3.n5086 vdd3p3.n5085 23.051
R6516 vdd3p3.n4903 vdd3p3.n4902 23.051
R6517 vdd3p3.n8531 vdd3p3.n8530 23.051
R6518 vdd3p3.n8876 vdd3p3.n8875 23.051
R6519 vdd3p3.n8793 vdd3p3.n8792 23.051
R6520 vdd3p3.n8721 vdd3p3.n8720 22.709
R6521 vdd3p3.n8646 vdd3p3.t73 22.288
R6522 vdd3p3.n3041 vdd3p3.t0 21.794
R6523 vdd3p3.t133 vdd3p3.n2665 21.794
R6524 vdd3p3.n3344 vdd3p3.t133 21.794
R6525 vdd3p3.n2195 vdd3p3.t75 21.794
R6526 vdd3p3.t169 vdd3p3.n1819 21.794
R6527 vdd3p3.n2498 vdd3p3.t169 21.794
R6528 vdd3p3.n1350 vdd3p3.t22 21.794
R6529 vdd3p3.t117 vdd3p3.n974 21.794
R6530 vdd3p3.n1653 vdd3p3.t117 21.794
R6531 vdd3p3.n504 vdd3p3.t18 21.794
R6532 vdd3p3.t19 vdd3p3.n128 21.794
R6533 vdd3p3.n807 vdd3p3.t19 21.794
R6534 vdd3p3.n36 vdd3p3.n31 21.134
R6535 vdd3p3.n889 vdd3p3.n885 21.134
R6536 vdd3p3.n1727 vdd3p3.n1722 21.134
R6537 vdd3p3.n2580 vdd3p3.n2576 21.134
R6538 vdd3p3.n8029 vdd3p3.n8028 20.718
R6539 vdd3p3.n7522 vdd3p3.n7521 20.718
R6540 vdd3p3.n7522 vdd3p3.n7518 20.718
R6541 vdd3p3.n7522 vdd3p3.n7515 20.718
R6542 vdd3p3.n7522 vdd3p3.n7512 20.718
R6543 vdd3p3.n7522 vdd3p3.n7511 20.718
R6544 vdd3p3.n3290 vdd3p3.n3289 20.603
R6545 vdd3p3.n2444 vdd3p3.n2443 20.603
R6546 vdd3p3.n1599 vdd3p3.n1598 20.603
R6547 vdd3p3.n753 vdd3p3.n752 20.603
R6548 vdd3p3.n3147 vdd3p3.n3049 20.512
R6549 vdd3p3.n3373 vdd3p3.n2611 20.512
R6550 vdd3p3.n3357 vdd3p3.n2629 20.512
R6551 vdd3p3.n2301 vdd3p3.n2203 20.512
R6552 vdd3p3.n2527 vdd3p3.n1765 20.512
R6553 vdd3p3.n2511 vdd3p3.n1783 20.512
R6554 vdd3p3.n1456 vdd3p3.n1358 20.512
R6555 vdd3p3.n1682 vdd3p3.n920 20.512
R6556 vdd3p3.n1666 vdd3p3.n938 20.512
R6557 vdd3p3.n610 vdd3p3.n512 20.512
R6558 vdd3p3.n836 vdd3p3.n74 20.512
R6559 vdd3p3.n820 vdd3p3.n92 20.512
R6560 vdd3p3.n4241 vdd3p3.n4240 19.758
R6561 vdd3p3.n5101 vdd3p3.n5100 19.758
R6562 vdd3p3.n4931 vdd3p3.n4930 19.758
R6563 vdd3p3.n3216 vdd3p3.n3215 18.742
R6564 vdd3p3.n2370 vdd3p3.n2369 18.742
R6565 vdd3p3.n1525 vdd3p3.n1524 18.742
R6566 vdd3p3.n679 vdd3p3.n678 18.742
R6567 vdd3p3.n40 vdd3p3.t116 17.826
R6568 vdd3p3.n900 vdd3p3.t147 17.826
R6569 vdd3p3.n1731 vdd3p3.t29 17.826
R6570 vdd3p3.n2591 vdd3p3.t127 17.826
R6571 vdd3p3.n4718 vdd3p3.n4716 17.824
R6572 vdd3p3.n4036 vdd3p3.n4035 17.62
R6573 vdd3p3.n46 vdd3p3.n32 17.248
R6574 vdd3p3.n898 vdd3p3.n897 17.248
R6575 vdd3p3.n1737 vdd3p3.n1723 17.248
R6576 vdd3p3.n2589 vdd3p3.n2588 17.248
R6577 vdd3p3.n5343 vdd3p3.n5279 17.242
R6578 vdd3p3.n4220 vdd3p3.n4219 16.465
R6579 vdd3p3.n5072 vdd3p3.n5071 16.465
R6580 vdd3p3.n3502 vdd3p3.n3501 16.465
R6581 vdd3p3.n4984 vdd3p3.n4983 16.465
R6582 vdd3p3.n8494 vdd3p3.n8493 16.465
R6583 vdd3p3.n8838 vdd3p3.n8837 16.465
R6584 vdd3p3.n8780 vdd3p3.n8779 16.465
R6585 vdd3p3.n3127 vdd3p3.n2614 15.616
R6586 vdd3p3.n2662 vdd3p3.n2661 15.616
R6587 vdd3p3.n2281 vdd3p3.n1768 15.616
R6588 vdd3p3.n1816 vdd3p3.n1815 15.616
R6589 vdd3p3.n1436 vdd3p3.n923 15.616
R6590 vdd3p3.n971 vdd3p3.n970 15.616
R6591 vdd3p3.n590 vdd3p3.n77 15.616
R6592 vdd3p3.n125 vdd3p3.n124 15.616
R6593 vdd3p3.n4718 vdd3p3.n4717 15.079
R6594 vdd3p3.t0 vdd3p3.n3035 14.743
R6595 vdd3p3.n3147 vdd3p3.t2 14.743
R6596 vdd3p3.n3373 vdd3p3.t162 14.743
R6597 vdd3p3.t130 vdd3p3.n2619 14.743
R6598 vdd3p3.n3364 vdd3p3.t130 14.743
R6599 vdd3p3.n3357 vdd3p3.t128 14.743
R6600 vdd3p3.t75 vdd3p3.n2189 14.743
R6601 vdd3p3.n2301 vdd3p3.t77 14.743
R6602 vdd3p3.n2527 vdd3p3.t110 14.743
R6603 vdd3p3.t15 vdd3p3.n1773 14.743
R6604 vdd3p3.n2518 vdd3p3.t15 14.743
R6605 vdd3p3.n2511 vdd3p3.t170 14.743
R6606 vdd3p3.t22 vdd3p3.n1344 14.743
R6607 vdd3p3.n1456 vdd3p3.t31 14.743
R6608 vdd3p3.n1682 vdd3p3.t165 14.743
R6609 vdd3p3.t118 vdd3p3.n928 14.743
R6610 vdd3p3.n1673 vdd3p3.t118 14.743
R6611 vdd3p3.n1666 vdd3p3.t23 14.743
R6612 vdd3p3.t18 vdd3p3.n498 14.743
R6613 vdd3p3.n610 vdd3p3.t135 14.743
R6614 vdd3p3.n836 vdd3p3.t159 14.743
R6615 vdd3p3.t16 vdd3p3.n82 14.743
R6616 vdd3p3.n827 vdd3p3.t16 14.743
R6617 vdd3p3.n820 vdd3p3.t20 14.743
R6618 vdd3p3.n8028 vdd3p3.n8027 14.25
R6619 vdd3p3.n3127 vdd3p3.n3126 14.208
R6620 vdd3p3.n3348 vdd3p3.n2662 14.208
R6621 vdd3p3.n2281 vdd3p3.n2280 14.208
R6622 vdd3p3.n2502 vdd3p3.n1816 14.208
R6623 vdd3p3.n1436 vdd3p3.n1435 14.208
R6624 vdd3p3.n1657 vdd3p3.n971 14.208
R6625 vdd3p3.n590 vdd3p3.n589 14.208
R6626 vdd3p3.n811 vdd3p3.n125 14.208
R6627 vdd3p3.n2618 vdd3p3.n2617 14.102
R6628 vdd3p3.n3367 vdd3p3.n2619 14.102
R6629 vdd3p3.n3364 vdd3p3.n3363 14.102
R6630 vdd3p3.n2630 vdd3p3.n2622 14.102
R6631 vdd3p3.n1772 vdd3p3.n1771 14.102
R6632 vdd3p3.n2521 vdd3p3.n1773 14.102
R6633 vdd3p3.n2518 vdd3p3.n2517 14.102
R6634 vdd3p3.n1784 vdd3p3.n1776 14.102
R6635 vdd3p3.n927 vdd3p3.n926 14.102
R6636 vdd3p3.n1676 vdd3p3.n928 14.102
R6637 vdd3p3.n1673 vdd3p3.n1672 14.102
R6638 vdd3p3.n939 vdd3p3.n931 14.102
R6639 vdd3p3.n81 vdd3p3.n80 14.102
R6640 vdd3p3.n830 vdd3p3.n82 14.102
R6641 vdd3p3.n827 vdd3p3.n826 14.102
R6642 vdd3p3.n93 vdd3p3.n85 14.102
R6643 vdd3p3.t92 vdd3p3.n6554 13.877
R6644 vdd3p3.n8727 vdd3p3.n8726 13.877
R6645 vdd3p3.n2665 vdd3p3.n2641 13.461
R6646 vdd3p3.n1819 vdd3p3.n1795 13.461
R6647 vdd3p3.n974 vdd3p3.n950 13.461
R6648 vdd3p3.n128 vdd3p3.n104 13.461
R6649 vdd3p3.t106 vdd3p3.n6561 13.036
R6650 vdd3p3.t120 vdd3p3.n6 12.788
R6651 vdd3p3.n867 vdd3p3.t155 12.788
R6652 vdd3p3.t11 vdd3p3.n1697 12.788
R6653 vdd3p3.n2558 vdd3p3.t81 12.788
R6654 vdd3p3.n4687 vdd3p3.n4684 12.688
R6655 vdd3p3.n7523 vdd3p3.n7522 12.666
R6656 vdd3p3.n3393 vdd3p3.n3392 12.134
R6657 vdd3p3.n5729 vdd3p3.n5728 12.063
R6658 vdd3p3.n3121 vdd3p3.n2753 12.032
R6659 vdd3p3.n3314 vdd3p3.n2663 12.032
R6660 vdd3p3.n2275 vdd3p3.n1907 12.032
R6661 vdd3p3.n2468 vdd3p3.n1817 12.032
R6662 vdd3p3.n1430 vdd3p3.n1062 12.032
R6663 vdd3p3.n1623 vdd3p3.n972 12.032
R6664 vdd3p3.n584 vdd3p3.n216 12.032
R6665 vdd3p3.n777 vdd3p3.n126 12.032
R6666 vdd3p3.n5274 vdd3p3.t145 11.897
R6667 vdd3p3.n3840 vdd3p3.n3839 11.67
R6668 vdd3p3.n5343 vdd3p3.n5272 11.354
R6669 vdd3p3.n6663 vdd3p3.t97 11.354
R6670 vdd3p3.n3387 vdd3p3.n3386 11.118
R6671 vdd3p3.n5022 vdd3p3.n5021 10.892
R6672 vdd3p3.n4721 vdd3p3.n4720 10.892
R6673 vdd3p3.n3053 vdd3p3.n3046 10.41
R6674 vdd3p3.n3054 vdd3p3.n3053 10.41
R6675 vdd3p3.n2207 vdd3p3.n2200 10.41
R6676 vdd3p3.n2208 vdd3p3.n2207 10.41
R6677 vdd3p3.n1362 vdd3p3.n1355 10.41
R6678 vdd3p3.n1363 vdd3p3.n1362 10.41
R6679 vdd3p3.n516 vdd3p3.n509 10.41
R6680 vdd3p3.n517 vdd3p3.n516 10.41
R6681 vdd3p3.n4209 vdd3p3.n4208 9.879
R6682 vdd3p3.n5061 vdd3p3.n5060 9.879
R6683 vdd3p3.n3486 vdd3p3.n3485 9.879
R6684 vdd3p3.n4968 vdd3p3.n4967 9.879
R6685 vdd3p3.n8515 vdd3p3.n8514 9.879
R6686 vdd3p3.n8859 vdd3p3.n8858 9.879
R6687 vdd3p3.n8770 vdd3p3.n8769 9.879
R6688 vdd3p3.n6633 vdd3p3.t8 9.672
R6689 vdd3p3.n8722 vdd3p3.n8721 9.672
R6690 vdd3p3.n4202 vdd3p3.n4201 9.3
R6691 vdd3p3.n4213 vdd3p3.n4212 9.3
R6692 vdd3p3.n4226 vdd3p3.n4225 9.3
R6693 vdd3p3.n4200 vdd3p3.n4199 9.3
R6694 vdd3p3.n4199 vdd3p3.n4198 9.3
R6695 vdd3p3.n4204 vdd3p3.n4203 9.3
R6696 vdd3p3.n4211 vdd3p3.n4210 9.3
R6697 vdd3p3.n4210 vdd3p3.n4209 9.3
R6698 vdd3p3.n4215 vdd3p3.n4214 9.3
R6699 vdd3p3.n4222 vdd3p3.n4221 9.3
R6700 vdd3p3.n4221 vdd3p3.n4220 9.3
R6701 vdd3p3.n4224 vdd3p3.n4223 9.3
R6702 vdd3p3.n4183 vdd3p3.n4182 9.3
R6703 vdd3p3.n4191 vdd3p3.n4190 9.3
R6704 vdd3p3.n4281 vdd3p3.n4280 9.3
R6705 vdd3p3.n4283 vdd3p3.n4282 9.3
R6706 vdd3p3.n4279 vdd3p3.n4278 9.3
R6707 vdd3p3.n4278 vdd3p3.n4277 9.3
R6708 vdd3p3.n4267 vdd3p3.n4266 9.3
R6709 vdd3p3.n4265 vdd3p3.n4264 9.3
R6710 vdd3p3.n4263 vdd3p3.n4262 9.3
R6711 vdd3p3.n4262 vdd3p3.n4261 9.3
R6712 vdd3p3.n4291 vdd3p3.n4290 9.3
R6713 vdd3p3.n4298 vdd3p3.n4297 9.3
R6714 vdd3p3.n4305 vdd3p3.n4304 9.3
R6715 vdd3p3.n4312 vdd3p3.n4311 9.3
R6716 vdd3p3.n4319 vdd3p3.n4318 9.3
R6717 vdd3p3.n4326 vdd3p3.n4325 9.3
R6718 vdd3p3.n4332 vdd3p3.n4331 9.3
R6719 vdd3p3.n4339 vdd3p3.n4338 9.3
R6720 vdd3p3.n4346 vdd3p3.n4345 9.3
R6721 vdd3p3.n4348 vdd3p3.n4347 9.3
R6722 vdd3p3.n4344 vdd3p3.n4343 9.3
R6723 vdd3p3.n4341 vdd3p3.n4340 9.3
R6724 vdd3p3.n4337 vdd3p3.n4336 9.3
R6725 vdd3p3.n4334 vdd3p3.n4333 9.3
R6726 vdd3p3.n4330 vdd3p3.n4329 9.3
R6727 vdd3p3.n4328 vdd3p3.n4327 9.3
R6728 vdd3p3.n4324 vdd3p3.n4323 9.3
R6729 vdd3p3.n4322 vdd3p3.n4321 9.3
R6730 vdd3p3.n4317 vdd3p3.n4316 9.3
R6731 vdd3p3.n4315 vdd3p3.n4314 9.3
R6732 vdd3p3.n4310 vdd3p3.n4309 9.3
R6733 vdd3p3.n4308 vdd3p3.n4307 9.3
R6734 vdd3p3.n4303 vdd3p3.n4302 9.3
R6735 vdd3p3.n4301 vdd3p3.n4300 9.3
R6736 vdd3p3.n4296 vdd3p3.n4295 9.3
R6737 vdd3p3.n4294 vdd3p3.n4293 9.3
R6738 vdd3p3.n4289 vdd3p3.n4288 9.3
R6739 vdd3p3.n4601 vdd3p3.n4600 9.3
R6740 vdd3p3.n4603 vdd3p3.n4602 9.3
R6741 vdd3p3.n4599 vdd3p3.n4598 9.3
R6742 vdd3p3.n4598 vdd3p3.n4597 9.3
R6743 vdd3p3.n4587 vdd3p3.n4586 9.3
R6744 vdd3p3.n4585 vdd3p3.n4584 9.3
R6745 vdd3p3.n4583 vdd3p3.n4582 9.3
R6746 vdd3p3.n4582 vdd3p3.n4581 9.3
R6747 vdd3p3.n4611 vdd3p3.n4610 9.3
R6748 vdd3p3.n4618 vdd3p3.n4617 9.3
R6749 vdd3p3.n4625 vdd3p3.n4624 9.3
R6750 vdd3p3.n4632 vdd3p3.n4631 9.3
R6751 vdd3p3.n4639 vdd3p3.n4638 9.3
R6752 vdd3p3.n4646 vdd3p3.n4645 9.3
R6753 vdd3p3.n4652 vdd3p3.n4651 9.3
R6754 vdd3p3.n4659 vdd3p3.n4658 9.3
R6755 vdd3p3.n4666 vdd3p3.n4665 9.3
R6756 vdd3p3.n4668 vdd3p3.n4667 9.3
R6757 vdd3p3.n4664 vdd3p3.n4663 9.3
R6758 vdd3p3.n4661 vdd3p3.n4660 9.3
R6759 vdd3p3.n4657 vdd3p3.n4656 9.3
R6760 vdd3p3.n4654 vdd3p3.n4653 9.3
R6761 vdd3p3.n4650 vdd3p3.n4649 9.3
R6762 vdd3p3.n4648 vdd3p3.n4647 9.3
R6763 vdd3p3.n4644 vdd3p3.n4643 9.3
R6764 vdd3p3.n4642 vdd3p3.n4641 9.3
R6765 vdd3p3.n4637 vdd3p3.n4636 9.3
R6766 vdd3p3.n4635 vdd3p3.n4634 9.3
R6767 vdd3p3.n4630 vdd3p3.n4629 9.3
R6768 vdd3p3.n4628 vdd3p3.n4627 9.3
R6769 vdd3p3.n4623 vdd3p3.n4622 9.3
R6770 vdd3p3.n4621 vdd3p3.n4620 9.3
R6771 vdd3p3.n4616 vdd3p3.n4615 9.3
R6772 vdd3p3.n4614 vdd3p3.n4613 9.3
R6773 vdd3p3.n4609 vdd3p3.n4608 9.3
R6774 vdd3p3.n5076 vdd3p3.n5075 9.3
R6775 vdd3p3.n5065 vdd3p3.n5064 9.3
R6776 vdd3p3.n5054 vdd3p3.n5053 9.3
R6777 vdd3p3.n5052 vdd3p3.n5051 9.3
R6778 vdd3p3.n5051 vdd3p3.n5050 9.3
R6779 vdd3p3.n5056 vdd3p3.n5055 9.3
R6780 vdd3p3.n5063 vdd3p3.n5062 9.3
R6781 vdd3p3.n5062 vdd3p3.n5061 9.3
R6782 vdd3p3.n5067 vdd3p3.n5066 9.3
R6783 vdd3p3.n5074 vdd3p3.n5073 9.3
R6784 vdd3p3.n5073 vdd3p3.n5072 9.3
R6785 vdd3p3.n5078 vdd3p3.n5077 9.3
R6786 vdd3p3.n5043 vdd3p3.n5042 9.3
R6787 vdd3p3.n5087 vdd3p3.n5086 9.3
R6788 vdd3p3.n3664 vdd3p3.n3663 9.3
R6789 vdd3p3.n3657 vdd3p3.n3656 9.3
R6790 vdd3p3.n3650 vdd3p3.n3649 9.3
R6791 vdd3p3.n3648 vdd3p3.n3647 9.3
R6792 vdd3p3.n3653 vdd3p3.n3652 9.3
R6793 vdd3p3.n3655 vdd3p3.n3654 9.3
R6794 vdd3p3.n3660 vdd3p3.n3659 9.3
R6795 vdd3p3.n3662 vdd3p3.n3661 9.3
R6796 vdd3p3.n3735 vdd3p3.n3734 9.3
R6797 vdd3p3.n3733 vdd3p3.n3732 9.3
R6798 vdd3p3.n3721 vdd3p3.n3720 9.3
R6799 vdd3p3.n3731 vdd3p3.n3730 9.3
R6800 vdd3p3.n3724 vdd3p3.n3723 9.3
R6801 vdd3p3.n3719 vdd3p3.n3718 9.3
R6802 vdd3p3.n3726 vdd3p3.n3725 9.3
R6803 vdd3p3.n3728 vdd3p3.n3727 9.3
R6804 vdd3p3.n3640 vdd3p3.n3639 9.3
R6805 vdd3p3.n3621 vdd3p3.n3620 9.3
R6806 vdd3p3.n3642 vdd3p3.n3641 9.3
R6807 vdd3p3.n3638 vdd3p3.n3637 9.3
R6808 vdd3p3.n3637 vdd3p3.n3636 9.3
R6809 vdd3p3.n3628 vdd3p3.n3627 9.3
R6810 vdd3p3.n3627 vdd3p3.n3626 9.3
R6811 vdd3p3.n3619 vdd3p3.n3618 9.3
R6812 vdd3p3.n3711 vdd3p3.n3710 9.3
R6813 vdd3p3.n3713 vdd3p3.n3712 9.3
R6814 vdd3p3.n3709 vdd3p3.n3708 9.3
R6815 vdd3p3.n3708 vdd3p3.n3707 9.3
R6816 vdd3p3.n3614 vdd3p3.n3613 9.3
R6817 vdd3p3.n3545 vdd3p3.n3544 9.3
R6818 vdd3p3.n3529 vdd3p3.n3528 9.3
R6819 vdd3p3.n3527 vdd3p3.n3526 9.3
R6820 vdd3p3.n3525 vdd3p3.n3524 9.3
R6821 vdd3p3.n3524 vdd3p3.n3523 9.3
R6822 vdd3p3.n3543 vdd3p3.n3542 9.3
R6823 vdd3p3.n3541 vdd3p3.n3540 9.3
R6824 vdd3p3.n3540 vdd3p3.n3539 9.3
R6825 vdd3p3.n3612 vdd3p3.n3611 9.3
R6826 vdd3p3.n3610 vdd3p3.n3609 9.3
R6827 vdd3p3.n3609 vdd3p3.n3608 9.3
R6828 vdd3p3.n3554 vdd3p3.n3553 9.3
R6829 vdd3p3.n3561 vdd3p3.n3560 9.3
R6830 vdd3p3.n3568 vdd3p3.n3567 9.3
R6831 vdd3p3.n3552 vdd3p3.n3551 9.3
R6832 vdd3p3.n3557 vdd3p3.n3556 9.3
R6833 vdd3p3.n3559 vdd3p3.n3558 9.3
R6834 vdd3p3.n3564 vdd3p3.n3563 9.3
R6835 vdd3p3.n3566 vdd3p3.n3565 9.3
R6836 vdd3p3.n3479 vdd3p3.n3478 9.3
R6837 vdd3p3.n3481 vdd3p3.n3480 9.3
R6838 vdd3p3.n3477 vdd3p3.n3476 9.3
R6839 vdd3p3.n3476 vdd3p3.n3475 9.3
R6840 vdd3p3.n3503 vdd3p3.n3502 9.3
R6841 vdd3p3.n3487 vdd3p3.n3486 9.3
R6842 vdd3p3.n4776 vdd3p3.n4775 9.3
R6843 vdd3p3.n4774 vdd3p3.n4773 9.3
R6844 vdd3p3.n4773 vdd3p3.n4772 9.3
R6845 vdd3p3.n4778 vdd3p3.n4777 9.3
R6846 vdd3p3.n4800 vdd3p3.n4799 9.3
R6847 vdd3p3.n4798 vdd3p3.n4797 9.3
R6848 vdd3p3.n4786 vdd3p3.n4785 9.3
R6849 vdd3p3.n4796 vdd3p3.n4795 9.3
R6850 vdd3p3.n4789 vdd3p3.n4788 9.3
R6851 vdd3p3.n4784 vdd3p3.n4783 9.3
R6852 vdd3p3.n4791 vdd3p3.n4790 9.3
R6853 vdd3p3.n4793 vdd3p3.n4792 9.3
R6854 vdd3p3.n4961 vdd3p3.n4960 9.3
R6855 vdd3p3.n4959 vdd3p3.n4958 9.3
R6856 vdd3p3.n4958 vdd3p3.n4957 9.3
R6857 vdd3p3.n4963 vdd3p3.n4962 9.3
R6858 vdd3p3.n4917 vdd3p3.n4916 9.3
R6859 vdd3p3.n4915 vdd3p3.n4914 9.3
R6860 vdd3p3.n4914 vdd3p3.n4913 9.3
R6861 vdd3p3.n4919 vdd3p3.n4918 9.3
R6862 vdd3p3.n4927 vdd3p3.n4926 9.3
R6863 vdd3p3.n4938 vdd3p3.n4937 9.3
R6864 vdd3p3.n4949 vdd3p3.n4948 9.3
R6865 vdd3p3.n4947 vdd3p3.n4946 9.3
R6866 vdd3p3.n4945 vdd3p3.n4944 9.3
R6867 vdd3p3.n4944 vdd3p3.n4943 9.3
R6868 vdd3p3.n4936 vdd3p3.n4935 9.3
R6869 vdd3p3.n4934 vdd3p3.n4933 9.3
R6870 vdd3p3.n4933 vdd3p3.n4932 9.3
R6871 vdd3p3.n4925 vdd3p3.n4924 9.3
R6872 vdd3p3.n4904 vdd3p3.n4903 9.3
R6873 vdd3p3.n4969 vdd3p3.n4968 9.3
R6874 vdd3p3.n4985 vdd3p3.n4984 9.3
R6875 vdd3p3.n8508 vdd3p3.n8507 9.3
R6876 vdd3p3.n8506 vdd3p3.n8505 9.3
R6877 vdd3p3.n8505 vdd3p3.n8504 9.3
R6878 vdd3p3.n8510 vdd3p3.n8509 9.3
R6879 vdd3p3.n8517 vdd3p3.n8516 9.3
R6880 vdd3p3.n8516 vdd3p3.n8515 9.3
R6881 vdd3p3.n8519 vdd3p3.n8518 9.3
R6882 vdd3p3.n8532 vdd3p3.n8531 9.3
R6883 vdd3p3.n8551 vdd3p3.n8550 9.3
R6884 vdd3p3.n8521 vdd3p3.n8520 9.3
R6885 vdd3p3.n8495 vdd3p3.n8494 9.3
R6886 vdd3p3.n8852 vdd3p3.n8851 9.3
R6887 vdd3p3.n8850 vdd3p3.n8849 9.3
R6888 vdd3p3.n8849 vdd3p3.n8848 9.3
R6889 vdd3p3.n8854 vdd3p3.n8853 9.3
R6890 vdd3p3.n8861 vdd3p3.n8860 9.3
R6891 vdd3p3.n8860 vdd3p3.n8859 9.3
R6892 vdd3p3.n8863 vdd3p3.n8862 9.3
R6893 vdd3p3.n8877 vdd3p3.n8876 9.3
R6894 vdd3p3.n8630 vdd3p3.n8629 9.3
R6895 vdd3p3.n8865 vdd3p3.n8864 9.3
R6896 vdd3p3.n8839 vdd3p3.n8838 9.3
R6897 vdd3p3.n8774 vdd3p3.n8773 9.3
R6898 vdd3p3.n8763 vdd3p3.n8762 9.3
R6899 vdd3p3.n8772 vdd3p3.n8771 9.3
R6900 vdd3p3.n8771 vdd3p3.n8770 9.3
R6901 vdd3p3.n8761 vdd3p3.n8760 9.3
R6902 vdd3p3.n8760 vdd3p3.n8759 9.3
R6903 vdd3p3.n8765 vdd3p3.n8764 9.3
R6904 vdd3p3.n8776 vdd3p3.n8775 9.3
R6905 vdd3p3.n8813 vdd3p3.n8812 9.3
R6906 vdd3p3.n8794 vdd3p3.n8793 9.3
R6907 vdd3p3.n8781 vdd3p3.n8780 9.3
R6908 vdd3p3.n3844 vdd3p3.n3843 9.3
R6909 vdd3p3.n3847 vdd3p3.n3846 9.3
R6910 vdd3p3.n3835 vdd3p3.n3834 9.3
R6911 vdd3p3.n3184 vdd3p3.n3018 8.96
R6912 vdd3p3.n2840 vdd3p3.n2627 8.96
R6913 vdd3p3.n2338 vdd3p3.n2172 8.96
R6914 vdd3p3.n1994 vdd3p3.n1781 8.96
R6915 vdd3p3.n1493 vdd3p3.n1327 8.96
R6916 vdd3p3.n1149 vdd3p3.n936 8.96
R6917 vdd3p3.n647 vdd3p3.n481 8.96
R6918 vdd3p3.n303 vdd3p3.n90 8.96
R6919 vdd3p3.n35 vdd3p3.n34 8.855
R6920 vdd3p3.n52 vdd3p3.n51 8.855
R6921 vdd3p3.n50 vdd3p3.n33 8.855
R6922 vdd3p3.n39 vdd3p3.n38 8.855
R6923 vdd3p3.n16 vdd3p3.n15 8.855
R6924 vdd3p3.n8 vdd3p3.n7 8.855
R6925 vdd3p3.n7 vdd3p3.n6 8.855
R6926 vdd3p3.n28 vdd3p3.n27 8.855
R6927 vdd3p3.n29 vdd3p3.n28 8.855
R6928 vdd3p3.n5 vdd3p3.n4 8.855
R6929 vdd3p3.n30 vdd3p3.n5 8.855
R6930 vdd3p3.n58 vdd3p3.n57 8.855
R6931 vdd3p3.n57 vdd3p3.n56 8.855
R6932 vdd3p3.n888 vdd3p3.n887 8.855
R6933 vdd3p3.n894 vdd3p3.n893 8.855
R6934 vdd3p3.n892 vdd3p3.n886 8.855
R6935 vdd3p3.n848 vdd3p3.n847 8.855
R6936 vdd3p3.n866 vdd3p3.n865 8.855
R6937 vdd3p3.n857 vdd3p3.n856 8.855
R6938 vdd3p3.n867 vdd3p3.n857 8.855
R6939 vdd3p3.n870 vdd3p3.n869 8.855
R6940 vdd3p3.n869 vdd3p3.n868 8.855
R6941 vdd3p3.n851 vdd3p3.n850 8.855
R6942 vdd3p3.n850 vdd3p3.n849 8.855
R6943 vdd3p3.n882 vdd3p3.n881 8.855
R6944 vdd3p3.n883 vdd3p3.n882 8.855
R6945 vdd3p3.n1726 vdd3p3.n1725 8.855
R6946 vdd3p3.n1743 vdd3p3.n1742 8.855
R6947 vdd3p3.n1741 vdd3p3.n1724 8.855
R6948 vdd3p3.n1730 vdd3p3.n1729 8.855
R6949 vdd3p3.n1707 vdd3p3.n1706 8.855
R6950 vdd3p3.n1699 vdd3p3.n1698 8.855
R6951 vdd3p3.n1698 vdd3p3.n1697 8.855
R6952 vdd3p3.n1719 vdd3p3.n1718 8.855
R6953 vdd3p3.n1720 vdd3p3.n1719 8.855
R6954 vdd3p3.n1696 vdd3p3.n1695 8.855
R6955 vdd3p3.n1721 vdd3p3.n1696 8.855
R6956 vdd3p3.n1749 vdd3p3.n1748 8.855
R6957 vdd3p3.n1748 vdd3p3.n1747 8.855
R6958 vdd3p3.n2579 vdd3p3.n2578 8.855
R6959 vdd3p3.n2585 vdd3p3.n2584 8.855
R6960 vdd3p3.n2583 vdd3p3.n2577 8.855
R6961 vdd3p3.n2539 vdd3p3.n2538 8.855
R6962 vdd3p3.n2557 vdd3p3.n2556 8.855
R6963 vdd3p3.n2548 vdd3p3.n2547 8.855
R6964 vdd3p3.n2558 vdd3p3.n2548 8.855
R6965 vdd3p3.n2561 vdd3p3.n2560 8.855
R6966 vdd3p3.n2560 vdd3p3.n2559 8.855
R6967 vdd3p3.n2542 vdd3p3.n2541 8.855
R6968 vdd3p3.n2541 vdd3p3.n2540 8.855
R6969 vdd3p3.n2573 vdd3p3.n2572 8.855
R6970 vdd3p3.n2574 vdd3p3.n2573 8.855
R6971 vdd3p3.n3630 vdd3p3.n3629 8.764
R6972 vdd3p3.n3533 vdd3p3.n3532 8.764
R6973 vdd3p3.n3122 vdd3p3.n3121 8.704
R6974 vdd3p3.n3123 vdd3p3.n3122 8.704
R6975 vdd3p3.n3126 vdd3p3.n3123 8.704
R6976 vdd3p3.n3371 vdd3p3.n2614 8.704
R6977 vdd3p3.n3371 vdd3p3.n3370 8.704
R6978 vdd3p3.n3370 vdd3p3.n3369 8.704
R6979 vdd3p3.n3369 vdd3p3.n2615 8.704
R6980 vdd3p3.n2661 vdd3p3.n2615 8.704
R6981 vdd3p3.n3348 vdd3p3.n3347 8.704
R6982 vdd3p3.n3347 vdd3p3.n3346 8.704
R6983 vdd3p3.n3346 vdd3p3.n2663 8.704
R6984 vdd3p3.n2276 vdd3p3.n2275 8.704
R6985 vdd3p3.n2277 vdd3p3.n2276 8.704
R6986 vdd3p3.n2280 vdd3p3.n2277 8.704
R6987 vdd3p3.n2525 vdd3p3.n1768 8.704
R6988 vdd3p3.n2525 vdd3p3.n2524 8.704
R6989 vdd3p3.n2524 vdd3p3.n2523 8.704
R6990 vdd3p3.n2523 vdd3p3.n1769 8.704
R6991 vdd3p3.n1815 vdd3p3.n1769 8.704
R6992 vdd3p3.n2502 vdd3p3.n2501 8.704
R6993 vdd3p3.n2501 vdd3p3.n2500 8.704
R6994 vdd3p3.n2500 vdd3p3.n1817 8.704
R6995 vdd3p3.n1431 vdd3p3.n1430 8.704
R6996 vdd3p3.n1432 vdd3p3.n1431 8.704
R6997 vdd3p3.n1435 vdd3p3.n1432 8.704
R6998 vdd3p3.n1680 vdd3p3.n923 8.704
R6999 vdd3p3.n1680 vdd3p3.n1679 8.704
R7000 vdd3p3.n1679 vdd3p3.n1678 8.704
R7001 vdd3p3.n1678 vdd3p3.n924 8.704
R7002 vdd3p3.n970 vdd3p3.n924 8.704
R7003 vdd3p3.n1657 vdd3p3.n1656 8.704
R7004 vdd3p3.n1656 vdd3p3.n1655 8.704
R7005 vdd3p3.n1655 vdd3p3.n972 8.704
R7006 vdd3p3.n585 vdd3p3.n584 8.704
R7007 vdd3p3.n586 vdd3p3.n585 8.704
R7008 vdd3p3.n589 vdd3p3.n586 8.704
R7009 vdd3p3.n834 vdd3p3.n77 8.704
R7010 vdd3p3.n834 vdd3p3.n833 8.704
R7011 vdd3p3.n833 vdd3p3.n832 8.704
R7012 vdd3p3.n832 vdd3p3.n78 8.704
R7013 vdd3p3.n124 vdd3p3.n78 8.704
R7014 vdd3p3.n811 vdd3p3.n810 8.704
R7015 vdd3p3.n810 vdd3p3.n809 8.704
R7016 vdd3p3.n809 vdd3p3.n126 8.704
R7017 vdd3p3.n8455 vdd3p3.n8450 8.464
R7018 vdd3p3.n4730 vdd3p3.n4729 8.45
R7019 vdd3p3.n8698 vdd3p3.n8697 8.45
R7020 vdd3p3.n3990 vdd3p3.n3989 8.45
R7021 vdd3p3.n3995 vdd3p3.n3992 8.45
R7022 vdd3p3.n3461 vdd3p3.n3460 8.45
R7023 vdd3p3.n8653 vdd3p3.n8652 8.409
R7024 vdd3p3.n53 vdd3p3.n33 8.394
R7025 vdd3p3.n53 vdd3p3.n52 8.394
R7026 vdd3p3.n38 vdd3p3.n32 8.394
R7027 vdd3p3.n895 vdd3p3.n886 8.394
R7028 vdd3p3.n895 vdd3p3.n894 8.394
R7029 vdd3p3.n897 vdd3p3.n848 8.394
R7030 vdd3p3.n1744 vdd3p3.n1724 8.394
R7031 vdd3p3.n1744 vdd3p3.n1743 8.394
R7032 vdd3p3.n1729 vdd3p3.n1723 8.394
R7033 vdd3p3.n2586 vdd3p3.n2577 8.394
R7034 vdd3p3.n2586 vdd3p3.n2585 8.394
R7035 vdd3p3.n2588 vdd3p3.n2539 8.394
R7036 vdd3p3.n34 vdd3p3.n31 8.394
R7037 vdd3p3.n887 vdd3p3.n885 8.394
R7038 vdd3p3.n1725 vdd3p3.n1722 8.394
R7039 vdd3p3.n2578 vdd3p3.n2576 8.394
R7040 vdd3p3.n3915 vdd3p3.n3914 8.067
R7041 vdd3p3.n3965 vdd3p3.n3964 8.067
R7042 vdd3p3.n3969 vdd3p3.n3968 8.067
R7043 vdd3p3.n3894 vdd3p3.n3891 8.067
R7044 vdd3p3.n3890 vdd3p3.n3887 8.067
R7045 vdd3p3.n3886 vdd3p3.n3883 8.067
R7046 vdd3p3.n3882 vdd3p3.n3879 8.067
R7047 vdd3p3.n4011 vdd3p3.n4010 8.067
R7048 vdd3p3.n4015 vdd3p3.n4014 8.067
R7049 vdd3p3.n4033 vdd3p3.n4030 8.067
R7050 vdd3p3.n4029 vdd3p3.n4026 8.067
R7051 vdd3p3.n4025 vdd3p3.n4022 8.067
R7052 vdd3p3.n4041 vdd3p3.n4040 8.067
R7053 vdd3p3.n4045 vdd3p3.n4044 8.067
R7054 vdd3p3.n4049 vdd3p3.n4048 8.067
R7055 vdd3p3.n4053 vdd3p3.n4052 8.067
R7056 vdd3p3.n4144 vdd3p3.n4141 8.067
R7057 vdd3p3.n4140 vdd3p3.n4137 8.067
R7058 vdd3p3.n4136 vdd3p3.n4133 8.067
R7059 vdd3p3.n4132 vdd3p3.n4129 8.067
R7060 vdd3p3.n4128 vdd3p3.n4125 8.067
R7061 vdd3p3.n4120 vdd3p3.n4117 8.067
R7062 vdd3p3.n4116 vdd3p3.n4113 8.067
R7063 vdd3p3.n4112 vdd3p3.n4109 8.067
R7064 vdd3p3.n4108 vdd3p3.n4105 8.067
R7065 vdd3p3.n4104 vdd3p3.n4101 8.067
R7066 vdd3p3.n4100 vdd3p3.n4097 8.067
R7067 vdd3p3.n4096 vdd3p3.n4093 8.067
R7068 vdd3p3.n4092 vdd3p3.n4089 8.067
R7069 vdd3p3.n4088 vdd3p3.n4085 8.067
R7070 vdd3p3.n4084 vdd3p3.n4081 8.067
R7071 vdd3p3.n4080 vdd3p3.n4077 8.067
R7072 vdd3p3.n4076 vdd3p3.n4073 8.067
R7073 vdd3p3.n8450 vdd3p3.n8449 8.067
R7074 vdd3p3.n6555 vdd3p3.t100 7.99
R7075 vdd3p3.n4260 vdd3p3.n4259 7.453
R7076 vdd3p3.n4276 vdd3p3.n4275 7.453
R7077 vdd3p3.n4580 vdd3p3.n4579 7.453
R7078 vdd3p3.n4596 vdd3p3.n4595 7.453
R7079 vdd3p3.n3522 vdd3p3.n3521 7.453
R7080 vdd3p3.n3538 vdd3p3.n3537 7.453
R7081 vdd3p3.n3607 vdd3p3.n3606 7.453
R7082 vdd3p3.n3706 vdd3p3.n3705 7.453
R7083 vdd3p3.n3635 vdd3p3.n3634 7.453
R7084 vdd3p3.n3625 vdd3p3.n3624 7.453
R7085 vdd3p3.n4771 vdd3p3.n4770 7.453
R7086 vdd3p3.n4912 vdd3p3.n4911 7.453
R7087 vdd3p3.n3984 vdd3p3.n3983 7.424
R7088 vdd3p3.n4724 vdd3p3.n4723 7.389
R7089 vdd3p3.n5008 vdd3p3.n5007 7.172
R7090 vdd3p3.n6457 vdd3p3.t102 7.149
R7091 vdd3p3.n2606 vdd3p3.n2605 7.088
R7092 vdd3p3.n3378 vdd3p3.n2602 7.088
R7093 vdd3p3.n1760 vdd3p3.n1759 7.088
R7094 vdd3p3.n2532 vdd3p3.n1756 7.088
R7095 vdd3p3.n915 vdd3p3.n914 7.088
R7096 vdd3p3.n1687 vdd3p3.n911 7.088
R7097 vdd3p3.n69 vdd3p3.n68 7.088
R7098 vdd3p3.n841 vdd3p3.n65 7.088
R7099 vdd3p3.n2975 vdd3p3.n2793 7.076
R7100 vdd3p3.n2969 vdd3p3.n2793 7.076
R7101 vdd3p3.n2969 vdd3p3.n2968 7.076
R7102 vdd3p3.n2968 vdd3p3.n2967 7.076
R7103 vdd3p3.n2967 vdd3p3.n2797 7.076
R7104 vdd3p3.n2961 vdd3p3.n2797 7.076
R7105 vdd3p3.n2961 vdd3p3.n2960 7.076
R7106 vdd3p3.n2960 vdd3p3.n2959 7.076
R7107 vdd3p3.n2959 vdd3p3.n2801 7.076
R7108 vdd3p3.n2953 vdd3p3.n2801 7.076
R7109 vdd3p3.n2953 vdd3p3.n2952 7.076
R7110 vdd3p3.n2952 vdd3p3.n2951 7.076
R7111 vdd3p3.n2951 vdd3p3.n2805 7.076
R7112 vdd3p3.n2945 vdd3p3.n2805 7.076
R7113 vdd3p3.n2945 vdd3p3.n2944 7.076
R7114 vdd3p3.n2944 vdd3p3.n2943 7.076
R7115 vdd3p3.n2943 vdd3p3.n2809 7.076
R7116 vdd3p3.n2937 vdd3p3.n2809 7.076
R7117 vdd3p3.n2937 vdd3p3.n2936 7.076
R7118 vdd3p3.n2936 vdd3p3.n2935 7.076
R7119 vdd3p3.n2935 vdd3p3.n2813 7.076
R7120 vdd3p3.n2929 vdd3p3.n2813 7.076
R7121 vdd3p3.n2929 vdd3p3.n2928 7.076
R7122 vdd3p3.n2928 vdd3p3.n2927 7.076
R7123 vdd3p3.n2927 vdd3p3.n2817 7.076
R7124 vdd3p3.n2129 vdd3p3.n1947 7.076
R7125 vdd3p3.n2123 vdd3p3.n1947 7.076
R7126 vdd3p3.n2123 vdd3p3.n2122 7.076
R7127 vdd3p3.n2122 vdd3p3.n2121 7.076
R7128 vdd3p3.n2121 vdd3p3.n1951 7.076
R7129 vdd3p3.n2115 vdd3p3.n1951 7.076
R7130 vdd3p3.n2115 vdd3p3.n2114 7.076
R7131 vdd3p3.n2114 vdd3p3.n2113 7.076
R7132 vdd3p3.n2113 vdd3p3.n1955 7.076
R7133 vdd3p3.n2107 vdd3p3.n1955 7.076
R7134 vdd3p3.n2107 vdd3p3.n2106 7.076
R7135 vdd3p3.n2106 vdd3p3.n2105 7.076
R7136 vdd3p3.n2105 vdd3p3.n1959 7.076
R7137 vdd3p3.n2099 vdd3p3.n1959 7.076
R7138 vdd3p3.n2099 vdd3p3.n2098 7.076
R7139 vdd3p3.n2098 vdd3p3.n2097 7.076
R7140 vdd3p3.n2097 vdd3p3.n1963 7.076
R7141 vdd3p3.n2091 vdd3p3.n1963 7.076
R7142 vdd3p3.n2091 vdd3p3.n2090 7.076
R7143 vdd3p3.n2090 vdd3p3.n2089 7.076
R7144 vdd3p3.n2089 vdd3p3.n1967 7.076
R7145 vdd3p3.n2083 vdd3p3.n1967 7.076
R7146 vdd3p3.n2083 vdd3p3.n2082 7.076
R7147 vdd3p3.n2082 vdd3p3.n2081 7.076
R7148 vdd3p3.n2081 vdd3p3.n1971 7.076
R7149 vdd3p3.n1284 vdd3p3.n1102 7.076
R7150 vdd3p3.n1278 vdd3p3.n1102 7.076
R7151 vdd3p3.n1278 vdd3p3.n1277 7.076
R7152 vdd3p3.n1277 vdd3p3.n1276 7.076
R7153 vdd3p3.n1276 vdd3p3.n1106 7.076
R7154 vdd3p3.n1270 vdd3p3.n1106 7.076
R7155 vdd3p3.n1270 vdd3p3.n1269 7.076
R7156 vdd3p3.n1269 vdd3p3.n1268 7.076
R7157 vdd3p3.n1268 vdd3p3.n1110 7.076
R7158 vdd3p3.n1262 vdd3p3.n1110 7.076
R7159 vdd3p3.n1262 vdd3p3.n1261 7.076
R7160 vdd3p3.n1261 vdd3p3.n1260 7.076
R7161 vdd3p3.n1260 vdd3p3.n1114 7.076
R7162 vdd3p3.n1254 vdd3p3.n1114 7.076
R7163 vdd3p3.n1254 vdd3p3.n1253 7.076
R7164 vdd3p3.n1253 vdd3p3.n1252 7.076
R7165 vdd3p3.n1252 vdd3p3.n1118 7.076
R7166 vdd3p3.n1246 vdd3p3.n1118 7.076
R7167 vdd3p3.n1246 vdd3p3.n1245 7.076
R7168 vdd3p3.n1245 vdd3p3.n1244 7.076
R7169 vdd3p3.n1244 vdd3p3.n1122 7.076
R7170 vdd3p3.n1238 vdd3p3.n1122 7.076
R7171 vdd3p3.n1238 vdd3p3.n1237 7.076
R7172 vdd3p3.n1237 vdd3p3.n1236 7.076
R7173 vdd3p3.n1236 vdd3p3.n1126 7.076
R7174 vdd3p3.n438 vdd3p3.n256 7.076
R7175 vdd3p3.n432 vdd3p3.n256 7.076
R7176 vdd3p3.n432 vdd3p3.n431 7.076
R7177 vdd3p3.n431 vdd3p3.n430 7.076
R7178 vdd3p3.n430 vdd3p3.n260 7.076
R7179 vdd3p3.n424 vdd3p3.n260 7.076
R7180 vdd3p3.n424 vdd3p3.n423 7.076
R7181 vdd3p3.n423 vdd3p3.n422 7.076
R7182 vdd3p3.n422 vdd3p3.n264 7.076
R7183 vdd3p3.n416 vdd3p3.n264 7.076
R7184 vdd3p3.n416 vdd3p3.n415 7.076
R7185 vdd3p3.n415 vdd3p3.n414 7.076
R7186 vdd3p3.n414 vdd3p3.n268 7.076
R7187 vdd3p3.n408 vdd3p3.n268 7.076
R7188 vdd3p3.n408 vdd3p3.n407 7.076
R7189 vdd3p3.n407 vdd3p3.n406 7.076
R7190 vdd3p3.n406 vdd3p3.n272 7.076
R7191 vdd3p3.n400 vdd3p3.n272 7.076
R7192 vdd3p3.n400 vdd3p3.n399 7.076
R7193 vdd3p3.n399 vdd3p3.n398 7.076
R7194 vdd3p3.n398 vdd3p3.n276 7.076
R7195 vdd3p3.n392 vdd3p3.n276 7.076
R7196 vdd3p3.n392 vdd3p3.n391 7.076
R7197 vdd3p3.n391 vdd3p3.n390 7.076
R7198 vdd3p3.n390 vdd3p3.n280 7.076
R7199 vdd3p3.n3161 vdd3p3.n3023 7.051
R7200 vdd3p3.n3160 vdd3p3.n3035 7.051
R7201 vdd3p3.n3153 vdd3p3.n3041 7.051
R7202 vdd3p3.n3048 vdd3p3.n3042 7.051
R7203 vdd3p3.n2315 vdd3p3.n2177 7.051
R7204 vdd3p3.n2314 vdd3p3.n2189 7.051
R7205 vdd3p3.n2307 vdd3p3.n2195 7.051
R7206 vdd3p3.n2202 vdd3p3.n2196 7.051
R7207 vdd3p3.n1470 vdd3p3.n1332 7.051
R7208 vdd3p3.n1469 vdd3p3.n1344 7.051
R7209 vdd3p3.n1462 vdd3p3.n1350 7.051
R7210 vdd3p3.n1357 vdd3p3.n1351 7.051
R7211 vdd3p3.n624 vdd3p3.n486 7.051
R7212 vdd3p3.n623 vdd3p3.n498 7.051
R7213 vdd3p3.n616 vdd3p3.n504 7.051
R7214 vdd3p3.n511 vdd3p3.n505 7.051
R7215 vdd3p3.n4151 vdd3p3.n4148 6.894
R7216 vdd3p3.n4256 vdd3p3.n4255 6.803
R7217 vdd3p3.n4576 vdd3p3.n4575 6.803
R7218 vdd3p3.n3518 vdd3p3.n3517 6.803
R7219 vdd3p3.n4767 vdd3p3.n4766 6.8
R7220 vdd3p3.n4908 vdd3p3.n4907 6.8
R7221 vdd3p3.n4272 vdd3p3.n4271 6.8
R7222 vdd3p3.n4592 vdd3p3.n4591 6.8
R7223 vdd3p3.n3702 vdd3p3.n3701 6.8
R7224 vdd3p3.n8731 vdd3p3.n8730 6.599
R7225 vdd3p3.n2920 vdd3p3.n2919 6.593
R7226 vdd3p3.n2919 vdd3p3.n2821 6.593
R7227 vdd3p3.n2914 vdd3p3.n2821 6.593
R7228 vdd3p3.n2914 vdd3p3.n2913 6.593
R7229 vdd3p3.n2913 vdd3p3.n2912 6.593
R7230 vdd3p3.n2912 vdd3p3.n2825 6.593
R7231 vdd3p3.n2906 vdd3p3.n2825 6.593
R7232 vdd3p3.n2906 vdd3p3.n2905 6.593
R7233 vdd3p3.n2905 vdd3p3.n2904 6.593
R7234 vdd3p3.n2904 vdd3p3.n2830 6.593
R7235 vdd3p3.n2898 vdd3p3.n2830 6.593
R7236 vdd3p3.n2898 vdd3p3.n2897 6.593
R7237 vdd3p3.n2897 vdd3p3.n2896 6.593
R7238 vdd3p3.n2896 vdd3p3.n2834 6.593
R7239 vdd3p3.n2890 vdd3p3.n2834 6.593
R7240 vdd3p3.n2890 vdd3p3.n2889 6.593
R7241 vdd3p3.n2889 vdd3p3.n2888 6.593
R7242 vdd3p3.n2074 vdd3p3.n2073 6.593
R7243 vdd3p3.n2073 vdd3p3.n1975 6.593
R7244 vdd3p3.n2068 vdd3p3.n1975 6.593
R7245 vdd3p3.n2068 vdd3p3.n2067 6.593
R7246 vdd3p3.n2067 vdd3p3.n2066 6.593
R7247 vdd3p3.n2066 vdd3p3.n1979 6.593
R7248 vdd3p3.n2060 vdd3p3.n1979 6.593
R7249 vdd3p3.n2060 vdd3p3.n2059 6.593
R7250 vdd3p3.n2059 vdd3p3.n2058 6.593
R7251 vdd3p3.n2058 vdd3p3.n1984 6.593
R7252 vdd3p3.n2052 vdd3p3.n1984 6.593
R7253 vdd3p3.n2052 vdd3p3.n2051 6.593
R7254 vdd3p3.n2051 vdd3p3.n2050 6.593
R7255 vdd3p3.n2050 vdd3p3.n1988 6.593
R7256 vdd3p3.n2044 vdd3p3.n1988 6.593
R7257 vdd3p3.n2044 vdd3p3.n2043 6.593
R7258 vdd3p3.n2043 vdd3p3.n2042 6.593
R7259 vdd3p3.n1229 vdd3p3.n1228 6.593
R7260 vdd3p3.n1228 vdd3p3.n1130 6.593
R7261 vdd3p3.n1223 vdd3p3.n1130 6.593
R7262 vdd3p3.n1223 vdd3p3.n1222 6.593
R7263 vdd3p3.n1222 vdd3p3.n1221 6.593
R7264 vdd3p3.n1221 vdd3p3.n1134 6.593
R7265 vdd3p3.n1215 vdd3p3.n1134 6.593
R7266 vdd3p3.n1215 vdd3p3.n1214 6.593
R7267 vdd3p3.n1214 vdd3p3.n1213 6.593
R7268 vdd3p3.n1213 vdd3p3.n1139 6.593
R7269 vdd3p3.n1207 vdd3p3.n1139 6.593
R7270 vdd3p3.n1207 vdd3p3.n1206 6.593
R7271 vdd3p3.n1206 vdd3p3.n1205 6.593
R7272 vdd3p3.n1205 vdd3p3.n1143 6.593
R7273 vdd3p3.n1199 vdd3p3.n1143 6.593
R7274 vdd3p3.n1199 vdd3p3.n1198 6.593
R7275 vdd3p3.n1198 vdd3p3.n1197 6.593
R7276 vdd3p3.n383 vdd3p3.n382 6.593
R7277 vdd3p3.n382 vdd3p3.n284 6.593
R7278 vdd3p3.n377 vdd3p3.n284 6.593
R7279 vdd3p3.n377 vdd3p3.n376 6.593
R7280 vdd3p3.n376 vdd3p3.n375 6.593
R7281 vdd3p3.n375 vdd3p3.n288 6.593
R7282 vdd3p3.n369 vdd3p3.n288 6.593
R7283 vdd3p3.n369 vdd3p3.n368 6.593
R7284 vdd3p3.n368 vdd3p3.n367 6.593
R7285 vdd3p3.n367 vdd3p3.n293 6.593
R7286 vdd3p3.n361 vdd3p3.n293 6.593
R7287 vdd3p3.n361 vdd3p3.n360 6.593
R7288 vdd3p3.n360 vdd3p3.n359 6.593
R7289 vdd3p3.n359 vdd3p3.n297 6.593
R7290 vdd3p3.n353 vdd3p3.n297 6.593
R7291 vdd3p3.n353 vdd3p3.n352 6.593
R7292 vdd3p3.n352 vdd3p3.n351 6.593
R7293 vdd3p3.n4072 vdd3p3.t51 6.348
R7294 vdd3p3.n3826 vdd3p3.n3825 6.313
R7295 vdd3p3.t73 vdd3p3.n8645 6.308
R7296 vdd3p3.n3192 vdd3p3.n3191 6.173
R7297 vdd3p3.n3193 vdd3p3.n3192 6.173
R7298 vdd3p3.n3193 vdd3p3.n2749 6.173
R7299 vdd3p3.n3199 vdd3p3.n2749 6.173
R7300 vdd3p3.n3200 vdd3p3.n3199 6.173
R7301 vdd3p3.n3201 vdd3p3.n3200 6.173
R7302 vdd3p3.n3201 vdd3p3.n2745 6.173
R7303 vdd3p3.n3207 vdd3p3.n2745 6.173
R7304 vdd3p3.n3208 vdd3p3.n3207 6.173
R7305 vdd3p3.n3209 vdd3p3.n3208 6.173
R7306 vdd3p3.n3209 vdd3p3.n2741 6.173
R7307 vdd3p3.n3215 vdd3p3.n2741 6.173
R7308 vdd3p3.n2346 vdd3p3.n2345 6.173
R7309 vdd3p3.n2347 vdd3p3.n2346 6.173
R7310 vdd3p3.n2347 vdd3p3.n1903 6.173
R7311 vdd3p3.n2353 vdd3p3.n1903 6.173
R7312 vdd3p3.n2354 vdd3p3.n2353 6.173
R7313 vdd3p3.n2355 vdd3p3.n2354 6.173
R7314 vdd3p3.n2355 vdd3p3.n1899 6.173
R7315 vdd3p3.n2361 vdd3p3.n1899 6.173
R7316 vdd3p3.n2362 vdd3p3.n2361 6.173
R7317 vdd3p3.n2363 vdd3p3.n2362 6.173
R7318 vdd3p3.n2363 vdd3p3.n1895 6.173
R7319 vdd3p3.n2369 vdd3p3.n1895 6.173
R7320 vdd3p3.n1501 vdd3p3.n1500 6.173
R7321 vdd3p3.n1502 vdd3p3.n1501 6.173
R7322 vdd3p3.n1502 vdd3p3.n1058 6.173
R7323 vdd3p3.n1508 vdd3p3.n1058 6.173
R7324 vdd3p3.n1509 vdd3p3.n1508 6.173
R7325 vdd3p3.n1510 vdd3p3.n1509 6.173
R7326 vdd3p3.n1510 vdd3p3.n1054 6.173
R7327 vdd3p3.n1516 vdd3p3.n1054 6.173
R7328 vdd3p3.n1517 vdd3p3.n1516 6.173
R7329 vdd3p3.n1518 vdd3p3.n1517 6.173
R7330 vdd3p3.n1518 vdd3p3.n1050 6.173
R7331 vdd3p3.n1524 vdd3p3.n1050 6.173
R7332 vdd3p3.n655 vdd3p3.n654 6.173
R7333 vdd3p3.n656 vdd3p3.n655 6.173
R7334 vdd3p3.n656 vdd3p3.n212 6.173
R7335 vdd3p3.n662 vdd3p3.n212 6.173
R7336 vdd3p3.n663 vdd3p3.n662 6.173
R7337 vdd3p3.n664 vdd3p3.n663 6.173
R7338 vdd3p3.n664 vdd3p3.n208 6.173
R7339 vdd3p3.n670 vdd3p3.n208 6.173
R7340 vdd3p3.n671 vdd3p3.n670 6.173
R7341 vdd3p3.n672 vdd3p3.n671 6.173
R7342 vdd3p3.n672 vdd3p3.n204 6.173
R7343 vdd3p3.n678 vdd3p3.n204 6.173
R7344 vdd3p3.n3961 vdd3p3.n3960 6.083
R7345 vdd3p3.n4195 vdd3p3.n4194 6.023
R7346 vdd3p3.n5047 vdd3p3.n5046 6.023
R7347 vdd3p3.n3473 vdd3p3.n3472 6.023
R7348 vdd3p3.n4954 vdd3p3.n4953 6.023
R7349 vdd3p3.n8501 vdd3p3.n8500 6.023
R7350 vdd3p3.n8845 vdd3p3.n8844 6.023
R7351 vdd3p3.n8756 vdd3p3.n8755 6.023
R7352 vdd3p3.n7381 vdd3p3.n7380 5.967
R7353 vdd3p3.n4007 vdd3p3.t153 5.951
R7354 vdd3p3.t39 vdd3p3.n4121 5.951
R7355 vdd3p3.n3045 vdd3p3.n3018 5.802
R7356 vdd3p3.n3151 vdd3p3.n3045 5.802
R7357 vdd3p3.n3151 vdd3p3.n3150 5.802
R7358 vdd3p3.n3150 vdd3p3.n3149 5.802
R7359 vdd3p3.n3149 vdd3p3.n3046 5.802
R7360 vdd3p3.n3054 vdd3p3.n2626 5.802
R7361 vdd3p3.n3361 vdd3p3.n2626 5.802
R7362 vdd3p3.n3361 vdd3p3.n3360 5.802
R7363 vdd3p3.n3360 vdd3p3.n3359 5.802
R7364 vdd3p3.n3359 vdd3p3.n2627 5.802
R7365 vdd3p3.n2199 vdd3p3.n2172 5.802
R7366 vdd3p3.n2305 vdd3p3.n2199 5.802
R7367 vdd3p3.n2305 vdd3p3.n2304 5.802
R7368 vdd3p3.n2304 vdd3p3.n2303 5.802
R7369 vdd3p3.n2303 vdd3p3.n2200 5.802
R7370 vdd3p3.n2208 vdd3p3.n1780 5.802
R7371 vdd3p3.n2515 vdd3p3.n1780 5.802
R7372 vdd3p3.n2515 vdd3p3.n2514 5.802
R7373 vdd3p3.n2514 vdd3p3.n2513 5.802
R7374 vdd3p3.n2513 vdd3p3.n1781 5.802
R7375 vdd3p3.n1354 vdd3p3.n1327 5.802
R7376 vdd3p3.n1460 vdd3p3.n1354 5.802
R7377 vdd3p3.n1460 vdd3p3.n1459 5.802
R7378 vdd3p3.n1459 vdd3p3.n1458 5.802
R7379 vdd3p3.n1458 vdd3p3.n1355 5.802
R7380 vdd3p3.n1363 vdd3p3.n935 5.802
R7381 vdd3p3.n1670 vdd3p3.n935 5.802
R7382 vdd3p3.n1670 vdd3p3.n1669 5.802
R7383 vdd3p3.n1669 vdd3p3.n1668 5.802
R7384 vdd3p3.n1668 vdd3p3.n936 5.802
R7385 vdd3p3.n508 vdd3p3.n481 5.802
R7386 vdd3p3.n614 vdd3p3.n508 5.802
R7387 vdd3p3.n614 vdd3p3.n613 5.802
R7388 vdd3p3.n613 vdd3p3.n612 5.802
R7389 vdd3p3.n612 vdd3p3.n509 5.802
R7390 vdd3p3.n517 vdd3p3.n89 5.802
R7391 vdd3p3.n824 vdd3p3.n89 5.802
R7392 vdd3p3.n824 vdd3p3.n823 5.802
R7393 vdd3p3.n823 vdd3p3.n822 5.802
R7394 vdd3p3.n822 vdd3p3.n90 5.802
R7395 vdd3p3.n4923 vdd3p3.n4922 5.737
R7396 vdd3p3.n4258 vdd3p3.n4257 5.647
R7397 vdd3p3.n4274 vdd3p3.n4273 5.647
R7398 vdd3p3.n4578 vdd3p3.n4577 5.647
R7399 vdd3p3.n4594 vdd3p3.n4593 5.647
R7400 vdd3p3.n3520 vdd3p3.n3519 5.647
R7401 vdd3p3.n3536 vdd3p3.n3535 5.647
R7402 vdd3p3.n3605 vdd3p3.n3604 5.647
R7403 vdd3p3.n3704 vdd3p3.n3703 5.647
R7404 vdd3p3.n3633 vdd3p3.n3632 5.647
R7405 vdd3p3.n3623 vdd3p3.n3622 5.647
R7406 vdd3p3.n4769 vdd3p3.n4768 5.647
R7407 vdd3p3.n4910 vdd3p3.n4909 5.647
R7408 vdd3p3.n4365 vdd3p3.n4364 5.629
R7409 vdd3p3.n4429 vdd3p3.n4428 5.629
R7410 vdd3p3.n4459 vdd3p3.n4458 5.629
R7411 vdd3p3.n4519 vdd3p3.n4518 5.629
R7412 vdd3p3.n4687 vdd3p3.n4686 5.629
R7413 vdd3p3.n4399 vdd3p3.n4398 5.629
R7414 vdd3p3.n4489 vdd3p3.n4488 5.629
R7415 vdd3p3.n3315 vdd3p3.n3313 5.615
R7416 vdd3p3.n3313 vdd3p3.n3312 5.615
R7417 vdd3p3.n3312 vdd3p3.n2687 5.615
R7418 vdd3p3.n3306 vdd3p3.n2687 5.615
R7419 vdd3p3.n3306 vdd3p3.n3305 5.615
R7420 vdd3p3.n3305 vdd3p3.n3304 5.615
R7421 vdd3p3.n3304 vdd3p3.n2692 5.615
R7422 vdd3p3.n3298 vdd3p3.n2692 5.615
R7423 vdd3p3.n3298 vdd3p3.n3297 5.615
R7424 vdd3p3.n3297 vdd3p3.n3296 5.615
R7425 vdd3p3.n3296 vdd3p3.n2696 5.615
R7426 vdd3p3.n3290 vdd3p3.n2696 5.615
R7427 vdd3p3.n2469 vdd3p3.n2467 5.615
R7428 vdd3p3.n2467 vdd3p3.n2466 5.615
R7429 vdd3p3.n2466 vdd3p3.n1841 5.615
R7430 vdd3p3.n2460 vdd3p3.n1841 5.615
R7431 vdd3p3.n2460 vdd3p3.n2459 5.615
R7432 vdd3p3.n2459 vdd3p3.n2458 5.615
R7433 vdd3p3.n2458 vdd3p3.n1846 5.615
R7434 vdd3p3.n2452 vdd3p3.n1846 5.615
R7435 vdd3p3.n2452 vdd3p3.n2451 5.615
R7436 vdd3p3.n2451 vdd3p3.n2450 5.615
R7437 vdd3p3.n2450 vdd3p3.n1850 5.615
R7438 vdd3p3.n2444 vdd3p3.n1850 5.615
R7439 vdd3p3.n1624 vdd3p3.n1622 5.615
R7440 vdd3p3.n1622 vdd3p3.n1621 5.615
R7441 vdd3p3.n1621 vdd3p3.n996 5.615
R7442 vdd3p3.n1615 vdd3p3.n996 5.615
R7443 vdd3p3.n1615 vdd3p3.n1614 5.615
R7444 vdd3p3.n1614 vdd3p3.n1613 5.615
R7445 vdd3p3.n1613 vdd3p3.n1001 5.615
R7446 vdd3p3.n1607 vdd3p3.n1001 5.615
R7447 vdd3p3.n1607 vdd3p3.n1606 5.615
R7448 vdd3p3.n1606 vdd3p3.n1605 5.615
R7449 vdd3p3.n1605 vdd3p3.n1005 5.615
R7450 vdd3p3.n1599 vdd3p3.n1005 5.615
R7451 vdd3p3.n778 vdd3p3.n776 5.615
R7452 vdd3p3.n776 vdd3p3.n775 5.615
R7453 vdd3p3.n775 vdd3p3.n150 5.615
R7454 vdd3p3.n769 vdd3p3.n150 5.615
R7455 vdd3p3.n769 vdd3p3.n768 5.615
R7456 vdd3p3.n768 vdd3p3.n767 5.615
R7457 vdd3p3.n767 vdd3p3.n155 5.615
R7458 vdd3p3.n761 vdd3p3.n155 5.615
R7459 vdd3p3.n761 vdd3p3.n760 5.615
R7460 vdd3p3.n760 vdd3p3.n759 5.615
R7461 vdd3p3.n759 vdd3p3.n159 5.615
R7462 vdd3p3.n753 vdd3p3.n159 5.615
R7463 vdd3p3.n5103 vdd3p3.n5102 5.572
R7464 vdd3p3.n4243 vdd3p3.n4242 5.572
R7465 vdd3p3.n4380 vdd3p3.n4378 5.539
R7466 vdd3p3.n4381 vdd3p3.n4380 5.539
R7467 vdd3p3.n4382 vdd3p3.n4381 5.539
R7468 vdd3p3.n4382 vdd3p3.t89 5.539
R7469 vdd3p3.n4415 vdd3p3.t113 5.539
R7470 vdd3p3.n4415 vdd3p3.t148 5.539
R7471 vdd3p3.n4445 vdd3p3.t149 5.539
R7472 vdd3p3.n4445 vdd3p3.t160 5.539
R7473 vdd3p3.n4475 vdd3p3.t161 5.539
R7474 vdd3p3.n4475 vdd3p3.t168 5.539
R7475 vdd3p3.n4505 vdd3p3.t10 5.539
R7476 vdd3p3.n4505 vdd3p3.t90 5.539
R7477 vdd3p3.n3444 vdd3p3.t91 5.539
R7478 vdd3p3.n3444 vdd3p3.t7 5.539
R7479 vdd3p3.n4563 vdd3p3.t5 5.539
R7480 vdd3p3.n4563 vdd3p3.n4562 5.539
R7481 vdd3p3.n4684 vdd3p3.t57 5.539
R7482 vdd3p3.n3574 vdd3p3.n3572 5.539
R7483 vdd3p3.n3574 vdd3p3.n3573 5.539
R7484 vdd3p3.n3668 vdd3p3.n3667 5.539
R7485 vdd3p3.n3738 vdd3p3.t49 5.539
R7486 vdd3p3.n4803 vdd3p3.t72 5.539
R7487 vdd3p3.n4803 vdd3p3.t151 5.539
R7488 vdd3p3.n4734 vdd3p3.t150 5.539
R7489 vdd3p3.n4734 vdd3p3.t60 5.539
R7490 vdd3p3.n8570 vdd3p3.t101 5.539
R7491 vdd3p3.n8570 vdd3p3.t105 5.539
R7492 vdd3p3.n4057 vdd3p3.n4056 5.422
R7493 vdd3p3.n8734 vdd3p3.n8714 5.377
R7494 vdd3p3.n903 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 5.28
R7495 vdd3p3.n2594 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 5.28
R7496 vdd3p3.n8466 vdd3p3.t132 5.273
R7497 vdd3p3.n4206 vdd3p3.n4205 5.27
R7498 vdd3p3.n5058 vdd3p3.n5057 5.27
R7499 vdd3p3.n8512 vdd3p3.n8511 5.27
R7500 vdd3p3.n8856 vdd3p3.n8855 5.27
R7501 vdd3p3.n8767 vdd3p3.n8766 5.27
R7502 vdd3p3.n8541 vdd3p3.n8540 5.251
R7503 vdd3p3.n8620 vdd3p3.n8619 5.251
R7504 vdd3p3.n8803 vdd3p3.n8802 5.251
R7505 vdd3p3.n3088 vdd3p3.n3087 5.231
R7506 vdd3p3.n2242 vdd3p3.n2241 5.231
R7507 vdd3p3.n1397 vdd3p3.n1396 5.231
R7508 vdd3p3.n551 vdd3p3.n550 5.231
R7509 vdd3p3.n4035 vdd3p3.n4018 5.158
R7510 vdd3p3.n4782 vdd3p3.n4781 4.967
R7511 vdd3p3.n4287 vdd3p3.n4286 4.955
R7512 vdd3p3.n4607 vdd3p3.n4606 4.955
R7513 vdd3p3.n3550 vdd3p3.n3549 4.955
R7514 vdd3p3.n3646 vdd3p3.n3645 4.955
R7515 vdd3p3.n3717 vdd3p3.n3716 4.955
R7516 vdd3p3.n3489 vdd3p3.n3483 4.894
R7517 vdd3p3.n4971 vdd3p3.n4965 4.894
R7518 vdd3p3.n3973 vdd3p3.n3972 4.893
R7519 vdd3p3.n8704 vdd3p3.n8702 4.889
R7520 vdd3p3.n3143 vdd3p3.n3142 4.786
R7521 vdd3p3.n2297 vdd3p3.n2296 4.786
R7522 vdd3p3.n1452 vdd3p3.n1451 4.786
R7523 vdd3p3.n606 vdd3p3.n605 4.786
R7524 vdd3p3.n3900 vdd3p3.n3899 4.75
R7525 vdd3p3.n3902 vdd3p3.n3901 4.75
R7526 vdd3p3.n3907 vdd3p3.n3906 4.75
R7527 vdd3p3.n3905 vdd3p3.n3904 4.75
R7528 vdd3p3.n4284 vdd3p3.n4270 4.735
R7529 vdd3p3.n4604 vdd3p3.n4590 4.735
R7530 vdd3p3.n3714 vdd3p3.n3700 4.735
R7531 vdd3p3.n3643 vdd3p3.n3617 4.735
R7532 vdd3p3.n4269 vdd3p3.n4268 4.735
R7533 vdd3p3.n4589 vdd3p3.n4588 4.735
R7534 vdd3p3.n3531 vdd3p3.n3530 4.735
R7535 vdd3p3.n3547 vdd3p3.n3546 4.735
R7536 vdd3p3.n3616 vdd3p3.n3615 4.735
R7537 vdd3p3.n3699 vdd3p3.n3698 4.735
R7538 vdd3p3.n4780 vdd3p3.n4779 4.735
R7539 vdd3p3.n4921 vdd3p3.n4920 4.735
R7540 vdd3p3.n2983 vdd3p3.n2982 4.73
R7541 vdd3p3.n2982 vdd3p3.n2976 4.73
R7542 vdd3p3.n2976 vdd3p3.n2787 4.73
R7543 vdd3p3.n2991 vdd3p3.n2787 4.73
R7544 vdd3p3.n2992 vdd3p3.n2991 4.73
R7545 vdd3p3.n2993 vdd3p3.n2992 4.73
R7546 vdd3p3.n2993 vdd3p3.n2783 4.73
R7547 vdd3p3.n2999 vdd3p3.n2783 4.73
R7548 vdd3p3.n3000 vdd3p3.n2999 4.73
R7549 vdd3p3.n3001 vdd3p3.n3000 4.73
R7550 vdd3p3.n3001 vdd3p3.n2779 4.73
R7551 vdd3p3.n3007 vdd3p3.n2779 4.73
R7552 vdd3p3.n3008 vdd3p3.n3007 4.73
R7553 vdd3p3.n3009 vdd3p3.n3008 4.73
R7554 vdd3p3.n3009 vdd3p3.n2775 4.73
R7555 vdd3p3.n3016 vdd3p3.n2775 4.73
R7556 vdd3p3.n3017 vdd3p3.n3016 4.73
R7557 vdd3p3.n2137 vdd3p3.n2136 4.73
R7558 vdd3p3.n2136 vdd3p3.n2130 4.73
R7559 vdd3p3.n2130 vdd3p3.n1941 4.73
R7560 vdd3p3.n2145 vdd3p3.n1941 4.73
R7561 vdd3p3.n2146 vdd3p3.n2145 4.73
R7562 vdd3p3.n2147 vdd3p3.n2146 4.73
R7563 vdd3p3.n2147 vdd3p3.n1937 4.73
R7564 vdd3p3.n2153 vdd3p3.n1937 4.73
R7565 vdd3p3.n2154 vdd3p3.n2153 4.73
R7566 vdd3p3.n2155 vdd3p3.n2154 4.73
R7567 vdd3p3.n2155 vdd3p3.n1933 4.73
R7568 vdd3p3.n2161 vdd3p3.n1933 4.73
R7569 vdd3p3.n2162 vdd3p3.n2161 4.73
R7570 vdd3p3.n2163 vdd3p3.n2162 4.73
R7571 vdd3p3.n2163 vdd3p3.n1929 4.73
R7572 vdd3p3.n2170 vdd3p3.n1929 4.73
R7573 vdd3p3.n2171 vdd3p3.n2170 4.73
R7574 vdd3p3.n1292 vdd3p3.n1291 4.73
R7575 vdd3p3.n1291 vdd3p3.n1285 4.73
R7576 vdd3p3.n1285 vdd3p3.n1096 4.73
R7577 vdd3p3.n1300 vdd3p3.n1096 4.73
R7578 vdd3p3.n1301 vdd3p3.n1300 4.73
R7579 vdd3p3.n1302 vdd3p3.n1301 4.73
R7580 vdd3p3.n1302 vdd3p3.n1092 4.73
R7581 vdd3p3.n1308 vdd3p3.n1092 4.73
R7582 vdd3p3.n1309 vdd3p3.n1308 4.73
R7583 vdd3p3.n1310 vdd3p3.n1309 4.73
R7584 vdd3p3.n1310 vdd3p3.n1088 4.73
R7585 vdd3p3.n1316 vdd3p3.n1088 4.73
R7586 vdd3p3.n1317 vdd3p3.n1316 4.73
R7587 vdd3p3.n1318 vdd3p3.n1317 4.73
R7588 vdd3p3.n1318 vdd3p3.n1084 4.73
R7589 vdd3p3.n1325 vdd3p3.n1084 4.73
R7590 vdd3p3.n1326 vdd3p3.n1325 4.73
R7591 vdd3p3.n446 vdd3p3.n445 4.73
R7592 vdd3p3.n445 vdd3p3.n439 4.73
R7593 vdd3p3.n439 vdd3p3.n250 4.73
R7594 vdd3p3.n454 vdd3p3.n250 4.73
R7595 vdd3p3.n455 vdd3p3.n454 4.73
R7596 vdd3p3.n456 vdd3p3.n455 4.73
R7597 vdd3p3.n456 vdd3p3.n246 4.73
R7598 vdd3p3.n462 vdd3p3.n246 4.73
R7599 vdd3p3.n463 vdd3p3.n462 4.73
R7600 vdd3p3.n464 vdd3p3.n463 4.73
R7601 vdd3p3.n464 vdd3p3.n242 4.73
R7602 vdd3p3.n470 vdd3p3.n242 4.73
R7603 vdd3p3.n471 vdd3p3.n470 4.73
R7604 vdd3p3.n472 vdd3p3.n471 4.73
R7605 vdd3p3.n472 vdd3p3.n238 4.73
R7606 vdd3p3.n479 vdd3p3.n238 4.73
R7607 vdd3p3.n480 vdd3p3.n479 4.73
R7608 vdd3p3.n17 vdd3p3.n16 4.652
R7609 vdd3p3.n865 vdd3p3.n864 4.652
R7610 vdd3p3.n1708 vdd3p3.n1707 4.652
R7611 vdd3p3.n2556 vdd3p3.n2555 4.652
R7612 vdd3p3.n51 vdd3p3.n37 4.65
R7613 vdd3p3.n50 vdd3p3.n49 4.65
R7614 vdd3p3.n48 vdd3p3.n39 4.65
R7615 vdd3p3.n47 vdd3p3.n46 4.65
R7616 vdd3p3.n20 vdd3p3.n8 4.65
R7617 vdd3p3.n27 vdd3p3.n26 4.65
R7618 vdd3p3.n11 vdd3p3.n4 4.65
R7619 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n58 4.65
R7620 vdd3p3.n10 vdd3p3.n3 4.65
R7621 vdd3p3.n13 vdd3p3.n10 4.65
R7622 vdd3p3.n19 vdd3p3.n18 4.65
R7623 vdd3p3.n893 vdd3p3.n890 4.65
R7624 vdd3p3.n892 vdd3p3.n891 4.65
R7625 vdd3p3.n847 vdd3p3.n846 4.65
R7626 vdd3p3.n899 vdd3p3.n898 4.65
R7627 vdd3p3.n860 vdd3p3.n856 4.65
R7628 vdd3p3.n871 vdd3p3.n870 4.65
R7629 vdd3p3.n877 vdd3p3.n851 4.65
R7630 vdd3p3.n881 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.vdd3p3 4.65
R7631 vdd3p3.n880 vdd3p3.n879 4.65
R7632 vdd3p3.n879 vdd3p3.n853 4.65
R7633 vdd3p3.n859 vdd3p3.n858 4.65
R7634 vdd3p3.n1742 vdd3p3.n1728 4.65
R7635 vdd3p3.n1741 vdd3p3.n1740 4.65
R7636 vdd3p3.n1739 vdd3p3.n1730 4.65
R7637 vdd3p3.n1738 vdd3p3.n1737 4.65
R7638 vdd3p3.n1711 vdd3p3.n1699 4.65
R7639 vdd3p3.n1718 vdd3p3.n1717 4.65
R7640 vdd3p3.n1702 vdd3p3.n1695 4.65
R7641 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n1749 4.65
R7642 vdd3p3.n1701 vdd3p3.n1694 4.65
R7643 vdd3p3.n1704 vdd3p3.n1701 4.65
R7644 vdd3p3.n1710 vdd3p3.n1709 4.65
R7645 vdd3p3.n2584 vdd3p3.n2581 4.65
R7646 vdd3p3.n2583 vdd3p3.n2582 4.65
R7647 vdd3p3.n2538 vdd3p3.n2537 4.65
R7648 vdd3p3.n2590 vdd3p3.n2589 4.65
R7649 vdd3p3.n2551 vdd3p3.n2547 4.65
R7650 vdd3p3.n2562 vdd3p3.n2561 4.65
R7651 vdd3p3.n2568 vdd3p3.n2542 4.65
R7652 vdd3p3.n2572 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.vdd3p3 4.65
R7653 vdd3p3.n2571 vdd3p3.n2570 4.65
R7654 vdd3p3.n2570 vdd3p3.n2544 4.65
R7655 vdd3p3.n2550 vdd3p3.n2549 4.65
R7656 vdd3p3.n3631 vdd3p3.n3630 4.65
R7657 vdd3p3.n3534 vdd3p3.n3533 4.65
R7658 vdd3p3.n3395 vdd3p3.n3385 4.65
R7659 vdd3p3.n6715 vdd3p3.n6714 4.65
R7660 vdd3p3.n6711 vdd3p3.n6710 4.65
R7661 vdd3p3.n6707 vdd3p3.n6706 4.65
R7662 vdd3p3.n6703 vdd3p3.n6702 4.65
R7663 vdd3p3.n6699 vdd3p3.n6698 4.65
R7664 vdd3p3.n6695 vdd3p3.n6694 4.65
R7665 vdd3p3.n6690 vdd3p3.n6689 4.65
R7666 vdd3p3.n6685 vdd3p3.n6684 4.65
R7667 vdd3p3.n6677 vdd3p3.n6676 4.65
R7668 vdd3p3.n6672 vdd3p3.n6671 4.65
R7669 vdd3p3.n6667 vdd3p3.n6666 4.65
R7670 vdd3p3.n6662 vdd3p3.n6661 4.65
R7671 vdd3p3.n6657 vdd3p3.n6656 4.65
R7672 vdd3p3.n6652 vdd3p3.n6651 4.65
R7673 vdd3p3.n6647 vdd3p3.n6646 4.65
R7674 vdd3p3.n6642 vdd3p3.n6641 4.65
R7675 vdd3p3.n6637 vdd3p3.n6636 4.65
R7676 vdd3p3.n6632 vdd3p3.n6631 4.65
R7677 vdd3p3.n6627 vdd3p3.n6626 4.65
R7678 vdd3p3.n6622 vdd3p3.n6621 4.65
R7679 vdd3p3.n6617 vdd3p3.n6616 4.65
R7680 vdd3p3.n6612 vdd3p3.n6611 4.65
R7681 vdd3p3.n6607 vdd3p3.n6606 4.65
R7682 vdd3p3.n6602 vdd3p3.n6601 4.65
R7683 vdd3p3.n6597 vdd3p3.n6596 4.65
R7684 vdd3p3.n6589 vdd3p3.n6588 4.65
R7685 vdd3p3.n6585 vdd3p3.n6584 4.65
R7686 vdd3p3.n6581 vdd3p3.n6580 4.65
R7687 vdd3p3.n6577 vdd3p3.n6576 4.65
R7688 vdd3p3.n6573 vdd3p3.n6572 4.65
R7689 vdd3p3.n6569 vdd3p3.n6568 4.65
R7690 vdd3p3.n6565 vdd3p3.n6564 4.65
R7691 vdd3p3.n6548 vdd3p3.n6547 4.65
R7692 vdd3p3.n6544 vdd3p3.n6543 4.65
R7693 vdd3p3.n6540 vdd3p3.n6539 4.65
R7694 vdd3p3.n6536 vdd3p3.n6535 4.65
R7695 vdd3p3.n6532 vdd3p3.n6531 4.65
R7696 vdd3p3.n6528 vdd3p3.n6527 4.65
R7697 vdd3p3.n6524 vdd3p3.n6523 4.65
R7698 vdd3p3.n6519 vdd3p3.n6518 4.65
R7699 vdd3p3.n6514 vdd3p3.n6513 4.65
R7700 vdd3p3.n6509 vdd3p3.n6508 4.65
R7701 vdd3p3.n6501 vdd3p3.n6500 4.65
R7702 vdd3p3.n6496 vdd3p3.n6495 4.65
R7703 vdd3p3.n6491 vdd3p3.n6490 4.65
R7704 vdd3p3.n6486 vdd3p3.n6485 4.65
R7705 vdd3p3.n6481 vdd3p3.n6480 4.65
R7706 vdd3p3.n6476 vdd3p3.n6475 4.65
R7707 vdd3p3.n6471 vdd3p3.n6470 4.65
R7708 vdd3p3.n6466 vdd3p3.n6465 4.65
R7709 vdd3p3.n6461 vdd3p3.n6460 4.65
R7710 vdd3p3.n6456 vdd3p3.n6455 4.65
R7711 vdd3p3.n6451 vdd3p3.n6450 4.65
R7712 vdd3p3.n6446 vdd3p3.n6445 4.65
R7713 vdd3p3.n6441 vdd3p3.n6440 4.65
R7714 vdd3p3.n6436 vdd3p3.n6435 4.65
R7715 vdd3p3.n6431 vdd3p3.n6430 4.65
R7716 vdd3p3.n6426 vdd3p3.n6425 4.65
R7717 vdd3p3.n6421 vdd3p3.n6420 4.65
R7718 vdd3p3.n6415 vdd3p3.n6414 4.65
R7719 vdd3p3.n6411 vdd3p3.n6410 4.65
R7720 vdd3p3.n6407 vdd3p3.n6406 4.65
R7721 vdd3p3.n6403 vdd3p3.n6402 4.65
R7722 vdd3p3.n7949 vdd3p3.n7948 4.65
R7723 vdd3p3.n7957 vdd3p3.n7956 4.65
R7724 vdd3p3.n7965 vdd3p3.n7964 4.65
R7725 vdd3p3.n7973 vdd3p3.n7972 4.65
R7726 vdd3p3.n7981 vdd3p3.n7980 4.65
R7727 vdd3p3.n7989 vdd3p3.n7988 4.65
R7728 vdd3p3.n7995 vdd3p3.n7994 4.65
R7729 vdd3p3.n8003 vdd3p3.n8002 4.65
R7730 vdd3p3.n8009 vdd3p3.n8008 4.65
R7731 vdd3p3.n8017 vdd3p3.n8016 4.65
R7732 vdd3p3.n8024 vdd3p3.n8023 4.65
R7733 vdd3p3.n8033 vdd3p3.n8032 4.65
R7734 vdd3p3.n8038 vdd3p3.n8037 4.65
R7735 vdd3p3.n8044 vdd3p3.n8043 4.65
R7736 vdd3p3.n8050 vdd3p3.n8049 4.65
R7737 vdd3p3.n8056 vdd3p3.n8055 4.65
R7738 vdd3p3.n8062 vdd3p3.n8061 4.65
R7739 vdd3p3.n8068 vdd3p3.n8067 4.65
R7740 vdd3p3.n8074 vdd3p3.n8073 4.65
R7741 vdd3p3.n8082 vdd3p3.n8081 4.65
R7742 vdd3p3.n8088 vdd3p3.n8087 4.65
R7743 vdd3p3.n8096 vdd3p3.n8095 4.65
R7744 vdd3p3.n8102 vdd3p3.n8101 4.65
R7745 vdd3p3.n8108 vdd3p3.n8107 4.65
R7746 vdd3p3.n8114 vdd3p3.n8113 4.65
R7747 vdd3p3.n8120 vdd3p3.n8119 4.65
R7748 vdd3p3.n8126 vdd3p3.n8125 4.65
R7749 vdd3p3.n8132 vdd3p3.n8131 4.65
R7750 vdd3p3.n8138 vdd3p3.n8137 4.65
R7751 vdd3p3.n8143 vdd3p3.n8142 4.65
R7752 vdd3p3.n8149 vdd3p3.n8148 4.65
R7753 vdd3p3.n8155 vdd3p3.n8154 4.65
R7754 vdd3p3.n8161 vdd3p3.n8160 4.65
R7755 vdd3p3.n8167 vdd3p3.n8166 4.65
R7756 vdd3p3.n8173 vdd3p3.n8172 4.65
R7757 vdd3p3.n8179 vdd3p3.n8178 4.65
R7758 vdd3p3.n8187 vdd3p3.n8186 4.65
R7759 vdd3p3.n8193 vdd3p3.n8192 4.65
R7760 vdd3p3.n8201 vdd3p3.n8200 4.65
R7761 vdd3p3.n8207 vdd3p3.n8206 4.65
R7762 vdd3p3.n8213 vdd3p3.n8212 4.65
R7763 vdd3p3.n8219 vdd3p3.n8218 4.65
R7764 vdd3p3.n8225 vdd3p3.n8224 4.65
R7765 vdd3p3.n8231 vdd3p3.n8230 4.65
R7766 vdd3p3.n8237 vdd3p3.n8236 4.65
R7767 vdd3p3.n8243 vdd3p3.n8242 4.65
R7768 vdd3p3.n8248 vdd3p3.n8247 4.65
R7769 vdd3p3.n8254 vdd3p3.n8253 4.65
R7770 vdd3p3.n8260 vdd3p3.n8259 4.65
R7771 vdd3p3.n8266 vdd3p3.n8265 4.65
R7772 vdd3p3.n8272 vdd3p3.n8271 4.65
R7773 vdd3p3.n8278 vdd3p3.n8277 4.65
R7774 vdd3p3.n8284 vdd3p3.n8283 4.65
R7775 vdd3p3.n8292 vdd3p3.n8291 4.65
R7776 vdd3p3.n8298 vdd3p3.n8297 4.65
R7777 vdd3p3.n8310 vdd3p3.n8309 4.65
R7778 vdd3p3.n8320 vdd3p3.n8319 4.65
R7779 vdd3p3.n8330 vdd3p3.n8329 4.65
R7780 vdd3p3.n8340 vdd3p3.n8339 4.65
R7781 vdd3p3.n8350 vdd3p3.n8349 4.65
R7782 vdd3p3.n8359 vdd3p3.n8358 4.65
R7783 vdd3p3.n8368 vdd3p3.n8367 4.65
R7784 vdd3p3.n8377 vdd3p3.n8376 4.65
R7785 vdd3p3.n8385 vdd3p3.n8384 4.65
R7786 vdd3p3.n8394 vdd3p3.n8393 4.65
R7787 vdd3p3.n8403 vdd3p3.n8402 4.65
R7788 vdd3p3.n8412 vdd3p3.n8411 4.65
R7789 vdd3p3.n8420 vdd3p3.n8419 4.65
R7790 vdd3p3.n8428 vdd3p3.n8427 4.65
R7791 vdd3p3.n8434 vdd3p3.n8433 4.65
R7792 vdd3p3.n7924 vdd3p3.n7923 4.65
R7793 vdd3p3.n7916 vdd3p3.n7915 4.65
R7794 vdd3p3.n7908 vdd3p3.n7907 4.65
R7795 vdd3p3.n7900 vdd3p3.n7899 4.65
R7796 vdd3p3.n7892 vdd3p3.n7891 4.65
R7797 vdd3p3.n7884 vdd3p3.n7883 4.65
R7798 vdd3p3.n7876 vdd3p3.n7875 4.65
R7799 vdd3p3.n7868 vdd3p3.n7867 4.65
R7800 vdd3p3.n7857 vdd3p3.n7856 4.65
R7801 vdd3p3.n7849 vdd3p3.n7848 4.65
R7802 vdd3p3.n7838 vdd3p3.n7837 4.65
R7803 vdd3p3.n7830 vdd3p3.n7829 4.65
R7804 vdd3p3.n7822 vdd3p3.n7821 4.65
R7805 vdd3p3.n7814 vdd3p3.n7813 4.65
R7806 vdd3p3.n7806 vdd3p3.n7805 4.65
R7807 vdd3p3.n7798 vdd3p3.n7797 4.65
R7808 vdd3p3.n7790 vdd3p3.n7789 4.65
R7809 vdd3p3.n7782 vdd3p3.n7781 4.65
R7810 vdd3p3.n7774 vdd3p3.n7773 4.65
R7811 vdd3p3.n7766 vdd3p3.n7765 4.65
R7812 vdd3p3.n7758 vdd3p3.n7757 4.65
R7813 vdd3p3.n7750 vdd3p3.n7749 4.65
R7814 vdd3p3.n7742 vdd3p3.n7741 4.65
R7815 vdd3p3.n7734 vdd3p3.n7733 4.65
R7816 vdd3p3.n7726 vdd3p3.n7725 4.65
R7817 vdd3p3.n7716 vdd3p3.n7715 4.65
R7818 vdd3p3.n7710 vdd3p3.n7709 4.65
R7819 vdd3p3.n7702 vdd3p3.n7701 4.65
R7820 vdd3p3.n7696 vdd3p3.n7695 4.65
R7821 vdd3p3.n7690 vdd3p3.n7689 4.65
R7822 vdd3p3.n7682 vdd3p3.n7681 4.65
R7823 vdd3p3.n7674 vdd3p3.n7673 4.65
R7824 vdd3p3.n7666 vdd3p3.n7665 4.65
R7825 vdd3p3.n7658 vdd3p3.n7657 4.65
R7826 vdd3p3.n7650 vdd3p3.n7649 4.65
R7827 vdd3p3.n7642 vdd3p3.n7641 4.65
R7828 vdd3p3.n7634 vdd3p3.n7633 4.65
R7829 vdd3p3.n7626 vdd3p3.n7625 4.65
R7830 vdd3p3.n7618 vdd3p3.n7617 4.65
R7831 vdd3p3.n7610 vdd3p3.n7609 4.65
R7832 vdd3p3.n7602 vdd3p3.n7601 4.65
R7833 vdd3p3.n7594 vdd3p3.n7593 4.65
R7834 vdd3p3.n7583 vdd3p3.n7582 4.65
R7835 vdd3p3.n7575 vdd3p3.n7574 4.65
R7836 vdd3p3.n7564 vdd3p3.n7563 4.65
R7837 vdd3p3.n7556 vdd3p3.n7555 4.65
R7838 vdd3p3.n7548 vdd3p3.n7547 4.65
R7839 vdd3p3.n7540 vdd3p3.n7539 4.65
R7840 vdd3p3.n7532 vdd3p3.n7531 4.65
R7841 vdd3p3.n7527 vdd3p3.n7526 4.65
R7842 vdd3p3.n7935 vdd3p3.n7934 4.65
R7843 vdd3p3.n7492 vdd3p3.n7491 4.65
R7844 vdd3p3.n7487 vdd3p3.n7486 4.65
R7845 vdd3p3.n7482 vdd3p3.n7481 4.65
R7846 vdd3p3.n7477 vdd3p3.n7476 4.65
R7847 vdd3p3.n7472 vdd3p3.n7471 4.65
R7848 vdd3p3.n7455 vdd3p3.n7454 4.65
R7849 vdd3p3.n7448 vdd3p3.n7447 4.65
R7850 vdd3p3.n7443 vdd3p3.n7442 4.65
R7851 vdd3p3.n7438 vdd3p3.n7437 4.65
R7852 vdd3p3.n7433 vdd3p3.n7432 4.65
R7853 vdd3p3.n7428 vdd3p3.n7427 4.65
R7854 vdd3p3.n7422 vdd3p3.n7421 4.65
R7855 vdd3p3.n7417 vdd3p3.n7416 4.65
R7856 vdd3p3.n7412 vdd3p3.n7411 4.65
R7857 vdd3p3.n7407 vdd3p3.n7406 4.65
R7858 vdd3p3.n7402 vdd3p3.n7401 4.65
R7859 vdd3p3.n7397 vdd3p3.n7396 4.65
R7860 vdd3p3.n7393 vdd3p3.n7392 4.65
R7861 vdd3p3.n7387 vdd3p3.n7386 4.65
R7862 vdd3p3.n7383 vdd3p3.n7382 4.65
R7863 vdd3p3.n7379 vdd3p3.n7378 4.65
R7864 vdd3p3.n7377 vdd3p3.n7376 4.65
R7865 vdd3p3.n7371 vdd3p3.n7370 4.65
R7866 vdd3p3.n7367 vdd3p3.n7366 4.65
R7867 vdd3p3.n7363 vdd3p3.n7362 4.65
R7868 vdd3p3.n7359 vdd3p3.n7358 4.65
R7869 vdd3p3.n7355 vdd3p3.n7354 4.65
R7870 vdd3p3.n7351 vdd3p3.n7350 4.65
R7871 vdd3p3.n7347 vdd3p3.n7346 4.65
R7872 vdd3p3.n7343 vdd3p3.n7342 4.65
R7873 vdd3p3.n7339 vdd3p3.n7338 4.65
R7874 vdd3p3.n7336 vdd3p3.n7335 4.65
R7875 vdd3p3.n7332 vdd3p3.n7331 4.65
R7876 vdd3p3.n7328 vdd3p3.n7327 4.65
R7877 vdd3p3.n7324 vdd3p3.n7323 4.65
R7878 vdd3p3.n7320 vdd3p3.n7319 4.65
R7879 vdd3p3.n7316 vdd3p3.n7315 4.65
R7880 vdd3p3.n7312 vdd3p3.n7311 4.65
R7881 vdd3p3.n7308 vdd3p3.n7307 4.65
R7882 vdd3p3.n7302 vdd3p3.n7301 4.65
R7883 vdd3p3.n7298 vdd3p3.n7297 4.65
R7884 vdd3p3.n7294 vdd3p3.n7293 4.65
R7885 vdd3p3.n7290 vdd3p3.n7289 4.65
R7886 vdd3p3.n7286 vdd3p3.n7285 4.65
R7887 vdd3p3.n7282 vdd3p3.n7281 4.65
R7888 vdd3p3.n7278 vdd3p3.n7277 4.65
R7889 vdd3p3.n7274 vdd3p3.n7273 4.65
R7890 vdd3p3.n7270 vdd3p3.n7269 4.65
R7891 vdd3p3.n7267 vdd3p3.n7266 4.65
R7892 vdd3p3.n7263 vdd3p3.n7262 4.65
R7893 vdd3p3.n7259 vdd3p3.n7258 4.65
R7894 vdd3p3.n7255 vdd3p3.n7254 4.65
R7895 vdd3p3.n7251 vdd3p3.n7250 4.65
R7896 vdd3p3.n7247 vdd3p3.n7246 4.65
R7897 vdd3p3.n7243 vdd3p3.n7242 4.65
R7898 vdd3p3.n7239 vdd3p3.n7238 4.65
R7899 vdd3p3.n7233 vdd3p3.n7232 4.65
R7900 vdd3p3.n7228 vdd3p3.n7227 4.65
R7901 vdd3p3.n7223 vdd3p3.n7222 4.65
R7902 vdd3p3.n7218 vdd3p3.n7217 4.65
R7903 vdd3p3.n7213 vdd3p3.n7212 4.65
R7904 vdd3p3.n7208 vdd3p3.n7207 4.65
R7905 vdd3p3.n7203 vdd3p3.n7202 4.65
R7906 vdd3p3.n7198 vdd3p3.n7197 4.65
R7907 vdd3p3.n7193 vdd3p3.n7192 4.65
R7908 vdd3p3.n7189 vdd3p3.n7188 4.65
R7909 vdd3p3.n7184 vdd3p3.n7183 4.65
R7910 vdd3p3.n7179 vdd3p3.n7178 4.65
R7911 vdd3p3.n7174 vdd3p3.n7173 4.65
R7912 vdd3p3.n7169 vdd3p3.n7168 4.65
R7913 vdd3p3.n7164 vdd3p3.n7163 4.65
R7914 vdd3p3.n7159 vdd3p3.n7158 4.65
R7915 vdd3p3.n7154 vdd3p3.n7153 4.65
R7916 vdd3p3.n7146 vdd3p3.n7145 4.65
R7917 vdd3p3.n7141 vdd3p3.n7140 4.65
R7918 vdd3p3.n7136 vdd3p3.n7135 4.65
R7919 vdd3p3.n7131 vdd3p3.n7130 4.65
R7920 vdd3p3.n7126 vdd3p3.n7125 4.65
R7921 vdd3p3.n7121 vdd3p3.n7120 4.65
R7922 vdd3p3.n7116 vdd3p3.n7115 4.65
R7923 vdd3p3.n7111 vdd3p3.n7110 4.65
R7924 vdd3p3.n7106 vdd3p3.n7105 4.65
R7925 vdd3p3.n7102 vdd3p3.n7101 4.65
R7926 vdd3p3.n7097 vdd3p3.n7096 4.65
R7927 vdd3p3.n7092 vdd3p3.n7091 4.65
R7928 vdd3p3.n7087 vdd3p3.n7086 4.65
R7929 vdd3p3.n7082 vdd3p3.n7081 4.65
R7930 vdd3p3.n7077 vdd3p3.n7076 4.65
R7931 vdd3p3.n7072 vdd3p3.n7071 4.65
R7932 vdd3p3.n7067 vdd3p3.n7066 4.65
R7933 vdd3p3.n7059 vdd3p3.n7058 4.65
R7934 vdd3p3.n7054 vdd3p3.n7053 4.65
R7935 vdd3p3.n7049 vdd3p3.n7048 4.65
R7936 vdd3p3.n7044 vdd3p3.n7043 4.65
R7937 vdd3p3.n7039 vdd3p3.n7038 4.65
R7938 vdd3p3.n7034 vdd3p3.n7033 4.65
R7939 vdd3p3.n7029 vdd3p3.n7028 4.65
R7940 vdd3p3.n7024 vdd3p3.n7023 4.65
R7941 vdd3p3.n5727 vdd3p3.n5726 4.65
R7942 vdd3p3.n5722 vdd3p3.n5721 4.65
R7943 vdd3p3.n5717 vdd3p3.n5716 4.65
R7944 vdd3p3.n5712 vdd3p3.n5711 4.65
R7945 vdd3p3.n5707 vdd3p3.n5706 4.65
R7946 vdd3p3.n5702 vdd3p3.n5701 4.65
R7947 vdd3p3.n5697 vdd3p3.n5696 4.65
R7948 vdd3p3.n5692 vdd3p3.n5691 4.65
R7949 vdd3p3.n5687 vdd3p3.n5686 4.65
R7950 vdd3p3.n5682 vdd3p3.n5681 4.65
R7951 vdd3p3.n5677 vdd3p3.n5676 4.65
R7952 vdd3p3.n5669 vdd3p3.n5668 4.65
R7953 vdd3p3.n5664 vdd3p3.n5663 4.65
R7954 vdd3p3.n5659 vdd3p3.n5658 4.65
R7955 vdd3p3.n5654 vdd3p3.n5653 4.65
R7956 vdd3p3.n5649 vdd3p3.n5648 4.65
R7957 vdd3p3.n5644 vdd3p3.n5643 4.65
R7958 vdd3p3.n5639 vdd3p3.n5638 4.65
R7959 vdd3p3.n5634 vdd3p3.n5633 4.65
R7960 vdd3p3.n5629 vdd3p3.n5628 4.65
R7961 vdd3p3.n5624 vdd3p3.n5623 4.65
R7962 vdd3p3.n5619 vdd3p3.n5618 4.65
R7963 vdd3p3.n5614 vdd3p3.n5613 4.65
R7964 vdd3p3.n5609 vdd3p3.n5608 4.65
R7965 vdd3p3.n5604 vdd3p3.n5603 4.65
R7966 vdd3p3.n5599 vdd3p3.n5598 4.65
R7967 vdd3p3.n5594 vdd3p3.n5593 4.65
R7968 vdd3p3.n5589 vdd3p3.n5588 4.65
R7969 vdd3p3.n5581 vdd3p3.n5580 4.65
R7970 vdd3p3.n5576 vdd3p3.n5575 4.65
R7971 vdd3p3.n5571 vdd3p3.n5570 4.65
R7972 vdd3p3.n5566 vdd3p3.n5565 4.65
R7973 vdd3p3.n5561 vdd3p3.n5560 4.65
R7974 vdd3p3.n5556 vdd3p3.n5555 4.65
R7975 vdd3p3.n5551 vdd3p3.n5550 4.65
R7976 vdd3p3.n5546 vdd3p3.n5545 4.65
R7977 vdd3p3.n5541 vdd3p3.n5540 4.65
R7978 vdd3p3.n5536 vdd3p3.n5535 4.65
R7979 vdd3p3.n5531 vdd3p3.n5530 4.65
R7980 vdd3p3.n5526 vdd3p3.n5525 4.65
R7981 vdd3p3.n5521 vdd3p3.n5520 4.65
R7982 vdd3p3.n5516 vdd3p3.n5515 4.65
R7983 vdd3p3.n5511 vdd3p3.n5510 4.65
R7984 vdd3p3.n5506 vdd3p3.n5505 4.65
R7985 vdd3p3.n5501 vdd3p3.n5500 4.65
R7986 vdd3p3.n5493 vdd3p3.n5492 4.65
R7987 vdd3p3.n5488 vdd3p3.n5487 4.65
R7988 vdd3p3.n5483 vdd3p3.n5482 4.65
R7989 vdd3p3.n5478 vdd3p3.n5477 4.65
R7990 vdd3p3.n5473 vdd3p3.n5472 4.65
R7991 vdd3p3.n5468 vdd3p3.n5467 4.65
R7992 vdd3p3.n5463 vdd3p3.n5462 4.65
R7993 vdd3p3.n5458 vdd3p3.n5457 4.65
R7994 vdd3p3.n5453 vdd3p3.n5452 4.65
R7995 vdd3p3.n5448 vdd3p3.n5447 4.65
R7996 vdd3p3.n5443 vdd3p3.n5442 4.65
R7997 vdd3p3.n5438 vdd3p3.n5437 4.65
R7998 vdd3p3.n5433 vdd3p3.n5432 4.65
R7999 vdd3p3.n5428 vdd3p3.n5427 4.65
R8000 vdd3p3.n5423 vdd3p3.n5422 4.65
R8001 vdd3p3.n5418 vdd3p3.n5417 4.65
R8002 vdd3p3.n5413 vdd3p3.n5412 4.65
R8003 vdd3p3.n5405 vdd3p3.n5404 4.65
R8004 vdd3p3.n5400 vdd3p3.n5399 4.65
R8005 vdd3p3.n5395 vdd3p3.n5394 4.65
R8006 vdd3p3.n5390 vdd3p3.n5389 4.65
R8007 vdd3p3.n5385 vdd3p3.n5384 4.65
R8008 vdd3p3.n5380 vdd3p3.n5379 4.65
R8009 vdd3p3.n5375 vdd3p3.n5374 4.65
R8010 vdd3p3.n5370 vdd3p3.n5369 4.65
R8011 vdd3p3.n5365 vdd3p3.n5364 4.65
R8012 vdd3p3.n5360 vdd3p3.n5359 4.65
R8013 vdd3p3.n5355 vdd3p3.n5354 4.65
R8014 vdd3p3.n5350 vdd3p3.n5349 4.65
R8015 vdd3p3.n6722 vdd3p3.n6721 4.65
R8016 vdd3p3.n6727 vdd3p3.n6726 4.65
R8017 vdd3p3.n6732 vdd3p3.n6731 4.65
R8018 vdd3p3.n6737 vdd3p3.n6736 4.65
R8019 vdd3p3.n6745 vdd3p3.n6744 4.65
R8020 vdd3p3.n6750 vdd3p3.n6749 4.65
R8021 vdd3p3.n6755 vdd3p3.n6754 4.65
R8022 vdd3p3.n6760 vdd3p3.n6759 4.65
R8023 vdd3p3.n6765 vdd3p3.n6764 4.65
R8024 vdd3p3.n6770 vdd3p3.n6769 4.65
R8025 vdd3p3.n6775 vdd3p3.n6774 4.65
R8026 vdd3p3.n6780 vdd3p3.n6779 4.65
R8027 vdd3p3.n6785 vdd3p3.n6784 4.65
R8028 vdd3p3.n6790 vdd3p3.n6789 4.65
R8029 vdd3p3.n6795 vdd3p3.n6794 4.65
R8030 vdd3p3.n6800 vdd3p3.n6799 4.65
R8031 vdd3p3.n6805 vdd3p3.n6804 4.65
R8032 vdd3p3.n6810 vdd3p3.n6809 4.65
R8033 vdd3p3.n6815 vdd3p3.n6814 4.65
R8034 vdd3p3.n6820 vdd3p3.n6819 4.65
R8035 vdd3p3.n6825 vdd3p3.n6824 4.65
R8036 vdd3p3.n6833 vdd3p3.n6832 4.65
R8037 vdd3p3.n6838 vdd3p3.n6837 4.65
R8038 vdd3p3.n6843 vdd3p3.n6842 4.65
R8039 vdd3p3.n6848 vdd3p3.n6847 4.65
R8040 vdd3p3.n6853 vdd3p3.n6852 4.65
R8041 vdd3p3.n6858 vdd3p3.n6857 4.65
R8042 vdd3p3.n6863 vdd3p3.n6862 4.65
R8043 vdd3p3.n6868 vdd3p3.n6867 4.65
R8044 vdd3p3.n6873 vdd3p3.n6872 4.65
R8045 vdd3p3.n6878 vdd3p3.n6877 4.65
R8046 vdd3p3.n6883 vdd3p3.n6882 4.65
R8047 vdd3p3.n6888 vdd3p3.n6887 4.65
R8048 vdd3p3.n6893 vdd3p3.n6892 4.65
R8049 vdd3p3.n6898 vdd3p3.n6897 4.65
R8050 vdd3p3.n6903 vdd3p3.n6902 4.65
R8051 vdd3p3.n6908 vdd3p3.n6907 4.65
R8052 vdd3p3.n6913 vdd3p3.n6912 4.65
R8053 vdd3p3.n6921 vdd3p3.n6920 4.65
R8054 vdd3p3.n6926 vdd3p3.n6925 4.65
R8055 vdd3p3.n6931 vdd3p3.n6930 4.65
R8056 vdd3p3.n6936 vdd3p3.n6935 4.65
R8057 vdd3p3.n6941 vdd3p3.n6940 4.65
R8058 vdd3p3.n6946 vdd3p3.n6945 4.65
R8059 vdd3p3.n6951 vdd3p3.n6950 4.65
R8060 vdd3p3.n6956 vdd3p3.n6955 4.65
R8061 vdd3p3.n6961 vdd3p3.n6960 4.65
R8062 vdd3p3.n6966 vdd3p3.n6965 4.65
R8063 vdd3p3.n6971 vdd3p3.n6970 4.65
R8064 vdd3p3.n6976 vdd3p3.n6975 4.65
R8065 vdd3p3.n6981 vdd3p3.n6980 4.65
R8066 vdd3p3.n6986 vdd3p3.n6985 4.65
R8067 vdd3p3.n6991 vdd3p3.n6990 4.65
R8068 vdd3p3.n6996 vdd3p3.n6995 4.65
R8069 vdd3p3.n7001 vdd3p3.n7000 4.65
R8070 vdd3p3.n7016 vdd3p3.n7015 4.65
R8071 vdd3p3.n6388 vdd3p3.n6387 4.65
R8072 vdd3p3.n6383 vdd3p3.n6382 4.65
R8073 vdd3p3.n6379 vdd3p3.n6378 4.65
R8074 vdd3p3.n6374 vdd3p3.n6373 4.65
R8075 vdd3p3.n6370 vdd3p3.n6369 4.65
R8076 vdd3p3.n6365 vdd3p3.n6364 4.65
R8077 vdd3p3.n6361 vdd3p3.n6360 4.65
R8078 vdd3p3.n6354 vdd3p3.n6353 4.65
R8079 vdd3p3.n6350 vdd3p3.n6349 4.65
R8080 vdd3p3.n6345 vdd3p3.n6344 4.65
R8081 vdd3p3.n6341 vdd3p3.n6340 4.65
R8082 vdd3p3.n6336 vdd3p3.n6335 4.65
R8083 vdd3p3.n6332 vdd3p3.n6331 4.65
R8084 vdd3p3.n6327 vdd3p3.n6326 4.65
R8085 vdd3p3.n6323 vdd3p3.n6322 4.65
R8086 vdd3p3.n6318 vdd3p3.n6317 4.65
R8087 vdd3p3.n6313 vdd3p3.n6312 4.65
R8088 vdd3p3.n6309 vdd3p3.n6308 4.65
R8089 vdd3p3.n6304 vdd3p3.n6303 4.65
R8090 vdd3p3.n6300 vdd3p3.n6299 4.65
R8091 vdd3p3.n6295 vdd3p3.n6294 4.65
R8092 vdd3p3.n6291 vdd3p3.n6290 4.65
R8093 vdd3p3.n6286 vdd3p3.n6285 4.65
R8094 vdd3p3.n6282 vdd3p3.n6281 4.65
R8095 vdd3p3.n6275 vdd3p3.n6274 4.65
R8096 vdd3p3.n6271 vdd3p3.n6270 4.65
R8097 vdd3p3.n6266 vdd3p3.n6265 4.65
R8098 vdd3p3.n6261 vdd3p3.n6260 4.65
R8099 vdd3p3.n6256 vdd3p3.n6255 4.65
R8100 vdd3p3.n6251 vdd3p3.n6250 4.65
R8101 vdd3p3.n6246 vdd3p3.n6245 4.65
R8102 vdd3p3.n6241 vdd3p3.n6240 4.65
R8103 vdd3p3.n6236 vdd3p3.n6235 4.65
R8104 vdd3p3.n6231 vdd3p3.n6230 4.65
R8105 vdd3p3.n6226 vdd3p3.n6225 4.65
R8106 vdd3p3.n6221 vdd3p3.n6220 4.65
R8107 vdd3p3.n6216 vdd3p3.n6215 4.65
R8108 vdd3p3.n6211 vdd3p3.n6210 4.65
R8109 vdd3p3.n6206 vdd3p3.n6205 4.65
R8110 vdd3p3.n6201 vdd3p3.n6200 4.65
R8111 vdd3p3.n6196 vdd3p3.n6195 4.65
R8112 vdd3p3.n6188 vdd3p3.n6187 4.65
R8113 vdd3p3.n6183 vdd3p3.n6182 4.65
R8114 vdd3p3.n6178 vdd3p3.n6177 4.65
R8115 vdd3p3.n6173 vdd3p3.n6172 4.65
R8116 vdd3p3.n6168 vdd3p3.n6167 4.65
R8117 vdd3p3.n6163 vdd3p3.n6162 4.65
R8118 vdd3p3.n6158 vdd3p3.n6157 4.65
R8119 vdd3p3.n6153 vdd3p3.n6152 4.65
R8120 vdd3p3.n6148 vdd3p3.n6147 4.65
R8121 vdd3p3.n6143 vdd3p3.n6142 4.65
R8122 vdd3p3.n6138 vdd3p3.n6137 4.65
R8123 vdd3p3.n6133 vdd3p3.n6132 4.65
R8124 vdd3p3.n6128 vdd3p3.n6127 4.65
R8125 vdd3p3.n6123 vdd3p3.n6122 4.65
R8126 vdd3p3.n6118 vdd3p3.n6117 4.65
R8127 vdd3p3.n6114 vdd3p3.n6113 4.65
R8128 vdd3p3.n6110 vdd3p3.n6109 4.65
R8129 vdd3p3.n6104 vdd3p3.n6103 4.65
R8130 vdd3p3.n6100 vdd3p3.n6099 4.65
R8131 vdd3p3.n6096 vdd3p3.n6095 4.65
R8132 vdd3p3.n6092 vdd3p3.n6091 4.65
R8133 vdd3p3.n6088 vdd3p3.n6087 4.65
R8134 vdd3p3.n6084 vdd3p3.n6083 4.65
R8135 vdd3p3.n6080 vdd3p3.n6079 4.65
R8136 vdd3p3.n6076 vdd3p3.n6075 4.65
R8137 vdd3p3.n6072 vdd3p3.n6071 4.65
R8138 vdd3p3.n6068 vdd3p3.n6067 4.65
R8139 vdd3p3.n6064 vdd3p3.n6063 4.65
R8140 vdd3p3.n6060 vdd3p3.n6059 4.65
R8141 vdd3p3.n6056 vdd3p3.n6055 4.65
R8142 vdd3p3.n6052 vdd3p3.n6051 4.65
R8143 vdd3p3.n6048 vdd3p3.n6047 4.65
R8144 vdd3p3.n6044 vdd3p3.n6043 4.65
R8145 vdd3p3.n6040 vdd3p3.n6039 4.65
R8146 vdd3p3.n6034 vdd3p3.n6033 4.65
R8147 vdd3p3.n6030 vdd3p3.n6029 4.65
R8148 vdd3p3.n6026 vdd3p3.n6025 4.65
R8149 vdd3p3.n6022 vdd3p3.n6021 4.65
R8150 vdd3p3.n6018 vdd3p3.n6017 4.65
R8151 vdd3p3.n6014 vdd3p3.n6013 4.65
R8152 vdd3p3.n6010 vdd3p3.n6009 4.65
R8153 vdd3p3.n6006 vdd3p3.n6005 4.65
R8154 vdd3p3.n6002 vdd3p3.n6001 4.65
R8155 vdd3p3.n5998 vdd3p3.n5997 4.65
R8156 vdd3p3.n5994 vdd3p3.n5993 4.65
R8157 vdd3p3.n5990 vdd3p3.n5989 4.65
R8158 vdd3p3.n5986 vdd3p3.n5985 4.65
R8159 vdd3p3.n5982 vdd3p3.n5981 4.65
R8160 vdd3p3.n5978 vdd3p3.n5977 4.65
R8161 vdd3p3.n5974 vdd3p3.n5973 4.65
R8162 vdd3p3.n5970 vdd3p3.n5969 4.65
R8163 vdd3p3.n5964 vdd3p3.n5963 4.65
R8164 vdd3p3.n5960 vdd3p3.n5959 4.65
R8165 vdd3p3.n5956 vdd3p3.n5955 4.65
R8166 vdd3p3.n5952 vdd3p3.n5951 4.65
R8167 vdd3p3.n5947 vdd3p3.n5946 4.65
R8168 vdd3p3.n5942 vdd3p3.n5941 4.65
R8169 vdd3p3.n5937 vdd3p3.n5936 4.65
R8170 vdd3p3.n5932 vdd3p3.n5931 4.65
R8171 vdd3p3.n5927 vdd3p3.n5926 4.65
R8172 vdd3p3.n5922 vdd3p3.n5921 4.65
R8173 vdd3p3.n5917 vdd3p3.n5916 4.65
R8174 vdd3p3.n5912 vdd3p3.n5911 4.65
R8175 vdd3p3.n5907 vdd3p3.n5906 4.65
R8176 vdd3p3.n5902 vdd3p3.n5901 4.65
R8177 vdd3p3.n5897 vdd3p3.n5896 4.65
R8178 vdd3p3.n5892 vdd3p3.n5891 4.65
R8179 vdd3p3.n5887 vdd3p3.n5886 4.65
R8180 vdd3p3.n5879 vdd3p3.n5878 4.65
R8181 vdd3p3.n5874 vdd3p3.n5873 4.65
R8182 vdd3p3.n5869 vdd3p3.n5868 4.65
R8183 vdd3p3.n5864 vdd3p3.n5863 4.65
R8184 vdd3p3.n5859 vdd3p3.n5858 4.65
R8185 vdd3p3.n5854 vdd3p3.n5853 4.65
R8186 vdd3p3.n5849 vdd3p3.n5848 4.65
R8187 vdd3p3.n5844 vdd3p3.n5843 4.65
R8188 vdd3p3.n5839 vdd3p3.n5838 4.65
R8189 vdd3p3.n5834 vdd3p3.n5833 4.65
R8190 vdd3p3.n5829 vdd3p3.n5828 4.65
R8191 vdd3p3.n5824 vdd3p3.n5823 4.65
R8192 vdd3p3.n5819 vdd3p3.n5818 4.65
R8193 vdd3p3.n5814 vdd3p3.n5813 4.65
R8194 vdd3p3.n5809 vdd3p3.n5808 4.65
R8195 vdd3p3.n5804 vdd3p3.n5803 4.65
R8196 vdd3p3.n5799 vdd3p3.n5798 4.65
R8197 vdd3p3.n5791 vdd3p3.n5790 4.65
R8198 vdd3p3.n5786 vdd3p3.n5785 4.65
R8199 vdd3p3.n5781 vdd3p3.n5780 4.65
R8200 vdd3p3.n5776 vdd3p3.n5775 4.65
R8201 vdd3p3.n5771 vdd3p3.n5770 4.65
R8202 vdd3p3.n5766 vdd3p3.n5765 4.65
R8203 vdd3p3.n5761 vdd3p3.n5760 4.65
R8204 vdd3p3.n6398 vdd3p3.n6397 4.65
R8205 vdd3p3.n5751 vdd3p3.n5750 4.65
R8206 vdd3p3.n5746 vdd3p3.n5745 4.65
R8207 vdd3p3.n5741 vdd3p3.n5740 4.65
R8208 vdd3p3.n5756 vdd3p3.n5755 4.65
R8209 vdd3p3.n7022 vdd3p3.n7018 4.581
R8210 vdd3p3.n3456 vdd3p3.n3455 4.534
R8211 vdd3p3.n4217 vdd3p3.n4216 4.517
R8212 vdd3p3.n5069 vdd3p3.n5068 4.517
R8213 vdd3p3.n3597 vdd3p3.n3596 4.517
R8214 vdd3p3.n3691 vdd3p3.n3690 4.517
R8215 vdd3p3.n3761 vdd3p3.n3760 4.517
R8216 vdd3p3.n3510 vdd3p3.n3509 4.517
R8217 vdd3p3.n4826 vdd3p3.n4825 4.517
R8218 vdd3p3.n4757 vdd3p3.n4756 4.517
R8219 vdd3p3.n4992 vdd3p3.n4991 4.517
R8220 vdd3p3.n8488 vdd3p3.n8487 4.517
R8221 vdd3p3.n8497 vdd3p3.n8496 4.517
R8222 vdd3p3.n8566 vdd3p3.n8565 4.517
R8223 vdd3p3.n8617 vdd3p3.n8616 4.517
R8224 vdd3p3.n8841 vdd3p3.n8840 4.517
R8225 vdd3p3.n8750 vdd3p3.n8749 4.517
R8226 vdd3p3.n8783 vdd3p3.n8782 4.517
R8227 vdd3p3.n3666 vdd3p3.n3603 4.5
R8228 vdd3p3.n3737 vdd3p3.n3697 4.5
R8229 vdd3p3.n3570 vdd3p3.n3516 4.5
R8230 vdd3p3.n3751 vdd3p3.n3750 4.5
R8231 vdd3p3.n3757 vdd3p3.n3756 4.5
R8232 vdd3p3.n3674 vdd3p3.n3673 4.5
R8233 vdd3p3.n3744 vdd3p3.n3743 4.5
R8234 vdd3p3.n3587 vdd3p3.n3586 4.5
R8235 vdd3p3.n3497 vdd3p3.n3496 4.5
R8236 vdd3p3.n3506 vdd3p3.n3505 4.5
R8237 vdd3p3.n3593 vdd3p3.n3592 4.5
R8238 vdd3p3.n3580 vdd3p3.n3579 4.5
R8239 vdd3p3.n3681 vdd3p3.n3680 4.5
R8240 vdd3p3.n3687 vdd3p3.n3686 4.5
R8241 vdd3p3.n3490 vdd3p3.n3489 4.5
R8242 vdd3p3.n4802 vdd3p3.n4765 4.5
R8243 vdd3p3.n4951 vdd3p3.n4906 4.5
R8244 vdd3p3.n4972 vdd3p3.n4971 4.5
R8245 vdd3p3.n4747 vdd3p3.n4746 4.5
R8246 vdd3p3.n4753 vdd3p3.n4752 4.5
R8247 vdd3p3.n4809 vdd3p3.n4808 4.5
R8248 vdd3p3.n4816 vdd3p3.n4815 4.5
R8249 vdd3p3.n4822 vdd3p3.n4821 4.5
R8250 vdd3p3.n4740 vdd3p3.n4739 4.5
R8251 vdd3p3.n4979 vdd3p3.n4978 4.5
R8252 vdd3p3.n4988 vdd3p3.n4987 4.5
R8253 vdd3p3.n8545 vdd3p3.n8544 4.5
R8254 vdd3p3.n8593 vdd3p3.n8592 4.5
R8255 vdd3p3.n8624 vdd3p3.n8623 4.5
R8256 vdd3p3.n8807 vdd3p3.n8806 4.5
R8257 vdd3p3.n8867 vdd3p3.n8842 4.5
R8258 vdd3p3.n8871 vdd3p3.n8835 4.5
R8259 vdd3p3.n8881 vdd3p3.n8880 4.5
R8260 vdd3p3.n8523 vdd3p3.n8498 4.5
R8261 vdd3p3.n8527 vdd3p3.n8491 4.5
R8262 vdd3p3.n8536 vdd3p3.n8535 4.5
R8263 vdd3p3.n8600 vdd3p3.n8599 4.5
R8264 vdd3p3.n8635 vdd3p3.n8634 4.5
R8265 vdd3p3.n8818 vdd3p3.n8817 4.5
R8266 vdd3p3.n8798 vdd3p3.n8797 4.5
R8267 vdd3p3.n8556 vdd3p3.n8555 4.5
R8268 vdd3p3.n8575 vdd3p3.n8574 4.5
R8269 vdd3p3.n8579 vdd3p3.n8569 4.5
R8270 vdd3p3.n8584 vdd3p3.n8583 4.5
R8271 vdd3p3.n8785 vdd3p3.n8784 4.5
R8272 vdd3p3.n8789 vdd3p3.n8753 4.5
R8273 vdd3p3.n8742 vdd3p3.n8741 4.5
R8274 vdd3p3.n8694 vdd3p3.n8693 4.5
R8275 vdd3p3.n3832 vdd3p3.n3831 4.5
R8276 vdd3p3.n3850 vdd3p3.n3822 4.5
R8277 vdd3p3.n3841 vdd3p3.n3840 4.5
R8278 vdd3p3.n3859 vdd3p3.n3858 4.5
R8279 vdd3p3.n3862 vdd3p3.n3817 4.5
R8280 vdd3p3.n3869 vdd3p3.n3868 4.5
R8281 vdd3p3.n3872 vdd3p3.n3814 4.5
R8282 vdd3p3.n4671 vdd3p3.n4574 4.5
R8283 vdd3p3.n4560 vdd3p3.n4559 4.5
R8284 vdd3p3.n5121 vdd3p3.n5120 4.5
R8285 vdd3p3.n4515 vdd3p3.n4501 4.5
R8286 vdd3p3.n5095 vdd3p3.n5044 4.5
R8287 vdd3p3.n5089 vdd3p3.n5088 4.5
R8288 vdd3p3.n4681 vdd3p3.n4680 4.5
R8289 vdd3p3.n5128 vdd3p3.n5126 4.5
R8290 vdd3p3.n3436 vdd3p3.n3433 4.5
R8291 vdd3p3.n3429 vdd3p3.n3428 4.5
R8292 vdd3p3.n3448 vdd3p3.n3443 4.5
R8293 vdd3p3.n4479 vdd3p3.n4474 4.5
R8294 vdd3p3.n4509 vdd3p3.n4504 4.5
R8295 vdd3p3.n4449 vdd3p3.n4444 4.5
R8296 vdd3p3.n4455 vdd3p3.n4441 4.5
R8297 vdd3p3.n4485 vdd3p3.n4471 4.5
R8298 vdd3p3.n4425 vdd3p3.n4411 4.5
R8299 vdd3p3.n4351 vdd3p3.n4254 4.5
R8300 vdd3p3.n4229 vdd3p3.n4192 4.5
R8301 vdd3p3.n4235 vdd3p3.n4184 4.5
R8302 vdd3p3.n4395 vdd3p3.n4377 4.5
R8303 vdd3p3.n4419 vdd3p3.n4414 4.5
R8304 vdd3p3.n4389 vdd3p3.n4388 4.5
R8305 vdd3p3.n4361 vdd3p3.n4360 4.5
R8306 vdd3p3.n3394 vdd3p3.n3393 4.482
R8307 vdd3p3.n3956 vdd3p3.n3955 4.364
R8308 vdd3p3.n8674 vdd3p3.n8673 4.313
R8309 vdd3p3.n5027 vdd3p3.n5026 4.313
R8310 vdd3p3.n4693 vdd3p3.n4691 4.313
R8311 vdd3p3.n5016 vdd3p3.n5013 4.313
R8312 vdd3p3.n4163 vdd3p3.n4162 4.313
R8313 vdd3p3.n4160 vdd3p3.n4159 4.313
R8314 vdd3p3.n4167 vdd3p3.n4166 4.313
R8315 vdd3p3.n8742 vdd3p3.n8739 4.312
R8316 vdd3p3.n4200 vdd3p3.n4193 4.236
R8317 vdd3p3.n5052 vdd3p3.n5045 4.236
R8318 vdd3p3.n3477 vdd3p3.n3471 4.236
R8319 vdd3p3.n8761 vdd3p3.n8754 4.236
R8320 vdd3p3.n4959 vdd3p3.n4952 4.235
R8321 vdd3p3.n8506 vdd3p3.n8499 4.235
R8322 vdd3p3.n8850 vdd3p3.n8843 4.235
R8323 vdd3p3.n3897 vdd3p3.n3896 4.219
R8324 vdd3p3.n4147 vdd3p3.n4146 4.184
R8325 vdd3p3.n3353 vdd3p3.n3352 4.173
R8326 vdd3p3.n2507 vdd3p3.n2506 4.173
R8327 vdd3p3.n1662 vdd3p3.n1661 4.173
R8328 vdd3p3.n816 vdd3p3.n815 4.173
R8329 vdd3p3.n4239 vdd3p3.n4238 4.141
R8330 vdd3p3.n5099 vdd3p3.n5098 4.141
R8331 vdd3p3.n3592 vdd3p3.n3589 4.141
R8332 vdd3p3.n3686 vdd3p3.n3683 4.141
R8333 vdd3p3.n3756 vdd3p3.n3753 4.141
R8334 vdd3p3.n3505 vdd3p3.n3499 4.141
R8335 vdd3p3.n4821 vdd3p3.n4818 4.141
R8336 vdd3p3.n4752 vdd3p3.n4749 4.141
R8337 vdd3p3.n4987 vdd3p3.n4981 4.141
R8338 vdd3p3.n4933 vdd3p3.n4929 4.141
R8339 vdd3p3.n8364 vdd3p3.t48 4.099
R8340 vdd3p3.n6396 vdd3p3.n6394 4.049
R8341 vdd3p3.n3396 vdd3p3.n3382 4.035
R8342 vdd3p3.n3396 vdd3p3.n3383 4.035
R8343 vdd3p3.n7471 vdd3p3.n7470 3.943
R8344 vdd3p3.n7930 vdd3p3.n7927 3.928
R8345 vdd3p3.n3394 vdd3p3.n3387 3.788
R8346 vdd3p3.n3145 vdd3p3.n3076 3.784
R8347 vdd3p3.n3375 vdd3p3.n2608 3.784
R8348 vdd3p3.n3355 vdd3p3.n2635 3.784
R8349 vdd3p3.n2299 vdd3p3.n2230 3.784
R8350 vdd3p3.n2529 vdd3p3.n1762 3.784
R8351 vdd3p3.n2509 vdd3p3.n1789 3.784
R8352 vdd3p3.n1454 vdd3p3.n1385 3.784
R8353 vdd3p3.n1684 vdd3p3.n917 3.784
R8354 vdd3p3.n1664 vdd3p3.n944 3.784
R8355 vdd3p3.n608 vdd3p3.n539 3.784
R8356 vdd3p3.n838 vdd3p3.n71 3.784
R8357 vdd3p3.n818 vdd3p3.n98 3.784
R8358 vdd3p3.t96 vdd3p3.n5266 3.784
R8359 vdd3p3.n4192 vdd3p3.n4185 3.764
R8360 vdd3p3.n4187 vdd3p3.n4186 3.764
R8361 vdd3p3.n4254 vdd3p3.n4251 3.764
R8362 vdd3p3.n4388 vdd3p3.n4386 3.764
R8363 vdd3p3.n4414 vdd3p3.n4412 3.764
R8364 vdd3p3.n4444 vdd3p3.n4442 3.764
R8365 vdd3p3.n4474 vdd3p3.n4472 3.764
R8366 vdd3p3.n4504 vdd3p3.n4502 3.764
R8367 vdd3p3.n3443 vdd3p3.n3441 3.764
R8368 vdd3p3.n4559 vdd3p3.n4557 3.764
R8369 vdd3p3.n4574 vdd3p3.n4571 3.764
R8370 vdd3p3.n5088 vdd3p3.n5081 3.764
R8371 vdd3p3.n5083 vdd3p3.n5082 3.764
R8372 vdd3p3.n8534 vdd3p3.n8533 3.764
R8373 vdd3p3.n3393 vdd3p3.n3389 3.764
R8374 vdd3p3.n8879 vdd3p3.n8878 3.764
R8375 vdd3p3.n8796 vdd3p3.n8795 3.764
R8376 vdd3p3.n8666 vdd3p3.n8665 3.74
R8377 vdd3p3.n7945 vdd3p3.n7944 3.738
R8378 vdd3p3.n3955 vdd3p3.n3918 3.703
R8379 vdd3p3.n36 vdd3p3.n35 3.678
R8380 vdd3p3.n889 vdd3p3.n888 3.678
R8381 vdd3p3.n1727 vdd3p3.n1726 3.678
R8382 vdd3p3.n2580 vdd3p3.n2579 3.678
R8383 vdd3p3.n2984 vdd3p3.n2975 3.642
R8384 vdd3p3.n2138 vdd3p3.n2129 3.642
R8385 vdd3p3.n1293 vdd3p3.n1284 3.642
R8386 vdd3p3.n447 vdd3p3.n438 3.642
R8387 vdd3p3.n8654 vdd3p3.n8653 3.443
R8388 vdd3p3.n906 vdd3p3.n899 3.434
R8389 vdd3p3.n2597 vdd3p3.n2590 3.434
R8390 vdd3p3.n4774 vdd3p3.n4767 3.427
R8391 vdd3p3.n4915 vdd3p3.n4908 3.427
R8392 vdd3p3.n4279 vdd3p3.n4272 3.427
R8393 vdd3p3.n4599 vdd3p3.n4592 3.427
R8394 vdd3p3.n3709 vdd3p3.n3702 3.427
R8395 vdd3p3.n4263 vdd3p3.n4256 3.426
R8396 vdd3p3.n4583 vdd3p3.n4576 3.426
R8397 vdd3p3.n3525 vdd3p3.n3518 3.426
R8398 vdd3p3.n2888 vdd3p3.n2838 3.421
R8399 vdd3p3.n2042 vdd3p3.n1992 3.421
R8400 vdd3p3.n1197 vdd3p3.n1147 3.421
R8401 vdd3p3.n351 vdd3p3.n301 3.421
R8402 vdd3p3.n3185 vdd3p3.n3017 3.393
R8403 vdd3p3.n2339 vdd3p3.n2171 3.393
R8404 vdd3p3.n1494 vdd3p3.n1326 3.393
R8405 vdd3p3.n648 vdd3p3.n480 3.393
R8406 vdd3p3.n4184 vdd3p3.n4183 3.388
R8407 vdd3p3.n4183 vdd3p3.n4179 3.388
R8408 vdd3p3.n4360 vdd3p3.n4359 3.388
R8409 vdd3p3.n4377 vdd3p3.n4376 3.388
R8410 vdd3p3.n4411 vdd3p3.n4410 3.388
R8411 vdd3p3.n4441 vdd3p3.n4440 3.388
R8412 vdd3p3.n4471 vdd3p3.n4470 3.388
R8413 vdd3p3.n4501 vdd3p3.n4500 3.388
R8414 vdd3p3.n3428 vdd3p3.n3427 3.388
R8415 vdd3p3.n5120 vdd3p3.n5119 3.388
R8416 vdd3p3.n4680 vdd3p3.n4679 3.388
R8417 vdd3p3.n5044 vdd3p3.n5043 3.388
R8418 vdd3p3.n5043 vdd3p3.n5039 3.388
R8419 vdd3p3.n3516 vdd3p3.n3513 3.388
R8420 vdd3p3.n3603 vdd3p3.n3600 3.388
R8421 vdd3p3.n3697 vdd3p3.n3694 3.388
R8422 vdd3p3.n4765 vdd3p3.n4762 3.388
R8423 vdd3p3.n4906 vdd3p3.n4900 3.388
R8424 vdd3p3.n4944 vdd3p3.n4940 3.388
R8425 vdd3p3.n5017 vdd3p3.n5016 3.339
R8426 vdd3p3.n5025 vdd3p3.n4693 3.339
R8427 vdd3p3.n5027 vdd3p3.n5025 3.339
R8428 vdd3p3.n4727 vdd3p3.n4726 3.339
R8429 vdd3p3.n5010 vdd3p3.n5009 3.339
R8430 vdd3p3.n3995 vdd3p3.n3994 3.339
R8431 vdd3p3.n3985 vdd3p3.n3982 3.339
R8432 vdd3p3.n4160 vdd3p3.n4158 3.339
R8433 vdd3p3.n4198 vdd3p3.n4197 3.293
R8434 vdd3p3.n5050 vdd3p3.n5049 3.293
R8435 vdd3p3.n3475 vdd3p3.n3474 3.293
R8436 vdd3p3.n4957 vdd3p3.n4956 3.293
R8437 vdd3p3.n8504 vdd3p3.n8503 3.293
R8438 vdd3p3.n8848 vdd3p3.n8847 3.293
R8439 vdd3p3.n8759 vdd3p3.n8758 3.293
R8440 vdd3p3.n8707 vdd3p3.n8705 3.252
R8441 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_1.vdd3p3 3.22
R8442 vdd3p3.n47 vdd3p3.n45 3.206
R8443 vdd3p3.n1738 vdd3p3.n1736 3.206
R8444 vdd3p3.n3974 vdd3p3.n3973 3.174
R8445 vdd3p3.n3896 vdd3p3.n3895 3.174
R8446 vdd3p3.n3158 vdd3p3.n3034 3.172
R8447 vdd3p3.n3157 vdd3p3.n3156 3.172
R8448 vdd3p3.n3155 vdd3p3.n3039 3.172
R8449 vdd3p3.n2312 vdd3p3.n2188 3.172
R8450 vdd3p3.n2311 vdd3p3.n2310 3.172
R8451 vdd3p3.n2309 vdd3p3.n2193 3.172
R8452 vdd3p3.n1467 vdd3p3.n1343 3.172
R8453 vdd3p3.n1466 vdd3p3.n1465 3.172
R8454 vdd3p3.n1464 vdd3p3.n1348 3.172
R8455 vdd3p3.n621 vdd3p3.n497 3.172
R8456 vdd3p3.n620 vdd3p3.n619 3.172
R8457 vdd3p3.n618 vdd3p3.n502 3.172
R8458 vdd3p3.n3909 vdd3p3.n3903 3.166
R8459 vdd3p3.n8736 vdd3p3.n8735 3.118
R8460 vdd3p3.n5261 vdd3p3.n5258 3.108
R8461 vdd3p3.n5258 vdd3p3.n5255 3.108
R8462 vdd3p3.n5255 vdd3p3.n5252 3.108
R8463 vdd3p3.n5252 vdd3p3.n5249 3.108
R8464 vdd3p3.n5249 vdd3p3.n5246 3.108
R8465 vdd3p3.n5246 vdd3p3.n5243 3.108
R8466 vdd3p3.n5243 vdd3p3.n5240 3.108
R8467 vdd3p3.n5240 vdd3p3.n5237 3.108
R8468 vdd3p3.n5237 vdd3p3.n5234 3.108
R8469 vdd3p3.n5234 vdd3p3.n5231 3.108
R8470 vdd3p3.n5231 vdd3p3.n5228 3.108
R8471 vdd3p3.n5228 vdd3p3.n5225 3.108
R8472 vdd3p3.n5225 vdd3p3.n5222 3.108
R8473 vdd3p3.n5222 vdd3p3.n5219 3.108
R8474 vdd3p3.n5219 vdd3p3.n5216 3.108
R8475 vdd3p3.n5216 vdd3p3.n5213 3.108
R8476 vdd3p3.n5213 vdd3p3.n5210 3.108
R8477 vdd3p3.n5210 vdd3p3.n5207 3.108
R8478 vdd3p3.n5207 vdd3p3.n5204 3.108
R8479 vdd3p3.n5204 vdd3p3.n5202 3.108
R8480 vdd3p3.n5202 vdd3p3.n5200 3.108
R8481 vdd3p3.n5200 vdd3p3.n5198 3.108
R8482 vdd3p3.n5198 vdd3p3.n5196 3.108
R8483 vdd3p3.n5196 vdd3p3.n5194 3.108
R8484 vdd3p3.n18 vdd3p3.n17 3.101
R8485 vdd3p3.n864 vdd3p3.n858 3.101
R8486 vdd3p3.n1709 vdd3p3.n1708 3.101
R8487 vdd3p3.n2555 vdd3p3.n2549 3.101
R8488 vdd3p3.n10 vdd3p3.n2 3.098
R8489 vdd3p3.n879 vdd3p3.n878 3.098
R8490 vdd3p3.n1701 vdd3p3.n1693 3.098
R8491 vdd3p3.n2570 vdd3p3.n2569 3.098
R8492 vdd3p3.n3511 vdd3p3.n3510 3.033
R8493 vdd3p3.n3598 vdd3p3.n3597 3.033
R8494 vdd3p3.n3692 vdd3p3.n3691 3.033
R8495 vdd3p3.n3762 vdd3p3.n3761 3.033
R8496 vdd3p3.n4758 vdd3p3.n4757 3.033
R8497 vdd3p3.n4827 vdd3p3.n4826 3.033
R8498 vdd3p3.n4993 vdd3p3.n4992 3.033
R8499 vdd3p3.n8539 vdd3p3.n8488 3.033
R8500 vdd3p3.n8618 vdd3p3.n8617 3.033
R8501 vdd3p3.n8801 vdd3p3.n8750 3.033
R8502 vdd3p3.n8587 vdd3p3.n8566 3.033
R8503 vdd3p3.n8738 vdd3p3.n8737 3.033
R8504 vdd3p3.n8699 vdd3p3.n8698 3.033
R8505 vdd3p3.n8668 vdd3p3.n8667 3.033
R8506 vdd3p3.n8656 vdd3p3.n8655 3.033
R8507 vdd3p3.n8675 vdd3p3.n8674 3.033
R8508 vdd3p3.n3986 vdd3p3.n3985 3.033
R8509 vdd3p3.n5009 vdd3p3.n5006 3.033
R8510 vdd3p3.n4731 vdd3p3.n4730 3.033
R8511 vdd3p3.n5028 vdd3p3.n5027 3.033
R8512 vdd3p3.n4728 vdd3p3.n4727 3.033
R8513 vdd3p3.n3464 vdd3p3.n3463 3.033
R8514 vdd3p3.n3462 vdd3p3.n3461 3.033
R8515 vdd3p3.n3457 vdd3p3.n3456 3.033
R8516 vdd3p3.n4164 vdd3p3.n4163 3.033
R8517 vdd3p3.n3853 vdd3p3.n3820 3.033
R8518 vdd3p3.n4693 vdd3p3.n4692 3.033
R8519 vdd3p3.n4168 vdd3p3.n4167 3.033
R8520 vdd3p3.n3996 vdd3p3.n3995 3.033
R8521 vdd3p3.n3991 vdd3p3.n3990 3.033
R8522 vdd3p3.n4161 vdd3p3.n4160 3.033
R8523 vdd3p3.n5016 vdd3p3.n5015 3.033
R8524 vdd3p3.n4184 vdd3p3.n4177 3.011
R8525 vdd3p3.n4179 vdd3p3.n4178 3.011
R8526 vdd3p3.n4360 vdd3p3.n4357 3.011
R8527 vdd3p3.n4377 vdd3p3.n4374 3.011
R8528 vdd3p3.n4411 vdd3p3.n4408 3.011
R8529 vdd3p3.n4441 vdd3p3.n4438 3.011
R8530 vdd3p3.n4471 vdd3p3.n4468 3.011
R8531 vdd3p3.n4501 vdd3p3.n4498 3.011
R8532 vdd3p3.n3433 vdd3p3.n3432 3.011
R8533 vdd3p3.n3428 vdd3p3.n3425 3.011
R8534 vdd3p3.n5126 vdd3p3.n5125 3.011
R8535 vdd3p3.n5120 vdd3p3.n5117 3.011
R8536 vdd3p3.n4680 vdd3p3.n4677 3.011
R8537 vdd3p3.n5044 vdd3p3.n5037 3.011
R8538 vdd3p3.n5039 vdd3p3.n5038 3.011
R8539 vdd3p3.n4940 vdd3p3.n4939 3.011
R8540 vdd3p3.n8554 vdd3p3.n8553 3.011
R8541 vdd3p3.n8633 vdd3p3.n8632 3.011
R8542 vdd3p3.n8816 vdd3p3.n8815 3.011
R8543 vdd3p3.n3858 vdd3p3.n3857 3.011
R8544 vdd3p3.n3820 vdd3p3.n3819 3.011
R8545 vdd3p3.n3516 vdd3p3.n3515 2.959
R8546 vdd3p3.n3603 vdd3p3.n3602 2.959
R8547 vdd3p3.n3697 vdd3p3.n3696 2.959
R8548 vdd3p3.n4765 vdd3p3.n4764 2.959
R8549 vdd3p3.n4035 vdd3p3.n4034 2.909
R8550 vdd3p3.n7454 vdd3p3.n7450 2.886
R8551 vdd3p3.n3824 vdd3p3.t154 2.769
R8552 vdd3p3.n3824 vdd3p3.t86 2.769
R8553 vdd3p3.n3320 vdd3p3.n2684 2.645
R8554 vdd3p3.n2474 vdd3p3.n1838 2.645
R8555 vdd3p3.n1629 vdd3p3.n993 2.645
R8556 vdd3p3.n783 vdd3p3.n147 2.645
R8557 vdd3p3.n4058 vdd3p3.n4057 2.645
R8558 vdd3p3.n4146 vdd3p3.n4145 2.645
R8559 vdd3p3.n4192 vdd3p3.n4191 2.635
R8560 vdd3p3.n4191 vdd3p3.n4187 2.635
R8561 vdd3p3.n4254 vdd3p3.n4253 2.635
R8562 vdd3p3.n4388 vdd3p3.n4387 2.635
R8563 vdd3p3.n4414 vdd3p3.n4413 2.635
R8564 vdd3p3.n4444 vdd3p3.n4443 2.635
R8565 vdd3p3.n4474 vdd3p3.n4473 2.635
R8566 vdd3p3.n4504 vdd3p3.n4503 2.635
R8567 vdd3p3.n3443 vdd3p3.n3442 2.635
R8568 vdd3p3.n4559 vdd3p3.n4558 2.635
R8569 vdd3p3.n4574 vdd3p3.n4573 2.635
R8570 vdd3p3.n5088 vdd3p3.n5087 2.635
R8571 vdd3p3.n5087 vdd3p3.n5083 2.635
R8572 vdd3p3.n4905 vdd3p3.n4904 2.635
R8573 vdd3p3.n8555 vdd3p3.n8552 2.635
R8574 vdd3p3.n8599 vdd3p3.n8597 2.635
R8575 vdd3p3.n3389 vdd3p3.n3388 2.635
R8576 vdd3p3.n8634 vdd3p3.n8631 2.635
R8577 vdd3p3.n8817 vdd3p3.n8814 2.635
R8578 vdd3p3.n3868 vdd3p3.n3867 2.635
R8579 vdd3p3.n3183 vdd3p3.n3182 2.567
R8580 vdd3p3.n3090 vdd3p3.n3032 2.567
R8581 vdd3p3.n3091 vdd3p3.n3090 2.567
R8582 vdd3p3.n3096 vdd3p3.n3094 2.567
R8583 vdd3p3.n3098 vdd3p3.n3096 2.567
R8584 vdd3p3.n3117 vdd3p3.n3115 2.567
R8585 vdd3p3.n2337 vdd3p3.n2336 2.567
R8586 vdd3p3.n2244 vdd3p3.n2186 2.567
R8587 vdd3p3.n2245 vdd3p3.n2244 2.567
R8588 vdd3p3.n2250 vdd3p3.n2248 2.567
R8589 vdd3p3.n2252 vdd3p3.n2250 2.567
R8590 vdd3p3.n2271 vdd3p3.n2269 2.567
R8591 vdd3p3.n1492 vdd3p3.n1491 2.567
R8592 vdd3p3.n1399 vdd3p3.n1341 2.567
R8593 vdd3p3.n1400 vdd3p3.n1399 2.567
R8594 vdd3p3.n1405 vdd3p3.n1403 2.567
R8595 vdd3p3.n1407 vdd3p3.n1405 2.567
R8596 vdd3p3.n1426 vdd3p3.n1424 2.567
R8597 vdd3p3.n646 vdd3p3.n645 2.567
R8598 vdd3p3.n553 vdd3p3.n495 2.567
R8599 vdd3p3.n554 vdd3p3.n553 2.567
R8600 vdd3p3.n559 vdd3p3.n557 2.567
R8601 vdd3p3.n561 vdd3p3.n559 2.567
R8602 vdd3p3.n580 vdd3p3.n578 2.567
R8603 vdd3p3.n8589 vdd3p3.n8588 2.565
R8604 vdd3p3.n3069 vdd3p3.n2621 2.56
R8605 vdd3p3.n2634 vdd3p3.n2633 2.56
R8606 vdd3p3.n2223 vdd3p3.n1775 2.56
R8607 vdd3p3.n1788 vdd3p3.n1787 2.56
R8608 vdd3p3.n1378 vdd3p3.n930 2.56
R8609 vdd3p3.n943 vdd3p3.n942 2.56
R8610 vdd3p3.n532 vdd3p3.n84 2.56
R8611 vdd3p3.n97 vdd3p3.n96 2.56
R8612 vdd3p3.n6360 vdd3p3.n6356 2.531
R8613 vdd3p3.n6281 vdd3p3.n6277 2.531
R8614 vdd3p3.n6195 vdd3p3.n6191 2.531
R8615 vdd3p3.n6109 vdd3p3.n6106 2.531
R8616 vdd3p3.n6039 vdd3p3.n6036 2.531
R8617 vdd3p3.n5969 vdd3p3.n5966 2.531
R8618 vdd3p3.n5886 vdd3p3.n5882 2.531
R8619 vdd3p3.n5798 vdd3p3.n5794 2.531
R8620 comparator_top_0.VDD vdd3p3 2.509
R8621 vdd3p3.n7980 vdd3p3.n7975 2.438
R8622 vdd3p3.n8095 vdd3p3.n8090 2.438
R8623 vdd3p3.n8200 vdd3p3.n8195 2.438
R8624 vdd3p3.n8309 vdd3p3.n8300 2.438
R8625 vdd3p3.n3340 vdd3p3.n2670 2.435
R8626 vdd3p3.n2494 vdd3p3.n1824 2.435
R8627 vdd3p3.n1649 vdd3p3.n979 2.435
R8628 vdd3p3.n803 vdd3p3.n133 2.435
R8629 vdd3p3.n7376 vdd3p3.n7375 2.425
R8630 vdd3p3.n7307 vdd3p3.n7306 2.425
R8631 vdd3p3.n7238 vdd3p3.n7237 2.425
R8632 vdd3p3.n7153 vdd3p3.n7152 2.425
R8633 vdd3p3.n7066 vdd3p3.n7065 2.425
R8634 vdd3p3.n902 vdd3p3.n901 2.423
R8635 vdd3p3.n2593 vdd3p3.n2592 2.423
R8636 vdd3p3.n6360 vdd3p3.n6359 2.386
R8637 vdd3p3.n6281 vdd3p3.n6280 2.386
R8638 vdd3p3.n6195 vdd3p3.n6194 2.386
R8639 vdd3p3.n6109 vdd3p3.n6108 2.386
R8640 vdd3p3.n6039 vdd3p3.n6038 2.386
R8641 vdd3p3.n5969 vdd3p3.n5968 2.386
R8642 vdd3p3.n5886 vdd3p3.n5885 2.386
R8643 vdd3p3.n5798 vdd3p3.n5797 2.386
R8644 vdd3p3.n5740 vdd3p3.n5739 2.386
R8645 vdd3p3.n3824 vdd3p3.n3823 2.379
R8646 vdd3p3.n3396 vdd3p3.n3395 2.375
R8647 vdd3p3.n8462 vdd3p3.n8461 2.37
R8648 vdd3p3.n22 vdd3p3.n14 2.306
R8649 vdd3p3.n863 vdd3p3.n862 2.306
R8650 vdd3p3.n1713 vdd3p3.n1705 2.306
R8651 vdd3p3.n2554 vdd3p3.n2553 2.306
R8652 vdd3p3.n7015 vdd3p3.n7014 2.302
R8653 vdd3p3.n6920 vdd3p3.n6916 2.302
R8654 vdd3p3.n6920 vdd3p3.n6919 2.302
R8655 vdd3p3.n6832 vdd3p3.n6828 2.302
R8656 vdd3p3.n6832 vdd3p3.n6831 2.302
R8657 vdd3p3.n6744 vdd3p3.n6740 2.302
R8658 vdd3p3.n6744 vdd3p3.n6743 2.302
R8659 vdd3p3.n5412 vdd3p3.n5408 2.302
R8660 vdd3p3.n5412 vdd3p3.n5411 2.302
R8661 vdd3p3.n5500 vdd3p3.n5496 2.302
R8662 vdd3p3.n5500 vdd3p3.n5499 2.302
R8663 vdd3p3.n5588 vdd3p3.n5584 2.302
R8664 vdd3p3.n5588 vdd3p3.n5587 2.302
R8665 vdd3p3.n5676 vdd3p3.n5672 2.302
R8666 vdd3p3.n5676 vdd3p3.n5675 2.302
R8667 vdd3p3.n4238 vdd3p3.n4237 2.258
R8668 vdd3p3.n5098 vdd3p3.n5097 2.258
R8669 vdd3p3.n3585 vdd3p3.n3584 2.258
R8670 vdd3p3.n3679 vdd3p3.n3678 2.258
R8671 vdd3p3.n3749 vdd3p3.n3748 2.258
R8672 vdd3p3.n3495 vdd3p3.n3494 2.258
R8673 vdd3p3.n4814 vdd3p3.n4813 2.258
R8674 vdd3p3.n4745 vdd3p3.n4744 2.258
R8675 vdd3p3.n4977 vdd3p3.n4976 2.258
R8676 vdd3p3.n4929 vdd3p3.n4928 2.258
R8677 vdd3p3.n8535 vdd3p3.n8532 2.258
R8678 vdd3p3.n8490 vdd3p3.n8489 2.258
R8679 vdd3p3.n8583 vdd3p3.n8581 2.258
R8680 vdd3p3.n8568 vdd3p3.n8567 2.258
R8681 vdd3p3.n8880 vdd3p3.n8877 2.258
R8682 vdd3p3.n8834 vdd3p3.n8833 2.258
R8683 vdd3p3.n8797 vdd3p3.n8794 2.258
R8684 vdd3p3.n8752 vdd3p3.n8751 2.258
R8685 vdd3p3.n3822 vdd3p3.n3821 2.258
R8686 vdd3p3.n8583 vdd3p3.n8582 2.252
R8687 vdd3p3.n5131 vdd3p3.n4565 2.25
R8688 vdd3p3.n22 vdd3p3.n21 2.25
R8689 vdd3p3.n23 vdd3p3.n9 2.25
R8690 vdd3p3.n25 vdd3p3.n24 2.25
R8691 vdd3p3.n12 vdd3p3.n1 2.25
R8692 vdd3p3.n60 vdd3p3.n59 2.25
R8693 vdd3p3.n862 vdd3p3.n861 2.25
R8694 vdd3p3.n855 vdd3p3.n854 2.25
R8695 vdd3p3.n873 vdd3p3.n872 2.25
R8696 vdd3p3.n876 vdd3p3.n875 2.25
R8697 vdd3p3.n874 vdd3p3.n852 2.25
R8698 vdd3p3.n1713 vdd3p3.n1712 2.25
R8699 vdd3p3.n1714 vdd3p3.n1700 2.25
R8700 vdd3p3.n1716 vdd3p3.n1715 2.25
R8701 vdd3p3.n1703 vdd3p3.n1692 2.25
R8702 vdd3p3.n1751 vdd3p3.n1750 2.25
R8703 vdd3p3.n2553 vdd3p3.n2552 2.25
R8704 vdd3p3.n2546 vdd3p3.n2545 2.25
R8705 vdd3p3.n2564 vdd3p3.n2563 2.25
R8706 vdd3p3.n2567 vdd3p3.n2566 2.25
R8707 vdd3p3.n2565 vdd3p3.n2543 2.25
R8708 vdd3p3.n5131 vdd3p3.n5130 2.249
R8709 vdd3p3.n6364 vdd3p3.n6363 2.241
R8710 vdd3p3.n6285 vdd3p3.n6284 2.241
R8711 vdd3p3.n6200 vdd3p3.n6199 2.241
R8712 vdd3p3.n6113 vdd3p3.n6112 2.241
R8713 vdd3p3.n6043 vdd3p3.n6042 2.241
R8714 vdd3p3.n5973 vdd3p3.n5972 2.241
R8715 vdd3p3.n5891 vdd3p3.n5890 2.241
R8716 vdd3p3.n5803 vdd3p3.n5802 2.241
R8717 vdd3p3.n5131 vdd3p3.n4570 2.239
R8718 vdd3p3.n5131 vdd3p3.n5123 2.239
R8719 vdd3p3.n7964 vdd3p3.n7963 2.234
R8720 vdd3p3.n8081 vdd3p3.n8080 2.234
R8721 vdd3p3.n8186 vdd3p3.n8185 2.234
R8722 vdd3p3.n8291 vdd3p3.n8290 2.234
R8723 vdd3p3.n3592 vdd3p3.n3591 2.223
R8724 vdd3p3.n3686 vdd3p3.n3685 2.223
R8725 vdd3p3.n3756 vdd3p3.n3755 2.223
R8726 vdd3p3.n4821 vdd3p3.n4820 2.223
R8727 vdd3p3.n4752 vdd3p3.n4751 2.223
R8728 vdd3p3.n7867 vdd3p3.n7866 2.217
R8729 vdd3p3.n7848 vdd3p3.n7841 2.217
R8730 vdd3p3.n7725 vdd3p3.n7724 2.217
R8731 vdd3p3.n7709 vdd3p3.n7704 2.217
R8732 vdd3p3.n7593 vdd3p3.n7592 2.217
R8733 vdd3p3.n7574 vdd3p3.n7567 2.217
R8734 vdd3p3.n904 vdd3p3.n903 2.196
R8735 vdd3p3.n2595 vdd3p3.n2594 2.196
R8736 vdd3p3.n8711 vdd3p3.n8710 2.183
R8737 vdd3p3.n7972 vdd3p3.n7968 2.167
R8738 vdd3p3.n8087 vdd3p3.n8084 2.167
R8739 vdd3p3.n8192 vdd3p3.n8189 2.167
R8740 vdd3p3.n8297 vdd3p3.n8294 2.167
R8741 vdd3p3.n7376 vdd3p3.n7373 2.155
R8742 vdd3p3.n7370 vdd3p3.n7369 2.155
R8743 vdd3p3.n7307 vdd3p3.n7304 2.155
R8744 vdd3p3.n7301 vdd3p3.n7300 2.155
R8745 vdd3p3.n7238 vdd3p3.n7235 2.155
R8746 vdd3p3.n7232 vdd3p3.n7231 2.155
R8747 vdd3p3.n7153 vdd3p3.n7149 2.155
R8748 vdd3p3.n7145 vdd3p3.n7144 2.155
R8749 vdd3p3.n7066 vdd3p3.n7062 2.155
R8750 vdd3p3.n7058 vdd3p3.n7057 2.155
R8751 vdd3p3.t153 vdd3p3.n4006 2.116
R8752 vdd3p3.n4124 vdd3p3.t39 2.116
R8753 vdd3p3.n3512 vdd3p3.n3470 2.103
R8754 vdd3p3.n6598 vdd3p3.t95 2.102
R8755 vdd3p3.n6353 vdd3p3.n6352 2.097
R8756 vdd3p3.n6274 vdd3p3.n6273 2.097
R8757 vdd3p3.n6187 vdd3p3.n6186 2.097
R8758 vdd3p3.n6103 vdd3p3.n6102 2.097
R8759 vdd3p3.n6033 vdd3p3.n6032 2.097
R8760 vdd3p3.n5963 vdd3p3.n5962 2.097
R8761 vdd3p3.n5878 vdd3p3.n5877 2.097
R8762 vdd3p3.n5790 vdd3p3.n5789 2.097
R8763 vdd3p3.n5265 vdd3p3.n5261 2.076
R8764 vdd3p3.n45 vdd3p3.n41 2.07
R8765 vdd3p3.n1736 vdd3p3.n1732 2.07
R8766 vdd3p3.n7000 vdd3p3.n6999 2.031
R8767 vdd3p3.n6925 vdd3p3.n6924 2.031
R8768 vdd3p3.n6912 vdd3p3.n6911 2.031
R8769 vdd3p3.n6837 vdd3p3.n6836 2.031
R8770 vdd3p3.n6824 vdd3p3.n6823 2.031
R8771 vdd3p3.n6749 vdd3p3.n6748 2.031
R8772 vdd3p3.n6736 vdd3p3.n6735 2.031
R8773 vdd3p3.n5404 vdd3p3.n5403 2.031
R8774 vdd3p3.n5417 vdd3p3.n5416 2.031
R8775 vdd3p3.n5492 vdd3p3.n5491 2.031
R8776 vdd3p3.n5505 vdd3p3.n5504 2.031
R8777 vdd3p3.n5580 vdd3p3.n5579 2.031
R8778 vdd3p3.n5593 vdd3p3.n5592 2.031
R8779 vdd3p3.n5668 vdd3p3.n5667 2.031
R8780 vdd3p3.n5681 vdd3p3.n5680 2.031
R8781 vdd3p3.n3144 vdd3p3.n3143 2.003
R8782 vdd3p3.n3142 vdd3p3.n2607 2.003
R8783 vdd3p3.n3354 vdd3p3.n3353 2.003
R8784 vdd3p3.n2298 vdd3p3.n2297 2.003
R8785 vdd3p3.n2296 vdd3p3.n1761 2.003
R8786 vdd3p3.n2508 vdd3p3.n2507 2.003
R8787 vdd3p3.n1453 vdd3p3.n1452 2.003
R8788 vdd3p3.n1451 vdd3p3.n916 2.003
R8789 vdd3p3.n1663 vdd3p3.n1662 2.003
R8790 vdd3p3.n607 vdd3p3.n606 2.003
R8791 vdd3p3.n605 vdd3p3.n70 2.003
R8792 vdd3p3.n817 vdd3p3.n816 2.003
R8793 vdd3p3.n3455 vdd3p3.n3454 1.998
R8794 vdd3p3.n3960 vdd3p3.n3959 1.983
R8795 vdd3p3.n2921 vdd3p3.n2817 1.977
R8796 vdd3p3.n2075 vdd3p3.n1971 1.977
R8797 vdd3p3.n1230 vdd3p3.n1126 1.977
R8798 vdd3p3.n384 vdd3p3.n280 1.977
R8799 vdd3p3.n7972 vdd3p3.n7971 1.964
R8800 vdd3p3.n8087 vdd3p3.n8086 1.964
R8801 vdd3p3.n8192 vdd3p3.n8191 1.964
R8802 vdd3p3.n8297 vdd3p3.n8296 1.964
R8803 vdd3p3.n7856 vdd3p3.n7852 1.964
R8804 vdd3p3.n7856 vdd3p3.n7855 1.964
R8805 vdd3p3.n7715 vdd3p3.n7712 1.964
R8806 vdd3p3.n7715 vdd3p3.n7714 1.964
R8807 vdd3p3.n7582 vdd3p3.n7578 1.964
R8808 vdd3p3.n7582 vdd3p3.n7581 1.964
R8809 vdd3p3.n3182 vdd3p3.n3180 1.963
R8810 vdd3p3.n3029 vdd3p3.n3020 1.963
R8811 vdd3p3.n3174 vdd3p3.n3031 1.963
R8812 vdd3p3.n3173 vdd3p3.n3171 1.963
R8813 vdd3p3.n3170 vdd3p3.n3168 1.963
R8814 vdd3p3.n3166 vdd3p3.n3164 1.963
R8815 vdd3p3.n2336 vdd3p3.n2334 1.963
R8816 vdd3p3.n2183 vdd3p3.n2174 1.963
R8817 vdd3p3.n2328 vdd3p3.n2185 1.963
R8818 vdd3p3.n2327 vdd3p3.n2325 1.963
R8819 vdd3p3.n2324 vdd3p3.n2322 1.963
R8820 vdd3p3.n2320 vdd3p3.n2318 1.963
R8821 vdd3p3.n1491 vdd3p3.n1489 1.963
R8822 vdd3p3.n1338 vdd3p3.n1329 1.963
R8823 vdd3p3.n1483 vdd3p3.n1340 1.963
R8824 vdd3p3.n1482 vdd3p3.n1480 1.963
R8825 vdd3p3.n1479 vdd3p3.n1477 1.963
R8826 vdd3p3.n1475 vdd3p3.n1473 1.963
R8827 vdd3p3.n645 vdd3p3.n643 1.963
R8828 vdd3p3.n492 vdd3p3.n483 1.963
R8829 vdd3p3.n637 vdd3p3.n494 1.963
R8830 vdd3p3.n636 vdd3p3.n634 1.963
R8831 vdd3p3.n633 vdd3p3.n631 1.963
R8832 vdd3p3.n629 vdd3p3.n627 1.963
R8833 vdd3p3.n6369 vdd3p3.n6368 1.952
R8834 vdd3p3.n6290 vdd3p3.n6289 1.952
R8835 vdd3p3.n6205 vdd3p3.n6204 1.952
R8836 vdd3p3.n6117 vdd3p3.n6116 1.952
R8837 vdd3p3.n6047 vdd3p3.n6046 1.952
R8838 vdd3p3.n5977 vdd3p3.n5976 1.952
R8839 vdd3p3.n5896 vdd3p3.n5895 1.952
R8840 vdd3p3.n5808 vdd3p3.n5807 1.952
R8841 vdd3p3.n3315 vdd3p3.n3314 1.945
R8842 vdd3p3.n2469 vdd3p3.n2468 1.945
R8843 vdd3p3.n1624 vdd3p3.n1623 1.945
R8844 vdd3p3.n778 vdd3p3.n777 1.945
R8845 vdd3p3.n5343 vdd3p3.n5342 1.899
R8846 vdd3p3.n7947 vdd3p3.n7945 1.896
R8847 vdd3p3.n7964 vdd3p3.n7961 1.896
R8848 vdd3p3.n8081 vdd3p3.n8078 1.896
R8849 vdd3p3.n8186 vdd3p3.n8183 1.896
R8850 vdd3p3.n8291 vdd3p3.n8288 1.896
R8851 vdd3p3.n3191 vdd3p3.n2753 1.887
R8852 vdd3p3.n2345 vdd3p3.n1907 1.887
R8853 vdd3p3.n1500 vdd3p3.n1062 1.887
R8854 vdd3p3.n654 vdd3p3.n216 1.887
R8855 vdd3p3.n7366 vdd3p3.n7365 1.886
R8856 vdd3p3.n7311 vdd3p3.n7310 1.886
R8857 vdd3p3.n7297 vdd3p3.n7296 1.886
R8858 vdd3p3.n7242 vdd3p3.n7241 1.886
R8859 vdd3p3.n7227 vdd3p3.n7226 1.886
R8860 vdd3p3.n7158 vdd3p3.n7157 1.886
R8861 vdd3p3.n7140 vdd3p3.n7139 1.886
R8862 vdd3p3.n7071 vdd3p3.n7070 1.886
R8863 vdd3p3.n7053 vdd3p3.n7052 1.886
R8864 vdd3p3.n4221 vdd3p3.n4217 1.882
R8865 vdd3p3.n5073 vdd3p3.n5069 1.882
R8866 vdd3p3.n3504 vdd3p3.n3503 1.882
R8867 vdd3p3.n4986 vdd3p3.n4985 1.882
R8868 vdd3p3.n7386 vdd3p3.n7385 1.882
R8869 vdd3p3.n8599 vdd3p3.n8598 1.878
R8870 vdd3p3.n8463 vdd3p3.n8459 1.852
R8871 vdd3p3.n7948 vdd3p3.n7947 1.828
R8872 vdd3p3.n4380 vdd3p3.n4379 1.813
R8873 vdd3p3.n4684 vdd3p3.n4683 1.813
R8874 vdd3p3.n6349 vdd3p3.n6348 1.807
R8875 vdd3p3.n6270 vdd3p3.n6269 1.807
R8876 vdd3p3.n6182 vdd3p3.n6181 1.807
R8877 vdd3p3.n6099 vdd3p3.n6098 1.807
R8878 vdd3p3.n6029 vdd3p3.n6028 1.807
R8879 vdd3p3.n5959 vdd3p3.n5958 1.807
R8880 vdd3p3.n5873 vdd3p3.n5872 1.807
R8881 vdd3p3.n5785 vdd3p3.n5784 1.807
R8882 vdd3p3.n3145 vdd3p3.n3144 1.78
R8883 vdd3p3.n3355 vdd3p3.n3354 1.78
R8884 vdd3p3.n2299 vdd3p3.n2298 1.78
R8885 vdd3p3.n2509 vdd3p3.n2508 1.78
R8886 vdd3p3.n1454 vdd3p3.n1453 1.78
R8887 vdd3p3.n1664 vdd3p3.n1663 1.78
R8888 vdd3p3.n608 vdd3p3.n607 1.78
R8889 vdd3p3.n818 vdd3p3.n817 1.78
R8890 vdd3p3.n6995 vdd3p3.n6994 1.76
R8891 vdd3p3.n6930 vdd3p3.n6929 1.76
R8892 vdd3p3.n6907 vdd3p3.n6906 1.76
R8893 vdd3p3.n6842 vdd3p3.n6841 1.76
R8894 vdd3p3.n6819 vdd3p3.n6818 1.76
R8895 vdd3p3.n6754 vdd3p3.n6753 1.76
R8896 vdd3p3.n6731 vdd3p3.n6730 1.76
R8897 vdd3p3.n5399 vdd3p3.n5398 1.76
R8898 vdd3p3.n5422 vdd3p3.n5421 1.76
R8899 vdd3p3.n5487 vdd3p3.n5486 1.76
R8900 vdd3p3.n5510 vdd3p3.n5509 1.76
R8901 vdd3p3.n5575 vdd3p3.n5574 1.76
R8902 vdd3p3.n5598 vdd3p3.n5597 1.76
R8903 vdd3p3.n5663 vdd3p3.n5662 1.76
R8904 vdd3p3.n5686 vdd3p3.n5685 1.76
R8905 vdd3p3.n2921 vdd3p3.n2920 1.745
R8906 vdd3p3.n2075 vdd3p3.n2074 1.745
R8907 vdd3p3.n1230 vdd3p3.n1229 1.745
R8908 vdd3p3.n384 vdd3p3.n383 1.745
R8909 vdd3p3.t51 vdd3p3.n4069 1.719
R8910 vdd3p3.n3335 vdd3p3.n2674 1.711
R8911 vdd3p3.n3334 vdd3p3.n2675 1.711
R8912 vdd3p3.n3331 vdd3p3.n3330 1.711
R8913 vdd3p3.n3326 vdd3p3.n2678 1.711
R8914 vdd3p3.n3325 vdd3p3.n2681 1.711
R8915 vdd3p3.n3321 vdd3p3.n3320 1.711
R8916 vdd3p3.n2489 vdd3p3.n1828 1.711
R8917 vdd3p3.n2488 vdd3p3.n1829 1.711
R8918 vdd3p3.n2485 vdd3p3.n2484 1.711
R8919 vdd3p3.n2480 vdd3p3.n1832 1.711
R8920 vdd3p3.n2479 vdd3p3.n1835 1.711
R8921 vdd3p3.n2475 vdd3p3.n2474 1.711
R8922 vdd3p3.n1644 vdd3p3.n983 1.711
R8923 vdd3p3.n1643 vdd3p3.n984 1.711
R8924 vdd3p3.n1640 vdd3p3.n1639 1.711
R8925 vdd3p3.n1635 vdd3p3.n987 1.711
R8926 vdd3p3.n1634 vdd3p3.n990 1.711
R8927 vdd3p3.n1630 vdd3p3.n1629 1.711
R8928 vdd3p3.n798 vdd3p3.n137 1.711
R8929 vdd3p3.n797 vdd3p3.n138 1.711
R8930 vdd3p3.n794 vdd3p3.n793 1.711
R8931 vdd3p3.n789 vdd3p3.n141 1.711
R8932 vdd3p3.n788 vdd3p3.n144 1.711
R8933 vdd3p3.n784 vdd3p3.n783 1.711
R8934 vdd3p3.n7867 vdd3p3.n7863 1.71
R8935 vdd3p3.n7848 vdd3p3.n7847 1.71
R8936 vdd3p3.n7725 vdd3p3.n7722 1.71
R8937 vdd3p3.n7709 vdd3p3.n7708 1.71
R8938 vdd3p3.n7593 vdd3p3.n7589 1.71
R8939 vdd3p3.n7574 vdd3p3.n7573 1.71
R8940 vdd3p3.n62 vdd3p3.n0 1.705
R8941 vdd3p3.n908 vdd3p3.n907 1.705
R8942 vdd3p3.n1753 vdd3p3.n1691 1.705
R8943 vdd3p3.n2599 vdd3p3.n2598 1.705
R8944 vdd3p3.n7980 vdd3p3.n7979 1.693
R8945 vdd3p3.n8095 vdd3p3.n8094 1.693
R8946 vdd3p3.n8200 vdd3p3.n8199 1.693
R8947 vdd3p3.n8309 vdd3p3.n8308 1.693
R8948 vdd3p3.t106 vdd3p3.t92 1.682
R8949 vdd3p3.n3352 vdd3p3.n2637 1.669
R8950 vdd3p3.n2506 vdd3p3.n1791 1.669
R8951 vdd3p3.n1661 vdd3p3.n946 1.669
R8952 vdd3p3.n815 vdd3p3.n100 1.669
R8953 vdd3p3.n6373 vdd3p3.n6372 1.663
R8954 vdd3p3.n6294 vdd3p3.n6293 1.663
R8955 vdd3p3.n6210 vdd3p3.n6209 1.663
R8956 vdd3p3.n6122 vdd3p3.n6121 1.663
R8957 vdd3p3.n6051 vdd3p3.n6050 1.663
R8958 vdd3p3.n5981 vdd3p3.n5980 1.663
R8959 vdd3p3.n5901 vdd3p3.n5900 1.663
R8960 vdd3p3.n5813 vdd3p3.n5812 1.663
R8961 vdd3p3.n3102 vdd3p3.n3100 1.661
R8962 vdd3p3.n3103 vdd3p3.n3086 1.661
R8963 vdd3p3.n3108 vdd3p3.n3106 1.661
R8964 vdd3p3.n3109 vdd3p3.n3084 1.661
R8965 vdd3p3.n3114 vdd3p3.n3112 1.661
R8966 vdd3p3.n3118 vdd3p3.n3117 1.661
R8967 vdd3p3.n2256 vdd3p3.n2254 1.661
R8968 vdd3p3.n2257 vdd3p3.n2240 1.661
R8969 vdd3p3.n2262 vdd3p3.n2260 1.661
R8970 vdd3p3.n2263 vdd3p3.n2238 1.661
R8971 vdd3p3.n2268 vdd3p3.n2266 1.661
R8972 vdd3p3.n2272 vdd3p3.n2271 1.661
R8973 vdd3p3.n1411 vdd3p3.n1409 1.661
R8974 vdd3p3.n1412 vdd3p3.n1395 1.661
R8975 vdd3p3.n1417 vdd3p3.n1415 1.661
R8976 vdd3p3.n1418 vdd3p3.n1393 1.661
R8977 vdd3p3.n1423 vdd3p3.n1421 1.661
R8978 vdd3p3.n1427 vdd3p3.n1426 1.661
R8979 vdd3p3.n565 vdd3p3.n563 1.661
R8980 vdd3p3.n566 vdd3p3.n549 1.661
R8981 vdd3p3.n571 vdd3p3.n569 1.661
R8982 vdd3p3.n572 vdd3p3.n547 1.661
R8983 vdd3p3.n577 vdd3p3.n575 1.661
R8984 vdd3p3.n581 vdd3p3.n580 1.661
R8985 vdd3p3.n3669 vdd3p3.n3668 1.642
R8986 vdd3p3.n3739 vdd3p3.n3738 1.642
R8987 vdd3p3.n3575 vdd3p3.n3574 1.642
R8988 vdd3p3.n4804 vdd3p3.n4803 1.642
R8989 vdd3p3.n4735 vdd3p3.n4734 1.642
R8990 vdd3p3.n7392 vdd3p3.n7391 1.631
R8991 vdd3p3.n7956 vdd3p3.n7955 1.625
R8992 vdd3p3.n8073 vdd3p3.n8072 1.625
R8993 vdd3p3.n8178 vdd3p3.n8177 1.625
R8994 vdd3p3.n8283 vdd3p3.n8282 1.625
R8995 vdd3p3.n8433 vdd3p3.n8432 1.625
R8996 vdd3p3.n3397 vdd3p3.n3396 1.618
R8997 vdd3p3.n7362 vdd3p3.n7361 1.616
R8998 vdd3p3.n7315 vdd3p3.n7314 1.616
R8999 vdd3p3.n7293 vdd3p3.n7292 1.616
R9000 vdd3p3.n7246 vdd3p3.n7245 1.616
R9001 vdd3p3.n7222 vdd3p3.n7221 1.616
R9002 vdd3p3.n7163 vdd3p3.n7162 1.616
R9003 vdd3p3.n7135 vdd3p3.n7134 1.616
R9004 vdd3p3.n7076 vdd3p3.n7075 1.616
R9005 vdd3p3.n7048 vdd3p3.n7047 1.616
R9006 vdd3p3.n5338 vdd3p3.n5335 1.614
R9007 vdd3p3.n5335 vdd3p3.n5332 1.614
R9008 vdd3p3.n5332 vdd3p3.n5329 1.614
R9009 vdd3p3.n5329 vdd3p3.n5326 1.614
R9010 vdd3p3.n5326 vdd3p3.n5323 1.614
R9011 vdd3p3.n5284 vdd3p3.n5281 1.614
R9012 vdd3p3.n5287 vdd3p3.n5284 1.614
R9013 vdd3p3.n5290 vdd3p3.n5287 1.614
R9014 vdd3p3.n5293 vdd3p3.n5290 1.614
R9015 vdd3p3.n5296 vdd3p3.n5293 1.614
R9016 vdd3p3.n5300 vdd3p3.n5296 1.614
R9017 vdd3p3.n5320 vdd3p3.n5317 1.614
R9018 vdd3p3.n5317 vdd3p3.n5314 1.614
R9019 vdd3p3.n5314 vdd3p3.n5311 1.614
R9020 vdd3p3.n5311 vdd3p3.n5308 1.614
R9021 vdd3p3.n5308 vdd3p3.n5305 1.614
R9022 vdd3p3.n5305 vdd3p3.n5302 1.614
R9023 vdd3p3.n5167 vdd3p3.n5164 1.614
R9024 vdd3p3.n5170 vdd3p3.n5167 1.614
R9025 vdd3p3.n5173 vdd3p3.n5170 1.614
R9026 vdd3p3.n5176 vdd3p3.n5173 1.614
R9027 vdd3p3.n5179 vdd3p3.n5176 1.614
R9028 vdd3p3.n3376 vdd3p3.n3375 1.613
R9029 vdd3p3.n2530 vdd3p3.n2529 1.613
R9030 vdd3p3.n1685 vdd3p3.n1684 1.613
R9031 vdd3p3.n839 vdd3p3.n838 1.613
R9032 vdd3p3.n8416 vdd3p3.t144 1.587
R9033 vdd3p3.n6684 vdd3p3.n6683 1.583
R9034 vdd3p3.n6596 vdd3p3.n6595 1.583
R9035 vdd3p3.n6508 vdd3p3.n6507 1.583
R9036 vdd3p3.n6420 vdd3p3.n6419 1.583
R9037 vdd3p3.n3909 vdd3p3.n3908 1.583
R9038 vdd3p3.n7015 vdd3p3.n7011 1.557
R9039 vdd3p3.n8465 vdd3p3.n8464 1.55
R9040 vdd3p3.n6344 vdd3p3.n6343 1.518
R9041 vdd3p3.n6265 vdd3p3.n6264 1.518
R9042 vdd3p3.n6177 vdd3p3.n6176 1.518
R9043 vdd3p3.n6095 vdd3p3.n6094 1.518
R9044 vdd3p3.n6025 vdd3p3.n6024 1.518
R9045 vdd3p3.n5955 vdd3p3.n5954 1.518
R9046 vdd3p3.n5868 vdd3p3.n5867 1.518
R9047 vdd3p3.n5780 vdd3p3.n5779 1.518
R9048 vdd3p3.n8737 vdd3p3.n8736 1.512
R9049 vdd3p3.n8498 vdd3p3.n8495 1.505
R9050 vdd3p3.n8574 vdd3p3.n8573 1.505
R9051 vdd3p3.n8842 vdd3p3.n8839 1.505
R9052 vdd3p3.n8784 vdd3p3.n8781 1.505
R9053 vdd3p3.n3814 vdd3p3.n3813 1.505
R9054 vdd3p3.n3840 vdd3p3.n3838 1.505
R9055 vdd3p3.n3873 vdd3p3.n3872 1.5
R9056 vdd3p3.n8571 vdd3p3.n8570 1.5
R9057 vdd3p3.n6990 vdd3p3.n6989 1.489
R9058 vdd3p3.n6935 vdd3p3.n6934 1.489
R9059 vdd3p3.n6902 vdd3p3.n6901 1.489
R9060 vdd3p3.n6847 vdd3p3.n6846 1.489
R9061 vdd3p3.n6814 vdd3p3.n6813 1.489
R9062 vdd3p3.n6759 vdd3p3.n6758 1.489
R9063 vdd3p3.n6726 vdd3p3.n6725 1.489
R9064 vdd3p3.n5394 vdd3p3.n5393 1.489
R9065 vdd3p3.n5427 vdd3p3.n5426 1.489
R9066 vdd3p3.n5482 vdd3p3.n5481 1.489
R9067 vdd3p3.n5515 vdd3p3.n5514 1.489
R9068 vdd3p3.n5570 vdd3p3.n5569 1.489
R9069 vdd3p3.n5603 vdd3p3.n5602 1.489
R9070 vdd3p3.n5658 vdd3p3.n5657 1.489
R9071 vdd3p3.n5691 vdd3p3.n5690 1.489
R9072 vdd3p3.n3579 vdd3p3.n3578 1.486
R9073 vdd3p3.n3673 vdd3p3.n3672 1.486
R9074 vdd3p3.n3743 vdd3p3.n3742 1.486
R9075 vdd3p3.n4808 vdd3p3.n4807 1.486
R9076 vdd3p3.n4739 vdd3p3.n4738 1.486
R9077 vdd3p3.n5106 vdd3p3.n5105 1.484
R9078 vdd3p3.n4493 vdd3p3.n4492 1.484
R9079 vdd3p3.n4403 vdd3p3.n4402 1.484
R9080 vdd3p3.n5111 vdd3p3.n4690 1.484
R9081 vdd3p3.n4463 vdd3p3.n4462 1.484
R9082 vdd3p3.n4369 vdd3p3.n4368 1.484
R9083 vdd3p3.n4246 vdd3p3.n4245 1.484
R9084 vdd3p3.n4433 vdd3p3.n4432 1.484
R9085 vdd3p3.n4523 vdd3p3.n4522 1.484
R9086 vdd3p3.n3446 vdd3p3.n3445 1.472
R9087 vdd3p3.n4565 vdd3p3.n4564 1.472
R9088 vdd3p3.n4384 vdd3p3.n4383 1.464
R9089 vdd3p3.n4417 vdd3p3.n4416 1.464
R9090 vdd3p3.n4507 vdd3p3.n4506 1.464
R9091 vdd3p3.n4447 vdd3p3.n4446 1.464
R9092 vdd3p3.n4477 vdd3p3.n4476 1.464
R9093 vdd3p3.n2881 vdd3p3.n2880 1.457
R9094 vdd3p3.n2862 vdd3p3.n2853 1.457
R9095 vdd3p3.n2857 vdd3p3.n2853 1.457
R9096 vdd3p3.n2035 vdd3p3.n2034 1.457
R9097 vdd3p3.n2016 vdd3p3.n2007 1.457
R9098 vdd3p3.n2011 vdd3p3.n2007 1.457
R9099 vdd3p3.n1190 vdd3p3.n1189 1.457
R9100 vdd3p3.n1171 vdd3p3.n1162 1.457
R9101 vdd3p3.n1166 vdd3p3.n1162 1.457
R9102 vdd3p3.n344 vdd3p3.n343 1.457
R9103 vdd3p3.n325 vdd3p3.n316 1.457
R9104 vdd3p3.n320 vdd3p3.n316 1.457
R9105 vdd3p3.n7875 vdd3p3.n7874 1.457
R9106 vdd3p3.n7837 vdd3p3.n7836 1.457
R9107 vdd3p3.n7733 vdd3p3.n7732 1.457
R9108 vdd3p3.n7701 vdd3p3.n7700 1.457
R9109 vdd3p3.n7601 vdd3p3.n7600 1.457
R9110 vdd3p3.n7563 vdd3p3.n7562 1.457
R9111 vdd3p3.n5274 vdd3p3.n5273 1.454
R9112 vdd3p3.n7988 vdd3p3.n7987 1.422
R9113 vdd3p3.n8101 vdd3p3.n8100 1.422
R9114 vdd3p3.n8206 vdd3p3.n8205 1.422
R9115 vdd3p3.n8319 vdd3p3.n8318 1.422
R9116 vdd3p3.n6676 vdd3p3.n6675 1.412
R9117 vdd3p3.n6588 vdd3p3.n6587 1.412
R9118 vdd3p3.n6500 vdd3p3.n6499 1.412
R9119 vdd3p3.n6414 vdd3p3.n6413 1.412
R9120 vdd3p3.n8734 vdd3p3.n8713 1.412
R9121 vdd3p3.n8692 vdd3p3.n8691 1.391
R9122 vdd3p3.n7454 vdd3p3.n7453 1.38
R9123 vdd3p3.n7396 vdd3p3.n7395 1.38
R9124 vdd3p3.n6378 vdd3p3.n6377 1.374
R9125 vdd3p3.n6299 vdd3p3.n6298 1.374
R9126 vdd3p3.n6215 vdd3p3.n6214 1.374
R9127 vdd3p3.n6127 vdd3p3.n6126 1.374
R9128 vdd3p3.n6055 vdd3p3.n6054 1.374
R9129 vdd3p3.n5985 vdd3p3.n5984 1.374
R9130 vdd3p3.n5906 vdd3p3.n5905 1.374
R9131 vdd3p3.n5818 vdd3p3.n5817 1.374
R9132 vdd3p3.n8067 vdd3p3.n8066 1.354
R9133 vdd3p3.n8172 vdd3p3.n8171 1.354
R9134 vdd3p3.n8277 vdd3p3.n8276 1.354
R9135 vdd3p3.n8427 vdd3p3.n8426 1.354
R9136 vdd3p3.n3341 vdd3p3.n2669 1.35
R9137 vdd3p3.n2495 vdd3p3.n1823 1.35
R9138 vdd3p3.n1650 vdd3p3.n978 1.35
R9139 vdd3p3.n804 vdd3p3.n132 1.35
R9140 vdd3p3.n7358 vdd3p3.n7357 1.347
R9141 vdd3p3.n7319 vdd3p3.n7318 1.347
R9142 vdd3p3.n7289 vdd3p3.n7288 1.347
R9143 vdd3p3.n7250 vdd3p3.n7249 1.347
R9144 vdd3p3.n7217 vdd3p3.n7216 1.347
R9145 vdd3p3.n7168 vdd3p3.n7167 1.347
R9146 vdd3p3.n7130 vdd3p3.n7129 1.347
R9147 vdd3p3.n7081 vdd3p3.n7080 1.347
R9148 vdd3p3.n7043 vdd3p3.n7042 1.347
R9149 vdd3p3.n4541 vdd3p3.n3438 1.344
R9150 vdd3p3.n4541 vdd3p3.n3450 1.342
R9151 vdd3p3.n3377 vdd3p3.n2603 1.335
R9152 vdd3p3.n2531 vdd3p3.n1757 1.335
R9153 vdd3p3.n1686 vdd3p3.n912 1.335
R9154 vdd3p3.n840 vdd3p3.n66 1.335
R9155 vdd3p3.n6684 vdd3p3.n6680 1.327
R9156 vdd3p3.n6596 vdd3p3.n6592 1.327
R9157 vdd3p3.n6508 vdd3p3.n6504 1.327
R9158 vdd3p3.n6420 vdd3p3.n6417 1.327
R9159 vdd3p3.n3184 vdd3p3.n3183 1.321
R9160 vdd3p3.n3094 vdd3p3.n3088 1.321
R9161 vdd3p3.n2338 vdd3p3.n2337 1.321
R9162 vdd3p3.n2248 vdd3p3.n2242 1.321
R9163 vdd3p3.n1493 vdd3p3.n1492 1.321
R9164 vdd3p3.n1403 vdd3p3.n1397 1.321
R9165 vdd3p3.n647 vdd3p3.n646 1.321
R9166 vdd3p3.n557 vdd3p3.n551 1.321
R9167 vdd3p3.n5343 vdd3p3.n5338 1.282
R9168 vdd3p3.n3827 vdd3p3.n3826 1.265
R9169 vdd3p3.n2984 vdd3p3.n2983 1.252
R9170 vdd3p3.n2138 vdd3p3.n2137 1.252
R9171 vdd3p3.n1293 vdd3p3.n1292 1.252
R9172 vdd3p3.n447 vdd3p3.n446 1.252
R9173 vdd3p3.n3185 vdd3p3.n3184 1.246
R9174 vdd3p3.n3091 vdd3p3.n3088 1.246
R9175 vdd3p3.n2339 vdd3p3.n2338 1.246
R9176 vdd3p3.n2245 vdd3p3.n2242 1.246
R9177 vdd3p3.n1494 vdd3p3.n1493 1.246
R9178 vdd3p3.n1400 vdd3p3.n1397 1.246
R9179 vdd3p3.n648 vdd3p3.n647 1.246
R9180 vdd3p3.n554 vdd3p3.n551 1.246
R9181 vdd3p3.n6671 vdd3p3.n6670 1.241
R9182 vdd3p3.n6584 vdd3p3.n6583 1.241
R9183 vdd3p3.n6495 vdd3p3.n6494 1.241
R9184 vdd3p3.n6410 vdd3p3.n6409 1.241
R9185 vdd3p3.n8736 vdd3p3.n8734 1.235
R9186 vdd3p3.n6340 vdd3p3.n6339 1.229
R9187 vdd3p3.n6260 vdd3p3.n6259 1.229
R9188 vdd3p3.n6172 vdd3p3.n6171 1.229
R9189 vdd3p3.n6091 vdd3p3.n6090 1.229
R9190 vdd3p3.n6021 vdd3p3.n6020 1.229
R9191 vdd3p3.n5951 vdd3p3.n5950 1.229
R9192 vdd3p3.n5863 vdd3p3.n5862 1.229
R9193 vdd3p3.n5775 vdd3p3.n5774 1.229
R9194 vdd3p3.n2608 vdd3p3.n2604 1.224
R9195 vdd3p3.n3377 vdd3p3.n2604 1.224
R9196 vdd3p3.n3069 vdd3p3.n2603 1.224
R9197 vdd3p3.n2633 vdd3p3.n2621 1.224
R9198 vdd3p3.n2635 vdd3p3.n2634 1.224
R9199 vdd3p3.n1762 vdd3p3.n1758 1.224
R9200 vdd3p3.n2531 vdd3p3.n1758 1.224
R9201 vdd3p3.n2223 vdd3p3.n1757 1.224
R9202 vdd3p3.n1787 vdd3p3.n1775 1.224
R9203 vdd3p3.n1789 vdd3p3.n1788 1.224
R9204 vdd3p3.n917 vdd3p3.n913 1.224
R9205 vdd3p3.n1686 vdd3p3.n913 1.224
R9206 vdd3p3.n1378 vdd3p3.n912 1.224
R9207 vdd3p3.n942 vdd3p3.n930 1.224
R9208 vdd3p3.n944 vdd3p3.n943 1.224
R9209 vdd3p3.n71 vdd3p3.n67 1.224
R9210 vdd3p3.n840 vdd3p3.n67 1.224
R9211 vdd3p3.n532 vdd3p3.n66 1.224
R9212 vdd3p3.n96 vdd3p3.n84 1.224
R9213 vdd3p3.n98 vdd3p3.n97 1.224
R9214 vdd3p3.n6985 vdd3p3.n6984 1.219
R9215 vdd3p3.n6940 vdd3p3.n6939 1.219
R9216 vdd3p3.n6897 vdd3p3.n6896 1.219
R9217 vdd3p3.n6852 vdd3p3.n6851 1.219
R9218 vdd3p3.n6809 vdd3p3.n6808 1.219
R9219 vdd3p3.n6764 vdd3p3.n6763 1.219
R9220 vdd3p3.n6721 vdd3p3.n6720 1.219
R9221 vdd3p3.n5389 vdd3p3.n5388 1.219
R9222 vdd3p3.n5432 vdd3p3.n5431 1.219
R9223 vdd3p3.n5477 vdd3p3.n5476 1.219
R9224 vdd3p3.n5520 vdd3p3.n5519 1.219
R9225 vdd3p3.n5565 vdd3p3.n5564 1.219
R9226 vdd3p3.n5608 vdd3p3.n5607 1.219
R9227 vdd3p3.n5653 vdd3p3.n5652 1.219
R9228 vdd3p3.n5696 vdd3p3.n5695 1.219
R9229 vdd3p3.n7883 vdd3p3.n7882 1.203
R9230 vdd3p3.n7829 vdd3p3.n7828 1.203
R9231 vdd3p3.n7741 vdd3p3.n7740 1.203
R9232 vdd3p3.n7695 vdd3p3.n7694 1.203
R9233 vdd3p3.n7609 vdd3p3.n7608 1.203
R9234 vdd3p3.n7555 vdd3p3.n7554 1.203
R9235 vdd3p3.n874 vdd3p3.n845 1.195
R9236 vdd3p3.n2565 vdd3p3.n2536 1.195
R9237 vdd3p3.n61 vdd3p3.n60 1.19
R9238 vdd3p3.n1752 vdd3p3.n1751 1.19
R9239 vdd3p3.n6689 vdd3p3.n6688 1.155
R9240 vdd3p3.n6601 vdd3p3.n6600 1.155
R9241 vdd3p3.n6513 vdd3p3.n6512 1.155
R9242 vdd3p3.n6425 vdd3p3.n6424 1.155
R9243 vdd3p3.n7994 vdd3p3.n7993 1.151
R9244 vdd3p3.n8107 vdd3p3.n8106 1.151
R9245 vdd3p3.n8212 vdd3p3.n8211 1.151
R9246 vdd3p3.n8329 vdd3p3.n8328 1.151
R9247 vdd3p3.n4171 vdd3p3.n4170 1.142
R9248 vdd3p3.n8657 vdd3p3.n8641 1.142
R9249 vdd3p3.n5148 vdd3p3.n3403 1.137
R9250 vdd3p3.n5148 vdd3p3.n5146 1.137
R9251 vdd3p3.n5148 vdd3p3.n5147 1.137
R9252 vdd3p3.n5148 vdd3p3.n3405 1.137
R9253 vdd3p3.n4172 vdd3p3.n3792 1.135
R9254 vdd3p3.n4210 vdd3p3.n4206 1.129
R9255 vdd3p3.n5062 vdd3p3.n5058 1.129
R9256 vdd3p3.n3488 vdd3p3.n3487 1.129
R9257 vdd3p3.n4970 vdd3p3.n4969 1.129
R9258 vdd3p3.n8516 vdd3p3.n8512 1.129
R9259 vdd3p3.n8860 vdd3p3.n8856 1.129
R9260 vdd3p3.n8771 vdd3p3.n8767 1.129
R9261 vdd3p3.n7447 vdd3p3.n7446 1.129
R9262 vdd3p3.n7401 vdd3p3.n7400 1.129
R9263 vdd3p3.n3867 vdd3p3.n3866 1.129
R9264 vdd3p3.n3857 vdd3p3.n3856 1.129
R9265 vdd3p3.n8657 vdd3p3.n8656 1.127
R9266 vdd3p3.n2880 vdd3p3.n2841 1.114
R9267 vdd3p3.n2877 vdd3p3.n2876 1.114
R9268 vdd3p3.n2872 vdd3p3.n2843 1.114
R9269 vdd3p3.n2871 vdd3p3.n2847 1.114
R9270 vdd3p3.n2867 vdd3p3.n2866 1.114
R9271 vdd3p3.n2863 vdd3p3.n2850 1.114
R9272 vdd3p3.n2034 vdd3p3.n1995 1.114
R9273 vdd3p3.n2031 vdd3p3.n2030 1.114
R9274 vdd3p3.n2026 vdd3p3.n1997 1.114
R9275 vdd3p3.n2025 vdd3p3.n2001 1.114
R9276 vdd3p3.n2021 vdd3p3.n2020 1.114
R9277 vdd3p3.n2017 vdd3p3.n2004 1.114
R9278 vdd3p3.n1189 vdd3p3.n1150 1.114
R9279 vdd3p3.n1186 vdd3p3.n1185 1.114
R9280 vdd3p3.n1181 vdd3p3.n1152 1.114
R9281 vdd3p3.n1180 vdd3p3.n1156 1.114
R9282 vdd3p3.n1176 vdd3p3.n1175 1.114
R9283 vdd3p3.n1172 vdd3p3.n1159 1.114
R9284 vdd3p3.n343 vdd3p3.n304 1.114
R9285 vdd3p3.n340 vdd3p3.n339 1.114
R9286 vdd3p3.n335 vdd3p3.n306 1.114
R9287 vdd3p3.n334 vdd3p3.n310 1.114
R9288 vdd3p3.n330 vdd3p3.n329 1.114
R9289 vdd3p3.n326 vdd3p3.n313 1.114
R9290 vdd3p3.n8602 vdd3p3.n8601 1.109
R9291 vdd3p3.n8820 vdd3p3.n8819 1.109
R9292 vdd3p3.n8560 vdd3p3.n8557 1.109
R9293 vdd3p3.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPB 1.097
R9294 vdd3p3.n1736 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPB 1.097
R9295 vdd3p3.n8467 vdd3p3.n8466 1.095
R9296 vdd3p3.n6382 vdd3p3.n6381 1.084
R9297 vdd3p3.n6303 vdd3p3.n6302 1.084
R9298 vdd3p3.n6220 vdd3p3.n6219 1.084
R9299 vdd3p3.n6132 vdd3p3.n6131 1.084
R9300 vdd3p3.n6059 vdd3p3.n6058 1.084
R9301 vdd3p3.n5989 vdd3p3.n5988 1.084
R9302 vdd3p3.n5911 vdd3p3.n5910 1.084
R9303 vdd3p3.n5823 vdd3p3.n5822 1.084
R9304 vdd3p3.n8061 vdd3p3.n8060 1.083
R9305 vdd3p3.n8166 vdd3p3.n8165 1.083
R9306 vdd3p3.n8271 vdd3p3.n8270 1.083
R9307 vdd3p3.n8419 vdd3p3.n8418 1.083
R9308 vdd3p3.n7354 vdd3p3.n7353 1.077
R9309 vdd3p3.n7323 vdd3p3.n7322 1.077
R9310 vdd3p3.n7285 vdd3p3.n7284 1.077
R9311 vdd3p3.n7254 vdd3p3.n7253 1.077
R9312 vdd3p3.n7212 vdd3p3.n7211 1.077
R9313 vdd3p3.n7173 vdd3p3.n7172 1.077
R9314 vdd3p3.n7125 vdd3p3.n7124 1.077
R9315 vdd3p3.n7086 vdd3p3.n7085 1.077
R9316 vdd3p3.n7038 vdd3p3.n7037 1.077
R9317 vdd3p3.n5342 vdd3p3.n5341 1.07
R9318 vdd3p3.n6666 vdd3p3.n6665 1.07
R9319 vdd3p3.n6580 vdd3p3.n6579 1.07
R9320 vdd3p3.n6490 vdd3p3.n6489 1.07
R9321 vdd3p3.n6406 vdd3p3.n6405 1.07
R9322 vdd3p3.n8676 vdd3p3.n8675 1.042
R9323 vdd3p3.n8883 vdd3p3.n8882 1.027
R9324 vdd3p3.n8883 vdd3p3.n8636 1.026
R9325 vdd3p3.n5344 vdd3p3.n5179 1.021
R9326 vdd3p3.n4261 vdd3p3.n4260 0.993
R9327 vdd3p3.n4277 vdd3p3.n4276 0.993
R9328 vdd3p3.n4581 vdd3p3.n4580 0.993
R9329 vdd3p3.n4597 vdd3p3.n4596 0.993
R9330 vdd3p3.n3523 vdd3p3.n3522 0.993
R9331 vdd3p3.n3539 vdd3p3.n3538 0.993
R9332 vdd3p3.n3608 vdd3p3.n3607 0.993
R9333 vdd3p3.n3707 vdd3p3.n3706 0.993
R9334 vdd3p3.n3636 vdd3p3.n3635 0.993
R9335 vdd3p3.n3626 vdd3p3.n3625 0.993
R9336 vdd3p3.n4772 vdd3p3.n4771 0.993
R9337 vdd3p3.n4913 vdd3p3.n4912 0.993
R9338 vdd3p3.n6694 vdd3p3.n6693 0.984
R9339 vdd3p3.n6606 vdd3p3.n6605 0.984
R9340 vdd3p3.n6518 vdd3p3.n6517 0.984
R9341 vdd3p3.n6430 vdd3p3.n6429 0.984
R9342 vdd3p3.n7891 vdd3p3.n7890 0.95
R9343 vdd3p3.n7821 vdd3p3.n7820 0.95
R9344 vdd3p3.n7749 vdd3p3.n7748 0.95
R9345 vdd3p3.n7689 vdd3p3.n7688 0.95
R9346 vdd3p3.n7617 vdd3p3.n7616 0.95
R9347 vdd3p3.n7547 vdd3p3.n7546 0.95
R9348 vdd3p3.n6980 vdd3p3.n6979 0.948
R9349 vdd3p3.n6945 vdd3p3.n6944 0.948
R9350 vdd3p3.n6892 vdd3p3.n6891 0.948
R9351 vdd3p3.n6857 vdd3p3.n6856 0.948
R9352 vdd3p3.n6804 vdd3p3.n6803 0.948
R9353 vdd3p3.n6769 vdd3p3.n6768 0.948
R9354 vdd3p3.n5349 vdd3p3.n5348 0.948
R9355 vdd3p3.n5384 vdd3p3.n5383 0.948
R9356 vdd3p3.n5437 vdd3p3.n5436 0.948
R9357 vdd3p3.n5472 vdd3p3.n5471 0.948
R9358 vdd3p3.n5525 vdd3p3.n5524 0.948
R9359 vdd3p3.n5560 vdd3p3.n5559 0.948
R9360 vdd3p3.n5613 vdd3p3.n5612 0.948
R9361 vdd3p3.n5648 vdd3p3.n5647 0.948
R9362 vdd3p3.n5701 vdd3p3.n5700 0.948
R9363 vdd3p3.n6564 vdd3p3.t106 0.941
R9364 vdd3p3.n8734 vdd3p3.n8708 0.941
R9365 vdd3p3.n6335 vdd3p3.n6334 0.94
R9366 vdd3p3.n6255 vdd3p3.n6254 0.94
R9367 vdd3p3.n6167 vdd3p3.n6166 0.94
R9368 vdd3p3.n6087 vdd3p3.n6086 0.94
R9369 vdd3p3.n6017 vdd3p3.n6016 0.94
R9370 vdd3p3.n5946 vdd3p3.n5945 0.94
R9371 vdd3p3.n5858 vdd3p3.n5857 0.94
R9372 vdd3p3.n5770 vdd3p3.n5769 0.94
R9373 vdd3p3.n2674 vdd3p3.n2670 0.933
R9374 vdd3p3.n3335 vdd3p3.n3334 0.933
R9375 vdd3p3.n3331 vdd3p3.n2675 0.933
R9376 vdd3p3.n3330 vdd3p3.n2678 0.933
R9377 vdd3p3.n3326 vdd3p3.n3325 0.933
R9378 vdd3p3.n3321 vdd3p3.n2681 0.933
R9379 vdd3p3.n1828 vdd3p3.n1824 0.933
R9380 vdd3p3.n2489 vdd3p3.n2488 0.933
R9381 vdd3p3.n2485 vdd3p3.n1829 0.933
R9382 vdd3p3.n2484 vdd3p3.n1832 0.933
R9383 vdd3p3.n2480 vdd3p3.n2479 0.933
R9384 vdd3p3.n2475 vdd3p3.n1835 0.933
R9385 vdd3p3.n983 vdd3p3.n979 0.933
R9386 vdd3p3.n1644 vdd3p3.n1643 0.933
R9387 vdd3p3.n1640 vdd3p3.n984 0.933
R9388 vdd3p3.n1639 vdd3p3.n987 0.933
R9389 vdd3p3.n1635 vdd3p3.n1634 0.933
R9390 vdd3p3.n1630 vdd3p3.n990 0.933
R9391 vdd3p3.n137 vdd3p3.n133 0.933
R9392 vdd3p3.n798 vdd3p3.n797 0.933
R9393 vdd3p3.n794 vdd3p3.n138 0.933
R9394 vdd3p3.n793 vdd3p3.n141 0.933
R9395 vdd3p3.n789 vdd3p3.n788 0.933
R9396 vdd3p3.n784 vdd3p3.n144 0.933
R9397 vdd3p3.n3985 vdd3p3.n3984 0.931
R9398 vdd3p3.n4727 vdd3p3.n4724 0.926
R9399 vdd3p3.n3914 vdd3p3.n3909 0.925
R9400 vdd3p3.n3918 vdd3p3.n3915 0.925
R9401 vdd3p3.n3959 vdd3p3.n3956 0.925
R9402 vdd3p3.n3964 vdd3p3.n3961 0.925
R9403 vdd3p3.n3968 vdd3p3.n3965 0.925
R9404 vdd3p3.n3972 vdd3p3.n3969 0.925
R9405 vdd3p3.n3977 vdd3p3.n3974 0.925
R9406 vdd3p3.n3895 vdd3p3.n3894 0.925
R9407 vdd3p3.n3891 vdd3p3.n3890 0.925
R9408 vdd3p3.n3887 vdd3p3.n3886 0.925
R9409 vdd3p3.n3883 vdd3p3.n3882 0.925
R9410 vdd3p3.n3879 vdd3p3.n3878 0.925
R9411 vdd3p3.n4006 vdd3p3.n4003 0.925
R9412 vdd3p3.n4010 vdd3p3.n4007 0.925
R9413 vdd3p3.n4014 vdd3p3.n4011 0.925
R9414 vdd3p3.n4018 vdd3p3.n4015 0.925
R9415 vdd3p3.n4034 vdd3p3.n4033 0.925
R9416 vdd3p3.n4030 vdd3p3.n4029 0.925
R9417 vdd3p3.n4026 vdd3p3.n4025 0.925
R9418 vdd3p3.n4040 vdd3p3.n4037 0.925
R9419 vdd3p3.n4044 vdd3p3.n4041 0.925
R9420 vdd3p3.n4048 vdd3p3.n4045 0.925
R9421 vdd3p3.n4052 vdd3p3.n4049 0.925
R9422 vdd3p3.n4056 vdd3p3.n4053 0.925
R9423 vdd3p3.n4061 vdd3p3.n4058 0.925
R9424 vdd3p3.n4145 vdd3p3.n4144 0.925
R9425 vdd3p3.n4141 vdd3p3.n4140 0.925
R9426 vdd3p3.n4137 vdd3p3.n4136 0.925
R9427 vdd3p3.n4133 vdd3p3.n4132 0.925
R9428 vdd3p3.n4129 vdd3p3.n4128 0.925
R9429 vdd3p3.n4125 vdd3p3.n4124 0.925
R9430 vdd3p3.n4121 vdd3p3.n4120 0.925
R9431 vdd3p3.n4117 vdd3p3.n4116 0.925
R9432 vdd3p3.n4113 vdd3p3.n4112 0.925
R9433 vdd3p3.n4109 vdd3p3.n4108 0.925
R9434 vdd3p3.n4105 vdd3p3.n4104 0.925
R9435 vdd3p3.n4101 vdd3p3.n4100 0.925
R9436 vdd3p3.n4093 vdd3p3.n4092 0.925
R9437 vdd3p3.n4089 vdd3p3.n4088 0.925
R9438 vdd3p3.n4085 vdd3p3.n4084 0.925
R9439 vdd3p3.n4081 vdd3p3.n4080 0.925
R9440 vdd3p3.n4077 vdd3p3.n4076 0.925
R9441 vdd3p3.n4073 vdd3p3.n4072 0.925
R9442 vdd3p3.n4069 vdd3p3.n4068 0.925
R9443 vdd3p3.n8449 vdd3p3.n8448 0.925
R9444 vdd3p3.n3100 vdd3p3.n3098 0.906
R9445 vdd3p3.n3103 vdd3p3.n3102 0.906
R9446 vdd3p3.n3106 vdd3p3.n3086 0.906
R9447 vdd3p3.n3109 vdd3p3.n3108 0.906
R9448 vdd3p3.n3112 vdd3p3.n3084 0.906
R9449 vdd3p3.n3118 vdd3p3.n3114 0.906
R9450 vdd3p3.n2254 vdd3p3.n2252 0.906
R9451 vdd3p3.n2257 vdd3p3.n2256 0.906
R9452 vdd3p3.n2260 vdd3p3.n2240 0.906
R9453 vdd3p3.n2263 vdd3p3.n2262 0.906
R9454 vdd3p3.n2266 vdd3p3.n2238 0.906
R9455 vdd3p3.n2272 vdd3p3.n2268 0.906
R9456 vdd3p3.n1409 vdd3p3.n1407 0.906
R9457 vdd3p3.n1412 vdd3p3.n1411 0.906
R9458 vdd3p3.n1415 vdd3p3.n1395 0.906
R9459 vdd3p3.n1418 vdd3p3.n1417 0.906
R9460 vdd3p3.n1421 vdd3p3.n1393 0.906
R9461 vdd3p3.n1427 vdd3p3.n1423 0.906
R9462 vdd3p3.n563 vdd3p3.n561 0.906
R9463 vdd3p3.n566 vdd3p3.n565 0.906
R9464 vdd3p3.n569 vdd3p3.n549 0.906
R9465 vdd3p3.n572 vdd3p3.n571 0.906
R9466 vdd3p3.n575 vdd3p3.n547 0.906
R9467 vdd3p3.n581 vdd3p3.n577 0.906
R9468 vdd3p3.n3766 vdd3p3.n3763 0.903
R9469 vdd3p3.n3780 vdd3p3.n3512 0.903
R9470 vdd3p3.n5343 vdd3p3.n5320 0.902
R9471 vdd3p3.n5009 vdd3p3.n5008 0.899
R9472 vdd3p3.n7470 vdd3p3.n7467 0.899
R9473 vdd3p3.n6661 vdd3p3.n6660 0.898
R9474 vdd3p3.n6576 vdd3p3.n6575 0.898
R9475 vdd3p3.n6485 vdd3p3.n6484 0.898
R9476 vdd3p3.n5005 vdd3p3.n5004 0.884
R9477 vdd3p3.n5004 vdd3p3.n4732 0.883
R9478 vdd3p3.n8002 vdd3p3.n8001 0.88
R9479 vdd3p3.n8113 vdd3p3.n8112 0.88
R9480 vdd3p3.n8218 vdd3p3.n8217 0.88
R9481 vdd3p3.n8339 vdd3p3.n8338 0.88
R9482 vdd3p3.n5739 vdd3p3.n5734 0.88
R9483 vdd3p3.n7442 vdd3p3.n7441 0.878
R9484 vdd3p3.n7406 vdd3p3.n7405 0.878
R9485 vdd3p3.n4857 vdd3p3.n4856 0.853
R9486 vdd3p3.n3786 vdd3p3.n3785 0.849
R9487 vdd3p3.n44 vdd3p3.n42 0.84
R9488 vdd3p3.n42 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.84
R9489 vdd3p3.n1735 vdd3p3.n1733 0.84
R9490 vdd3p3.n1733 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.84
R9491 vdd3p3.n3785 vdd3p3.n3458 0.828
R9492 vdd3p3.n3785 vdd3p3.n3465 0.825
R9493 vdd3p3.n7531 vdd3p3.n7530 0.823
R9494 vdd3p3.n6698 vdd3p3.n6697 0.813
R9495 vdd3p3.n6611 vdd3p3.n6610 0.813
R9496 vdd3p3.n6523 vdd3p3.n6522 0.813
R9497 vdd3p3.n6435 vdd3p3.n6434 0.813
R9498 vdd3p3.n8055 vdd3p3.n8054 0.812
R9499 vdd3p3.n8160 vdd3p3.n8159 0.812
R9500 vdd3p3.n8265 vdd3p3.n8264 0.812
R9501 vdd3p3.n8411 vdd3p3.n8410 0.812
R9502 vdd3p3.n8463 vdd3p3.n8462 0.812
R9503 vdd3p3.n7350 vdd3p3.n7349 0.808
R9504 vdd3p3.n7327 vdd3p3.n7326 0.808
R9505 vdd3p3.n7281 vdd3p3.n7280 0.808
R9506 vdd3p3.n7258 vdd3p3.n7257 0.808
R9507 vdd3p3.n7207 vdd3p3.n7206 0.808
R9508 vdd3p3.n7178 vdd3p3.n7177 0.808
R9509 vdd3p3.n7120 vdd3p3.n7119 0.808
R9510 vdd3p3.n7091 vdd3p3.n7090 0.808
R9511 vdd3p3.n7033 vdd3p3.n7032 0.808
R9512 vdd3p3.n6387 vdd3p3.n6386 0.795
R9513 vdd3p3.n6308 vdd3p3.n6307 0.795
R9514 vdd3p3.n6225 vdd3p3.n6224 0.795
R9515 vdd3p3.n6137 vdd3p3.n6136 0.795
R9516 vdd3p3.n6063 vdd3p3.n6062 0.795
R9517 vdd3p3.n5993 vdd3p3.n5992 0.795
R9518 vdd3p3.n5916 vdd3p3.n5915 0.795
R9519 vdd3p3.n5828 vdd3p3.n5827 0.795
R9520 vdd3p3.n5740 vdd3p3.n5731 0.795
R9521 vdd3p3.n4062 vdd3p3.n4061 0.793
R9522 vdd3p3.n3435 vdd3p3.n3434 0.774
R9523 vdd3p3.n5130 vdd3p3.n5129 0.774
R9524 vdd3p3.n7471 vdd3p3.n7458 0.761
R9525 vdd3p3.n37 vdd3p3.n36 0.76
R9526 vdd3p3.n890 vdd3p3.n889 0.76
R9527 vdd3p3.n1728 vdd3p3.n1727 0.76
R9528 vdd3p3.n2581 vdd3p3.n2580 0.76
R9529 vdd3p3.n4262 vdd3p3.n4258 0.752
R9530 vdd3p3.n4278 vdd3p3.n4274 0.752
R9531 vdd3p3.n4582 vdd3p3.n4578 0.752
R9532 vdd3p3.n4598 vdd3p3.n4594 0.752
R9533 vdd3p3.n3586 vdd3p3.n3585 0.752
R9534 vdd3p3.n3524 vdd3p3.n3520 0.752
R9535 vdd3p3.n3540 vdd3p3.n3536 0.752
R9536 vdd3p3.n3609 vdd3p3.n3605 0.752
R9537 vdd3p3.n3708 vdd3p3.n3704 0.752
R9538 vdd3p3.n3637 vdd3p3.n3633 0.752
R9539 vdd3p3.n3627 vdd3p3.n3623 0.752
R9540 vdd3p3.n3680 vdd3p3.n3679 0.752
R9541 vdd3p3.n3750 vdd3p3.n3749 0.752
R9542 vdd3p3.n3496 vdd3p3.n3495 0.752
R9543 vdd3p3.n4815 vdd3p3.n4814 0.752
R9544 vdd3p3.n4773 vdd3p3.n4769 0.752
R9545 vdd3p3.n4746 vdd3p3.n4745 0.752
R9546 vdd3p3.n4978 vdd3p3.n4977 0.752
R9547 vdd3p3.n4914 vdd3p3.n4910 0.752
R9548 vdd3p3.n8544 vdd3p3.n8543 0.752
R9549 vdd3p3.n8491 vdd3p3.n8490 0.752
R9550 vdd3p3.n8592 vdd3p3.n8591 0.752
R9551 vdd3p3.n8569 vdd3p3.n8568 0.752
R9552 vdd3p3.n8623 vdd3p3.n8622 0.752
R9553 vdd3p3.n8835 vdd3p3.n8834 0.752
R9554 vdd3p3.n8806 vdd3p3.n8805 0.752
R9555 vdd3p3.n8753 vdd3p3.n8752 0.752
R9556 vdd3p3.n3817 vdd3p3.n3816 0.752
R9557 vdd3p3.n3831 vdd3p3.n3830 0.752
R9558 vdd3p3.n2881 vdd3p3.n2840 0.75
R9559 vdd3p3.n2669 vdd3p3.n2637 0.75
R9560 vdd3p3.n2035 vdd3p3.n1994 0.75
R9561 vdd3p3.n1823 vdd3p3.n1791 0.75
R9562 vdd3p3.n1190 vdd3p3.n1149 0.75
R9563 vdd3p3.n978 vdd3p3.n946 0.75
R9564 vdd3p3.n344 vdd3p3.n303 0.75
R9565 vdd3p3.n132 vdd3p3.n100 0.75
R9566 vdd3p3.n3770 vdd3p3.n3693 0.743
R9567 vdd3p3.n4831 vdd3p3.n4828 0.743
R9568 vdd3p3.n3775 vdd3p3.n3599 0.743
R9569 vdd3p3.n6656 vdd3p3.n6655 0.727
R9570 vdd3p3.n6572 vdd3p3.n6571 0.727
R9571 vdd3p3.n6480 vdd3p3.n6479 0.727
R9572 vdd3p3.n8713 vdd3p3.n8711 0.727
R9573 vdd3p3.n3998 vdd3p3.n3987 0.725
R9574 vdd3p3.n3998 vdd3p3.n3997 0.724
R9575 vdd3p3.n5343 vdd3p3.n5300 0.712
R9576 vdd3p3.n2840 vdd3p3.n2838 0.707
R9577 vdd3p3.n1994 vdd3p3.n1992 0.707
R9578 vdd3p3.n1149 vdd3p3.n1147 0.707
R9579 vdd3p3.n303 vdd3p3.n301 0.707
R9580 vdd3p3.n3314 vdd3p3.n2684 0.7
R9581 vdd3p3.n2468 vdd3p3.n1838 0.7
R9582 vdd3p3.n1623 vdd3p3.n993 0.7
R9583 vdd3p3.n777 vdd3p3.n147 0.7
R9584 vdd3p3.n5149 vdd3p3.n3397 0.698
R9585 vdd3p3.n7899 vdd3p3.n7898 0.697
R9586 vdd3p3.n7813 vdd3p3.n7812 0.697
R9587 vdd3p3.n7757 vdd3p3.n7756 0.697
R9588 vdd3p3.n7681 vdd3p3.n7680 0.697
R9589 vdd3p3.n7625 vdd3p3.n7624 0.697
R9590 vdd3p3.n7539 vdd3p3.n7538 0.697
R9591 vdd3p3.n4172 vdd3p3.n4169 0.692
R9592 vdd3p3.n4863 vdd3p3.n4841 0.682
R9593 vdd3p3.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.682
R9594 vdd3p3.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.682
R9595 vdd3p3.n1736 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.682
R9596 vdd3p3.n1736 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.682
R9597 vdd3p3.n8563 vdd3p3.n8562 0.682
R9598 vdd3p3.n4406 vdd3p3.n4405 0.682
R9599 vdd3p3.n4436 vdd3p3.n4435 0.682
R9600 vdd3p3.n4466 vdd3p3.n4465 0.682
R9601 vdd3p3.n4496 vdd3p3.n4495 0.682
R9602 vdd3p3.n5143 vdd3p3.n5142 0.682
R9603 vdd3p3.n4548 vdd3p3.n4547 0.682
R9604 vdd3p3.n4885 vdd3p3.n4884 0.682
R9605 vdd3p3.n3115 vdd3p3.n2753 0.679
R9606 vdd3p3.n2269 vdd3p3.n1907 0.679
R9607 vdd3p3.n1424 vdd3p3.n1062 0.679
R9608 vdd3p3.n578 vdd3p3.n216 0.679
R9609 vdd3p3.n6975 vdd3p3.n6974 0.677
R9610 vdd3p3.n6950 vdd3p3.n6949 0.677
R9611 vdd3p3.n6887 vdd3p3.n6886 0.677
R9612 vdd3p3.n6862 vdd3p3.n6861 0.677
R9613 vdd3p3.n6799 vdd3p3.n6798 0.677
R9614 vdd3p3.n6774 vdd3p3.n6773 0.677
R9615 vdd3p3.n5354 vdd3p3.n5353 0.677
R9616 vdd3p3.n5379 vdd3p3.n5378 0.677
R9617 vdd3p3.n5442 vdd3p3.n5441 0.677
R9618 vdd3p3.n5467 vdd3p3.n5466 0.677
R9619 vdd3p3.n5530 vdd3p3.n5529 0.677
R9620 vdd3p3.n5555 vdd3p3.n5554 0.677
R9621 vdd3p3.n5618 vdd3p3.n5617 0.677
R9622 vdd3p3.n5643 vdd3p3.n5642 0.677
R9623 vdd3p3.n5706 vdd3p3.n5705 0.677
R9624 vdd3p3.n4022 vdd3p3.t85 0.661
R9625 vdd3p3.n4097 vdd3p3.t34 0.661
R9626 vdd3p3.n6331 vdd3p3.n6330 0.65
R9627 vdd3p3.n6250 vdd3p3.n6249 0.65
R9628 vdd3p3.n6162 vdd3p3.n6161 0.65
R9629 vdd3p3.n6083 vdd3p3.n6082 0.65
R9630 vdd3p3.n6013 vdd3p3.n6012 0.65
R9631 vdd3p3.n5941 vdd3p3.n5940 0.65
R9632 vdd3p3.n5853 vdd3p3.n5852 0.65
R9633 vdd3p3.n5765 vdd3p3.n5764 0.65
R9634 vdd3p3.n8705 vdd3p3.n8704 0.647
R9635 vdd3p3.n6702 vdd3p3.n6701 0.642
R9636 vdd3p3.n6616 vdd3p3.n6615 0.642
R9637 vdd3p3.n6527 vdd3p3.n6526 0.642
R9638 vdd3p3.n6440 vdd3p3.n6439 0.642
R9639 vdd3p3.n8744 vdd3p3.n8743 0.63
R9640 vdd3p3.n7437 vdd3p3.n7436 0.627
R9641 vdd3p3.n7411 vdd3p3.n7410 0.627
R9642 vdd3p3.n5032 vdd3p3.n5029 0.614
R9643 vdd3p3.n3087 vdd3p3.n3034 0.612
R9644 vdd3p3.n3158 vdd3p3.n3157 0.612
R9645 vdd3p3.n3156 vdd3p3.n3155 0.612
R9646 vdd3p3.n3076 vdd3p3.n3039 0.612
R9647 vdd3p3.n2241 vdd3p3.n2188 0.612
R9648 vdd3p3.n2312 vdd3p3.n2311 0.612
R9649 vdd3p3.n2310 vdd3p3.n2309 0.612
R9650 vdd3p3.n2230 vdd3p3.n2193 0.612
R9651 vdd3p3.n1396 vdd3p3.n1343 0.612
R9652 vdd3p3.n1467 vdd3p3.n1466 0.612
R9653 vdd3p3.n1465 vdd3p3.n1464 0.612
R9654 vdd3p3.n1385 vdd3p3.n1348 0.612
R9655 vdd3p3.n550 vdd3p3.n497 0.612
R9656 vdd3p3.n621 vdd3p3.n620 0.612
R9657 vdd3p3.n619 vdd3p3.n618 0.612
R9658 vdd3p3.n539 vdd3p3.n502 0.612
R9659 vdd3p3.n8008 vdd3p3.n8007 0.609
R9660 vdd3p3.n8119 vdd3p3.n8118 0.609
R9661 vdd3p3.n8224 vdd3p3.n8223 0.609
R9662 vdd3p3.n8349 vdd3p3.n8348 0.609
R9663 vdd3p3.n3180 vdd3p3.n3020 0.604
R9664 vdd3p3.n3031 vdd3p3.n3029 0.604
R9665 vdd3p3.n3174 vdd3p3.n3173 0.604
R9666 vdd3p3.n3171 vdd3p3.n3170 0.604
R9667 vdd3p3.n3168 vdd3p3.n3166 0.604
R9668 vdd3p3.n3164 vdd3p3.n3032 0.604
R9669 vdd3p3.n2334 vdd3p3.n2174 0.604
R9670 vdd3p3.n2185 vdd3p3.n2183 0.604
R9671 vdd3p3.n2328 vdd3p3.n2327 0.604
R9672 vdd3p3.n2325 vdd3p3.n2324 0.604
R9673 vdd3p3.n2322 vdd3p3.n2320 0.604
R9674 vdd3p3.n2318 vdd3p3.n2186 0.604
R9675 vdd3p3.n1489 vdd3p3.n1329 0.604
R9676 vdd3p3.n1340 vdd3p3.n1338 0.604
R9677 vdd3p3.n1483 vdd3p3.n1482 0.604
R9678 vdd3p3.n1480 vdd3p3.n1479 0.604
R9679 vdd3p3.n1477 vdd3p3.n1475 0.604
R9680 vdd3p3.n1473 vdd3p3.n1341 0.604
R9681 vdd3p3.n643 vdd3p3.n483 0.604
R9682 vdd3p3.n494 vdd3p3.n492 0.604
R9683 vdd3p3.n637 vdd3p3.n636 0.604
R9684 vdd3p3.n634 vdd3p3.n633 0.604
R9685 vdd3p3.n631 vdd3p3.n629 0.604
R9686 vdd3p3.n627 vdd3p3.n495 0.604
R9687 vdd3p3.n4995 vdd3p3.n4994 0.604
R9688 vdd3p3.n4886 vdd3p3.n4759 0.604
R9689 vdd3p3.n4759 vdd3p3.n4733 0.575
R9690 vdd3p3.n7945 vdd3p3.n7942 0.57
R9691 vdd3p3.n7526 vdd3p3.n7525 0.57
R9692 vdd3p3.n8888 vdd3p3.n8887 0.568
R9693 vdd3p3.n6651 vdd3p3.n6650 0.556
R9694 vdd3p3.n6568 vdd3p3.n6567 0.556
R9695 vdd3p3.n6475 vdd3p3.n6474 0.556
R9696 vdd3p3.n8708 vdd3p3.n8707 0.556
R9697 vdd3p3.n43 vdd3p3.n0 0.543
R9698 vdd3p3.n907 vdd3p3.n906 0.543
R9699 vdd3p3.n1734 vdd3p3.n1691 0.543
R9700 vdd3p3.n2598 vdd3p3.n2597 0.543
R9701 vdd3p3.n8049 vdd3p3.n8048 0.541
R9702 vdd3p3.n8154 vdd3p3.n8153 0.541
R9703 vdd3p3.n8259 vdd3p3.n8258 0.541
R9704 vdd3p3.n8402 vdd3p3.n8401 0.541
R9705 vdd3p3.n7346 vdd3p3.n7345 0.538
R9706 vdd3p3.n7331 vdd3p3.n7330 0.538
R9707 vdd3p3.n7277 vdd3p3.n7276 0.538
R9708 vdd3p3.n7262 vdd3p3.n7261 0.538
R9709 vdd3p3.n7202 vdd3p3.n7201 0.538
R9710 vdd3p3.n7183 vdd3p3.n7182 0.538
R9711 vdd3p3.n7115 vdd3p3.n7114 0.538
R9712 vdd3p3.n7096 vdd3p3.n7095 0.538
R9713 vdd3p3.n7028 vdd3p3.n7027 0.538
R9714 vdd3p3.n905 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPB 0.529
R9715 vdd3p3.n2596 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPB 0.529
R9716 vdd3p3.n8456 vdd3p3.n8455 0.529
R9717 vdd3p3.n8466 vdd3p3.n5345 0.522
R9718 vdd3p3.n5343 vdd3p3.n5265 0.522
R9719 vdd3p3.n8655 vdd3p3.n8654 0.515
R9720 vdd3p3.n2857 vdd3p3.n2601 0.514
R9721 vdd3p3.n2011 vdd3p3.n1755 0.514
R9722 vdd3p3.n1166 vdd3p3.n910 0.514
R9723 vdd3p3.n320 vdd3p3.n64 0.514
R9724 vdd3p3.n6397 vdd3p3.n6396 0.506
R9725 vdd3p3.n6312 vdd3p3.n6311 0.506
R9726 vdd3p3.n6230 vdd3p3.n6229 0.506
R9727 vdd3p3.n6142 vdd3p3.n6141 0.506
R9728 vdd3p3.n6067 vdd3p3.n6066 0.506
R9729 vdd3p3.n5997 vdd3p3.n5996 0.506
R9730 vdd3p3.n5921 vdd3p3.n5920 0.506
R9731 vdd3p3.n5833 vdd3p3.n5832 0.506
R9732 vdd3p3.n5745 vdd3p3.n5744 0.506
R9733 vdd3p3.n7467 vdd3p3.n7466 0.501
R9734 vdd3p3.n904 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.497
R9735 vdd3p3.n2595 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.497
R9736 vdd3p3.n3789 vdd3p3.n3788 0.491
R9737 vdd3p3.n4000 vdd3p3.n3999 0.49
R9738 vdd3p3.n4001 vdd3p3.n4000 0.487
R9739 vdd3p3.n7476 vdd3p3.n7475 0.484
R9740 vdd3p3.n3670 vdd3p3.n3669 0.481
R9741 vdd3p3.n4805 vdd3p3.n4804 0.481
R9742 vdd3p3.n8572 vdd3p3.n8571 0.475
R9743 vdd3p3.n7955 vdd3p3.n7952 0.474
R9744 vdd3p3.n7961 vdd3p3.n7959 0.474
R9745 vdd3p3.n7979 vdd3p3.n7977 0.474
R9746 vdd3p3.n7987 vdd3p3.n7984 0.474
R9747 vdd3p3.n7993 vdd3p3.n7991 0.474
R9748 vdd3p3.n8001 vdd3p3.n7998 0.474
R9749 vdd3p3.n8007 vdd3p3.n8005 0.474
R9750 vdd3p3.n8015 vdd3p3.n8012 0.474
R9751 vdd3p3.n8022 vdd3p3.n8019 0.474
R9752 vdd3p3.n8037 vdd3p3.n8035 0.474
R9753 vdd3p3.n8042 vdd3p3.n8040 0.474
R9754 vdd3p3.n8048 vdd3p3.n8046 0.474
R9755 vdd3p3.n8054 vdd3p3.n8052 0.474
R9756 vdd3p3.n8060 vdd3p3.n8058 0.474
R9757 vdd3p3.n8066 vdd3p3.n8064 0.474
R9758 vdd3p3.n8072 vdd3p3.n8070 0.474
R9759 vdd3p3.n8078 vdd3p3.n8076 0.474
R9760 vdd3p3.n8094 vdd3p3.n8092 0.474
R9761 vdd3p3.n8100 vdd3p3.n8098 0.474
R9762 vdd3p3.n8106 vdd3p3.n8104 0.474
R9763 vdd3p3.n8112 vdd3p3.n8110 0.474
R9764 vdd3p3.n8118 vdd3p3.n8116 0.474
R9765 vdd3p3.n8124 vdd3p3.n8122 0.474
R9766 vdd3p3.n8130 vdd3p3.n8128 0.474
R9767 vdd3p3.n8142 vdd3p3.n8140 0.474
R9768 vdd3p3.n8147 vdd3p3.n8145 0.474
R9769 vdd3p3.n8153 vdd3p3.n8151 0.474
R9770 vdd3p3.n8159 vdd3p3.n8157 0.474
R9771 vdd3p3.n8165 vdd3p3.n8163 0.474
R9772 vdd3p3.n8171 vdd3p3.n8169 0.474
R9773 vdd3p3.n8177 vdd3p3.n8175 0.474
R9774 vdd3p3.n8183 vdd3p3.n8181 0.474
R9775 vdd3p3.n8199 vdd3p3.n8197 0.474
R9776 vdd3p3.n8205 vdd3p3.n8203 0.474
R9777 vdd3p3.n8211 vdd3p3.n8209 0.474
R9778 vdd3p3.n8217 vdd3p3.n8215 0.474
R9779 vdd3p3.n8223 vdd3p3.n8221 0.474
R9780 vdd3p3.n8229 vdd3p3.n8227 0.474
R9781 vdd3p3.n8235 vdd3p3.n8233 0.474
R9782 vdd3p3.n8247 vdd3p3.n8245 0.474
R9783 vdd3p3.n8252 vdd3p3.n8250 0.474
R9784 vdd3p3.n8258 vdd3p3.n8256 0.474
R9785 vdd3p3.n8264 vdd3p3.n8262 0.474
R9786 vdd3p3.n8270 vdd3p3.n8268 0.474
R9787 vdd3p3.n8276 vdd3p3.n8274 0.474
R9788 vdd3p3.n8282 vdd3p3.n8280 0.474
R9789 vdd3p3.n8288 vdd3p3.n8286 0.474
R9790 vdd3p3.n8308 vdd3p3.n8305 0.474
R9791 vdd3p3.n8318 vdd3p3.n8315 0.474
R9792 vdd3p3.n8328 vdd3p3.n8325 0.474
R9793 vdd3p3.n8338 vdd3p3.n8335 0.474
R9794 vdd3p3.n8348 vdd3p3.n8345 0.474
R9795 vdd3p3.n8357 vdd3p3.n8354 0.474
R9796 vdd3p3.n8366 vdd3p3.n8363 0.474
R9797 vdd3p3.n8384 vdd3p3.n8380 0.474
R9798 vdd3p3.n8392 vdd3p3.n8388 0.474
R9799 vdd3p3.n8401 vdd3p3.n8397 0.474
R9800 vdd3p3.n8410 vdd3p3.n8406 0.474
R9801 vdd3p3.n8418 vdd3p3.n8415 0.474
R9802 vdd3p3.n8426 vdd3p3.n8423 0.474
R9803 vdd3p3.n8432 vdd3p3.n8430 0.474
R9804 vdd3p3.n4736 vdd3p3.n4735 0.471
R9805 vdd3p3.n6706 vdd3p3.n6705 0.47
R9806 vdd3p3.n6621 vdd3p3.n6620 0.47
R9807 vdd3p3.n6531 vdd3p3.n6530 0.47
R9808 vdd3p3.n6445 vdd3p3.n6444 0.47
R9809 vdd3p3.n8667 vdd3p3.n8666 0.469
R9810 vdd3p3.n3740 vdd3p3.n3739 0.467
R9811 vdd3p3.n3576 vdd3p3.n3575 0.467
R9812 vdd3p3.n8686 vdd3p3.n8685 0.461
R9813 vdd3p3.n7907 vdd3p3.n7906 0.443
R9814 vdd3p3.n7805 vdd3p3.n7804 0.443
R9815 vdd3p3.n7765 vdd3p3.n7764 0.443
R9816 vdd3p3.n7673 vdd3p3.n7672 0.443
R9817 vdd3p3.n7633 vdd3p3.n7632 0.443
R9818 vdd3p3.n7526 vdd3p3.n7510 0.443
R9819 vdd3p3.n4923 vdd3p3.n4921 0.442
R9820 vdd3p3.n2600 EF_AMUX21m_1.array_1ls_1tgm_0.vdd3p3 0.434
R9821 vdd3p3.n6394 vdd3p3.n6390 0.431
R9822 vdd3p3.n7949 vdd3p3.n7935 0.427
R9823 vdd3p3.n909 EF_AMUX21m_2.array_1ls_1tgm_0.vdd3p3 0.426
R9824 vdd3p3.n6492 vdd3p3.t104 0.42
R9825 vdd3p3.n8652 vdd3p3.n8651 0.42
R9826 vdd3p3.n8734 vdd3p3.n8727 0.42
R9827 vdd3p3.n8726 vdd3p3.n8725 0.42
R9828 vdd3p3.n6970 vdd3p3.n6969 0.406
R9829 vdd3p3.n6955 vdd3p3.n6954 0.406
R9830 vdd3p3.n6882 vdd3p3.n6881 0.406
R9831 vdd3p3.n6867 vdd3p3.n6866 0.406
R9832 vdd3p3.n6794 vdd3p3.n6793 0.406
R9833 vdd3p3.n6779 vdd3p3.n6778 0.406
R9834 vdd3p3.n5359 vdd3p3.n5358 0.406
R9835 vdd3p3.n5374 vdd3p3.n5373 0.406
R9836 vdd3p3.n5447 vdd3p3.n5446 0.406
R9837 vdd3p3.n5462 vdd3p3.n5461 0.406
R9838 vdd3p3.n5535 vdd3p3.n5534 0.406
R9839 vdd3p3.n5550 vdd3p3.n5549 0.406
R9840 vdd3p3.n5623 vdd3p3.n5622 0.406
R9841 vdd3p3.n5638 vdd3p3.n5637 0.406
R9842 vdd3p3.n5711 vdd3p3.n5710 0.406
R9843 vdd3p3.n5726 vdd3p3.n5725 0.406
R9844 vdd3p3.n4383 vdd3p3.n4382 0.4
R9845 vdd3p3.n4416 vdd3p3.n4415 0.4
R9846 vdd3p3.n4506 vdd3p3.n4505 0.4
R9847 vdd3p3.n4446 vdd3p3.n4445 0.4
R9848 vdd3p3.n4476 vdd3p3.n4475 0.4
R9849 vdd3p3.n3445 vdd3p3.n3444 0.4
R9850 vdd3p3.n4564 vdd3p3.n4563 0.4
R9851 vdd3p3.n3979 vdd3p3.n3977 0.396
R9852 vdd3p3.n6646 vdd3p3.n6645 0.385
R9853 vdd3p3.n6564 vdd3p3.n6563 0.385
R9854 vdd3p3.n6470 vdd3p3.n6469 0.385
R9855 vdd3p3.n7914 vdd3p3.n7911 0.38
R9856 vdd3p3.n7906 vdd3p3.n7903 0.38
R9857 vdd3p3.n7898 vdd3p3.n7895 0.38
R9858 vdd3p3.n7890 vdd3p3.n7887 0.38
R9859 vdd3p3.n7882 vdd3p3.n7879 0.38
R9860 vdd3p3.n7874 vdd3p3.n7871 0.38
R9861 vdd3p3.n7863 vdd3p3.n7860 0.38
R9862 vdd3p3.n7847 vdd3p3.n7844 0.38
R9863 vdd3p3.n7836 vdd3p3.n7833 0.38
R9864 vdd3p3.n7828 vdd3p3.n7825 0.38
R9865 vdd3p3.n7820 vdd3p3.n7817 0.38
R9866 vdd3p3.n7812 vdd3p3.n7809 0.38
R9867 vdd3p3.n7804 vdd3p3.n7801 0.38
R9868 vdd3p3.n7796 vdd3p3.n7793 0.38
R9869 vdd3p3.n7772 vdd3p3.n7769 0.38
R9870 vdd3p3.n7764 vdd3p3.n7761 0.38
R9871 vdd3p3.n7756 vdd3p3.n7753 0.38
R9872 vdd3p3.n7748 vdd3p3.n7745 0.38
R9873 vdd3p3.n7740 vdd3p3.n7737 0.38
R9874 vdd3p3.n7732 vdd3p3.n7729 0.38
R9875 vdd3p3.n7722 vdd3p3.n7719 0.38
R9876 vdd3p3.n7708 vdd3p3.n7706 0.38
R9877 vdd3p3.n7700 vdd3p3.n7698 0.38
R9878 vdd3p3.n7694 vdd3p3.n7692 0.38
R9879 vdd3p3.n7688 vdd3p3.n7685 0.38
R9880 vdd3p3.n7680 vdd3p3.n7677 0.38
R9881 vdd3p3.n7672 vdd3p3.n7669 0.38
R9882 vdd3p3.n7664 vdd3p3.n7661 0.38
R9883 vdd3p3.n7640 vdd3p3.n7637 0.38
R9884 vdd3p3.n7632 vdd3p3.n7629 0.38
R9885 vdd3p3.n7624 vdd3p3.n7621 0.38
R9886 vdd3p3.n7616 vdd3p3.n7613 0.38
R9887 vdd3p3.n7608 vdd3p3.n7605 0.38
R9888 vdd3p3.n7600 vdd3p3.n7597 0.38
R9889 vdd3p3.n7589 vdd3p3.n7586 0.38
R9890 vdd3p3.n7573 vdd3p3.n7570 0.38
R9891 vdd3p3.n7562 vdd3p3.n7559 0.38
R9892 vdd3p3.n7554 vdd3p3.n7551 0.38
R9893 vdd3p3.n7546 vdd3p3.n7543 0.38
R9894 vdd3p3.n7538 vdd3p3.n7535 0.38
R9895 vdd3p3.n6399 vdd3p3.n6398 0.377
R9896 vdd3p3.n4199 vdd3p3.n4195 0.376
R9897 vdd3p3.n5051 vdd3p3.n5047 0.376
R9898 vdd3p3.n3476 vdd3p3.n3473 0.376
R9899 vdd3p3.n3489 vdd3p3.n3488 0.376
R9900 vdd3p3.n3505 vdd3p3.n3504 0.376
R9901 vdd3p3.n4958 vdd3p3.n4954 0.376
R9902 vdd3p3.n4971 vdd3p3.n4970 0.376
R9903 vdd3p3.n4987 vdd3p3.n4986 0.376
R9904 vdd3p3.n4906 vdd3p3.n4905 0.376
R9905 vdd3p3.n8552 vdd3p3.n8551 0.376
R9906 vdd3p3.n8555 vdd3p3.n8554 0.376
R9907 vdd3p3.n8535 vdd3p3.n8534 0.376
R9908 vdd3p3.n8498 vdd3p3.n8497 0.376
R9909 vdd3p3.n8505 vdd3p3.n8501 0.376
R9910 vdd3p3.n8597 vdd3p3.n8596 0.376
R9911 vdd3p3.n8631 vdd3p3.n8630 0.376
R9912 vdd3p3.n8634 vdd3p3.n8633 0.376
R9913 vdd3p3.n8880 vdd3p3.n8879 0.376
R9914 vdd3p3.n8842 vdd3p3.n8841 0.376
R9915 vdd3p3.n8849 vdd3p3.n8845 0.376
R9916 vdd3p3.n8814 vdd3p3.n8813 0.376
R9917 vdd3p3.n8817 vdd3p3.n8816 0.376
R9918 vdd3p3.n8797 vdd3p3.n8796 0.376
R9919 vdd3p3.n8784 vdd3p3.n8783 0.376
R9920 vdd3p3.n8760 vdd3p3.n8756 0.376
R9921 vdd3p3.n7432 vdd3p3.n7431 0.376
R9922 vdd3p3.n7416 vdd3p3.n7415 0.376
R9923 vdd3p3.n6326 vdd3p3.n6325 0.361
R9924 vdd3p3.n6245 vdd3p3.n6244 0.361
R9925 vdd3p3.n6157 vdd3p3.n6156 0.361
R9926 vdd3p3.n6079 vdd3p3.n6078 0.361
R9927 vdd3p3.n6009 vdd3p3.n6008 0.361
R9928 vdd3p3.n5936 vdd3p3.n5935 0.361
R9929 vdd3p3.n5848 vdd3p3.n5847 0.361
R9930 vdd3p3.n5760 vdd3p3.n5759 0.361
R9931 vdd3p3.n3826 vdd3p3.n3824 0.356
R9932 vdd3p3.n7491 vdd3p3.n7490 0.345
R9933 vdd3p3.n2877 vdd3p3.n2841 0.343
R9934 vdd3p3.n2876 vdd3p3.n2843 0.343
R9935 vdd3p3.n2872 vdd3p3.n2871 0.343
R9936 vdd3p3.n2867 vdd3p3.n2847 0.343
R9937 vdd3p3.n2866 vdd3p3.n2850 0.343
R9938 vdd3p3.n2863 vdd3p3.n2862 0.343
R9939 vdd3p3.n2031 vdd3p3.n1995 0.343
R9940 vdd3p3.n2030 vdd3p3.n1997 0.343
R9941 vdd3p3.n2026 vdd3p3.n2025 0.343
R9942 vdd3p3.n2021 vdd3p3.n2001 0.343
R9943 vdd3p3.n2020 vdd3p3.n2004 0.343
R9944 vdd3p3.n2017 vdd3p3.n2016 0.343
R9945 vdd3p3.n1186 vdd3p3.n1150 0.343
R9946 vdd3p3.n1185 vdd3p3.n1152 0.343
R9947 vdd3p3.n1181 vdd3p3.n1180 0.343
R9948 vdd3p3.n1176 vdd3p3.n1156 0.343
R9949 vdd3p3.n1175 vdd3p3.n1159 0.343
R9950 vdd3p3.n1172 vdd3p3.n1171 0.343
R9951 vdd3p3.n340 vdd3p3.n304 0.343
R9952 vdd3p3.n339 vdd3p3.n306 0.343
R9953 vdd3p3.n335 vdd3p3.n334 0.343
R9954 vdd3p3.n330 vdd3p3.n310 0.343
R9955 vdd3p3.n329 vdd3p3.n313 0.343
R9956 vdd3p3.n326 vdd3p3.n325 0.343
R9957 vdd3p3.n4782 vdd3p3.n4780 0.339
R9958 vdd3p3.n8016 vdd3p3.n8015 0.338
R9959 vdd3p3.n8125 vdd3p3.n8124 0.338
R9960 vdd3p3.n8230 vdd3p3.n8229 0.338
R9961 vdd3p3.n8358 vdd3p3.n8357 0.338
R9962 vdd3p3.n7011 vdd3p3.n7010 0.336
R9963 vdd3p3.n5021 vdd3p3.n5020 0.33
R9964 vdd3p3.n5022 vdd3p3.n4721 0.33
R9965 vdd3p3.n4720 vdd3p3.n4719 0.33
R9966 vdd3p3.n902 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.329
R9967 vdd3p3.n2593 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.329
R9968 vdd3p3.n3778 vdd3p3.n3777 0.324
R9969 vdd3p3.n3773 vdd3p3.n3772 0.324
R9970 vdd3p3.n3769 vdd3p3.n3768 0.324
R9971 vdd3p3.n4249 vdd3p3.n4248 0.324
R9972 vdd3p3.n4372 vdd3p3.n4371 0.324
R9973 vdd3p3.n5114 vdd3p3.n5113 0.324
R9974 vdd3p3.n5109 vdd3p3.n5108 0.324
R9975 vdd3p3.n7934 vdd3p3.n7933 0.316
R9976 vdd3p3.n7923 vdd3p3.n7919 0.316
R9977 vdd3p3.n7789 vdd3p3.n7788 0.316
R9978 vdd3p3.n7781 vdd3p3.n7777 0.316
R9979 vdd3p3.n7657 vdd3p3.n7656 0.316
R9980 vdd3p3.n7649 vdd3p3.n7645 0.316
R9981 vdd3p3.n7472 vdd3p3.n7455 0.313
R9982 vdd3p3.n8464 vdd3p3.n8463 0.308
R9983 vdd3p3.n6710 vdd3p3.n6709 0.299
R9984 vdd3p3.n6626 vdd3p3.n6625 0.299
R9985 vdd3p3.n6535 vdd3p3.n6534 0.299
R9986 vdd3p3.n6450 vdd3p3.n6449 0.299
R9987 vdd3p3.n906 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd3p3 0.298
R9988 vdd3p3.n2597 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd3p3 0.298
R9989 vdd3p3.n908 vdd3p3.n845 0.293
R9990 vdd3p3.n2599 vdd3p3.n2536 0.293
R9991 vdd3p3.n62 vdd3p3.n61 0.292
R9992 vdd3p3.n1753 vdd3p3.n1752 0.292
R9993 vdd3p3.n4520 vdd3p3.n4519 0.278
R9994 vdd3p3.n4430 vdd3p3.n4429 0.278
R9995 vdd3p3.n4688 vdd3p3.n4687 0.278
R9996 vdd3p3.n4460 vdd3p3.n4459 0.278
R9997 vdd3p3.n4366 vdd3p3.n4365 0.278
R9998 vdd3p3.n4400 vdd3p3.n4399 0.278
R9999 vdd3p3.n4490 vdd3p3.n4489 0.278
R10000 vdd3p3.n63 EF_AMUX21m_2.vdd3p3 0.276
R10001 vdd3p3.n1754 EF_AMUX21m_1.vdd3p3 0.276
R10002 vdd3p3.n7024 vdd3p3.n7016 0.272
R10003 vdd3p3.n8032 vdd3p3.n8031 0.27
R10004 vdd3p3.n8043 vdd3p3.n8042 0.27
R10005 vdd3p3.n8137 vdd3p3.n8136 0.27
R10006 vdd3p3.n8148 vdd3p3.n8147 0.27
R10007 vdd3p3.n8242 vdd3p3.n8241 0.27
R10008 vdd3p3.n8253 vdd3p3.n8252 0.27
R10009 vdd3p3.n8376 vdd3p3.n8375 0.27
R10010 vdd3p3.n8393 vdd3p3.n8392 0.27
R10011 vdd3p3.n7342 vdd3p3.n7341 0.269
R10012 vdd3p3.n7335 vdd3p3.n7334 0.269
R10013 vdd3p3.n7273 vdd3p3.n7272 0.269
R10014 vdd3p3.n7266 vdd3p3.n7265 0.269
R10015 vdd3p3.n7197 vdd3p3.n7196 0.269
R10016 vdd3p3.n7188 vdd3p3.n7187 0.269
R10017 vdd3p3.n7110 vdd3p3.n7109 0.269
R10018 vdd3p3.n7101 vdd3p3.n7100 0.269
R10019 vdd3p3.n7023 vdd3p3.n7022 0.269
R10020 vdd3p3.n4833 vdd3p3.n4832 0.268
R10021 vdd3p3.n3379 vdd3p3.n3378 0.266
R10022 vdd3p3.n2533 vdd3p3.n2532 0.266
R10023 vdd3p3.n1688 vdd3p3.n1687 0.266
R10024 vdd3p3.n842 vdd3p3.n841 0.266
R10025 vdd3p3.t85 vdd3p3.n4021 0.264
R10026 vdd3p3.t34 vdd3p3.n4096 0.264
R10027 vdd3p3.n49 vdd3p3.n37 0.26
R10028 vdd3p3.n49 vdd3p3.n48 0.26
R10029 vdd3p3.n48 vdd3p3.n47 0.26
R10030 vdd3p3.n891 vdd3p3.n890 0.26
R10031 vdd3p3.n891 vdd3p3.n846 0.26
R10032 vdd3p3.n899 vdd3p3.n846 0.26
R10033 vdd3p3.n1740 vdd3p3.n1728 0.26
R10034 vdd3p3.n1740 vdd3p3.n1739 0.26
R10035 vdd3p3.n1739 vdd3p3.n1738 0.26
R10036 vdd3p3.n2582 vdd3p3.n2581 0.26
R10037 vdd3p3.n2582 vdd3p3.n2537 0.26
R10038 vdd3p3.n2590 vdd3p3.n2537 0.26
R10039 vdd3p3.n3387 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VPB 0.259
R10040 vdd3p3.n3395 vdd3p3.n3394 0.254
R10041 vdd3p3.n5741 vdd3p3.n5727 0.235
R10042 vdd3p3.n54 vdd3p3.n31 0.231
R10043 vdd3p3.n896 vdd3p3.n885 0.231
R10044 vdd3p3.n1745 vdd3p3.n1722 0.231
R10045 vdd3p3.n2587 vdd3p3.n2576 0.231
R10046 vdd3p3.n54 vdd3p3.n53 0.231
R10047 vdd3p3.n54 vdd3p3.n32 0.231
R10048 vdd3p3.n896 vdd3p3.n895 0.231
R10049 vdd3p3.n897 vdd3p3.n896 0.231
R10050 vdd3p3.n1745 vdd3p3.n1744 0.231
R10051 vdd3p3.n1745 vdd3p3.n1723 0.231
R10052 vdd3p3.n2587 vdd3p3.n2586 0.231
R10053 vdd3p3.n2588 vdd3p3.n2587 0.231
R10054 vdd3p3.n4285 vdd3p3.n4269 0.228
R10055 vdd3p3.n4285 vdd3p3.n4284 0.228
R10056 vdd3p3.n4605 vdd3p3.n4589 0.228
R10057 vdd3p3.n4605 vdd3p3.n4604 0.228
R10058 vdd3p3.n3548 vdd3p3.n3531 0.228
R10059 vdd3p3.n3548 vdd3p3.n3547 0.228
R10060 vdd3p3.n3644 vdd3p3.n3616 0.228
R10061 vdd3p3.n3644 vdd3p3.n3643 0.228
R10062 vdd3p3.n3715 vdd3p3.n3699 0.228
R10063 vdd3p3.n3715 vdd3p3.n3714 0.228
R10064 vdd3p3.n909 vdd3p3.n908 0.222
R10065 vdd3p3.n2600 vdd3p3.n2599 0.222
R10066 vdd3p3.n63 vdd3p3.n62 0.221
R10067 vdd3p3.n1754 vdd3p3.n1753 0.221
R10068 vdd3p3.n6317 vdd3p3.n6316 0.216
R10069 vdd3p3.n6235 vdd3p3.n6234 0.216
R10070 vdd3p3.n6147 vdd3p3.n6146 0.216
R10071 vdd3p3.n6071 vdd3p3.n6070 0.216
R10072 vdd3p3.n6001 vdd3p3.n6000 0.216
R10073 vdd3p3.n5926 vdd3p3.n5925 0.216
R10074 vdd3p3.n5838 vdd3p3.n5837 0.216
R10075 vdd3p3.n5750 vdd3p3.n5749 0.216
R10076 vdd3p3.n6717 vdd3p3.n6716 0.215
R10077 vdd3p3.n4287 vdd3p3.n4285 0.214
R10078 vdd3p3.n4607 vdd3p3.n4605 0.214
R10079 vdd3p3.n3646 vdd3p3.n3644 0.214
R10080 vdd3p3.n3717 vdd3p3.n3715 0.214
R10081 vdd3p3.n3550 vdd3p3.n3548 0.214
R10082 vdd3p3.n2606 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.vdd 0.214
R10083 vdd3p3.n1760 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.vdd 0.214
R10084 vdd3p3.n915 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.vdd 0.214
R10085 vdd3p3.n69 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.vdd 0.214
R10086 vdd3p3.n6641 vdd3p3.n6640 0.214
R10087 vdd3p3.n6547 vdd3p3.n6546 0.214
R10088 vdd3p3.n6465 vdd3p3.n6464 0.214
R10089 vdd3p3.n7383 vdd3p3.n7381 0.213
R10090 vdd3p3.n4155 vdd3p3.n4147 0.211
R10091 vdd3p3.n8437 vdd3p3.n6717 0.21
R10092 vdd3p3.n8605 vdd3p3.n8604 0.21
R10093 vdd3p3.n4242 vdd3p3.n4239 0.21
R10094 vdd3p3.n5102 vdd3p3.n5099 0.21
R10095 vdd3p3.n7481 vdd3p3.n7480 0.207
R10096 vdd3p3.n8032 vdd3p3.n8026 0.203
R10097 vdd3p3.n8137 vdd3p3.n8134 0.203
R10098 vdd3p3.n8242 vdd3p3.n8239 0.203
R10099 vdd3p3.n8376 vdd3p3.n8371 0.203
R10100 vdd3p3.n4526 vdd3p3.n4525 0.202
R10101 vdd3p3.n8897 vdd3p3.n5161 0.202
R10102 vdd3p3.n2637 vdd3p3.n2601 0.192
R10103 vdd3p3.n1791 vdd3p3.n1755 0.192
R10104 vdd3p3.n946 vdd3p3.n910 0.192
R10105 vdd3p3.n100 vdd3p3.n64 0.192
R10106 vdd3p3.n4330 vdd3p3.n4328 0.19
R10107 vdd3p3.n4650 vdd3p3.n4648 0.19
R10108 vdd3p3.n3541 vdd3p3.n3534 0.19
R10109 vdd3p3.n3638 vdd3p3.n3631 0.19
R10110 vdd3p3.n3631 vdd3p3.n3628 0.19
R10111 vdd3p3.n7915 vdd3p3.n7914 0.19
R10112 vdd3p3.n7797 vdd3p3.n7796 0.19
R10113 vdd3p3.n7773 vdd3p3.n7772 0.19
R10114 vdd3p3.n7665 vdd3p3.n7664 0.19
R10115 vdd3p3.n7641 vdd3p3.n7640 0.19
R10116 vdd3p3.n3846 vdd3p3.n3845 0.189
R10117 vdd3p3.n8693 vdd3p3.n8692 0.185
R10118 vdd3p3.n3820 vdd3p3.n3818 0.178
R10119 vdd3p3.n3979 vdd3p3.n3897 0.176
R10120 vdd3p3.n61 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vdd3p3 0.172
R10121 vdd3p3.n1752 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vdd3p3 0.172
R10122 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vdd3p3 vdd3p3.n845 0.172
R10123 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vdd3p3 vdd3p3.n2536 0.172
R10124 vdd3p3.n44 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.167
R10125 vdd3p3.n1735 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.167
R10126 vdd3p3.n3816 vdd3p3.n3815 0.166
R10127 vdd3p3.n3376 vdd3p3.n2607 0.166
R10128 vdd3p3.n2530 vdd3p3.n1761 0.166
R10129 vdd3p3.n1685 vdd3p3.n916 0.166
R10130 vdd3p3.n839 vdd3p3.n70 0.166
R10131 vdd3p3.n4289 vdd3p3.n4287 0.164
R10132 vdd3p3.n4609 vdd3p3.n4607 0.164
R10133 vdd3p3.n3648 vdd3p3.n3646 0.164
R10134 vdd3p3.n3719 vdd3p3.n3717 0.164
R10135 vdd3p3.n3552 vdd3p3.n3550 0.164
R10136 vdd3p3.n4925 vdd3p3.n4923 0.164
R10137 vdd3p3.n4364 vdd3p3.n4363 0.161
R10138 vdd3p3.n4293 vdd3p3.n4292 0.161
R10139 vdd3p3.n4398 vdd3p3.n4397 0.161
R10140 vdd3p3.n4428 vdd3p3.n4427 0.161
R10141 vdd3p3.n4458 vdd3p3.n4457 0.161
R10142 vdd3p3.n4488 vdd3p3.n4487 0.161
R10143 vdd3p3.n4518 vdd3p3.n4517 0.161
R10144 vdd3p3.n3432 vdd3p3.n3431 0.161
R10145 vdd3p3.n5125 vdd3p3.n5124 0.161
R10146 vdd3p3.n4686 vdd3p3.n4685 0.161
R10147 vdd3p3.n4613 vdd3p3.n4612 0.161
R10148 vdd3p3.n3556 vdd3p3.n3555 0.161
R10149 vdd3p3.n3652 vdd3p3.n3651 0.161
R10150 vdd3p3.n3723 vdd3p3.n3722 0.161
R10151 vdd3p3.n4788 vdd3p3.n4787 0.161
R10152 vdd3p3.n4269 vdd3p3.n4267 0.158
R10153 vdd3p3.n4284 vdd3p3.n4283 0.158
R10154 vdd3p3.n4589 vdd3p3.n4587 0.158
R10155 vdd3p3.n4604 vdd3p3.n4603 0.158
R10156 vdd3p3.n3531 vdd3p3.n3529 0.158
R10157 vdd3p3.n3547 vdd3p3.n3545 0.158
R10158 vdd3p3.n3616 vdd3p3.n3614 0.158
R10159 vdd3p3.n3643 vdd3p3.n3642 0.158
R10160 vdd3p3.n3714 vdd3p3.n3713 0.158
R10161 vdd3p3.n4780 vdd3p3.n4778 0.158
R10162 vdd3p3.n4921 vdd3p3.n4919 0.158
R10163 vdd3p3.n8466 vdd3p3.n8465 0.157
R10164 vdd3p3.n4359 vdd3p3.n4358 0.15
R10165 vdd3p3.n4300 vdd3p3.n4299 0.15
R10166 vdd3p3.n4376 vdd3p3.n4375 0.15
R10167 vdd3p3.n4410 vdd3p3.n4409 0.15
R10168 vdd3p3.n4440 vdd3p3.n4439 0.15
R10169 vdd3p3.n4470 vdd3p3.n4469 0.15
R10170 vdd3p3.n4500 vdd3p3.n4499 0.15
R10171 vdd3p3.n3427 vdd3p3.n3426 0.15
R10172 vdd3p3.n5119 vdd3p3.n5118 0.15
R10173 vdd3p3.n4679 vdd3p3.n4678 0.15
R10174 vdd3p3.n4620 vdd3p3.n4619 0.15
R10175 vdd3p3.n3563 vdd3p3.n3562 0.15
R10176 vdd3p3.n3659 vdd3p3.n3658 0.15
R10177 vdd3p3.n3730 vdd3p3.n3729 0.15
R10178 vdd3p3.n4795 vdd3p3.n4794 0.15
R10179 vdd3p3.n3381 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.vdd3p3 0.145
R10180 vdd3p3.n2535 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.vdd3p3 0.145
R10181 vdd3p3.n1690 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.vdd3p3 0.145
R10182 vdd3p3.n844 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.vdd3p3 0.145
R10183 vdd3p3.n4222 vdd3p3.n4215 0.144
R10184 vdd3p3.n4211 vdd3p3.n4204 0.144
R10185 vdd3p3.n4344 vdd3p3.n4341 0.144
R10186 vdd3p3.n4337 vdd3p3.n4334 0.144
R10187 vdd3p3.n4324 vdd3p3.n4322 0.144
R10188 vdd3p3.n4317 vdd3p3.n4315 0.144
R10189 vdd3p3.n4310 vdd3p3.n4308 0.144
R10190 vdd3p3.n4303 vdd3p3.n4301 0.144
R10191 vdd3p3.n4296 vdd3p3.n4294 0.144
R10192 vdd3p3.n4664 vdd3p3.n4661 0.144
R10193 vdd3p3.n4657 vdd3p3.n4654 0.144
R10194 vdd3p3.n4644 vdd3p3.n4642 0.144
R10195 vdd3p3.n4637 vdd3p3.n4635 0.144
R10196 vdd3p3.n4630 vdd3p3.n4628 0.144
R10197 vdd3p3.n4623 vdd3p3.n4621 0.144
R10198 vdd3p3.n4616 vdd3p3.n4614 0.144
R10199 vdd3p3.n5074 vdd3p3.n5067 0.144
R10200 vdd3p3.n5063 vdd3p3.n5056 0.144
R10201 vdd3p3.n3662 vdd3p3.n3660 0.144
R10202 vdd3p3.n3655 vdd3p3.n3653 0.144
R10203 vdd3p3.n3733 vdd3p3.n3731 0.144
R10204 vdd3p3.n3726 vdd3p3.n3724 0.144
R10205 vdd3p3.n3566 vdd3p3.n3564 0.144
R10206 vdd3p3.n3559 vdd3p3.n3557 0.144
R10207 vdd3p3.n4798 vdd3p3.n4796 0.144
R10208 vdd3p3.n4791 vdd3p3.n4789 0.144
R10209 vdd3p3.n4947 vdd3p3.n4945 0.144
R10210 vdd3p3.n4936 vdd3p3.n4934 0.144
R10211 vdd3p3.n8517 vdd3p3.n8510 0.144
R10212 vdd3p3.n8861 vdd3p3.n8854 0.144
R10213 vdd3p3.n8772 vdd3p3.n8765 0.144
R10214 vdd3p3.n4784 vdd3p3.n4782 0.141
R10215 vdd3p3.n4253 vdd3p3.n4252 0.138
R10216 vdd3p3.n4307 vdd3p3.n4306 0.138
R10217 vdd3p3.n4573 vdd3p3.n4572 0.138
R10218 vdd3p3.n4627 vdd3p3.n4626 0.138
R10219 vdd3p3.n6965 vdd3p3.n6964 0.135
R10220 vdd3p3.n6960 vdd3p3.n6959 0.135
R10221 vdd3p3.n6877 vdd3p3.n6876 0.135
R10222 vdd3p3.n6872 vdd3p3.n6871 0.135
R10223 vdd3p3.n6789 vdd3p3.n6788 0.135
R10224 vdd3p3.n6784 vdd3p3.n6783 0.135
R10225 vdd3p3.n5364 vdd3p3.n5363 0.135
R10226 vdd3p3.n5369 vdd3p3.n5368 0.135
R10227 vdd3p3.n5452 vdd3p3.n5451 0.135
R10228 vdd3p3.n5457 vdd3p3.n5456 0.135
R10229 vdd3p3.n5540 vdd3p3.n5539 0.135
R10230 vdd3p3.n5545 vdd3p3.n5544 0.135
R10231 vdd3p3.n5628 vdd3p3.n5627 0.135
R10232 vdd3p3.n5633 vdd3p3.n5632 0.135
R10233 vdd3p3.n5716 vdd3p3.n5715 0.135
R10234 vdd3p3.n5721 vdd3p3.n5720 0.135
R10235 vdd3p3.n3376 vdd3p3.n2606 0.134
R10236 vdd3p3.n2530 vdd3p3.n1760 0.134
R10237 vdd3p3.n1685 vdd3p3.n915 0.134
R10238 vdd3p3.n839 vdd3p3.n69 0.134
R10239 EF_AMUX21m_1.vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_1.vdd3p3 0.132
R10240 vdd3p3.n4155 vdd3p3.n4062 0.132
R10241 vdd3p3.n6714 vdd3p3.n6713 0.128
R10242 vdd3p3.n6631 vdd3p3.n6630 0.128
R10243 vdd3p3.n6539 vdd3p3.n6538 0.128
R10244 vdd3p3.n6455 vdd3p3.n6454 0.128
R10245 vdd3p3.n4343 vdd3p3.n4342 0.127
R10246 vdd3p3.n4314 vdd3p3.n4313 0.127
R10247 vdd3p3.n4663 vdd3p3.n4662 0.127
R10248 vdd3p3.n4634 vdd3p3.n4633 0.127
R10249 vdd3p3.n8896 vdd3p3.n8895 0.126
R10250 vdd3p3.n7427 vdd3p3.n7426 0.125
R10251 vdd3p3.n7421 vdd3p3.n7420 0.125
R10252 vdd3p3.n8898 vdd3p3.n8897 0.12
R10253 vdd3p3.n8897 vdd3p3.n8896 0.119
R10254 vdd3p3.n5150 vdd3p3.n5149 0.116
R10255 vdd3p3.n4336 vdd3p3.n4335 0.116
R10256 vdd3p3.n4321 vdd3p3.n4320 0.116
R10257 vdd3p3.n4656 vdd3p3.n4655 0.116
R10258 vdd3p3.n4641 vdd3p3.n4640 0.116
R10259 vdd3p3.n3382 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VPWR 0.115
R10260 vdd3p3.n3383 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VPWR 0.115
R10261 vdd3p3.n4175 vdd3p3.n4174 0.109
R10262 vdd3p3.n4849 vdd3p3.n4848 0.109
R10263 vdd3p3.n3783 vdd3p3.n3782 0.108
R10264 vdd3p3.n7935 vdd3p3.n7924 0.108
R10265 vdd3p3.n7924 vdd3p3.n7916 0.108
R10266 vdd3p3.n7916 vdd3p3.n7908 0.108
R10267 vdd3p3.n7908 vdd3p3.n7900 0.108
R10268 vdd3p3.n7900 vdd3p3.n7892 0.108
R10269 vdd3p3.n7892 vdd3p3.n7884 0.108
R10270 vdd3p3.n7884 vdd3p3.n7876 0.108
R10271 vdd3p3.n7876 vdd3p3.n7868 0.108
R10272 vdd3p3.n7868 vdd3p3.n7857 0.108
R10273 vdd3p3.n7857 vdd3p3.n7849 0.108
R10274 vdd3p3.n7849 vdd3p3.n7838 0.108
R10275 vdd3p3.n7838 vdd3p3.n7830 0.108
R10276 vdd3p3.n7830 vdd3p3.n7822 0.108
R10277 vdd3p3.n7822 vdd3p3.n7814 0.108
R10278 vdd3p3.n7814 vdd3p3.n7806 0.108
R10279 vdd3p3.n7806 vdd3p3.n7798 0.108
R10280 vdd3p3.n7798 vdd3p3.n7790 0.108
R10281 vdd3p3.n7790 vdd3p3.n7782 0.108
R10282 vdd3p3.n7782 vdd3p3.n7774 0.108
R10283 vdd3p3.n7774 vdd3p3.n7766 0.108
R10284 vdd3p3.n7766 vdd3p3.n7758 0.108
R10285 vdd3p3.n7758 vdd3p3.n7750 0.108
R10286 vdd3p3.n7750 vdd3p3.n7742 0.108
R10287 vdd3p3.n7742 vdd3p3.n7734 0.108
R10288 vdd3p3.n7734 vdd3p3.n7726 0.108
R10289 vdd3p3.n7726 vdd3p3.n7716 0.108
R10290 vdd3p3.n7716 vdd3p3.n7710 0.108
R10291 vdd3p3.n7710 vdd3p3.n7702 0.108
R10292 vdd3p3.n7702 vdd3p3.n7696 0.108
R10293 vdd3p3.n7696 vdd3p3.n7690 0.108
R10294 vdd3p3.n7690 vdd3p3.n7682 0.108
R10295 vdd3p3.n7682 vdd3p3.n7674 0.108
R10296 vdd3p3.n7674 vdd3p3.n7666 0.108
R10297 vdd3p3.n7666 vdd3p3.n7658 0.108
R10298 vdd3p3.n7658 vdd3p3.n7650 0.108
R10299 vdd3p3.n7650 vdd3p3.n7642 0.108
R10300 vdd3p3.n7642 vdd3p3.n7634 0.108
R10301 vdd3p3.n7634 vdd3p3.n7626 0.108
R10302 vdd3p3.n7626 vdd3p3.n7618 0.108
R10303 vdd3p3.n7618 vdd3p3.n7610 0.108
R10304 vdd3p3.n7610 vdd3p3.n7602 0.108
R10305 vdd3p3.n7602 vdd3p3.n7594 0.108
R10306 vdd3p3.n7594 vdd3p3.n7583 0.108
R10307 vdd3p3.n7583 vdd3p3.n7575 0.108
R10308 vdd3p3.n7575 vdd3p3.n7564 0.108
R10309 vdd3p3.n7564 vdd3p3.n7556 0.108
R10310 vdd3p3.n7556 vdd3p3.n7548 0.108
R10311 vdd3p3.n7548 vdd3p3.n7540 0.108
R10312 vdd3p3.n7540 vdd3p3.n7532 0.108
R10313 vdd3p3.n7532 vdd3p3.n7527 0.108
R10314 vdd3p3.n7527 vdd3p3.n7492 0.108
R10315 vdd3p3.n7492 vdd3p3.n7487 0.108
R10316 vdd3p3.n7487 vdd3p3.n7482 0.108
R10317 vdd3p3.n7482 vdd3p3.n7477 0.108
R10318 vdd3p3.n7477 vdd3p3.n7472 0.108
R10319 vdd3p3.n7455 vdd3p3.n7448 0.108
R10320 vdd3p3.n7448 vdd3p3.n7443 0.108
R10321 vdd3p3.n7443 vdd3p3.n7438 0.108
R10322 vdd3p3.n7438 vdd3p3.n7433 0.108
R10323 vdd3p3.n7433 vdd3p3.n7428 0.108
R10324 vdd3p3.n7428 vdd3p3.n7422 0.108
R10325 vdd3p3.n7422 vdd3p3.n7417 0.108
R10326 vdd3p3.n7417 vdd3p3.n7412 0.108
R10327 vdd3p3.n7412 vdd3p3.n7407 0.108
R10328 vdd3p3.n7407 vdd3p3.n7402 0.108
R10329 vdd3p3.n7402 vdd3p3.n7397 0.108
R10330 vdd3p3.n7397 vdd3p3.n7393 0.108
R10331 vdd3p3.n7393 vdd3p3.n7387 0.108
R10332 vdd3p3.n7387 vdd3p3.n7383 0.108
R10333 vdd3p3.n7381 vdd3p3.n7379 0.108
R10334 vdd3p3.n7379 vdd3p3.n7377 0.108
R10335 vdd3p3.n7377 vdd3p3.n7371 0.108
R10336 vdd3p3.n7371 vdd3p3.n7367 0.108
R10337 vdd3p3.n7367 vdd3p3.n7363 0.108
R10338 vdd3p3.n7363 vdd3p3.n7359 0.108
R10339 vdd3p3.n7359 vdd3p3.n7355 0.108
R10340 vdd3p3.n7355 vdd3p3.n7351 0.108
R10341 vdd3p3.n7351 vdd3p3.n7347 0.108
R10342 vdd3p3.n7347 vdd3p3.n7343 0.108
R10343 vdd3p3.n7343 vdd3p3.n7339 0.108
R10344 vdd3p3.n7339 vdd3p3.n7336 0.108
R10345 vdd3p3.n7336 vdd3p3.n7332 0.108
R10346 vdd3p3.n7332 vdd3p3.n7328 0.108
R10347 vdd3p3.n7328 vdd3p3.n7324 0.108
R10348 vdd3p3.n7324 vdd3p3.n7320 0.108
R10349 vdd3p3.n7320 vdd3p3.n7316 0.108
R10350 vdd3p3.n7316 vdd3p3.n7312 0.108
R10351 vdd3p3.n7312 vdd3p3.n7308 0.108
R10352 vdd3p3.n7308 vdd3p3.n7302 0.108
R10353 vdd3p3.n7302 vdd3p3.n7298 0.108
R10354 vdd3p3.n7298 vdd3p3.n7294 0.108
R10355 vdd3p3.n7294 vdd3p3.n7290 0.108
R10356 vdd3p3.n7290 vdd3p3.n7286 0.108
R10357 vdd3p3.n7286 vdd3p3.n7282 0.108
R10358 vdd3p3.n7282 vdd3p3.n7278 0.108
R10359 vdd3p3.n7278 vdd3p3.n7274 0.108
R10360 vdd3p3.n7274 vdd3p3.n7270 0.108
R10361 vdd3p3.n7270 vdd3p3.n7267 0.108
R10362 vdd3p3.n7267 vdd3p3.n7263 0.108
R10363 vdd3p3.n7263 vdd3p3.n7259 0.108
R10364 vdd3p3.n7259 vdd3p3.n7255 0.108
R10365 vdd3p3.n7255 vdd3p3.n7251 0.108
R10366 vdd3p3.n7251 vdd3p3.n7247 0.108
R10367 vdd3p3.n7247 vdd3p3.n7243 0.108
R10368 vdd3p3.n7243 vdd3p3.n7239 0.108
R10369 vdd3p3.n7239 vdd3p3.n7233 0.108
R10370 vdd3p3.n7233 vdd3p3.n7228 0.108
R10371 vdd3p3.n7228 vdd3p3.n7223 0.108
R10372 vdd3p3.n7223 vdd3p3.n7218 0.108
R10373 vdd3p3.n7218 vdd3p3.n7213 0.108
R10374 vdd3p3.n7213 vdd3p3.n7208 0.108
R10375 vdd3p3.n7208 vdd3p3.n7203 0.108
R10376 vdd3p3.n7203 vdd3p3.n7198 0.108
R10377 vdd3p3.n7198 vdd3p3.n7193 0.108
R10378 vdd3p3.n7193 vdd3p3.n7189 0.108
R10379 vdd3p3.n7189 vdd3p3.n7184 0.108
R10380 vdd3p3.n7184 vdd3p3.n7179 0.108
R10381 vdd3p3.n7179 vdd3p3.n7174 0.108
R10382 vdd3p3.n7174 vdd3p3.n7169 0.108
R10383 vdd3p3.n7169 vdd3p3.n7164 0.108
R10384 vdd3p3.n7164 vdd3p3.n7159 0.108
R10385 vdd3p3.n7159 vdd3p3.n7154 0.108
R10386 vdd3p3.n7154 vdd3p3.n7146 0.108
R10387 vdd3p3.n7146 vdd3p3.n7141 0.108
R10388 vdd3p3.n7141 vdd3p3.n7136 0.108
R10389 vdd3p3.n7136 vdd3p3.n7131 0.108
R10390 vdd3p3.n7131 vdd3p3.n7126 0.108
R10391 vdd3p3.n7126 vdd3p3.n7121 0.108
R10392 vdd3p3.n7121 vdd3p3.n7116 0.108
R10393 vdd3p3.n7116 vdd3p3.n7111 0.108
R10394 vdd3p3.n7111 vdd3p3.n7106 0.108
R10395 vdd3p3.n7106 vdd3p3.n7102 0.108
R10396 vdd3p3.n7102 vdd3p3.n7097 0.108
R10397 vdd3p3.n7097 vdd3p3.n7092 0.108
R10398 vdd3p3.n7092 vdd3p3.n7087 0.108
R10399 vdd3p3.n7087 vdd3p3.n7082 0.108
R10400 vdd3p3.n7082 vdd3p3.n7077 0.108
R10401 vdd3p3.n7077 vdd3p3.n7072 0.108
R10402 vdd3p3.n7072 vdd3p3.n7067 0.108
R10403 vdd3p3.n7067 vdd3p3.n7059 0.108
R10404 vdd3p3.n7059 vdd3p3.n7054 0.108
R10405 vdd3p3.n7054 vdd3p3.n7049 0.108
R10406 vdd3p3.n7049 vdd3p3.n7044 0.108
R10407 vdd3p3.n7044 vdd3p3.n7039 0.108
R10408 vdd3p3.n7039 vdd3p3.n7034 0.108
R10409 vdd3p3.n7034 vdd3p3.n7029 0.108
R10410 vdd3p3.n7029 vdd3p3.n7024 0.108
R10411 vdd3p3.n7016 vdd3p3.n7001 0.108
R10412 vdd3p3.n7001 vdd3p3.n6996 0.108
R10413 vdd3p3.n6996 vdd3p3.n6991 0.108
R10414 vdd3p3.n6991 vdd3p3.n6986 0.108
R10415 vdd3p3.n6986 vdd3p3.n6981 0.108
R10416 vdd3p3.n6981 vdd3p3.n6976 0.108
R10417 vdd3p3.n6976 vdd3p3.n6971 0.108
R10418 vdd3p3.n6971 vdd3p3.n6966 0.108
R10419 vdd3p3.n6966 vdd3p3.n6961 0.108
R10420 vdd3p3.n6961 vdd3p3.n6956 0.108
R10421 vdd3p3.n6956 vdd3p3.n6951 0.108
R10422 vdd3p3.n6951 vdd3p3.n6946 0.108
R10423 vdd3p3.n6946 vdd3p3.n6941 0.108
R10424 vdd3p3.n6941 vdd3p3.n6936 0.108
R10425 vdd3p3.n6936 vdd3p3.n6931 0.108
R10426 vdd3p3.n6931 vdd3p3.n6926 0.108
R10427 vdd3p3.n6926 vdd3p3.n6921 0.108
R10428 vdd3p3.n6921 vdd3p3.n6913 0.108
R10429 vdd3p3.n6913 vdd3p3.n6908 0.108
R10430 vdd3p3.n6908 vdd3p3.n6903 0.108
R10431 vdd3p3.n6903 vdd3p3.n6898 0.108
R10432 vdd3p3.n6898 vdd3p3.n6893 0.108
R10433 vdd3p3.n6893 vdd3p3.n6888 0.108
R10434 vdd3p3.n6888 vdd3p3.n6883 0.108
R10435 vdd3p3.n6883 vdd3p3.n6878 0.108
R10436 vdd3p3.n6878 vdd3p3.n6873 0.108
R10437 vdd3p3.n6873 vdd3p3.n6868 0.108
R10438 vdd3p3.n6868 vdd3p3.n6863 0.108
R10439 vdd3p3.n6863 vdd3p3.n6858 0.108
R10440 vdd3p3.n6858 vdd3p3.n6853 0.108
R10441 vdd3p3.n6853 vdd3p3.n6848 0.108
R10442 vdd3p3.n6848 vdd3p3.n6843 0.108
R10443 vdd3p3.n6843 vdd3p3.n6838 0.108
R10444 vdd3p3.n6838 vdd3p3.n6833 0.108
R10445 vdd3p3.n6833 vdd3p3.n6825 0.108
R10446 vdd3p3.n6825 vdd3p3.n6820 0.108
R10447 vdd3p3.n6820 vdd3p3.n6815 0.108
R10448 vdd3p3.n6815 vdd3p3.n6810 0.108
R10449 vdd3p3.n6810 vdd3p3.n6805 0.108
R10450 vdd3p3.n6805 vdd3p3.n6800 0.108
R10451 vdd3p3.n6800 vdd3p3.n6795 0.108
R10452 vdd3p3.n6795 vdd3p3.n6790 0.108
R10453 vdd3p3.n6790 vdd3p3.n6785 0.108
R10454 vdd3p3.n6785 vdd3p3.n6780 0.108
R10455 vdd3p3.n6780 vdd3p3.n6775 0.108
R10456 vdd3p3.n6775 vdd3p3.n6770 0.108
R10457 vdd3p3.n6770 vdd3p3.n6765 0.108
R10458 vdd3p3.n6765 vdd3p3.n6760 0.108
R10459 vdd3p3.n6760 vdd3p3.n6755 0.108
R10460 vdd3p3.n6755 vdd3p3.n6750 0.108
R10461 vdd3p3.n6750 vdd3p3.n6745 0.108
R10462 vdd3p3.n6745 vdd3p3.n6737 0.108
R10463 vdd3p3.n6737 vdd3p3.n6732 0.108
R10464 vdd3p3.n6732 vdd3p3.n6727 0.108
R10465 vdd3p3.n6727 vdd3p3.n6722 0.108
R10466 vdd3p3.n5355 vdd3p3.n5350 0.108
R10467 vdd3p3.n5360 vdd3p3.n5355 0.108
R10468 vdd3p3.n5365 vdd3p3.n5360 0.108
R10469 vdd3p3.n5370 vdd3p3.n5365 0.108
R10470 vdd3p3.n5375 vdd3p3.n5370 0.108
R10471 vdd3p3.n5380 vdd3p3.n5375 0.108
R10472 vdd3p3.n5385 vdd3p3.n5380 0.108
R10473 vdd3p3.n5390 vdd3p3.n5385 0.108
R10474 vdd3p3.n5395 vdd3p3.n5390 0.108
R10475 vdd3p3.n5400 vdd3p3.n5395 0.108
R10476 vdd3p3.n5405 vdd3p3.n5400 0.108
R10477 vdd3p3.n5413 vdd3p3.n5405 0.108
R10478 vdd3p3.n5418 vdd3p3.n5413 0.108
R10479 vdd3p3.n5423 vdd3p3.n5418 0.108
R10480 vdd3p3.n5428 vdd3p3.n5423 0.108
R10481 vdd3p3.n5433 vdd3p3.n5428 0.108
R10482 vdd3p3.n5438 vdd3p3.n5433 0.108
R10483 vdd3p3.n5443 vdd3p3.n5438 0.108
R10484 vdd3p3.n5448 vdd3p3.n5443 0.108
R10485 vdd3p3.n5453 vdd3p3.n5448 0.108
R10486 vdd3p3.n5458 vdd3p3.n5453 0.108
R10487 vdd3p3.n5463 vdd3p3.n5458 0.108
R10488 vdd3p3.n5468 vdd3p3.n5463 0.108
R10489 vdd3p3.n5473 vdd3p3.n5468 0.108
R10490 vdd3p3.n5478 vdd3p3.n5473 0.108
R10491 vdd3p3.n5483 vdd3p3.n5478 0.108
R10492 vdd3p3.n5488 vdd3p3.n5483 0.108
R10493 vdd3p3.n5493 vdd3p3.n5488 0.108
R10494 vdd3p3.n5501 vdd3p3.n5493 0.108
R10495 vdd3p3.n5506 vdd3p3.n5501 0.108
R10496 vdd3p3.n5511 vdd3p3.n5506 0.108
R10497 vdd3p3.n5516 vdd3p3.n5511 0.108
R10498 vdd3p3.n5521 vdd3p3.n5516 0.108
R10499 vdd3p3.n5526 vdd3p3.n5521 0.108
R10500 vdd3p3.n5531 vdd3p3.n5526 0.108
R10501 vdd3p3.n5536 vdd3p3.n5531 0.108
R10502 vdd3p3.n5541 vdd3p3.n5536 0.108
R10503 vdd3p3.n5546 vdd3p3.n5541 0.108
R10504 vdd3p3.n5551 vdd3p3.n5546 0.108
R10505 vdd3p3.n5556 vdd3p3.n5551 0.108
R10506 vdd3p3.n5561 vdd3p3.n5556 0.108
R10507 vdd3p3.n5566 vdd3p3.n5561 0.108
R10508 vdd3p3.n5571 vdd3p3.n5566 0.108
R10509 vdd3p3.n5576 vdd3p3.n5571 0.108
R10510 vdd3p3.n5581 vdd3p3.n5576 0.108
R10511 vdd3p3.n5589 vdd3p3.n5581 0.108
R10512 vdd3p3.n5594 vdd3p3.n5589 0.108
R10513 vdd3p3.n5599 vdd3p3.n5594 0.108
R10514 vdd3p3.n5604 vdd3p3.n5599 0.108
R10515 vdd3p3.n5609 vdd3p3.n5604 0.108
R10516 vdd3p3.n5614 vdd3p3.n5609 0.108
R10517 vdd3p3.n5619 vdd3p3.n5614 0.108
R10518 vdd3p3.n5624 vdd3p3.n5619 0.108
R10519 vdd3p3.n5629 vdd3p3.n5624 0.108
R10520 vdd3p3.n5634 vdd3p3.n5629 0.108
R10521 vdd3p3.n5639 vdd3p3.n5634 0.108
R10522 vdd3p3.n5644 vdd3p3.n5639 0.108
R10523 vdd3p3.n5649 vdd3p3.n5644 0.108
R10524 vdd3p3.n5654 vdd3p3.n5649 0.108
R10525 vdd3p3.n5659 vdd3p3.n5654 0.108
R10526 vdd3p3.n5664 vdd3p3.n5659 0.108
R10527 vdd3p3.n5669 vdd3p3.n5664 0.108
R10528 vdd3p3.n5677 vdd3p3.n5669 0.108
R10529 vdd3p3.n5682 vdd3p3.n5677 0.108
R10530 vdd3p3.n5687 vdd3p3.n5682 0.108
R10531 vdd3p3.n5692 vdd3p3.n5687 0.108
R10532 vdd3p3.n5697 vdd3p3.n5692 0.108
R10533 vdd3p3.n5702 vdd3p3.n5697 0.108
R10534 vdd3p3.n5707 vdd3p3.n5702 0.108
R10535 vdd3p3.n5712 vdd3p3.n5707 0.108
R10536 vdd3p3.n5717 vdd3p3.n5712 0.108
R10537 vdd3p3.n5722 vdd3p3.n5717 0.108
R10538 vdd3p3.n5727 vdd3p3.n5722 0.108
R10539 vdd3p3.n6398 vdd3p3.n6388 0.108
R10540 vdd3p3.n6388 vdd3p3.n6383 0.108
R10541 vdd3p3.n6383 vdd3p3.n6379 0.108
R10542 vdd3p3.n6379 vdd3p3.n6374 0.108
R10543 vdd3p3.n6374 vdd3p3.n6370 0.108
R10544 vdd3p3.n6370 vdd3p3.n6365 0.108
R10545 vdd3p3.n6365 vdd3p3.n6361 0.108
R10546 vdd3p3.n6361 vdd3p3.n6354 0.108
R10547 vdd3p3.n6354 vdd3p3.n6350 0.108
R10548 vdd3p3.n6350 vdd3p3.n6345 0.108
R10549 vdd3p3.n6345 vdd3p3.n6341 0.108
R10550 vdd3p3.n6341 vdd3p3.n6336 0.108
R10551 vdd3p3.n6336 vdd3p3.n6332 0.108
R10552 vdd3p3.n6332 vdd3p3.n6327 0.108
R10553 vdd3p3.n6327 vdd3p3.n6323 0.108
R10554 vdd3p3.n6323 vdd3p3.n6318 0.108
R10555 vdd3p3.n6318 vdd3p3.n6313 0.108
R10556 vdd3p3.n6313 vdd3p3.n6309 0.108
R10557 vdd3p3.n6309 vdd3p3.n6304 0.108
R10558 vdd3p3.n6304 vdd3p3.n6300 0.108
R10559 vdd3p3.n6300 vdd3p3.n6295 0.108
R10560 vdd3p3.n6295 vdd3p3.n6291 0.108
R10561 vdd3p3.n6291 vdd3p3.n6286 0.108
R10562 vdd3p3.n6286 vdd3p3.n6282 0.108
R10563 vdd3p3.n6282 vdd3p3.n6275 0.108
R10564 vdd3p3.n6275 vdd3p3.n6271 0.108
R10565 vdd3p3.n6271 vdd3p3.n6266 0.108
R10566 vdd3p3.n6266 vdd3p3.n6261 0.108
R10567 vdd3p3.n6261 vdd3p3.n6256 0.108
R10568 vdd3p3.n6256 vdd3p3.n6251 0.108
R10569 vdd3p3.n6251 vdd3p3.n6246 0.108
R10570 vdd3p3.n6246 vdd3p3.n6241 0.108
R10571 vdd3p3.n6241 vdd3p3.n6236 0.108
R10572 vdd3p3.n6236 vdd3p3.n6231 0.108
R10573 vdd3p3.n6231 vdd3p3.n6226 0.108
R10574 vdd3p3.n6226 vdd3p3.n6221 0.108
R10575 vdd3p3.n6221 vdd3p3.n6216 0.108
R10576 vdd3p3.n6216 vdd3p3.n6211 0.108
R10577 vdd3p3.n6211 vdd3p3.n6206 0.108
R10578 vdd3p3.n6206 vdd3p3.n6201 0.108
R10579 vdd3p3.n6201 vdd3p3.n6196 0.108
R10580 vdd3p3.n6196 vdd3p3.n6188 0.108
R10581 vdd3p3.n6188 vdd3p3.n6183 0.108
R10582 vdd3p3.n6183 vdd3p3.n6178 0.108
R10583 vdd3p3.n6178 vdd3p3.n6173 0.108
R10584 vdd3p3.n6173 vdd3p3.n6168 0.108
R10585 vdd3p3.n6168 vdd3p3.n6163 0.108
R10586 vdd3p3.n6163 vdd3p3.n6158 0.108
R10587 vdd3p3.n6158 vdd3p3.n6153 0.108
R10588 vdd3p3.n6153 vdd3p3.n6148 0.108
R10589 vdd3p3.n6148 vdd3p3.n6143 0.108
R10590 vdd3p3.n6143 vdd3p3.n6138 0.108
R10591 vdd3p3.n6138 vdd3p3.n6133 0.108
R10592 vdd3p3.n6133 vdd3p3.n6128 0.108
R10593 vdd3p3.n6128 vdd3p3.n6123 0.108
R10594 vdd3p3.n6123 vdd3p3.n6118 0.108
R10595 vdd3p3.n6118 vdd3p3.n6114 0.108
R10596 vdd3p3.n6114 vdd3p3.n6110 0.108
R10597 vdd3p3.n6110 vdd3p3.n6104 0.108
R10598 vdd3p3.n6104 vdd3p3.n6100 0.108
R10599 vdd3p3.n6100 vdd3p3.n6096 0.108
R10600 vdd3p3.n6096 vdd3p3.n6092 0.108
R10601 vdd3p3.n6092 vdd3p3.n6088 0.108
R10602 vdd3p3.n6088 vdd3p3.n6084 0.108
R10603 vdd3p3.n6084 vdd3p3.n6080 0.108
R10604 vdd3p3.n6080 vdd3p3.n6076 0.108
R10605 vdd3p3.n6076 vdd3p3.n6072 0.108
R10606 vdd3p3.n6072 vdd3p3.n6068 0.108
R10607 vdd3p3.n6068 vdd3p3.n6064 0.108
R10608 vdd3p3.n6064 vdd3p3.n6060 0.108
R10609 vdd3p3.n6060 vdd3p3.n6056 0.108
R10610 vdd3p3.n6056 vdd3p3.n6052 0.108
R10611 vdd3p3.n6052 vdd3p3.n6048 0.108
R10612 vdd3p3.n6048 vdd3p3.n6044 0.108
R10613 vdd3p3.n6044 vdd3p3.n6040 0.108
R10614 vdd3p3.n6040 vdd3p3.n6034 0.108
R10615 vdd3p3.n6034 vdd3p3.n6030 0.108
R10616 vdd3p3.n6030 vdd3p3.n6026 0.108
R10617 vdd3p3.n6026 vdd3p3.n6022 0.108
R10618 vdd3p3.n6022 vdd3p3.n6018 0.108
R10619 vdd3p3.n6018 vdd3p3.n6014 0.108
R10620 vdd3p3.n6014 vdd3p3.n6010 0.108
R10621 vdd3p3.n6010 vdd3p3.n6006 0.108
R10622 vdd3p3.n6006 vdd3p3.n6002 0.108
R10623 vdd3p3.n6002 vdd3p3.n5998 0.108
R10624 vdd3p3.n5998 vdd3p3.n5994 0.108
R10625 vdd3p3.n5994 vdd3p3.n5990 0.108
R10626 vdd3p3.n5990 vdd3p3.n5986 0.108
R10627 vdd3p3.n5986 vdd3p3.n5982 0.108
R10628 vdd3p3.n5982 vdd3p3.n5978 0.108
R10629 vdd3p3.n5978 vdd3p3.n5974 0.108
R10630 vdd3p3.n5974 vdd3p3.n5970 0.108
R10631 vdd3p3.n5970 vdd3p3.n5964 0.108
R10632 vdd3p3.n5964 vdd3p3.n5960 0.108
R10633 vdd3p3.n5960 vdd3p3.n5956 0.108
R10634 vdd3p3.n5956 vdd3p3.n5952 0.108
R10635 vdd3p3.n5952 vdd3p3.n5947 0.108
R10636 vdd3p3.n5947 vdd3p3.n5942 0.108
R10637 vdd3p3.n5942 vdd3p3.n5937 0.108
R10638 vdd3p3.n5937 vdd3p3.n5932 0.108
R10639 vdd3p3.n5932 vdd3p3.n5927 0.108
R10640 vdd3p3.n5927 vdd3p3.n5922 0.108
R10641 vdd3p3.n5922 vdd3p3.n5917 0.108
R10642 vdd3p3.n5917 vdd3p3.n5912 0.108
R10643 vdd3p3.n5912 vdd3p3.n5907 0.108
R10644 vdd3p3.n5907 vdd3p3.n5902 0.108
R10645 vdd3p3.n5902 vdd3p3.n5897 0.108
R10646 vdd3p3.n5897 vdd3p3.n5892 0.108
R10647 vdd3p3.n5892 vdd3p3.n5887 0.108
R10648 vdd3p3.n5887 vdd3p3.n5879 0.108
R10649 vdd3p3.n5879 vdd3p3.n5874 0.108
R10650 vdd3p3.n5874 vdd3p3.n5869 0.108
R10651 vdd3p3.n5869 vdd3p3.n5864 0.108
R10652 vdd3p3.n5864 vdd3p3.n5859 0.108
R10653 vdd3p3.n5859 vdd3p3.n5854 0.108
R10654 vdd3p3.n5854 vdd3p3.n5849 0.108
R10655 vdd3p3.n5849 vdd3p3.n5844 0.108
R10656 vdd3p3.n5844 vdd3p3.n5839 0.108
R10657 vdd3p3.n5839 vdd3p3.n5834 0.108
R10658 vdd3p3.n5834 vdd3p3.n5829 0.108
R10659 vdd3p3.n5829 vdd3p3.n5824 0.108
R10660 vdd3p3.n5824 vdd3p3.n5819 0.108
R10661 vdd3p3.n5819 vdd3p3.n5814 0.108
R10662 vdd3p3.n5814 vdd3p3.n5809 0.108
R10663 vdd3p3.n5809 vdd3p3.n5804 0.108
R10664 vdd3p3.n5804 vdd3p3.n5799 0.108
R10665 vdd3p3.n5799 vdd3p3.n5791 0.108
R10666 vdd3p3.n5791 vdd3p3.n5786 0.108
R10667 vdd3p3.n5786 vdd3p3.n5781 0.108
R10668 vdd3p3.n5781 vdd3p3.n5776 0.108
R10669 vdd3p3.n5776 vdd3p3.n5771 0.108
R10670 vdd3p3.n5771 vdd3p3.n5766 0.108
R10671 vdd3p3.n5766 vdd3p3.n5761 0.108
R10672 vdd3p3.n5761 vdd3p3.n5756 0.108
R10673 vdd3p3.n5756 vdd3p3.n5751 0.108
R10674 vdd3p3.n5751 vdd3p3.n5746 0.108
R10675 vdd3p3.n5746 vdd3p3.n5741 0.108
R10676 vdd3p3.n6716 vdd3p3.n6715 0.108
R10677 vdd3p3.n6715 vdd3p3.n6711 0.108
R10678 vdd3p3.n6711 vdd3p3.n6707 0.108
R10679 vdd3p3.n6707 vdd3p3.n6703 0.108
R10680 vdd3p3.n6703 vdd3p3.n6699 0.108
R10681 vdd3p3.n6699 vdd3p3.n6695 0.108
R10682 vdd3p3.n6695 vdd3p3.n6690 0.108
R10683 vdd3p3.n6690 vdd3p3.n6685 0.108
R10684 vdd3p3.n6685 vdd3p3.n6677 0.108
R10685 vdd3p3.n6677 vdd3p3.n6672 0.108
R10686 vdd3p3.n6672 vdd3p3.n6667 0.108
R10687 vdd3p3.n6667 vdd3p3.n6662 0.108
R10688 vdd3p3.n6662 vdd3p3.n6657 0.108
R10689 vdd3p3.n6657 vdd3p3.n6652 0.108
R10690 vdd3p3.n6652 vdd3p3.n6647 0.108
R10691 vdd3p3.n6647 vdd3p3.n6642 0.108
R10692 vdd3p3.n6642 vdd3p3.n6637 0.108
R10693 vdd3p3.n6637 vdd3p3.n6632 0.108
R10694 vdd3p3.n6632 vdd3p3.n6627 0.108
R10695 vdd3p3.n6627 vdd3p3.n6622 0.108
R10696 vdd3p3.n6622 vdd3p3.n6617 0.108
R10697 vdd3p3.n6617 vdd3p3.n6612 0.108
R10698 vdd3p3.n6612 vdd3p3.n6607 0.108
R10699 vdd3p3.n6607 vdd3p3.n6602 0.108
R10700 vdd3p3.n6602 vdd3p3.n6597 0.108
R10701 vdd3p3.n6597 vdd3p3.n6589 0.108
R10702 vdd3p3.n6589 vdd3p3.n6585 0.108
R10703 vdd3p3.n6585 vdd3p3.n6581 0.108
R10704 vdd3p3.n6581 vdd3p3.n6577 0.108
R10705 vdd3p3.n6577 vdd3p3.n6573 0.108
R10706 vdd3p3.n6573 vdd3p3.n6569 0.108
R10707 vdd3p3.n6569 vdd3p3.n6565 0.108
R10708 vdd3p3.n6565 vdd3p3.n6548 0.108
R10709 vdd3p3.n6548 vdd3p3.n6544 0.108
R10710 vdd3p3.n6544 vdd3p3.n6540 0.108
R10711 vdd3p3.n6540 vdd3p3.n6536 0.108
R10712 vdd3p3.n6536 vdd3p3.n6532 0.108
R10713 vdd3p3.n6532 vdd3p3.n6528 0.108
R10714 vdd3p3.n6528 vdd3p3.n6524 0.108
R10715 vdd3p3.n6524 vdd3p3.n6519 0.108
R10716 vdd3p3.n6519 vdd3p3.n6514 0.108
R10717 vdd3p3.n6514 vdd3p3.n6509 0.108
R10718 vdd3p3.n6509 vdd3p3.n6501 0.108
R10719 vdd3p3.n6501 vdd3p3.n6496 0.108
R10720 vdd3p3.n6496 vdd3p3.n6491 0.108
R10721 vdd3p3.n6491 vdd3p3.n6486 0.108
R10722 vdd3p3.n6486 vdd3p3.n6481 0.108
R10723 vdd3p3.n6481 vdd3p3.n6476 0.108
R10724 vdd3p3.n6476 vdd3p3.n6471 0.108
R10725 vdd3p3.n6471 vdd3p3.n6466 0.108
R10726 vdd3p3.n6466 vdd3p3.n6461 0.108
R10727 vdd3p3.n6461 vdd3p3.n6456 0.108
R10728 vdd3p3.n6456 vdd3p3.n6451 0.108
R10729 vdd3p3.n6451 vdd3p3.n6446 0.108
R10730 vdd3p3.n6446 vdd3p3.n6441 0.108
R10731 vdd3p3.n6441 vdd3p3.n6436 0.108
R10732 vdd3p3.n6436 vdd3p3.n6431 0.108
R10733 vdd3p3.n6431 vdd3p3.n6426 0.108
R10734 vdd3p3.n6426 vdd3p3.n6421 0.108
R10735 vdd3p3.n6421 vdd3p3.n6415 0.108
R10736 vdd3p3.n6415 vdd3p3.n6411 0.108
R10737 vdd3p3.n6411 vdd3p3.n6407 0.108
R10738 vdd3p3.n6407 vdd3p3.n6403 0.108
R10739 vdd3p3.n6403 vdd3p3.n6401 0.108
R10740 vdd3p3.n6401 vdd3p3.n6400 0.108
R10741 vdd3p3.n6400 vdd3p3.n6399 0.108
R10742 vdd3p3.n7957 vdd3p3.n7949 0.108
R10743 vdd3p3.n7965 vdd3p3.n7957 0.108
R10744 vdd3p3.n7973 vdd3p3.n7965 0.108
R10745 vdd3p3.n7981 vdd3p3.n7973 0.108
R10746 vdd3p3.n7989 vdd3p3.n7981 0.108
R10747 vdd3p3.n7995 vdd3p3.n7989 0.108
R10748 vdd3p3.n8003 vdd3p3.n7995 0.108
R10749 vdd3p3.n8009 vdd3p3.n8003 0.108
R10750 vdd3p3.n8017 vdd3p3.n8009 0.108
R10751 vdd3p3.n8024 vdd3p3.n8017 0.108
R10752 vdd3p3.n8033 vdd3p3.n8024 0.108
R10753 vdd3p3.n8038 vdd3p3.n8033 0.108
R10754 vdd3p3.n8044 vdd3p3.n8038 0.108
R10755 vdd3p3.n8050 vdd3p3.n8044 0.108
R10756 vdd3p3.n8056 vdd3p3.n8050 0.108
R10757 vdd3p3.n8062 vdd3p3.n8056 0.108
R10758 vdd3p3.n8068 vdd3p3.n8062 0.108
R10759 vdd3p3.n8074 vdd3p3.n8068 0.108
R10760 vdd3p3.n8082 vdd3p3.n8074 0.108
R10761 vdd3p3.n8088 vdd3p3.n8082 0.108
R10762 vdd3p3.n8096 vdd3p3.n8088 0.108
R10763 vdd3p3.n8102 vdd3p3.n8096 0.108
R10764 vdd3p3.n8108 vdd3p3.n8102 0.108
R10765 vdd3p3.n8114 vdd3p3.n8108 0.108
R10766 vdd3p3.n8120 vdd3p3.n8114 0.108
R10767 vdd3p3.n8126 vdd3p3.n8120 0.108
R10768 vdd3p3.n8132 vdd3p3.n8126 0.108
R10769 vdd3p3.n8138 vdd3p3.n8132 0.108
R10770 vdd3p3.n8143 vdd3p3.n8138 0.108
R10771 vdd3p3.n8149 vdd3p3.n8143 0.108
R10772 vdd3p3.n8155 vdd3p3.n8149 0.108
R10773 vdd3p3.n8161 vdd3p3.n8155 0.108
R10774 vdd3p3.n8167 vdd3p3.n8161 0.108
R10775 vdd3p3.n8173 vdd3p3.n8167 0.108
R10776 vdd3p3.n8179 vdd3p3.n8173 0.108
R10777 vdd3p3.n8187 vdd3p3.n8179 0.108
R10778 vdd3p3.n8193 vdd3p3.n8187 0.108
R10779 vdd3p3.n8201 vdd3p3.n8193 0.108
R10780 vdd3p3.n8207 vdd3p3.n8201 0.108
R10781 vdd3p3.n8213 vdd3p3.n8207 0.108
R10782 vdd3p3.n8219 vdd3p3.n8213 0.108
R10783 vdd3p3.n8225 vdd3p3.n8219 0.108
R10784 vdd3p3.n8231 vdd3p3.n8225 0.108
R10785 vdd3p3.n8237 vdd3p3.n8231 0.108
R10786 vdd3p3.n8243 vdd3p3.n8237 0.108
R10787 vdd3p3.n8248 vdd3p3.n8243 0.108
R10788 vdd3p3.n8254 vdd3p3.n8248 0.108
R10789 vdd3p3.n8260 vdd3p3.n8254 0.108
R10790 vdd3p3.n8266 vdd3p3.n8260 0.108
R10791 vdd3p3.n8272 vdd3p3.n8266 0.108
R10792 vdd3p3.n8278 vdd3p3.n8272 0.108
R10793 vdd3p3.n8284 vdd3p3.n8278 0.108
R10794 vdd3p3.n8292 vdd3p3.n8284 0.108
R10795 vdd3p3.n8298 vdd3p3.n8292 0.108
R10796 vdd3p3.n8310 vdd3p3.n8298 0.108
R10797 vdd3p3.n8320 vdd3p3.n8310 0.108
R10798 vdd3p3.n8330 vdd3p3.n8320 0.108
R10799 vdd3p3.n8340 vdd3p3.n8330 0.108
R10800 vdd3p3.n8350 vdd3p3.n8340 0.108
R10801 vdd3p3.n8359 vdd3p3.n8350 0.108
R10802 vdd3p3.n8368 vdd3p3.n8359 0.108
R10803 vdd3p3.n8377 vdd3p3.n8368 0.108
R10804 vdd3p3.n8385 vdd3p3.n8377 0.108
R10805 vdd3p3.n8394 vdd3p3.n8385 0.108
R10806 vdd3p3.n8403 vdd3p3.n8394 0.108
R10807 vdd3p3.n8412 vdd3p3.n8403 0.108
R10808 vdd3p3.n8420 vdd3p3.n8412 0.108
R10809 vdd3p3.n8428 vdd3p3.n8420 0.108
R10810 vdd3p3.n8434 vdd3p3.n8428 0.108
R10811 vdd3p3.n8435 vdd3p3.n8434 0.108
R10812 vdd3p3.n8436 vdd3p3.n8435 0.108
R10813 vdd3p3.n4732 vdd3p3.n4731 0.107
R10814 vdd3p3.n3341 vdd3p3.n3340 0.107
R10815 vdd3p3.n2495 vdd3p3.n2494 0.107
R10816 vdd3p3.n1650 vdd3p3.n1649 0.107
R10817 vdd3p3.n804 vdd3p3.n803 0.107
R10818 vdd3p3.n4227 vdd3p3.n4226 0.098
R10819 vdd3p3.n4349 vdd3p3.n4348 0.098
R10820 vdd3p3.n4669 vdd3p3.n4668 0.098
R10821 vdd3p3.n5079 vdd3p3.n5078 0.098
R10822 vdd3p3.n3465 vdd3p3.n3462 0.095
R10823 vdd3p3.n4165 vdd3p3.n4164 0.095
R10824 vdd3p3.n8741 vdd3p3.n8740 0.092
R10825 vdd3p3.n42 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.091
R10826 vdd3p3.n1733 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VPWR 0.091
R10827 vdd3p3.n4169 vdd3p3.n4168 0.089
R10828 vdd3p3.n8823 vdd3p3.n8822 0.089
R10829 vdd3p3.n3997 vdd3p3.n3991 0.088
R10830 vdd3p3.n5000 vdd3p3.n4999 0.085
R10831 vdd3p3.n3799 vdd3p3.n3798 0.082
R10832 vdd3p3.n3796 vdd3p3.n3795 0.082
R10833 comparator_top_0.comparator_0.VDD vdd3p3.n5034 0.073
R10834 vdd3p3.n3450 vdd3p3.n3440 0.072
R10835 vdd3p3.n6322 vdd3p3.n6321 0.072
R10836 vdd3p3.n6240 vdd3p3.n6239 0.072
R10837 vdd3p3.n6152 vdd3p3.n6151 0.072
R10838 vdd3p3.n6075 vdd3p3.n6074 0.072
R10839 vdd3p3.n6005 vdd3p3.n6004 0.072
R10840 vdd3p3.n5931 vdd3p3.n5930 0.072
R10841 vdd3p3.n5843 vdd3p3.n5842 0.072
R10842 vdd3p3.n5755 vdd3p3.n5754 0.072
R10843 vdd3p3.n5344 vdd3p3.n5343 0.071
R10844 vdd3p3.n3763 vdd3p3.n3762 0.07
R10845 vdd3p3.n3512 vdd3p3.n3511 0.07
R10846 vdd3p3.n7486 vdd3p3.n7485 0.069
R10847 vdd3p3.n3378 vdd3p3.n3377 0.068
R10848 vdd3p3.n2532 vdd3p3.n2531 0.068
R10849 vdd3p3.n1687 vdd3p3.n1686 0.068
R10850 vdd3p3.n841 vdd3p3.n840 0.068
R10851 vdd3p3.n3482 vdd3p3.n3481 0.067
R10852 vdd3p3.n8023 vdd3p3.n8022 0.067
R10853 vdd3p3.n8131 vdd3p3.n8130 0.067
R10854 vdd3p3.n8236 vdd3p3.n8235 0.067
R10855 vdd3p3.n8367 vdd3p3.n8366 0.067
R10856 vdd3p3.n4964 vdd3p3.n4963 0.067
R10857 vdd3p3.n8747 comparator_top_0.comparator_bias_0.VDD 0.064
R10858 vdd3p3.n3377 vdd3p3.n3376 0.063
R10859 vdd3p3.n2531 vdd3p3.n2530 0.063
R10860 vdd3p3.n1686 vdd3p3.n1685 0.063
R10861 vdd3p3.n840 vdd3p3.n839 0.063
R10862 vdd3p3.n7934 vdd3p3.n7930 0.063
R10863 vdd3p3.n7923 vdd3p3.n7922 0.063
R10864 vdd3p3.n7789 vdd3p3.n7785 0.063
R10865 vdd3p3.n7781 vdd3p3.n7780 0.063
R10866 vdd3p3.n7657 vdd3p3.n7653 0.063
R10867 vdd3p3.n7649 vdd3p3.n7648 0.063
R10868 vdd3p3.n5029 vdd3p3.n5028 0.062
R10869 vdd3p3.n4402 vdd3p3.n4396 0.061
R10870 vdd3p3.n4492 vdd3p3.n4486 0.061
R10871 vdd3p3.n5105 vdd3p3.n5096 0.061
R10872 vdd3p3.n4690 vdd3p3.n4682 0.061
R10873 vdd3p3.n4462 vdd3p3.n4456 0.061
R10874 vdd3p3.n4245 vdd3p3.n4236 0.061
R10875 vdd3p3.n4368 vdd3p3.n4362 0.061
R10876 vdd3p3.n4432 vdd3p3.n4426 0.061
R10877 vdd3p3.n4522 vdd3p3.n4516 0.061
R10878 vdd3p3.n43 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd3p3 0.06
R10879 vdd3p3.n1734 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd3p3 0.06
R10880 vdd3p3.n3687 vdd3p3.n3682 0.059
R10881 vdd3p3.n3593 vdd3p3.n3588 0.059
R10882 vdd3p3.n3506 vdd3p3.n3498 0.059
R10883 vdd3p3.n4822 vdd3p3.n4817 0.059
R10884 vdd3p3.n3458 vdd3p3.n3457 0.059
R10885 vdd3p3.n8528 vdd3p3.n8527 0.059
R10886 vdd3p3.n3599 vdd3p3.n3598 0.059
R10887 vdd3p3.n3693 vdd3p3.n3692 0.058
R10888 vdd3p3.n4828 vdd3p3.n4827 0.058
R10889 vdd3p3.n8798 vdd3p3.n8790 0.058
R10890 vdd3p3.n8584 vdd3p3.n8580 0.058
R10891 vdd3p3.n4988 vdd3p3.n4980 0.058
R10892 vdd3p3.n8743 vdd3p3.n8738 0.057
R10893 vdd3p3.n3438 vdd3p3.n3430 0.056
R10894 vdd3p3.n23 vdd3p3.n22 0.056
R10895 vdd3p3.n24 vdd3p3.n23 0.056
R10896 vdd3p3.n24 vdd3p3.n1 0.056
R10897 vdd3p3.n60 vdd3p3.n1 0.056
R10898 vdd3p3.n862 vdd3p3.n854 0.056
R10899 vdd3p3.n873 vdd3p3.n854 0.056
R10900 vdd3p3.n875 vdd3p3.n873 0.056
R10901 vdd3p3.n875 vdd3p3.n874 0.056
R10902 vdd3p3.n1714 vdd3p3.n1713 0.056
R10903 vdd3p3.n1715 vdd3p3.n1714 0.056
R10904 vdd3p3.n1715 vdd3p3.n1692 0.056
R10905 vdd3p3.n1751 vdd3p3.n1692 0.056
R10906 vdd3p3.n2553 vdd3p3.n2545 0.056
R10907 vdd3p3.n2564 vdd3p3.n2545 0.056
R10908 vdd3p3.n2566 vdd3p3.n2564 0.056
R10909 vdd3p3.n2566 vdd3p3.n2565 0.056
R10910 comparator_top_0.comparator_bias_0.VDD vdd3p3.n8746 0.056
R10911 vdd3p3.n4233 vdd3p3.n4232 0.055
R10912 vdd3p3.n4355 vdd3p3.n4354 0.055
R10913 vdd3p3.n4393 vdd3p3.n4392 0.055
R10914 vdd3p3.n4423 vdd3p3.n4422 0.055
R10915 vdd3p3.n4453 vdd3p3.n4452 0.055
R10916 vdd3p3.n4483 vdd3p3.n4482 0.055
R10917 vdd3p3.n4513 vdd3p3.n4512 0.055
R10918 vdd3p3.n4570 vdd3p3.n4569 0.055
R10919 vdd3p3.n4675 vdd3p3.n4674 0.055
R10920 vdd3p3.n5093 vdd3p3.n5092 0.055
R10921 vdd3p3.n5015 vdd3p3.n5014 0.055
R10922 vdd3p3.n4759 vdd3p3.n4758 0.055
R10923 vdd3p3.n4994 vdd3p3.n4993 0.054
R10924 vdd3p3.n8522 vdd3p3.n8521 0.053
R10925 vdd3p3.n8866 vdd3p3.n8865 0.053
R10926 vdd3p3.n8777 vdd3p3.n8776 0.053
R10927 EF_AMUX21m_1.array_1ls_1tgm_1.vdd3p3 vdd3p3.n3381 0.052
R10928 EF_AMUX21m_2.array_1ls_1tgm_1.vdd3p3 vdd3p3.n1690 0.051
R10929 vdd3p3.n8437 vdd3p3.n8436 0.051
R10930 vdd3p3.n3997 vdd3p3.n3996 0.051
R10931 vdd3p3.n4169 vdd3p3.n4161 0.051
R10932 vdd3p3.n3987 vdd3p3.n3986 0.05
R10933 vdd3p3.n3836 vdd3p3.n3835 0.048
R10934 vdd3p3.n3381 vdd3p3.n3380 0.047
R10935 vdd3p3.n4232 vdd3p3.n4231 0.047
R10936 vdd3p3.n4354 vdd3p3.n4353 0.047
R10937 vdd3p3.n4392 vdd3p3.n4391 0.047
R10938 vdd3p3.n4422 vdd3p3.n4421 0.047
R10939 vdd3p3.n4452 vdd3p3.n4451 0.047
R10940 vdd3p3.n4482 vdd3p3.n4481 0.047
R10941 vdd3p3.n4512 vdd3p3.n4511 0.047
R10942 vdd3p3.n4674 vdd3p3.n4673 0.047
R10943 vdd3p3.n5092 vdd3p3.n5091 0.047
R10944 EF_AMUX21m_2.array_1ls_1tgm_0.vdd3p3 vdd3p3.n844 0.047
R10945 EF_AMUX21m_1.array_1ls_1tgm_0.vdd3p3 vdd3p3.n2535 0.047
R10946 vdd3p3.n1690 vdd3p3.n1689 0.047
R10947 vdd3p3.n3438 vdd3p3.n3437 0.046
R10948 vdd3p3.n4855 vdd3p3.n4854 0.046
R10949 vdd3p3.n3757 vdd3p3.n3752 0.045
R10950 vdd3p3.n8557 vdd3p3.n8539 0.045
R10951 vdd3p3.n8819 vdd3p3.n8801 0.045
R10952 vdd3p3.n19 vdd3p3.n14 0.045
R10953 vdd3p3.n863 vdd3p3.n859 0.045
R10954 vdd3p3.n1710 vdd3p3.n1705 0.045
R10955 vdd3p3.n2554 vdd3p3.n2550 0.045
R10956 vdd3p3.n4841 vdd3p3.n4840 0.045
R10957 vdd3p3.n4753 vdd3p3.n4748 0.045
R10958 vdd3p3.n8601 vdd3p3.n8587 0.045
R10959 vdd3p3.n8636 vdd3p3.n8618 0.045
R10960 vdd3p3.n8882 vdd3p3.n8871 0.045
R10961 vdd3p3.n8636 vdd3p3.n8635 0.044
R10962 vdd3p3.n8601 vdd3p3.n8600 0.044
R10963 vdd3p3.n4748 vdd3p3.n4747 0.044
R10964 vdd3p3.n844 vdd3p3.n843 0.044
R10965 vdd3p3.n2535 vdd3p3.n2534 0.044
R10966 vdd3p3.n3752 vdd3p3.n3751 0.044
R10967 vdd3p3.n8557 vdd3p3.n8556 0.044
R10968 vdd3p3.n8819 vdd3p3.n8818 0.044
R10969 vdd3p3.n3873 vdd3p3.n3809 0.044
R10970 vdd3p3.n3806 vdd3p3.n3805 0.044
R10971 vdd3p3.n3802 vdd3p3.n3801 0.044
R10972 vdd3p3.n4168 vdd3p3.n4165 0.044
R10973 vdd3p3.n8828 vdd3p3.n8827 0.044
R10974 vdd3p3.n3465 vdd3p3.n3464 0.044
R10975 vdd3p3.n8882 vdd3p3.n8881 0.044
R10976 vdd3p3.n5123 vdd3p3.n5122 0.043
R10977 vdd3p3.n20 vdd3p3.n9 0.043
R10978 vdd3p3.n860 vdd3p3.n855 0.043
R10979 vdd3p3.n1711 vdd3p3.n1700 0.043
R10980 vdd3p3.n2551 vdd3p3.n2546 0.043
R10981 vdd3p3.n4204 vdd3p3.n4202 0.043
R10982 vdd3p3.n4334 vdd3p3.n4332 0.043
R10983 vdd3p3.n4326 vdd3p3.n4324 0.043
R10984 vdd3p3.n4654 vdd3p3.n4652 0.043
R10985 vdd3p3.n4646 vdd3p3.n4644 0.043
R10986 vdd3p3.n5056 vdd3p3.n5054 0.043
R10987 vdd3p3.n3481 vdd3p3.n3479 0.043
R10988 vdd3p3.n4963 vdd3p3.n4961 0.043
R10989 vdd3p3.n8510 vdd3p3.n8508 0.043
R10990 vdd3p3.n8854 vdd3p3.n8852 0.043
R10991 vdd3p3.n8765 vdd3p3.n8763 0.043
R10992 vdd3p3.n8700 vdd3p3.n8699 0.042
R10993 vdd3p3.n8827 vdd3p3.n8826 0.042
R10994 vdd3p3.n8738 vdd3p3.n8700 0.042
R10995 vdd3p3.n4835 vdd3p3.n4834 0.042
R10996 vdd3p3.n4836 vdd3p3.n4835 0.042
R10997 vdd3p3.n4837 vdd3p3.n4836 0.042
R10998 vdd3p3.n4840 vdd3p3.n4839 0.042
R10999 vdd3p3.n4839 vdd3p3.n4838 0.042
R11000 vdd3p3.n4890 vdd3p3.n4889 0.042
R11001 vdd3p3.n4891 vdd3p3.n4890 0.042
R11002 vdd3p3.n4892 vdd3p3.n4891 0.042
R11003 vdd3p3.n4895 vdd3p3.n4894 0.042
R11004 vdd3p3.n4896 vdd3p3.n4895 0.042
R11005 vdd3p3.n4897 vdd3p3.n4896 0.042
R11006 vdd3p3.n8607 vdd3p3.n8606 0.042
R11007 vdd3p3.n8608 vdd3p3.n8607 0.042
R11008 vdd3p3.n8609 vdd3p3.n8608 0.042
R11009 vdd3p3.n8610 vdd3p3.n8609 0.042
R11010 vdd3p3.n8613 vdd3p3.n8612 0.042
R11011 vdd3p3.n8614 vdd3p3.n8613 0.042
R11012 vdd3p3.n8615 vdd3p3.n8614 0.042
R11013 vdd3p3.n8887 vdd3p3.n8615 0.042
R11014 vdd3p3.n8887 vdd3p3.n8886 0.042
R11015 vdd3p3.n8830 vdd3p3.n8829 0.042
R11016 vdd3p3.n8829 vdd3p3.n8828 0.042
R11017 vdd3p3.n8826 vdd3p3.n8825 0.042
R11018 vdd3p3.n8825 vdd3p3.n8824 0.042
R11019 vdd3p3.n5341 vdd3p3.n5340 0.042
R11020 vdd3p3.n6636 vdd3p3.n6635 0.042
R11021 vdd3p3.n6543 vdd3p3.n6542 0.042
R11022 vdd3p3.n6460 vdd3p3.n6459 0.042
R11023 vdd3p3.n3854 vdd3p3.n3853 0.042
R11024 vdd3p3.n3803 vdd3p3.n3802 0.042
R11025 vdd3p3.n4528 vdd3p3.n4527 0.042
R11026 vdd3p3.n4529 vdd3p3.n4528 0.042
R11027 vdd3p3.n4530 vdd3p3.n4529 0.042
R11028 vdd3p3.n4531 vdd3p3.n4530 0.042
R11029 vdd3p3.n4534 vdd3p3.n4533 0.042
R11030 vdd3p3.n4535 vdd3p3.n4534 0.042
R11031 vdd3p3.n4536 vdd3p3.n4535 0.042
R11032 vdd3p3.n4537 vdd3p3.n4536 0.042
R11033 vdd3p3.n4538 vdd3p3.n4537 0.042
R11034 vdd3p3.n4547 vdd3p3.n4544 0.042
R11035 vdd3p3.n4547 vdd3p3.n4546 0.042
R11036 vdd3p3.n4546 vdd3p3.n4545 0.042
R11037 vdd3p3.n4555 vdd3p3.n4554 0.042
R11038 vdd3p3.n4556 vdd3p3.n4555 0.042
R11039 vdd3p3.n5142 vdd3p3.n4556 0.042
R11040 vdd3p3.n5142 vdd3p3.n5141 0.042
R11041 vdd3p3.n5141 vdd3p3.n5140 0.042
R11042 vdd3p3.n5140 vdd3p3.n5139 0.042
R11043 vdd3p3.n5139 vdd3p3.n5138 0.042
R11044 vdd3p3.n5138 vdd3p3.n5137 0.042
R11045 vdd3p3.n5137 vdd3p3.n5136 0.042
R11046 vdd3p3.n5136 vdd3p3.n5135 0.042
R11047 vdd3p3.n4841 vdd3p3.n4837 0.042
R11048 vdd3p3.n3744 vdd3p3.n3740 0.042
R11049 vdd3p3.n3580 vdd3p3.n3576 0.042
R11050 vdd3p3.n8523 vdd3p3.n8522 0.042
R11051 vdd3p3.n8575 vdd3p3.n8572 0.042
R11052 vdd3p3.n8867 vdd3p3.n8866 0.042
R11053 vdd3p3.n8785 vdd3p3.n8777 0.042
R11054 vdd3p3.n3515 vdd3p3.n3514 0.042
R11055 vdd3p3.n3602 vdd3p3.n3601 0.042
R11056 vdd3p3.n3696 vdd3p3.n3695 0.042
R11057 vdd3p3.n4764 vdd3p3.n4763 0.042
R11058 vdd3p3.n4570 vdd3p3.n4567 0.041
R11059 vdd3p3.n4432 vdd3p3.n4431 0.041
R11060 vdd3p3.n4522 vdd3p3.n4521 0.041
R11061 vdd3p3.n3859 vdd3p3.n3855 0.041
R11062 vdd3p3.n3848 vdd3p3.n3847 0.041
R11063 vdd3p3.n3805 vdd3p3.n3804 0.041
R11064 vdd3p3.n4402 vdd3p3.n4401 0.041
R11065 vdd3p3.n4492 vdd3p3.n4491 0.041
R11066 vdd3p3.n5105 vdd3p3.n5104 0.041
R11067 vdd3p3.n4245 vdd3p3.n4244 0.041
R11068 vdd3p3.n4368 vdd3p3.n4367 0.041
R11069 vdd3p3.n4462 vdd3p3.n4461 0.041
R11070 vdd3p3.n4690 vdd3p3.n4689 0.041
R11071 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd3p3 vdd3p3.n905 0.04
R11072 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd3p3 vdd3p3.n2596 0.04
R11073 vdd3p3.n4267 vdd3p3.n4265 0.04
R11074 vdd3p3.n4283 vdd3p3.n4281 0.04
R11075 vdd3p3.n4587 vdd3p3.n4585 0.04
R11076 vdd3p3.n4603 vdd3p3.n4601 0.04
R11077 vdd3p3.n3529 vdd3p3.n3527 0.04
R11078 vdd3p3.n3545 vdd3p3.n3543 0.04
R11079 vdd3p3.n3614 vdd3p3.n3612 0.04
R11080 vdd3p3.n3642 vdd3p3.n3640 0.04
R11081 vdd3p3.n3621 vdd3p3.n3619 0.04
R11082 vdd3p3.n3713 vdd3p3.n3711 0.04
R11083 vdd3p3.n4778 vdd3p3.n4776 0.04
R11084 vdd3p3.n4919 vdd3p3.n4917 0.04
R11085 vdd3p3.n5035 comparator_top_0.comparator_0.VDD 0.04
R11086 vdd3p3.n4761 vdd3p3.n4760 0.039
R11087 vdd3p3.n8831 vdd3p3.n8830 0.039
R11088 vdd3p3.n3807 vdd3p3.n3806 0.039
R11089 vdd3p3.n4544 vdd3p3.n4543 0.039
R11090 vdd3p3.n4740 vdd3p3.n4736 0.038
R11091 vdd3p3.n26 vdd3p3.n9 0.038
R11092 vdd3p3.n59 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.vdd3p3 0.038
R11093 vdd3p3.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VPWR 0.038
R11094 vdd3p3.n871 vdd3p3.n855 0.038
R11095 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n852 0.038
R11096 vdd3p3.n880 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VPWR 0.038
R11097 vdd3p3.n1717 vdd3p3.n1700 0.038
R11098 vdd3p3.n1750 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.vdd3p3 0.038
R11099 vdd3p3.n1694 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VPWR 0.038
R11100 vdd3p3.n2562 vdd3p3.n2546 0.038
R11101 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n2543 0.038
R11102 vdd3p3.n2571 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VPWR 0.038
R11103 vdd3p3.n4215 vdd3p3.n4213 0.038
R11104 vdd3p3.n4341 vdd3p3.n4339 0.038
R11105 vdd3p3.n4319 vdd3p3.n4317 0.038
R11106 vdd3p3.n4661 vdd3p3.n4659 0.038
R11107 vdd3p3.n4639 vdd3p3.n4637 0.038
R11108 vdd3p3.n5067 vdd3p3.n5065 0.038
R11109 vdd3p3.n8521 vdd3p3.n8519 0.038
R11110 vdd3p3.n8865 vdd3p3.n8863 0.038
R11111 vdd3p3.n8776 vdd3p3.n8774 0.038
R11112 vdd3p3.n3869 vdd3p3.n3865 0.037
R11113 vdd3p3.n3809 vdd3p3.n3808 0.037
R11114 vdd3p3.n4527 vdd3p3.n4526 0.037
R11115 vdd3p3.n5135 vdd3p3.n5134 0.037
R11116 vdd3p3.n8542 vdd3p3.n8541 0.037
R11117 vdd3p3.n8590 vdd3p3.n8589 0.037
R11118 vdd3p3.n8621 vdd3p3.n8620 0.037
R11119 vdd3p3.n8804 vdd3p3.n8803 0.037
R11120 vdd3p3.n8699 vdd3p3.n8696 0.037
R11121 vdd3p3.n3864 vdd3p3.n3863 0.035
R11122 vdd3p3.n4732 vdd3p3.n4728 0.034
R11123 vdd3p3.n4994 vdd3p3.n4951 0.034
R11124 vdd3p3.n45 vdd3p3.n44 0.033
R11125 vdd3p3.n1736 vdd3p3.n1735 0.033
R11126 vdd3p3.n3850 vdd3p3.n3849 0.033
R11127 vdd3p3.n3801 vdd3p3.n3800 0.033
R11128 vdd3p3.n8696 vdd3p3.n8695 0.033
R11129 vdd3p3.n5006 vdd3p3.n5005 0.033
R11130 vdd3p3.n8896 vdd3p3.n8467 0.033
R11131 vdd3p3.n4226 vdd3p3.n4224 0.032
R11132 vdd3p3.n4348 vdd3p3.n4346 0.032
R11133 vdd3p3.n4312 vdd3p3.n4310 0.032
R11134 vdd3p3.n4668 vdd3p3.n4666 0.032
R11135 vdd3p3.n4632 vdd3p3.n4630 0.032
R11136 vdd3p3.n5078 vdd3p3.n5076 0.032
R11137 vdd3p3.n5123 vdd3p3.n5116 0.031
R11138 vdd3p3.n4980 vdd3p3.n4979 0.031
R11139 vdd3p3.n3874 vdd3p3.n3873 0.031
R11140 vdd3p3.n3693 vdd3p3.n3666 0.031
R11141 vdd3p3.n4828 vdd3p3.n4802 0.031
R11142 vdd3p3.n3450 vdd3p3.n3449 0.03
R11143 vdd3p3.n3599 vdd3p3.n3570 0.03
R11144 vdd3p3.n8580 vdd3p3.n8579 0.03
R11145 vdd3p3.n4972 vdd3p3.n4964 0.03
R11146 vdd3p3.n3591 vdd3p3.n3590 0.03
R11147 vdd3p3.n3685 vdd3p3.n3684 0.03
R11148 vdd3p3.n3755 vdd3p3.n3754 0.03
R11149 vdd3p3.n4820 vdd3p3.n4819 0.03
R11150 vdd3p3.n4751 vdd3p3.n4750 0.03
R11151 vdd3p3.n8790 vdd3p3.n8789 0.03
R11152 vdd3p3.n3588 vdd3p3.n3587 0.029
R11153 vdd3p3.n3498 vdd3p3.n3497 0.029
R11154 vdd3p3.n3682 vdd3p3.n3681 0.029
R11155 vdd3p3.n4817 vdd3p3.n4816 0.029
R11156 vdd3p3.n4294 vdd3p3.n4291 0.029
R11157 vdd3p3.n4614 vdd3p3.n4611 0.029
R11158 vdd3p3.n3653 vdd3p3.n3650 0.029
R11159 vdd3p3.n3724 vdd3p3.n3721 0.029
R11160 vdd3p3.n3557 vdd3p3.n3554 0.029
R11161 vdd3p3.n4789 vdd3p3.n4786 0.029
R11162 vdd3p3.n4934 vdd3p3.n4927 0.029
R11163 vdd3p3.n4834 vdd3p3.n4833 0.029
R11164 vdd3p3.n8546 vdd3p3.n8545 0.029
R11165 vdd3p3.n8594 vdd3p3.n8593 0.029
R11166 vdd3p3.n8659 vdd3p3.n8658 0.029
R11167 vdd3p3.n8625 vdd3p3.n8624 0.029
R11168 vdd3p3.n8808 vdd3p3.n8807 0.029
R11169 vdd3p3.n8606 vdd3p3.n8605 0.029
R11170 vdd3p3.n8824 vdd3p3.n8823 0.029
R11171 vdd3p3.n8644 vdd3p3.n8643 0.029
R11172 vdd3p3.n3835 vdd3p3.n3833 0.029
R11173 vdd3p3.n8536 vdd3p3.n8528 0.029
R11174 vdd3p3.n3674 vdd3p3.n3670 0.028
R11175 vdd3p3.n3490 vdd3p3.n3482 0.028
R11176 vdd3p3.n4809 vdd3p3.n4805 0.028
R11177 vdd3p3.n8681 vdd3p3.n8680 0.028
R11178 vdd3p3.n8670 vdd3p3.n8669 0.028
R11179 vdd3p3.n25 vdd3p3.n13 0.027
R11180 vdd3p3.n13 vdd3p3.n12 0.027
R11181 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vdd3p3 vdd3p3.n0 0.027
R11182 vdd3p3.n872 vdd3p3.n853 0.027
R11183 vdd3p3.n876 vdd3p3.n853 0.027
R11184 vdd3p3.n907 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vdd3p3 0.027
R11185 vdd3p3.n1716 vdd3p3.n1704 0.027
R11186 vdd3p3.n1704 vdd3p3.n1703 0.027
R11187 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vdd3p3 vdd3p3.n1691 0.027
R11188 vdd3p3.n2563 vdd3p3.n2544 0.027
R11189 vdd3p3.n2567 vdd3p3.n2544 0.027
R11190 vdd3p3.n2598 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vdd3p3 0.027
R11191 vdd3p3.n4228 vdd3p3.n4227 0.027
R11192 vdd3p3.n4305 vdd3p3.n4303 0.027
R11193 vdd3p3.n4350 vdd3p3.n4349 0.027
R11194 vdd3p3.n4385 vdd3p3.n4384 0.027
R11195 vdd3p3.n4418 vdd3p3.n4417 0.027
R11196 vdd3p3.n4448 vdd3p3.n4447 0.027
R11197 vdd3p3.n4478 vdd3p3.n4477 0.027
R11198 vdd3p3.n4508 vdd3p3.n4507 0.027
R11199 vdd3p3.n4625 vdd3p3.n4623 0.027
R11200 vdd3p3.n4670 vdd3p3.n4669 0.027
R11201 vdd3p3.n5080 vdd3p3.n5079 0.027
R11202 vdd3p3.n8672 vdd3p3.n8671 0.027
R11203 vdd3p3.n8743 vdd3p3.n8742 0.027
R11204 vdd3p3.n8611 vdd3p3.n8610 0.026
R11205 vdd3p3.n8677 vdd3p3.n8676 0.025
R11206 vdd3p3.n8675 vdd3p3.n8672 0.025
R11207 vdd3p3.n3872 vdd3p3.n3871 0.025
R11208 vdd3p3.n3844 vdd3p3.n3842 0.025
R11209 vdd3p3.n3841 vdd3p3.n3837 0.025
R11210 vdd3p3.n3837 vdd3p3.n3836 0.025
R11211 vdd3p3.n3798 vdd3p3.n3797 0.025
R11212 vdd3p3.n3797 vdd3p3.n3796 0.025
R11213 vdd3p3.n4301 vdd3p3.n4298 0.024
R11214 vdd3p3.n4621 vdd3p3.n4618 0.024
R11215 vdd3p3.n3665 vdd3p3.n3664 0.024
R11216 vdd3p3.n3660 vdd3p3.n3657 0.024
R11217 vdd3p3.n3736 vdd3p3.n3735 0.024
R11218 vdd3p3.n3731 vdd3p3.n3728 0.024
R11219 vdd3p3.n3569 vdd3p3.n3568 0.024
R11220 vdd3p3.n3564 vdd3p3.n3561 0.024
R11221 vdd3p3.n4801 vdd3p3.n4800 0.024
R11222 vdd3p3.n4796 vdd3p3.n4793 0.024
R11223 vdd3p3.n4950 vdd3p3.n4949 0.024
R11224 vdd3p3.n4945 vdd3p3.n4938 0.024
R11225 vdd3p3.n8676 vdd3p3.n8662 0.024
R11226 vdd3p3.n8675 vdd3p3.n8663 0.024
R11227 vdd3p3.n4533 vdd3p3.n4532 0.024
R11228 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd3p3 vdd3p3.n42 0.023
R11229 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd3p3 vdd3p3.n1733 0.023
R11230 vdd3p3.n3692 vdd3p3.n3689 0.023
R11231 vdd3p3.n3762 vdd3p3.n3759 0.023
R11232 vdd3p3.n3598 vdd3p3.n3595 0.023
R11233 vdd3p3.n3511 vdd3p3.n3508 0.023
R11234 vdd3p3.n4827 vdd3p3.n4824 0.023
R11235 vdd3p3.n4758 vdd3p3.n4755 0.023
R11236 vdd3p3.n4993 vdd3p3.n4990 0.023
R11237 vdd3p3.n8539 vdd3p3.n8538 0.023
R11238 vdd3p3.n8587 vdd3p3.n8586 0.023
R11239 vdd3p3.n8801 vdd3p3.n8800 0.023
R11240 vdd3p3.n3812 vdd3p3.n3811 0.023
R11241 vdd3p3.n3862 vdd3p3.n3861 0.023
R11242 vdd3p3.n59 vdd3p3.n2 0.022
R11243 vdd3p3.n878 vdd3p3.n852 0.022
R11244 vdd3p3.n1750 vdd3p3.n1693 0.022
R11245 vdd3p3.n2569 vdd3p3.n2543 0.022
R11246 vdd3p3.n4894 vdd3p3.n4893 0.022
R11247 vdd3p3.n4298 vdd3p3.n4296 0.021
R11248 vdd3p3.n4618 vdd3p3.n4616 0.021
R11249 vdd3p3.n3676 vdd3p3.n3675 0.021
R11250 vdd3p3.n3664 vdd3p3.n3662 0.021
R11251 vdd3p3.n3657 vdd3p3.n3655 0.021
R11252 vdd3p3.n3746 vdd3p3.n3745 0.021
R11253 vdd3p3.n3735 vdd3p3.n3733 0.021
R11254 vdd3p3.n3728 vdd3p3.n3726 0.021
R11255 vdd3p3.n3568 vdd3p3.n3566 0.021
R11256 vdd3p3.n3561 vdd3p3.n3559 0.021
R11257 vdd3p3.n3582 vdd3p3.n3581 0.021
R11258 vdd3p3.n3492 vdd3p3.n3491 0.021
R11259 vdd3p3.n4800 vdd3p3.n4798 0.021
R11260 vdd3p3.n4793 vdd3p3.n4791 0.021
R11261 vdd3p3.n4811 vdd3p3.n4810 0.021
R11262 vdd3p3.n4742 vdd3p3.n4741 0.021
R11263 vdd3p3.n4949 vdd3p3.n4947 0.021
R11264 vdd3p3.n4938 vdd3p3.n4936 0.021
R11265 vdd3p3.n4974 vdd3p3.n4973 0.021
R11266 vdd3p3.n4998 vdd3p3.n4997 0.021
R11267 vdd3p3.n8525 vdd3p3.n8524 0.021
R11268 vdd3p3.n8577 vdd3p3.n8576 0.021
R11269 vdd3p3.n8661 vdd3p3.n8660 0.021
R11270 vdd3p3.n8679 vdd3p3.n8678 0.021
R11271 vdd3p3.n8869 vdd3p3.n8868 0.021
R11272 vdd3p3.n8787 vdd3p3.n8786 0.021
R11273 vdd3p3.n8668 vdd3p3.n8664 0.021
R11274 vdd3p3.n3828 vdd3p3.n3827 0.021
R11275 vdd3p3.n4893 vdd3p3.n4892 0.02
R11276 vdd3p3.n5149 vdd3p3.n5148 0.02
R11277 vdd3p3.n8898 vdd3p3.n5160 0.02
R11278 vdd3p3.n11 vdd3p3.n2 0.019
R11279 vdd3p3.n878 vdd3p3.n877 0.019
R11280 vdd3p3.n1702 vdd3p3.n1693 0.019
R11281 vdd3p3.n2569 vdd3p3.n2568 0.019
R11282 vdd3p3.n1689 vdd3p3.n909 0.019
R11283 vdd3p3.n3380 vdd3p3.n2600 0.019
R11284 vdd3p3.n4308 vdd3p3.n4305 0.019
R11285 vdd3p3.n3449 vdd3p3.n3448 0.019
R11286 vdd3p3.n4628 vdd3p3.n4625 0.019
R11287 vdd3p3.n3811 vdd3p3.n3810 0.019
R11288 vdd3p3.n3875 vdd3p3.n3874 0.019
R11289 vdd3p3.n3447 vdd3p3.n3446 0.019
R11290 vdd3p3.n4565 vdd3p3.n4561 0.019
R11291 vdd3p3.n3763 vdd3p3.n3737 0.019
R11292 vdd3p3.n3578 vdd3p3.n3577 0.018
R11293 vdd3p3.n3672 vdd3p3.n3671 0.018
R11294 vdd3p3.n3742 vdd3p3.n3741 0.018
R11295 vdd3p3.n4807 vdd3p3.n4806 0.018
R11296 vdd3p3.n4738 vdd3p3.n4737 0.018
R11297 vdd3p3.n843 vdd3p3.n63 0.018
R11298 vdd3p3.n2534 vdd3p3.n1754 0.018
R11299 vdd3p3.n8744 vdd3p3.n8687 0.018
R11300 vdd3p3.n4532 vdd3p3.n4531 0.018
R11301 vdd3p3.n3770 vdd3p3.n3769 0.017
R11302 vdd3p3.n4832 vdd3p3.n4831 0.017
R11303 vdd3p3.n8744 vdd3p3.n8688 0.017
R11304 vdd3p3.n8690 vdd3p3.n8689 0.017
R11305 vdd3p3.n3852 vdd3p3.n3851 0.017
R11306 vdd3p3.n3849 vdd3p3.n3848 0.017
R11307 vdd3p3.n3832 vdd3p3.n3829 0.017
R11308 vdd3p3.n3800 vdd3p3.n3799 0.017
R11309 vdd3p3.n3795 vdd3p3.n3794 0.017
R11310 vdd3p3.n3999 vdd3p3.n3998 0.017
R11311 vdd3p3.n4231 vdd3p3.n4230 0.017
R11312 vdd3p3.n4421 vdd3p3.n4420 0.017
R11313 vdd3p3.n4451 vdd3p3.n4450 0.017
R11314 vdd3p3.n4511 vdd3p3.n4510 0.017
R11315 vdd3p3.n3792 vdd3p3.n3791 0.016
R11316 vdd3p3.n26 vdd3p3.n25 0.016
R11317 vdd3p3.n872 vdd3p3.n871 0.016
R11318 vdd3p3.n1717 vdd3p3.n1716 0.016
R11319 vdd3p3.n2563 vdd3p3.n2562 0.016
R11320 vdd3p3.n4291 vdd3p3.n4289 0.016
R11321 vdd3p3.n4611 vdd3p3.n4609 0.016
R11322 vdd3p3.n3650 vdd3p3.n3648 0.016
R11323 vdd3p3.n3721 vdd3p3.n3719 0.016
R11324 vdd3p3.n3554 vdd3p3.n3552 0.016
R11325 vdd3p3.n3785 vdd3p3.n3784 0.016
R11326 vdd3p3.n4786 vdd3p3.n4784 0.016
R11327 vdd3p3.n4927 vdd3p3.n4925 0.016
R11328 vdd3p3.n8612 vdd3p3.n8611 0.016
R11329 vdd3p3.n3998 vdd3p3.n3988 0.016
R11330 vdd3p3.n3787 vdd3p3.n3786 0.016
R11331 vdd3p3.n4244 vdd3p3.n4243 0.015
R11332 vdd3p3.n4236 vdd3p3.n4235 0.015
R11333 vdd3p3.n4367 vdd3p3.n4366 0.015
R11334 vdd3p3.n4362 vdd3p3.n4361 0.015
R11335 vdd3p3.n4353 vdd3p3.n4352 0.015
R11336 vdd3p3.n4401 vdd3p3.n4400 0.015
R11337 vdd3p3.n4396 vdd3p3.n4395 0.015
R11338 vdd3p3.n4391 vdd3p3.n4390 0.015
R11339 vdd3p3.n4431 vdd3p3.n4430 0.015
R11340 vdd3p3.n4426 vdd3p3.n4425 0.015
R11341 vdd3p3.n4461 vdd3p3.n4460 0.015
R11342 vdd3p3.n4456 vdd3p3.n4455 0.015
R11343 vdd3p3.n4491 vdd3p3.n4490 0.015
R11344 vdd3p3.n4486 vdd3p3.n4485 0.015
R11345 vdd3p3.n4481 vdd3p3.n4480 0.015
R11346 vdd3p3.n4521 vdd3p3.n4520 0.015
R11347 vdd3p3.n4516 vdd3p3.n4515 0.015
R11348 vdd3p3.n3437 vdd3p3.n3436 0.015
R11349 vdd3p3.n3430 vdd3p3.n3429 0.015
R11350 vdd3p3.n5128 vdd3p3.n5127 0.015
R11351 vdd3p3.n5122 vdd3p3.n5121 0.015
R11352 vdd3p3.n4689 vdd3p3.n4688 0.015
R11353 vdd3p3.n4682 vdd3p3.n4681 0.015
R11354 vdd3p3.n4673 vdd3p3.n4672 0.015
R11355 vdd3p3.n5104 vdd3p3.n5103 0.015
R11356 vdd3p3.n5096 vdd3p3.n5095 0.015
R11357 vdd3p3.n5091 vdd3p3.n5090 0.015
R11358 vdd3p3.n3666 vdd3p3.n3665 0.015
R11359 vdd3p3.n3737 vdd3p3.n3736 0.015
R11360 vdd3p3.n3570 vdd3p3.n3569 0.015
R11361 vdd3p3.n4802 vdd3p3.n4801 0.015
R11362 vdd3p3.n4951 vdd3p3.n4950 0.015
R11363 vdd3p3.n4996 vdd3p3.n4995 0.015
R11364 vdd3p3.n3860 vdd3p3.n3859 0.015
R11365 vdd3p3.n3853 vdd3p3.n3852 0.015
R11366 vdd3p3.n4000 vdd3p3.n3875 0.015
R11367 vdd3p3.n4173 vdd3p3.n4172 0.015
R11368 vdd3p3.n8883 vdd3p3.n8832 0.014
R11369 vdd3p3.n4542 vdd3p3.n4541 0.014
R11370 vdd3p3.n17 vdd3p3.n14 0.014
R11371 vdd3p3.n864 vdd3p3.n863 0.014
R11372 vdd3p3.n1708 vdd3p3.n1705 0.014
R11373 vdd3p3.n2555 vdd3p3.n2554 0.014
R11374 vdd3p3.n4224 vdd3p3.n4222 0.013
R11375 vdd3p3.n4229 vdd3p3.n4228 0.013
R11376 vdd3p3.n4346 vdd3p3.n4344 0.013
R11377 vdd3p3.n4315 vdd3p3.n4312 0.013
R11378 vdd3p3.n4351 vdd3p3.n4350 0.013
R11379 vdd3p3.n4389 vdd3p3.n4385 0.013
R11380 vdd3p3.n4419 vdd3p3.n4418 0.013
R11381 vdd3p3.n4449 vdd3p3.n4448 0.013
R11382 vdd3p3.n4479 vdd3p3.n4478 0.013
R11383 vdd3p3.n4509 vdd3p3.n4508 0.013
R11384 vdd3p3.n3448 vdd3p3.n3447 0.013
R11385 vdd3p3.n4561 vdd3p3.n4560 0.013
R11386 vdd3p3.n4666 vdd3p3.n4664 0.013
R11387 vdd3p3.n4635 vdd3p3.n4632 0.013
R11388 vdd3p3.n4671 vdd3p3.n4670 0.013
R11389 vdd3p3.n5076 vdd3p3.n5074 0.013
R11390 vdd3p3.n5089 vdd3p3.n5080 0.013
R11391 vdd3p3.n4860 vdd3p3.n4859 0.013
R11392 vdd3p3.n4861 vdd3p3.n4860 0.013
R11393 vdd3p3.n4862 vdd3p3.n4861 0.013
R11394 vdd3p3.n4863 vdd3p3.n4862 0.013
R11395 vdd3p3.n4864 vdd3p3.n4863 0.013
R11396 vdd3p3.n4865 vdd3p3.n4864 0.013
R11397 vdd3p3.n4866 vdd3p3.n4865 0.013
R11398 vdd3p3.n4867 vdd3p3.n4866 0.013
R11399 vdd3p3.n4884 vdd3p3.n4867 0.013
R11400 vdd3p3.n4882 vdd3p3.n4881 0.013
R11401 vdd3p3.n4881 vdd3p3.n4880 0.013
R11402 vdd3p3.n4880 vdd3p3.n4879 0.013
R11403 vdd3p3.n4877 vdd3p3.n4876 0.013
R11404 vdd3p3.n4876 vdd3p3.n4875 0.013
R11405 vdd3p3.n4875 vdd3p3.n4874 0.013
R11406 vdd3p3.n4886 vdd3p3.n4885 0.013
R11407 vdd3p3.n8556 vdd3p3.n8547 0.013
R11408 vdd3p3.n8600 vdd3p3.n8595 0.013
R11409 vdd3p3.n8472 vdd3p3.n8471 0.013
R11410 vdd3p3.n8473 vdd3p3.n8472 0.013
R11411 vdd3p3.n8895 vdd3p3.n8473 0.013
R11412 vdd3p3.n8895 vdd3p3.n8894 0.013
R11413 vdd3p3.n8892 vdd3p3.n8891 0.013
R11414 vdd3p3.n8891 vdd3p3.n8890 0.013
R11415 vdd3p3.n8890 vdd3p3.n8889 0.013
R11416 vdd3p3.n8889 vdd3p3.n8888 0.013
R11417 vdd3p3.n8888 vdd3p3.n8486 0.013
R11418 vdd3p3.n8484 vdd3p3.n8483 0.013
R11419 vdd3p3.n8483 vdd3p3.n8482 0.013
R11420 vdd3p3.n8482 vdd3p3.n8481 0.013
R11421 vdd3p3.n8481 vdd3p3.n8480 0.013
R11422 vdd3p3.n8480 vdd3p3.n8479 0.013
R11423 vdd3p3.n8479 vdd3p3.n8478 0.013
R11424 vdd3p3.n8478 vdd3p3.n8477 0.013
R11425 vdd3p3.n8635 vdd3p3.n8626 0.013
R11426 vdd3p3.n8818 vdd3p3.n8809 0.013
R11427 vdd3p3.n3870 vdd3p3.n3869 0.013
R11428 vdd3p3.n3411 vdd3p3.n3410 0.013
R11429 vdd3p3.n3412 vdd3p3.n3411 0.013
R11430 vdd3p3.n3413 vdd3p3.n3412 0.013
R11431 vdd3p3.n3414 vdd3p3.n3413 0.013
R11432 vdd3p3.n3417 vdd3p3.n3416 0.013
R11433 vdd3p3.n3418 vdd3p3.n3417 0.013
R11434 vdd3p3.n3419 vdd3p3.n3418 0.013
R11435 vdd3p3.n3420 vdd3p3.n3419 0.013
R11436 vdd3p3.n3421 vdd3p3.n3420 0.013
R11437 vdd3p3.n3424 vdd3p3.n3423 0.013
R11438 vdd3p3.n4548 vdd3p3.n3424 0.013
R11439 vdd3p3.n4549 vdd3p3.n4548 0.013
R11440 vdd3p3.n4550 vdd3p3.n4549 0.013
R11441 vdd3p3.n4551 vdd3p3.n4550 0.013
R11442 vdd3p3.n4552 vdd3p3.n4551 0.013
R11443 vdd3p3.n4553 vdd3p3.n4552 0.013
R11444 vdd3p3.n5143 vdd3p3.n4553 0.013
R11445 vdd3p3.n5144 vdd3p3.n5143 0.013
R11446 vdd3p3.n5146 vdd3p3.n5144 0.013
R11447 vdd3p3.n5146 vdd3p3.n5145 0.013
R11448 vdd3p3.n3405 vdd3p3.n3404 0.013
R11449 vdd3p3.n3791 vdd3p3.n3790 0.013
R11450 vdd3p3.n4889 vdd3p3.n4888 0.012
R11451 vdd3p3.n8886 vdd3p3.n8885 0.012
R11452 vdd3p3.n4539 vdd3p3.n4538 0.012
R11453 vdd3p3.n3410 vdd3p3.n3409 0.012
R11454 vdd3p3.n3400 vdd3p3.n3399 0.012
R11455 vdd3p3.n3453 vdd3p3.n3452 0.012
R11456 vdd3p3.n3452 vdd3p3.n3451 0.012
R11457 vdd3p3.n4235 vdd3p3.n4234 0.011
R11458 vdd3p3.n4425 vdd3p3.n4424 0.011
R11459 vdd3p3.n4455 vdd3p3.n4454 0.011
R11460 vdd3p3.n4515 vdd3p3.n4514 0.011
R11461 vdd3p3.n3677 vdd3p3.n3676 0.011
R11462 vdd3p3.n3688 vdd3p3.n3687 0.011
R11463 vdd3p3.n3747 vdd3p3.n3746 0.011
R11464 vdd3p3.n3758 vdd3p3.n3757 0.011
R11465 vdd3p3.n3583 vdd3p3.n3582 0.011
R11466 vdd3p3.n3594 vdd3p3.n3593 0.011
R11467 vdd3p3.n3493 vdd3p3.n3492 0.011
R11468 vdd3p3.n3507 vdd3p3.n3506 0.011
R11469 vdd3p3.n4812 vdd3p3.n4811 0.011
R11470 vdd3p3.n4823 vdd3p3.n4822 0.011
R11471 vdd3p3.n4743 vdd3p3.n4742 0.011
R11472 vdd3p3.n4754 vdd3p3.n4753 0.011
R11473 vdd3p3.n4975 vdd3p3.n4974 0.011
R11474 vdd3p3.n4989 vdd3p3.n4988 0.011
R11475 vdd3p3.n8537 vdd3p3.n8536 0.011
R11476 vdd3p3.n8526 vdd3p3.n8525 0.011
R11477 vdd3p3.n8585 vdd3p3.n8584 0.011
R11478 vdd3p3.n8578 vdd3p3.n8577 0.011
R11479 vdd3p3.n8684 vdd3p3.n8683 0.011
R11480 vdd3p3.n8687 vdd3p3.n8686 0.011
R11481 vdd3p3.n8881 vdd3p3.n8873 0.011
R11482 vdd3p3.n8870 vdd3p3.n8869 0.011
R11483 vdd3p3.n8799 vdd3p3.n8798 0.011
R11484 vdd3p3.n8788 vdd3p3.n8787 0.011
R11485 vdd3p3.n8695 vdd3p3.n8694 0.011
R11486 vdd3p3.n3865 vdd3p3.n3864 0.011
R11487 vdd3p3.n3851 vdd3p3.n3850 0.011
R11488 vdd3p3.n3829 vdd3p3.n3828 0.011
R11489 vdd3p3.n3808 vdd3p3.n3807 0.011
R11490 vdd3p3.n4356 vdd3p3.n4355 0.011
R11491 vdd3p3.n4394 vdd3p3.n4393 0.011
R11492 vdd3p3.n4484 vdd3p3.n4483 0.011
R11493 vdd3p3.n4676 vdd3p3.n4675 0.011
R11494 vdd3p3.n5094 vdd3p3.n5093 0.011
R11495 vdd3p3.n21 vdd3p3.n20 0.01
R11496 vdd3p3.n12 vdd3p3.n11 0.01
R11497 vdd3p3.n861 vdd3p3.n860 0.01
R11498 vdd3p3.n877 vdd3p3.n876 0.01
R11499 vdd3p3.n1712 vdd3p3.n1711 0.01
R11500 vdd3p3.n1703 vdd3p3.n1702 0.01
R11501 vdd3p3.n2552 vdd3p3.n2551 0.01
R11502 vdd3p3.n2568 vdd3p3.n2567 0.01
R11503 vdd3p3.n4898 vdd3p3.n4897 0.01
R11504 vdd3p3.n8685 vdd3p3.n8684 0.01
R11505 vdd3p3.n5132 vdd3p3.n5131 0.01
R11506 vdd3p3.n5131 vdd3p3.n5115 0.01
R11507 vdd3p3.n3786 vdd3p3.n3453 0.009
R11508 vdd3p3.n3689 vdd3p3.n3688 0.009
R11509 vdd3p3.n3759 vdd3p3.n3758 0.009
R11510 vdd3p3.n3595 vdd3p3.n3594 0.009
R11511 vdd3p3.n3508 vdd3p3.n3507 0.009
R11512 vdd3p3.n4824 vdd3p3.n4823 0.009
R11513 vdd3p3.n4755 vdd3p3.n4754 0.009
R11514 vdd3p3.n4990 vdd3p3.n4989 0.009
R11515 vdd3p3.n4859 vdd3p3.n4858 0.009
R11516 vdd3p3.n4883 vdd3p3.n4882 0.009
R11517 vdd3p3.n8538 vdd3p3.n8537 0.009
R11518 vdd3p3.n8586 vdd3p3.n8585 0.009
R11519 vdd3p3.n8683 vdd3p3.n8682 0.009
R11520 vdd3p3.n8471 vdd3p3.n8470 0.009
R11521 vdd3p3.n8486 vdd3p3.n8485 0.009
R11522 vdd3p3.n8477 vdd3p3.n8476 0.009
R11523 vdd3p3.n8873 vdd3p3.n8872 0.009
R11524 vdd3p3.n8800 vdd3p3.n8799 0.009
R11525 vdd3p3.n4172 vdd3p3.n3793 0.009
R11526 vdd3p3.n3422 vdd3p3.n3421 0.009
R11527 vdd3p3.n3790 vdd3p3.n3789 0.009
R11528 vdd3p3.n3780 vdd3p3.n3779 0.009
R11529 vdd3p3.n3774 vdd3p3.n3773 0.009
R11530 vdd3p3.n3765 vdd3p3.n3764 0.009
R11531 vdd3p3.n3779 vdd3p3.n3778 0.009
R11532 vdd3p3.n3775 vdd3p3.n3774 0.009
R11533 vdd3p3.n3766 vdd3p3.n3765 0.009
R11534 vdd3p3.n4888 vdd3p3.n4887 0.009
R11535 vdd3p3.n5003 vdd3p3.n5002 0.009
R11536 vdd3p3.n4887 vdd3p3.n4886 0.009
R11537 vdd3p3.n5004 vdd3p3.n5003 0.009
R11538 vdd3p3.n8562 vdd3p3.n8561 0.009
R11539 vdd3p3.n8604 vdd3p3.n8603 0.009
R11540 vdd3p3.n8748 vdd3p3.n8747 0.009
R11541 vdd3p3.n8561 vdd3p3.n8560 0.009
R11542 vdd3p3.n8603 vdd3p3.n8602 0.009
R11543 vdd3p3.n8820 vdd3p3.n8748 0.009
R11544 vdd3p3.n4247 vdd3p3.n4246 0.009
R11545 vdd3p3.n4370 vdd3p3.n4369 0.009
R11546 vdd3p3.n4405 vdd3p3.n4404 0.009
R11547 vdd3p3.n4435 vdd3p3.n4434 0.009
R11548 vdd3p3.n4464 vdd3p3.n4463 0.009
R11549 vdd3p3.n4495 vdd3p3.n4494 0.009
R11550 vdd3p3.n4525 vdd3p3.n4524 0.009
R11551 vdd3p3.n5111 vdd3p3.n5110 0.009
R11552 vdd3p3.n5036 vdd3p3.n5035 0.009
R11553 vdd3p3.n5031 vdd3p3.n5030 0.009
R11554 vdd3p3.n5106 vdd3p3.n5036 0.009
R11555 vdd3p3.n4524 vdd3p3.n4523 0.009
R11556 vdd3p3.n4494 vdd3p3.n4493 0.009
R11557 vdd3p3.n4434 vdd3p3.n4433 0.009
R11558 vdd3p3.n4465 vdd3p3.n4464 0.009
R11559 vdd3p3.n4404 vdd3p3.n4403 0.009
R11560 vdd3p3.n4248 vdd3p3.n4247 0.009
R11561 vdd3p3.n4371 vdd3p3.n4370 0.009
R11562 vdd3p3.n5110 vdd3p3.n5109 0.009
R11563 vdd3p3.n5032 vdd3p3.n5031 0.009
R11564 vdd3p3.n5033 vdd3p3.n5032 0.009
R11565 vdd3p3.n3468 vdd3p3.n3467 0.008
R11566 vdd3p3.n3782 vdd3p3.n3781 0.008
R11567 vdd3p3.n3776 vdd3p3.n3775 0.008
R11568 vdd3p3.n3771 vdd3p3.n3770 0.008
R11569 vdd3p3.n3767 vdd3p3.n3766 0.008
R11570 vdd3p3.n3781 vdd3p3.n3780 0.008
R11571 vdd3p3.n3768 vdd3p3.n3767 0.008
R11572 vdd3p3.n3772 vdd3p3.n3771 0.008
R11573 vdd3p3.n3777 vdd3p3.n3776 0.008
R11574 vdd3p3.n4831 vdd3p3.n4830 0.008
R11575 vdd3p3.n4995 vdd3p3.n4899 0.008
R11576 vdd3p3.n5001 vdd3p3.n5000 0.008
R11577 vdd3p3.n4899 vdd3p3.n4898 0.008
R11578 vdd3p3.n5004 vdd3p3.n5001 0.008
R11579 vdd3p3.n4830 vdd3p3.n4829 0.008
R11580 vdd3p3.n8559 vdd3p3.n8558 0.008
R11581 vdd3p3.n8564 vdd3p3.n8563 0.008
R11582 vdd3p3.n8885 vdd3p3.n8884 0.008
R11583 vdd3p3.n8822 vdd3p3.n8821 0.008
R11584 vdd3p3.n8746 vdd3p3.n8745 0.008
R11585 vdd3p3.n8884 vdd3p3.n8883 0.008
R11586 vdd3p3.n8560 vdd3p3.n8559 0.008
R11587 vdd3p3.n8821 vdd3p3.n8820 0.008
R11588 vdd3p3.n8602 vdd3p3.n8564 0.008
R11589 vdd3p3.n8745 vdd3p3.n8744 0.008
R11590 vdd3p3.n3785 vdd3p3.n3468 0.008
R11591 vdd3p3.n4172 vdd3p3.n4002 0.008
R11592 vdd3p3.n4246 vdd3p3.n4176 0.008
R11593 vdd3p3.n4369 vdd3p3.n4250 0.008
R11594 vdd3p3.n4373 vdd3p3.n4372 0.008
R11595 vdd3p3.n4407 vdd3p3.n4406 0.008
R11596 vdd3p3.n4463 vdd3p3.n4437 0.008
R11597 vdd3p3.n4493 vdd3p3.n4467 0.008
R11598 vdd3p3.n4497 vdd3p3.n4496 0.008
R11599 vdd3p3.n4540 vdd3p3.n4539 0.008
R11600 vdd3p3.n5112 vdd3p3.n5111 0.008
R11601 vdd3p3.n5108 vdd3p3.n5107 0.008
R11602 vdd3p3.n4523 vdd3p3.n4497 0.008
R11603 vdd3p3.n5113 vdd3p3.n5112 0.008
R11604 vdd3p3.n5107 vdd3p3.n5106 0.008
R11605 vdd3p3.n4541 vdd3p3.n4540 0.008
R11606 vdd3p3.n4467 vdd3p3.n4466 0.008
R11607 vdd3p3.n4437 vdd3p3.n4436 0.008
R11608 vdd3p3.n4433 vdd3p3.n4407 0.008
R11609 vdd3p3.n4176 vdd3p3.n4175 0.008
R11610 vdd3p3.n4002 vdd3p3.n4001 0.008
R11611 vdd3p3.n4250 vdd3p3.n4249 0.008
R11612 vdd3p3.n4403 vdd3p3.n4373 0.008
R11613 vdd3p3.n5034 vdd3p3.n5033 0.008
R11614 vdd3p3.n44 vdd3p3.n43 0.008
R11615 vdd3p3.n21 vdd3p3.n19 0.008
R11616 vdd3p3.n905 vdd3p3.n902 0.008
R11617 vdd3p3.n905 vdd3p3.n904 0.008
R11618 vdd3p3.n861 vdd3p3.n859 0.008
R11619 vdd3p3.n1735 vdd3p3.n1734 0.008
R11620 vdd3p3.n1712 vdd3p3.n1710 0.008
R11621 vdd3p3.n2596 vdd3p3.n2593 0.008
R11622 vdd3p3.n2596 vdd3p3.n2595 0.008
R11623 vdd3p3.n2552 vdd3p3.n2550 0.008
R11624 vdd3p3.n4213 vdd3p3.n4211 0.008
R11625 vdd3p3.n4339 vdd3p3.n4337 0.008
R11626 vdd3p3.n4322 vdd3p3.n4319 0.008
R11627 vdd3p3.n4659 vdd3p3.n4657 0.008
R11628 vdd3p3.n4642 vdd3p3.n4639 0.008
R11629 vdd3p3.n5065 vdd3p3.n5063 0.008
R11630 vdd3p3.n4874 vdd3p3.n4873 0.008
R11631 vdd3p3.n8519 vdd3p3.n8517 0.008
R11632 vdd3p3.n8894 vdd3p3.n8893 0.008
R11633 vdd3p3.n8863 vdd3p3.n8861 0.008
R11634 vdd3p3.n8774 vdd3p3.n8772 0.008
R11635 vdd3p3.n3380 vdd3p3.n3379 0.008
R11636 vdd3p3.n2534 vdd3p3.n2533 0.008
R11637 vdd3p3.n1689 vdd3p3.n1688 0.008
R11638 vdd3p3.n843 vdd3p3.n842 0.008
R11639 vdd3p3.n3675 vdd3p3.n3674 0.007
R11640 vdd3p3.n3745 vdd3p3.n3744 0.007
R11641 vdd3p3.n3581 vdd3p3.n3580 0.007
R11642 vdd3p3.n3491 vdd3p3.n3490 0.007
R11643 vdd3p3.n4810 vdd3p3.n4809 0.007
R11644 vdd3p3.n4741 vdd3p3.n4740 0.007
R11645 vdd3p3.n4973 vdd3p3.n4972 0.007
R11646 vdd3p3.n4878 vdd3p3.n4877 0.007
R11647 vdd3p3.n4872 vdd3p3.n4871 0.007
R11648 vdd3p3.n8524 vdd3p3.n8523 0.007
R11649 vdd3p3.n8576 vdd3p3.n8575 0.007
R11650 vdd3p3.n8662 vdd3p3.n8661 0.007
R11651 vdd3p3.n8868 vdd3p3.n8867 0.007
R11652 vdd3p3.n8786 vdd3p3.n8785 0.007
R11653 vdd3p3.n3872 vdd3p3.n3812 0.007
R11654 vdd3p3.n3847 vdd3p3.n3844 0.007
R11655 vdd3p3.n3842 vdd3p3.n3841 0.007
R11656 vdd3p3.n5115 vdd3p3.n5114 0.007
R11657 vdd3p3.n3416 vdd3p3.n3415 0.007
R11658 vdd3p3.n3788 vdd3p3.n3787 0.007
R11659 vdd3p3.n4879 vdd3p3.n4878 0.006
R11660 vdd3p3.n4999 vdd3p3.n4998 0.006
R11661 vdd3p3.n5133 vdd3p3.n5132 0.006
R11662 vdd3p3.n3415 vdd3p3.n3414 0.006
R11663 vdd3p3.n5095 vdd3p3.n5094 0.006
R11664 vdd3p3.n4681 vdd3p3.n4676 0.006
R11665 vdd3p3.n4485 vdd3p3.n4484 0.006
R11666 vdd3p3.n4395 vdd3p3.n4394 0.006
R11667 vdd3p3.n4361 vdd3p3.n4356 0.006
R11668 vdd3p3.n4234 vdd3p3.n4233 0.005
R11669 vdd3p3.n4265 vdd3p3.n4263 0.005
R11670 vdd3p3.n4281 vdd3p3.n4279 0.005
R11671 vdd3p3.n4424 vdd3p3.n4423 0.005
R11672 vdd3p3.n4454 vdd3p3.n4453 0.005
R11673 vdd3p3.n4514 vdd3p3.n4513 0.005
R11674 vdd3p3.n3440 vdd3p3.n3439 0.005
R11675 vdd3p3.n4569 vdd3p3.n4568 0.005
R11676 vdd3p3.n4567 vdd3p3.n4566 0.005
R11677 vdd3p3.n4585 vdd3p3.n4583 0.005
R11678 vdd3p3.n4601 vdd3p3.n4599 0.005
R11679 vdd3p3.n3527 vdd3p3.n3525 0.005
R11680 vdd3p3.n3543 vdd3p3.n3541 0.005
R11681 vdd3p3.n3612 vdd3p3.n3610 0.005
R11682 vdd3p3.n3640 vdd3p3.n3638 0.005
R11683 vdd3p3.n3628 vdd3p3.n3621 0.005
R11684 vdd3p3.n3711 vdd3p3.n3709 0.005
R11685 vdd3p3.n4776 vdd3p3.n4774 0.005
R11686 vdd3p3.n4917 vdd3p3.n4915 0.005
R11687 vdd3p3.n4873 vdd3p3.n4872 0.005
R11688 vdd3p3.n8678 vdd3p3.n8677 0.005
R11689 vdd3p3.n8893 vdd3p3.n8892 0.005
R11690 vdd3p3.n3871 vdd3p3.n3870 0.005
R11691 vdd3p3.n3861 vdd3p3.n3860 0.005
R11692 vdd3p3.n3784 vdd3p3.n3783 0.004
R11693 vdd3p3.n4858 vdd3p3.n4857 0.004
R11694 vdd3p3.n4884 vdd3p3.n4883 0.004
R11695 vdd3p3.n4870 vdd3p3.n4869 0.004
R11696 vdd3p3.n8470 vdd3p3.n8469 0.004
R11697 vdd3p3.n8485 vdd3p3.n8484 0.004
R11698 vdd3p3.n8476 vdd3p3.n8475 0.004
R11699 vdd3p3.n4174 vdd3p3.n4173 0.004
R11700 vdd3p3.n3423 vdd3p3.n3422 0.004
R11701 vdd3p3.n5130 vdd3p3.n5128 0.004
R11702 vdd3p3.n3436 vdd3p3.n3435 0.004
R11703 vdd3p3.n8641 vdd3p3.n8637 0.004
R11704 vdd3p3.n8640 vdd3p3.n8639 0.004
R11705 vdd3p3.n8637 vdd3p3.n5161 0.004
R11706 vdd3p3.n8641 vdd3p3.n8640 0.004
R11707 vdd3p3.n8658 vdd3p3.n8657 0.004
R11708 vdd3p3.n3407 vdd3p3.n3406 0.003
R11709 vdd3p3.n3785 vdd3p3.n3469 0.003
R11710 vdd3p3.n4172 vdd3p3.n4171 0.003
R11711 vdd3p3.n4352 vdd3p3.n4351 0.003
R11712 vdd3p3.n4390 vdd3p3.n4389 0.003
R11713 vdd3p3.n4480 vdd3p3.n4479 0.003
R11714 vdd3p3.n4672 vdd3p3.n4671 0.003
R11715 vdd3p3.n5090 vdd3p3.n5089 0.003
R11716 vdd3p3.n3681 vdd3p3.n3677 0.003
R11717 vdd3p3.n3751 vdd3p3.n3747 0.003
R11718 vdd3p3.n3587 vdd3p3.n3583 0.003
R11719 vdd3p3.n3497 vdd3p3.n3493 0.003
R11720 vdd3p3.n3467 vdd3p3.n3466 0.003
R11721 vdd3p3.n4816 vdd3p3.n4812 0.003
R11722 vdd3p3.n4747 vdd3p3.n4743 0.003
R11723 vdd3p3.n4979 vdd3p3.n4975 0.003
R11724 vdd3p3.n4885 vdd3p3.n4761 0.003
R11725 vdd3p3.n8545 vdd3p3.n8542 0.003
R11726 vdd3p3.n8527 vdd3p3.n8526 0.003
R11727 vdd3p3.n8593 vdd3p3.n8590 0.003
R11728 vdd3p3.n8579 vdd3p3.n8578 0.003
R11729 vdd3p3.n8641 vdd3p3.n8638 0.003
R11730 vdd3p3.n8469 vdd3p3.n8468 0.003
R11731 vdd3p3.n8475 vdd3p3.n8474 0.003
R11732 vdd3p3.n8624 vdd3p3.n8621 0.003
R11733 vdd3p3.n8871 vdd3p3.n8870 0.003
R11734 vdd3p3.n8807 vdd3p3.n8804 0.003
R11735 vdd3p3.n8789 vdd3p3.n8788 0.003
R11736 vdd3p3.n8832 vdd3p3.n8831 0.003
R11737 vdd3p3.n3863 vdd3p3.n3862 0.003
R11738 vdd3p3.n3855 vdd3p3.n3854 0.003
R11739 vdd3p3.n3833 vdd3p3.n3832 0.003
R11740 vdd3p3.n3804 vdd3p3.n3803 0.003
R11741 vdd3p3.n4543 vdd3p3.n4542 0.003
R11742 vdd3p3.n5134 vdd3p3.n5133 0.003
R11743 vdd3p3.n4856 vdd3p3.n4853 0.003
R11744 vdd3p3.n3785 vdd3p3.n3459 0.003
R11745 vdd3p3.n8731 vdd3p3.n8729 0.002
R11746 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n3 0.002
R11747 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n880 0.002
R11748 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n1694 0.002
R11749 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.vdd3p3 vdd3p3.n2571 0.002
R11750 vdd3p3.n4202 vdd3p3.n4200 0.002
R11751 vdd3p3.n4332 vdd3p3.n4330 0.002
R11752 vdd3p3.n4328 vdd3p3.n4326 0.002
R11753 vdd3p3.n4652 vdd3p3.n4650 0.002
R11754 vdd3p3.n4648 vdd3p3.n4646 0.002
R11755 vdd3p3.n5054 vdd3p3.n5052 0.002
R11756 vdd3p3.n3479 vdd3p3.n3477 0.002
R11757 vdd3p3.n4961 vdd3p3.n4959 0.002
R11758 vdd3p3.n4871 vdd3p3.n4870 0.002
R11759 vdd3p3.n8508 vdd3p3.n8506 0.002
R11760 vdd3p3.n8465 vdd3p3.n8437 0.002
R11761 vdd3p3.n8680 vdd3p3.n8679 0.002
R11762 vdd3p3.n8852 vdd3p3.n8850 0.002
R11763 vdd3p3.n8763 vdd3p3.n8761 0.002
R11764 vdd3p3.n8671 vdd3p3.n8670 0.002
R11765 vdd3p3.n8694 vdd3p3.n8690 0.002
R11766 comparator_top_0.VDD vdd3p3.n8898 0.002
R11767 vdd3p3.n4230 vdd3p3.n4229 0.002
R11768 vdd3p3.n4420 vdd3p3.n4419 0.002
R11769 vdd3p3.n4450 vdd3p3.n4449 0.002
R11770 vdd3p3.n4510 vdd3p3.n4509 0.002
R11771 vdd3p3.n4845 vdd3p3.n4844 0.002
R11772 vdd3p3.n4846 vdd3p3.n4845 0.002
R11773 vdd3p3.n5155 vdd3p3.n5154 0.002
R11774 vdd3p3.n5156 vdd3p3.n5155 0.002
R11775 vdd3p3.n4854 vdd3p3.n3398 0.001
R11776 vdd3p3.n5148 vdd3p3.n3398 0.001
R11777 vdd3p3.n4869 vdd3p3.n4868 0.001
R11778 vdd3p3.n5023 vdd3p3.n5022 0.001
R11779 vdd3p3.n4156 vdd3p3.n4155 0.001
R11780 vdd3p3.n4155 vdd3p3.n4154 0.001
R11781 vdd3p3.n4856 vdd3p3.n4855 0.001
R11782 vdd3p3.n4151 vdd3p3.n4150 0.001
R11783 vdd3p3.n8719 vdd3p3.n8718 0.001
R11784 vdd3p3.n3981 vdd3p3.n3980 0.001
R11785 vdd3p3.n5012 vdd3p3.n5011 0.001
R11786 vdd3p3.n5022 vdd3p3.n5019 0.001
R11787 vdd3p3.n3403 vdd3p3.n3400 0.001
R11788 vdd3p3.n4155 vdd3p3.n4065 0.001
R11789 vdd3p3.n4997 vdd3p3.n4996 0.001
R11790 vdd3p3.n8547 vdd3p3.n8546 0.001
R11791 vdd3p3.n8595 vdd3p3.n8594 0.001
R11792 vdd3p3.n8660 vdd3p3.n8659 0.001
R11793 vdd3p3.n8682 vdd3p3.n8681 0.001
R11794 vdd3p3.n8626 vdd3p3.n8625 0.001
R11795 vdd3p3.n8809 vdd3p3.n8808 0.001
R11796 vdd3p3.n8656 vdd3p3.n8644 0.001
R11797 vdd3p3.n8643 vdd3p3.n8642 0.001
R11798 vdd3p3.n8669 vdd3p3.n8668 0.001
R11799 vdd3p3.n8716 vdd3p3.n8715 0.001
R11800 vdd3p3.n8734 vdd3p3.n8716 0.001
R11801 vdd3p3.n8733 vdd3p3.n8732 0.001
R11802 vdd3p3.n8734 vdd3p3.n8733 0.001
R11803 vdd3p3.n8729 vdd3p3.n8728 0.001
R11804 vdd3p3.n8718 vdd3p3.n8717 0.001
R11805 vdd3p3.n3982 vdd3p3.n3981 0.001
R11806 vdd3p3.n3994 vdd3p3.n3993 0.001
R11807 vdd3p3.n4726 vdd3p3.n4725 0.001
R11808 vdd3p3.n5011 vdd3p3.n5010 0.001
R11809 vdd3p3.n5025 vdd3p3.n5024 0.001
R11810 vdd3p3.n5018 vdd3p3.n5017 0.001
R11811 vdd3p3.n4150 vdd3p3.n4149 0.001
R11812 vdd3p3.n4153 vdd3p3.n4152 0.001
R11813 vdd3p3.n4158 vdd3p3.n4157 0.001
R11814 vdd3p3.n4064 vdd3p3.n4063 0.001
R11815 vdd3p3.n3402 vdd3p3.n3401 0.001
R11816 vdd3p3.n3408 vdd3p3.n3407 0.001
R11817 vdd3p3.n3409 vdd3p3.n3408 0.001
R11818 vdd3p3.n8734 vdd3p3.n8731 0.001
R11819 vdd3p3.n4065 vdd3p3.n4064 0.001
R11820 vdd3p3.n3403 vdd3p3.n3402 0.001
R11821 vdd3p3.n5019 vdd3p3.n5018 0.001
R11822 vdd3p3.n4155 vdd3p3.n4036 0.001
R11823 vdd3p3.n8734 vdd3p3.n8719 0.001
R11824 vdd3p3.n3980 vdd3p3.n3979 0.001
R11825 vdd3p3.n3979 vdd3p3.n3978 0.001
R11826 vdd3p3.n5022 vdd3p3.n4694 0.001
R11827 vdd3p3.n5022 vdd3p3.n5012 0.001
R11828 vdd3p3.n4155 vdd3p3.n4151 0.001
R11829 vdd3p3.n5345 vdd3p3.n5344 0.001
R11830 vdd3p3.n3379 vdd3p3.n2601 0.001
R11831 vdd3p3.n2533 vdd3p3.n1755 0.001
R11832 vdd3p3.n1688 vdd3p3.n910 0.001
R11833 vdd3p3.n842 vdd3p3.n64 0.001
R11834 vdd3p3.n4154 vdd3p3.n4153 0.001
R11835 vdd3p3.n4157 vdd3p3.n4156 0.001
R11836 vdd3p3.n5024 vdd3p3.n5023 0.001
R11837 vdd3p3.n4843 vdd3p3.n4842 0.001
R11838 vdd3p3.n4848 vdd3p3.n4847 0.001
R11839 vdd3p3.n4844 vdd3p3.n4843 0.001
R11840 vdd3p3.n4847 vdd3p3.n4846 0.001
R11841 vdd3p3.n4853 vdd3p3.n4852 0.001
R11842 vdd3p3.n4851 vdd3p3.n4850 0.001
R11843 vdd3p3.n4852 vdd3p3.n4851 0.001
R11844 vdd3p3.n4850 vdd3p3.n4849 0.001
R11845 vdd3p3.n5160 vdd3p3.n5159 0.001
R11846 vdd3p3.n5158 vdd3p3.n5157 0.001
R11847 vdd3p3.n5154 vdd3p3.n5153 0.001
R11848 vdd3p3.n5152 vdd3p3.n5151 0.001
R11849 vdd3p3.n5153 vdd3p3.n5152 0.001
R11850 vdd3p3.n5159 vdd3p3.n5158 0.001
R11851 vdd3p3.n5157 vdd3p3.n5156 0.001
R11852 vdd3p3.n5151 vdd3p3.n5150 0.001
R11853 vss.n1915 vss.t47 1304.5
R11854 vss.n1917 vss.t15 1299.15
R11855 vss.t61 vss.t63 1224.3
R11856 vss.t18 vss.t59 1224.3
R11857 vss.t35 vss.t30 720.228
R11858 vss.t30 vss.t21 720.228
R11859 vss.t0 vss.t12 720.228
R11860 vss.t68 vss.t0 720.228
R11861 vss.t72 vss.t68 720.228
R11862 vss.t4 vss.t3 720.228
R11863 vss.t3 vss.t2 720.228
R11864 vss.t2 vss.t5 720.228
R11865 vss.t66 vss.t40 720.228
R11866 vss.t7 vss.t66 720.228
R11867 vss.t26 vss.t7 720.228
R11868 vss.n1916 vss.t61 612.15
R11869 vss.n1916 vss.t18 612.15
R11870 vss.n401 vss.t35 602.287
R11871 vss.n163 vss.t26 602.287
R11872 vss.n738 vss.n737 388.348
R11873 vss.n734 vss.t74 360.114
R11874 vss.n734 vss.t4 360.114
R11875 vss.n735 vss.n734 332.425
R11876 vss.n737 vss.n736 271.139
R11877 vss.n717 vss.t57 212.294
R11878 vss.n718 vss.t81 91.223
R11879 vss.n1917 vss.n1916 68.662
R11880 vss.n778 vss.t51 68.231
R11881 vss.n190 vss.t28 68.231
R11882 vss.n1916 vss.n1915 67.106
R11883 vss.n737 vss.t72 61.329
R11884 vss.n1784 vss.t46 60.25
R11885 vss.n1511 vss.t17 60.25
R11886 vss.n1624 vss.t14 60.25
R11887 vss.n1166 vss.t42 60.25
R11888 vss.n1150 vss.t52 60.25
R11889 vss.n1268 vss.t20 60.25
R11890 vss.n1351 vss.t11 60.25
R11891 vss.n338 vss.t39 60.25
R11892 vss.n229 vss.t25 60.25
R11893 vss.n865 vss.t49 60.25
R11894 vss.n849 vss.t6 60.25
R11895 vss.n553 vss.t29 60.25
R11896 vss.n537 vss.t34 60.25
R11897 vss.n736 vss.n401 51.895
R11898 vss.n172 vss.n171 51.894
R11899 vss.n1868 vss.t48 35.379
R11900 vss.n1709 vss.t16 35.379
R11901 vss.n1215 vss.n1214 35.379
R11902 vss.n503 vss.n502 35.379
R11903 vss.n722 vss.n721 33.475
R11904 vss.n1862 vss.n1861 31.448
R11905 vss.n1869 vss.n1868 31.448
R11906 vss.n1703 vss.n1702 31.448
R11907 vss.n1710 vss.n1709 31.448
R11908 vss.n194 vss.n193 31.448
R11909 vss.n782 vss.n781 31.448
R11910 vss.n1753 vss.n1749 30.02
R11911 vss.n1746 vss.n1745 30.02
R11912 vss.n1851 vss.n1850 27.517
R11913 vss.n1880 vss.n1879 27.517
R11914 vss.n1692 vss.n1691 27.517
R11915 vss.n1721 vss.n1720 27.517
R11916 vss.n1081 vss.n1080 27.517
R11917 vss.n204 vss.n203 27.517
R11918 vss.n793 vss.n792 27.517
R11919 vss.n443 vss.n442 27.517
R11920 vss.n165 vss.n164 26.59
R11921 vss.n1840 vss.n1839 23.586
R11922 vss.n1893 vss.n1892 23.586
R11923 vss.n1681 vss.n1680 23.586
R11924 vss.n1734 vss.n1733 23.586
R11925 vss.n1106 vss.n1105 23.586
R11926 vss.n217 vss.n216 23.586
R11927 vss.n804 vss.n803 23.586
R11928 vss.n454 vss.n453 23.586
R11929 vss.n1808 vss.n1807 21.62
R11930 vss.n1649 vss.n1648 21.62
R11931 vss.n253 vss.n252 21.62
R11932 vss.n766 vss.n765 21.62
R11933 vss.n414 vss.n413 21.62
R11934 vss.n1829 vss.n1828 19.655
R11935 vss.n1774 vss.n1773 19.655
R11936 vss.n1670 vss.n1669 19.655
R11937 vss.n1615 vss.n1614 19.655
R11938 vss.n273 vss.n272 19.655
R11939 vss.n817 vss.n816 19.655
R11940 vss.n467 vss.n466 19.655
R11941 vss.n1819 vss.n1818 17.689
R11942 vss.n1759 vss.n1758 17.689
R11943 vss.n1660 vss.n1659 17.689
R11944 vss.n1603 vss.n1602 17.689
R11945 vss.n264 vss.n263 17.689
R11946 vss.n755 vss.n754 17.689
R11947 vss.n406 vss.n405 17.689
R11948 vss.n1818 vss.n1817 15.724
R11949 vss.n1758 vss.n1757 15.724
R11950 vss.n1659 vss.n1658 15.724
R11951 vss.n1602 vss.n1601 15.724
R11952 vss.n263 vss.n262 15.724
R11953 vss.n754 vss.n753 15.724
R11954 vss.n405 vss.n404 15.724
R11955 vss.n1830 vss.n1829 13.758
R11956 vss.n1775 vss.n1774 13.758
R11957 vss.n1671 vss.n1670 13.758
R11958 vss.n1616 vss.n1615 13.758
R11959 vss.n274 vss.n273 13.758
R11960 vss.n818 vss.n817 13.758
R11961 vss.n468 vss.n467 13.758
R11962 vss.n1594 vss.n1591 12.005
R11963 vss.n1807 vss.n1806 11.793
R11964 vss.n1749 vss.n1748 11.793
R11965 vss.n1648 vss.n1647 11.793
R11966 vss.n1745 vss.n1744 11.793
R11967 vss.n252 vss.n251 11.793
R11968 vss.n765 vss.n764 11.793
R11969 vss.n413 vss.n412 11.793
R11970 vss.n1841 vss.n1840 9.827
R11971 vss.n1894 vss.n1893 9.827
R11972 vss.n1682 vss.n1681 9.827
R11973 vss.n1735 vss.n1734 9.827
R11974 vss.n1107 vss.n1106 9.827
R11975 vss.n218 vss.n217 9.827
R11976 vss.n805 vss.n804 9.827
R11977 vss.n455 vss.n454 9.827
R11978 vss.n1794 vss.n1793 9.3
R11979 vss.n1796 vss.n1795 9.3
R11980 vss.n1792 vss.n1791 9.3
R11981 vss.n1791 vss.n1790 9.3
R11982 vss.n1885 vss.n1884 9.3
R11983 vss.n1874 vss.n1873 9.3
R11984 vss.n1858 vss.n1857 9.3
R11985 vss.n1847 vss.n1846 9.3
R11986 vss.n1836 vss.n1835 9.3
R11987 vss.n1825 vss.n1824 9.3
R11988 vss.n1814 vss.n1813 9.3
R11989 vss.n1803 vss.n1802 9.3
R11990 vss.n1801 vss.n1800 9.3
R11991 vss.n1810 vss.n1809 9.3
R11992 vss.n1809 vss.n1808 9.3
R11993 vss.n1812 vss.n1811 9.3
R11994 vss.n1821 vss.n1820 9.3
R11995 vss.n1820 vss.n1819 9.3
R11996 vss.n1823 vss.n1822 9.3
R11997 vss.n1832 vss.n1831 9.3
R11998 vss.n1831 vss.n1830 9.3
R11999 vss.n1834 vss.n1833 9.3
R12000 vss.n1843 vss.n1842 9.3
R12001 vss.n1842 vss.n1841 9.3
R12002 vss.n1845 vss.n1844 9.3
R12003 vss.n1854 vss.n1853 9.3
R12004 vss.n1853 vss.n1852 9.3
R12005 vss.n1856 vss.n1855 9.3
R12006 vss.n1865 vss.n1864 9.3
R12007 vss.n1864 vss.n1863 9.3
R12008 vss.n1872 vss.n1871 9.3
R12009 vss.n1871 vss.n1870 9.3
R12010 vss.n1876 vss.n1875 9.3
R12011 vss.n1883 vss.n1882 9.3
R12012 vss.n1882 vss.n1881 9.3
R12013 vss.n1887 vss.n1886 9.3
R12014 vss.n1895 vss.n1894 9.3
R12015 vss.n1776 vss.n1775 9.3
R12016 vss.n1760 vss.n1759 9.3
R12017 vss.n1521 vss.n1520 9.3
R12018 vss.n1523 vss.n1522 9.3
R12019 vss.n1519 vss.n1518 9.3
R12020 vss.n1518 vss.n1517 9.3
R12021 vss.n1579 vss.n1578 9.3
R12022 vss.n1572 vss.n1571 9.3
R12023 vss.n1566 vss.n1565 9.3
R12024 vss.n1559 vss.n1558 9.3
R12025 vss.n1552 vss.n1551 9.3
R12026 vss.n1545 vss.n1544 9.3
R12027 vss.n1538 vss.n1537 9.3
R12028 vss.n1531 vss.n1530 9.3
R12029 vss.n1529 vss.n1528 9.3
R12030 vss.n1534 vss.n1533 9.3
R12031 vss.n1536 vss.n1535 9.3
R12032 vss.n1541 vss.n1540 9.3
R12033 vss.n1543 vss.n1542 9.3
R12034 vss.n1548 vss.n1547 9.3
R12035 vss.n1550 vss.n1549 9.3
R12036 vss.n1555 vss.n1554 9.3
R12037 vss.n1557 vss.n1556 9.3
R12038 vss.n1562 vss.n1561 9.3
R12039 vss.n1564 vss.n1563 9.3
R12040 vss.n1568 vss.n1567 9.3
R12041 vss.n1570 vss.n1569 9.3
R12042 vss.n1574 vss.n1573 9.3
R12043 vss.n1577 vss.n1576 9.3
R12044 vss.n1581 vss.n1580 9.3
R12045 vss.n1634 vss.n1633 9.3
R12046 vss.n1636 vss.n1635 9.3
R12047 vss.n1632 vss.n1631 9.3
R12048 vss.n1631 vss.n1630 9.3
R12049 vss.n1726 vss.n1725 9.3
R12050 vss.n1715 vss.n1714 9.3
R12051 vss.n1699 vss.n1698 9.3
R12052 vss.n1688 vss.n1687 9.3
R12053 vss.n1677 vss.n1676 9.3
R12054 vss.n1666 vss.n1665 9.3
R12055 vss.n1655 vss.n1654 9.3
R12056 vss.n1644 vss.n1643 9.3
R12057 vss.n1642 vss.n1641 9.3
R12058 vss.n1651 vss.n1650 9.3
R12059 vss.n1650 vss.n1649 9.3
R12060 vss.n1653 vss.n1652 9.3
R12061 vss.n1662 vss.n1661 9.3
R12062 vss.n1661 vss.n1660 9.3
R12063 vss.n1664 vss.n1663 9.3
R12064 vss.n1673 vss.n1672 9.3
R12065 vss.n1672 vss.n1671 9.3
R12066 vss.n1675 vss.n1674 9.3
R12067 vss.n1684 vss.n1683 9.3
R12068 vss.n1683 vss.n1682 9.3
R12069 vss.n1686 vss.n1685 9.3
R12070 vss.n1695 vss.n1694 9.3
R12071 vss.n1694 vss.n1693 9.3
R12072 vss.n1697 vss.n1696 9.3
R12073 vss.n1706 vss.n1705 9.3
R12074 vss.n1705 vss.n1704 9.3
R12075 vss.n1713 vss.n1712 9.3
R12076 vss.n1712 vss.n1711 9.3
R12077 vss.n1717 vss.n1716 9.3
R12078 vss.n1724 vss.n1723 9.3
R12079 vss.n1723 vss.n1722 9.3
R12080 vss.n1728 vss.n1727 9.3
R12081 vss.n1604 vss.n1603 9.3
R12082 vss.n1736 vss.n1735 9.3
R12083 vss.n1617 vss.n1616 9.3
R12084 vss.n1371 vss.n1370 9.3
R12085 vss.n1378 vss.n1377 9.3
R12086 vss.n1385 vss.n1384 9.3
R12087 vss.n1383 vss.n1382 9.3
R12088 vss.n1381 vss.n1380 9.3
R12089 vss.n1376 vss.n1375 9.3
R12090 vss.n1374 vss.n1373 9.3
R12091 vss.n1369 vss.n1368 9.3
R12092 vss.n1292 vss.n1291 9.3
R12093 vss.n1296 vss.n1295 9.3
R12094 vss.n1294 vss.n1293 9.3
R12095 vss.n1299 vss.n1298 9.3
R12096 vss.n1301 vss.n1300 9.3
R12097 vss.n1303 vss.n1302 9.3
R12098 vss.n1289 vss.n1288 9.3
R12099 vss.n1287 vss.n1286 9.3
R12100 vss.n1279 vss.n1278 9.3
R12101 vss.n1260 vss.n1259 9.3
R12102 vss.n1361 vss.n1360 9.3
R12103 vss.n1363 vss.n1362 9.3
R12104 vss.n1359 vss.n1358 9.3
R12105 vss.n1358 vss.n1357 9.3
R12106 vss.n1281 vss.n1280 9.3
R12107 vss.n1277 vss.n1276 9.3
R12108 vss.n1276 vss.n1275 9.3
R12109 vss.n1267 vss.n1266 9.3
R12110 vss.n1266 vss.n1265 9.3
R12111 vss.n1348 vss.n1347 9.3
R12112 vss.n1162 vss.n1161 9.3
R12113 vss.n1160 vss.n1159 9.3
R12114 vss.n1158 vss.n1157 9.3
R12115 vss.n1157 vss.n1156 9.3
R12116 vss.n1179 vss.n1178 9.3
R12117 vss.n1175 vss.n1174 9.3
R12118 vss.n1174 vss.n1173 9.3
R12119 vss.n1177 vss.n1176 9.3
R12120 vss.n1252 vss.n1251 9.3
R12121 vss.n1251 vss.n1250 9.3
R12122 vss.n1256 vss.n1255 9.3
R12123 vss.n1254 vss.n1253 9.3
R12124 vss.n1187 vss.n1186 9.3
R12125 vss.n1194 vss.n1193 9.3
R12126 vss.n1201 vss.n1200 9.3
R12127 vss.n1199 vss.n1198 9.3
R12128 vss.n1197 vss.n1196 9.3
R12129 vss.n1192 vss.n1191 9.3
R12130 vss.n1190 vss.n1189 9.3
R12131 vss.n1185 vss.n1184 9.3
R12132 vss.n1093 vss.n1092 9.3
R12133 vss.n1092 vss.n1091 9.3
R12134 vss.n1095 vss.n1094 9.3
R12135 vss.n1108 vss.n1107 9.3
R12136 vss.n1097 vss.n1096 9.3
R12137 vss.n1083 vss.n1082 9.3
R12138 vss.n346 vss.n345 9.3
R12139 vss.n345 vss.n344 9.3
R12140 vss.n350 vss.n349 9.3
R12141 vss.n348 vss.n347 9.3
R12142 vss.n357 vss.n356 9.3
R12143 vss.n364 vss.n363 9.3
R12144 vss.n371 vss.n370 9.3
R12145 vss.n369 vss.n368 9.3
R12146 vss.n367 vss.n366 9.3
R12147 vss.n362 vss.n361 9.3
R12148 vss.n360 vss.n359 9.3
R12149 vss.n355 vss.n354 9.3
R12150 vss.n199 vss.n198 9.3
R12151 vss.n197 vss.n196 9.3
R12152 vss.n196 vss.n195 9.3
R12153 vss.n237 vss.n236 9.3
R12154 vss.n236 vss.n235 9.3
R12155 vss.n241 vss.n240 9.3
R12156 vss.n239 vss.n238 9.3
R12157 vss.n248 vss.n247 9.3
R12158 vss.n259 vss.n258 9.3
R12159 vss.n270 vss.n269 9.3
R12160 vss.n275 vss.n274 9.3
R12161 vss.n268 vss.n267 9.3
R12162 vss.n266 vss.n265 9.3
R12163 vss.n265 vss.n264 9.3
R12164 vss.n257 vss.n256 9.3
R12165 vss.n255 vss.n254 9.3
R12166 vss.n254 vss.n253 9.3
R12167 vss.n246 vss.n245 9.3
R12168 vss.n201 vss.n200 9.3
R12169 vss.n206 vss.n205 9.3
R12170 vss.n219 vss.n218 9.3
R12171 vss.n861 vss.n860 9.3
R12172 vss.n859 vss.n858 9.3
R12173 vss.n857 vss.n856 9.3
R12174 vss.n856 vss.n855 9.3
R12175 vss.n877 vss.n876 9.3
R12176 vss.n873 vss.n872 9.3
R12177 vss.n872 vss.n871 9.3
R12178 vss.n875 vss.n874 9.3
R12179 vss.n885 vss.n884 9.3
R12180 vss.n892 vss.n891 9.3
R12181 vss.n899 vss.n898 9.3
R12182 vss.n906 vss.n905 9.3
R12183 vss.n913 vss.n912 9.3
R12184 vss.n920 vss.n919 9.3
R12185 vss.n926 vss.n925 9.3
R12186 vss.n933 vss.n932 9.3
R12187 vss.n940 vss.n939 9.3
R12188 vss.n942 vss.n941 9.3
R12189 vss.n938 vss.n937 9.3
R12190 vss.n935 vss.n934 9.3
R12191 vss.n931 vss.n930 9.3
R12192 vss.n928 vss.n927 9.3
R12193 vss.n924 vss.n923 9.3
R12194 vss.n922 vss.n921 9.3
R12195 vss.n918 vss.n917 9.3
R12196 vss.n916 vss.n915 9.3
R12197 vss.n911 vss.n910 9.3
R12198 vss.n909 vss.n908 9.3
R12199 vss.n904 vss.n903 9.3
R12200 vss.n902 vss.n901 9.3
R12201 vss.n897 vss.n896 9.3
R12202 vss.n895 vss.n894 9.3
R12203 vss.n890 vss.n889 9.3
R12204 vss.n888 vss.n887 9.3
R12205 vss.n883 vss.n882 9.3
R12206 vss.n945 vss.n944 9.3
R12207 vss.n787 vss.n786 9.3
R12208 vss.n798 vss.n797 9.3
R12209 vss.n785 vss.n784 9.3
R12210 vss.n784 vss.n783 9.3
R12211 vss.n789 vss.n788 9.3
R12212 vss.n796 vss.n795 9.3
R12213 vss.n795 vss.n794 9.3
R12214 vss.n800 vss.n799 9.3
R12215 vss.n807 vss.n806 9.3
R12216 vss.n806 vss.n805 9.3
R12217 vss.n811 vss.n810 9.3
R12218 vss.n809 vss.n808 9.3
R12219 vss.n767 vss.n766 9.3
R12220 vss.n756 vss.n755 9.3
R12221 vss.n819 vss.n818 9.3
R12222 vss.n814 vss.n813 9.3
R12223 vss.n437 vss.n436 9.3
R12224 vss.n448 vss.n447 9.3
R12225 vss.n435 vss.n434 9.3
R12226 vss.n434 vss.n433 9.3
R12227 vss.n439 vss.n438 9.3
R12228 vss.n446 vss.n445 9.3
R12229 vss.n445 vss.n444 9.3
R12230 vss.n450 vss.n449 9.3
R12231 vss.n457 vss.n456 9.3
R12232 vss.n456 vss.n455 9.3
R12233 vss.n461 vss.n460 9.3
R12234 vss.n459 vss.n458 9.3
R12235 vss.n407 vss.n406 9.3
R12236 vss.n415 vss.n414 9.3
R12237 vss.n469 vss.n468 9.3
R12238 vss.n464 vss.n463 9.3
R12239 vss.n549 vss.n548 9.3
R12240 vss.n547 vss.n546 9.3
R12241 vss.n545 vss.n544 9.3
R12242 vss.n544 vss.n543 9.3
R12243 vss.n565 vss.n564 9.3
R12244 vss.n561 vss.n560 9.3
R12245 vss.n560 vss.n559 9.3
R12246 vss.n563 vss.n562 9.3
R12247 vss.n573 vss.n572 9.3
R12248 vss.n580 vss.n579 9.3
R12249 vss.n587 vss.n586 9.3
R12250 vss.n594 vss.n593 9.3
R12251 vss.n601 vss.n600 9.3
R12252 vss.n608 vss.n607 9.3
R12253 vss.n614 vss.n613 9.3
R12254 vss.n621 vss.n620 9.3
R12255 vss.n628 vss.n627 9.3
R12256 vss.n630 vss.n629 9.3
R12257 vss.n626 vss.n625 9.3
R12258 vss.n623 vss.n622 9.3
R12259 vss.n619 vss.n618 9.3
R12260 vss.n616 vss.n615 9.3
R12261 vss.n612 vss.n611 9.3
R12262 vss.n610 vss.n609 9.3
R12263 vss.n606 vss.n605 9.3
R12264 vss.n604 vss.n603 9.3
R12265 vss.n599 vss.n598 9.3
R12266 vss.n597 vss.n596 9.3
R12267 vss.n592 vss.n591 9.3
R12268 vss.n590 vss.n589 9.3
R12269 vss.n585 vss.n584 9.3
R12270 vss.n583 vss.n582 9.3
R12271 vss.n578 vss.n577 9.3
R12272 vss.n576 vss.n575 9.3
R12273 vss.n571 vss.n570 9.3
R12274 vss.n633 vss.n632 9.3
R12275 vss.n687 vss.n686 9.3
R12276 vss.n1269 vss.n1268 8.764
R12277 vss.n1167 vss.n1166 8.764
R12278 vss.n733 vss.n732 8.399
R12279 vss.n1789 vss.n1788 8.215
R12280 vss.n1516 vss.n1515 8.215
R12281 vss.n1629 vss.n1628 8.215
R12282 vss.n1155 vss.n1154 8.215
R12283 vss.n1356 vss.n1355 8.215
R12284 vss.n1274 vss.n1273 8.215
R12285 vss.n1264 vss.n1263 8.215
R12286 vss.n1172 vss.n1171 8.215
R12287 vss.n1249 vss.n1248 8.215
R12288 vss.n343 vss.n342 8.215
R12289 vss.n234 vss.n233 8.215
R12290 vss.n854 vss.n853 8.215
R12291 vss.n870 vss.n869 8.215
R12292 vss.n542 vss.n541 8.215
R12293 vss.n558 vss.n557 8.215
R12294 vss.n178 vss.n173 7.697
R12295 vss.n731 vss.n728 7.697
R12296 vss.n727 vss.n726 7.476
R12297 vss.n738 vss.n161 6.997
R12298 vss.n1151 vss.n1150 6.922
R12299 vss.n850 vss.n849 6.922
R12300 vss.n538 vss.n537 6.922
R12301 vss.n1512 vss.n1511 6.92
R12302 vss.n1625 vss.n1624 6.92
R12303 vss.n1352 vss.n1351 6.92
R12304 vss.n866 vss.n865 6.92
R12305 vss.n554 vss.n553 6.92
R12306 vss.n1785 vss.n1784 6.92
R12307 vss.n339 vss.n338 6.919
R12308 vss.n230 vss.n229 6.919
R12309 vss.n166 vss.n165 6.81
R12310 vss.n743 vss.n742 6.81
R12311 vss.n157 vss.n156 6.81
R12312 vss.n760 vss.n759 6.549
R12313 vss.n419 vss.n418 6.548
R12314 vss.n1799 vss.n1798 6.434
R12315 vss.n1640 vss.n1639 6.434
R12316 vss.n244 vss.n243 6.434
R12317 vss.n1860 vss.n1859 6.023
R12318 vss.n1867 vss.n1866 6.023
R12319 vss.n1701 vss.n1700 6.023
R12320 vss.n1708 vss.n1707 6.023
R12321 vss.n1089 vss.n1088 6.023
R12322 vss.n192 vss.n191 6.023
R12323 vss.n780 vss.n779 6.023
R12324 vss.n431 vss.n430 6.023
R12325 vss.n1852 vss.n1851 5.896
R12326 vss.n1881 vss.n1880 5.896
R12327 vss.n1693 vss.n1692 5.896
R12328 vss.n1722 vss.n1721 5.896
R12329 vss.n1082 vss.n1081 5.896
R12330 vss.n205 vss.n204 5.896
R12331 vss.n794 vss.n793 5.896
R12332 vss.n444 vss.n443 5.896
R12333 vss.n1787 vss.n1786 5.647
R12334 vss.n1514 vss.n1513 5.647
R12335 vss.n1627 vss.n1626 5.647
R12336 vss.n1153 vss.n1152 5.647
R12337 vss.n1354 vss.n1353 5.647
R12338 vss.n1272 vss.n1271 5.647
R12339 vss.n1262 vss.n1261 5.647
R12340 vss.n1170 vss.n1169 5.647
R12341 vss.n1247 vss.n1246 5.647
R12342 vss.n341 vss.n340 5.647
R12343 vss.n232 vss.n231 5.647
R12344 vss.n852 vss.n851 5.647
R12345 vss.n868 vss.n867 5.647
R12346 vss.n540 vss.n539 5.647
R12347 vss.n556 vss.n555 5.647
R12348 vss.n1489 vss.n1488 5.609
R12349 vss.n1594 vss.n1593 5.609
R12350 vss.n25 vss.n24 5.397
R12351 vss.n978 vss.n977 5.389
R12352 vss.n831 vss.n830 5.389
R12353 vss.n519 vss.n518 5.389
R12354 vss.n58 vss.n57 5.388
R12355 vss.n83 vss.n82 5.388
R12356 vss.n108 vss.n107 5.388
R12357 vss.n133 vss.n132 5.388
R12358 vss.n492 vss.n491 5.388
R12359 vss.n712 vss.n711 5.386
R12360 vss.n1754 vss.n1753 5.37
R12361 vss.n1747 vss.n1746 5.37
R12362 vss.n353 vss.n352 5.286
R12363 vss.n1527 vss.n1526 5.286
R12364 vss.n1183 vss.n1182 5.275
R12365 vss.n1367 vss.n1366 5.275
R12366 vss.n1285 vss.n1284 5.275
R12367 vss.n881 vss.n880 5.274
R12368 vss.n569 vss.n568 5.274
R12369 vss.n1849 vss.n1848 5.27
R12370 vss.n1878 vss.n1877 5.27
R12371 vss.n1690 vss.n1689 5.27
R12372 vss.n1719 vss.n1718 5.27
R12373 vss.n791 vss.n790 5.27
R12374 vss.n441 vss.n440 5.27
R12375 vss.n70 vss.n69 5.134
R12376 vss.n95 vss.n94 5.134
R12377 vss.n990 vss.n989 5.134
R12378 vss.n120 vss.n119 5.134
R12379 vss.n148 vss.n147 5.134
R12380 vss.n509 vss.n508 5.134
R12381 vss.n738 vss.n159 4.794
R12382 vss.n1797 vss.n1783 4.764
R12383 vss.n1364 vss.n1350 4.764
R12384 vss.n1282 vss.n1258 4.764
R12385 vss.n1349 vss.n1346 4.764
R12386 vss.n1180 vss.n1165 4.764
R12387 vss.n1257 vss.n1245 4.764
R12388 vss.n351 vss.n337 4.764
R12389 vss.n242 vss.n228 4.764
R12390 vss.n878 vss.n864 4.764
R12391 vss.n566 vss.n552 4.764
R12392 vss.n1525 vss.n1524 4.764
R12393 vss.n1638 vss.n1637 4.764
R12394 vss.n1164 vss.n1163 4.764
R12395 vss.n863 vss.n862 4.764
R12396 vss.n551 vss.n550 4.764
R12397 vss.n723 vss.n722 4.749
R12398 vss.n197 vss.n190 4.683
R12399 vss.n1093 vss.n1087 4.682
R12400 vss.n785 vss.n778 4.682
R12401 vss.n435 vss.n429 4.682
R12402 vss.n1270 vss.n1269 4.65
R12403 vss.n1168 vss.n1167 4.65
R12404 vss.n1484 vss.n1483 4.517
R12405 vss.n1838 vss.n1837 4.517
R12406 vss.n1891 vss.n1890 4.517
R12407 vss.n1897 vss.n1896 4.517
R12408 vss.n1587 vss.n1586 4.517
R12409 vss.n1679 vss.n1678 4.517
R12410 vss.n1732 vss.n1731 4.517
R12411 vss.n1738 vss.n1737 4.517
R12412 vss.n1086 vss.n1085 4.517
R12413 vss.n209 vss.n208 4.517
R12414 vss.n802 vss.n801 4.517
R12415 vss.n452 vss.n451 4.517
R12416 vss.n1485 vss.n1484 4.5
R12417 vss.n1898 vss.n1897 4.5
R12418 vss.n1588 vss.n1587 4.5
R12419 vss.n1739 vss.n1738 4.5
R12420 vss.n1498 vss.n1494 4.5
R12421 vss.n1507 vss.n1506 4.5
R12422 vss.n1620 vss.n1619 4.5
R12423 vss.n1766 vss.n1762 4.5
R12424 vss.n1779 vss.n1778 4.5
R12425 vss.n1465 vss.n1461 4.5
R12426 vss.n1474 vss.n1473 4.5
R12427 vss.n1607 vss.n1606 4.5
R12428 vss.n1391 vss.n1390 4.5
R12429 vss.n1309 vss.n1308 4.5
R12430 vss.n1207 vss.n1206 4.5
R12431 vss.n377 vss.n376 4.5
R12432 vss.n279 vss.n278 4.5
R12433 vss.n291 vss.n287 4.5
R12434 vss.n295 vss.n284 4.5
R12435 vss.n301 vss.n300 4.5
R12436 vss.n307 vss.n306 4.5
R12437 vss.n322 vss.n321 4.5
R12438 vss.n326 vss.n315 4.5
R12439 vss.n332 vss.n331 4.5
R12440 vss.n335 vss.n312 4.5
R12441 vss.n210 vss.n209 4.5
R12442 vss.n214 vss.n189 4.5
R12443 vss.n223 vss.n222 4.5
R12444 vss.n226 vss.n186 4.5
R12445 vss.n714 vss.n710 4.5
R12446 vss.n702 vss.n701 4.5
R12447 vss.n692 vss.n691 4.5
R12448 vss.n681 vss.n680 4.5
R12449 vss.n676 vss.n675 4.5
R12450 vss.n36 vss.n34 4.5
R12451 vss.n43 vss.n42 4.5
R12452 vss.n525 vss.n524 4.5
R12453 vss.n535 vss.n534 4.5
R12454 vss.n472 vss.n471 4.5
R12455 vss.n421 vss.n417 4.5
R12456 vss.n822 vss.n821 4.5
R12457 vss.n837 vss.n836 4.5
R12458 vss.n847 vss.n846 4.5
R12459 vss.n135 vss.n131 4.5
R12460 vss.n110 vss.n106 4.5
R12461 vss.n116 vss.n102 4.5
R12462 vss.n776 vss.n758 4.5
R12463 vss.n770 vss.n769 4.5
R12464 vss.n141 vss.n127 4.5
R12465 vss.n986 vss.n972 4.5
R12466 vss.n85 vss.n81 4.5
R12467 vss.n980 vss.n976 4.5
R12468 vss.n494 vss.n490 4.5
R12469 vss.n500 vss.n486 4.5
R12470 vss.n427 vss.n409 4.5
R12471 vss.n27 vss.n23 4.5
R12472 vss.n60 vss.n56 4.5
R12473 vss.n66 vss.n52 4.5
R12474 vss.n91 vss.n77 4.5
R12475 vss.n951 vss.n950 4.5
R12476 vss.n639 vss.n638 4.5
R12477 vss.n1099 vss.n1086 4.5
R12478 vss.n1103 vss.n1079 4.5
R12479 vss.n1112 vss.n1111 4.5
R12480 vss.n1118 vss.n1117 4.5
R12481 vss.n1336 vss.n1312 4.5
R12482 vss.n1404 vss.n1403 4.5
R12483 vss.n1408 vss.n1397 4.5
R12484 vss.n1414 vss.n1413 4.5
R12485 vss.n1417 vss.n1394 4.5
R12486 vss.n1236 vss.n1210 4.5
R12487 vss.n1233 vss.n1232 4.5
R12488 vss.n1223 vss.n1222 4.5
R12489 vss.n1227 vss.n1213 4.5
R12490 vss.n1333 vss.n1332 4.5
R12491 vss.n1323 vss.n1322 4.5
R12492 vss.n1327 vss.n1315 4.5
R12493 vss.n1809 vss.n1805 4.141
R12494 vss.n1752 vss.n1751 4.141
R12495 vss.n1650 vss.n1646 4.141
R12496 vss.n1743 vss.n1742 4.141
R12497 vss.n1210 vss.n1209 4.141
R12498 vss.n1394 vss.n1393 4.141
R12499 vss.n1312 vss.n1311 4.141
R12500 vss.n1117 vss.n1116 4.141
R12501 vss.n312 vss.n311 4.141
R12502 vss.n306 vss.n305 4.141
R12503 vss.n254 vss.n250 4.141
R12504 vss.n186 vss.n185 4.141
R12505 vss.n56 vss.n54 4.141
R12506 vss.n81 vss.n79 4.141
R12507 vss.n976 vss.n974 4.141
R12508 vss.n106 vss.n104 4.141
R12509 vss.n131 vss.n129 4.141
R12510 vss.n836 vss.n834 4.141
R12511 vss.n767 vss.n763 4.141
R12512 vss.n769 vss.n767 4.141
R12513 vss.n415 vss.n411 4.141
R12514 vss.n417 vss.n415 4.141
R12515 vss.n524 vss.n522 4.141
R12516 vss.n490 vss.n488 4.141
R12517 vss.n23 vss.n21 4.141
R12518 vss.n691 vss.n689 4.141
R12519 vss.n710 vss.n708 4.141
R12520 vss.n1473 vss.n1472 3.764
R12521 vss.n1827 vss.n1826 3.764
R12522 vss.n1772 vss.n1771 3.764
R12523 vss.n1778 vss.n1777 3.764
R12524 vss.n1506 vss.n1505 3.764
R12525 vss.n1668 vss.n1667 3.764
R12526 vss.n1613 vss.n1612 3.764
R12527 vss.n1619 vss.n1618 3.764
R12528 vss.n1232 vss.n1231 3.764
R12529 vss.n1413 vss.n1412 3.764
R12530 vss.n1332 vss.n1331 3.764
R12531 vss.n1111 vss.n1110 3.764
R12532 vss.n331 vss.n330 3.764
R12533 vss.n300 vss.n299 3.764
R12534 vss.n222 vss.n221 3.764
R12535 vss.n944 vss.n943 3.764
R12536 vss.n950 vss.n948 3.764
R12537 vss.n813 vss.n812 3.764
R12538 vss.n821 vss.n819 3.764
R12539 vss.n463 vss.n462 3.764
R12540 vss.n471 vss.n469 3.764
R12541 vss.n632 vss.n631 3.764
R12542 vss.n638 vss.n636 3.764
R12543 vss.n666 vss.n664 3.49
R12544 vss.n346 vss.n339 3.478
R12545 vss.n237 vss.n230 3.478
R12546 vss.n1519 vss.n1512 3.477
R12547 vss.n1632 vss.n1625 3.477
R12548 vss.n1359 vss.n1352 3.477
R12549 vss.n873 vss.n866 3.477
R12550 vss.n561 vss.n554 3.477
R12551 vss.n1792 vss.n1785 3.477
R12552 vss.n1158 vss.n1151 3.476
R12553 vss.n857 vss.n850 3.476
R12554 vss.n545 vss.n538 3.476
R12555 vss.n1461 vss.n1459 3.388
R12556 vss.n1820 vss.n1816 3.388
R12557 vss.n1760 vss.n1756 3.388
R12558 vss.n1762 vss.n1760 3.388
R12559 vss.n1494 vss.n1492 3.388
R12560 vss.n1661 vss.n1657 3.388
R12561 vss.n1604 vss.n1600 3.388
R12562 vss.n1606 vss.n1604 3.388
R12563 vss.n265 vss.n261 3.388
R12564 vss.n52 vss.n50 3.388
R12565 vss.n77 vss.n75 3.388
R12566 vss.n972 vss.n970 3.388
R12567 vss.n102 vss.n100 3.388
R12568 vss.n127 vss.n125 3.388
R12569 vss.n846 vss.n844 3.388
R12570 vss.n756 vss.n752 3.388
R12571 vss.n758 vss.n756 3.388
R12572 vss.n407 vss.n403 3.388
R12573 vss.n409 vss.n407 3.388
R12574 vss.n534 vss.n532 3.388
R12575 vss.n486 vss.n484 3.388
R12576 vss.n34 vss.n32 3.388
R12577 vss.n701 vss.n699 3.388
R12578 vss.n398 vss.n181 3.339
R12579 vss.n398 vss.n397 3.339
R12580 vss.n176 vss.n175 3.339
R12581 vss.n741 vss.n157 3.339
R12582 vss.n743 vss.n741 3.339
R12583 vss.n167 vss.n166 3.339
R12584 vss.n1478 vss.t64 3.306
R12585 vss.n1478 vss.t62 3.306
R12586 vss.n1591 vss.t19 3.306
R12587 vss.n1591 vss.t60 3.306
R12588 vss.n1217 vss.n1215 3.306
R12589 vss.n1217 vss.n1216 3.306
R12590 vss.n1398 vss.t13 3.306
R12591 vss.n1317 vss.n1316 3.306
R12592 vss.n316 vss.t41 3.306
R12593 vss.n316 vss.t67 3.306
R12594 vss.n288 vss.t65 3.306
R12595 vss.n288 vss.t27 3.306
R12596 vss.n68 vss.t69 3.306
R12597 vss.n68 vss.t73 3.306
R12598 vss.n93 vss.t75 3.306
R12599 vss.n93 vss.t71 3.306
R12600 vss.n988 vss.t70 3.306
R12601 vss.n988 vss.t56 3.306
R12602 vss.n118 vss.t79 3.306
R12603 vss.n118 vss.t80 3.306
R12604 vss.n146 vss.t78 3.306
R12605 vss.n146 vss.n145 3.306
R12606 vss.n145 vss.n144 3.306
R12607 vss.n144 vss.t50 3.306
R12608 vss.n505 vss.n503 3.306
R12609 vss.n506 vss.n505 3.306
R12610 vss.n507 vss.n506 3.306
R12611 vss.n507 vss.t76 3.306
R12612 vss.n38 vss.t77 3.306
R12613 vss.n38 vss.t1 3.306
R12614 vss.n665 vss.t82 3.306
R12615 vss.n665 vss.t58 3.306
R12616 vss.n1206 vss.n1204 3.228
R12617 vss.n1390 vss.n1388 3.228
R12618 vss.n1308 vss.n1306 3.228
R12619 vss.n376 vss.n374 3.228
R12620 vss.n719 vss.n718 3.211
R12621 vss.n157 vss.n155 3.033
R12622 vss.n181 vss.n180 3.033
R12623 vss.n166 vss.n162 3.033
R12624 vss.n744 vss.n743 3.033
R12625 vss.n175 vss.n174 3.033
R12626 vss.n397 vss.n396 3.033
R12627 vss.n1124 vss.n1123 3.033
R12628 vss.n1126 vss.n1125 3.033
R12629 vss.n1129 vss.n1128 3.033
R12630 vss.n1461 vss.n1460 3.011
R12631 vss.n1816 vss.n1815 3.011
R12632 vss.n1756 vss.n1755 3.011
R12633 vss.n1762 vss.n1761 3.011
R12634 vss.n1494 vss.n1493 3.011
R12635 vss.n1657 vss.n1656 3.011
R12636 vss.n1600 vss.n1599 3.011
R12637 vss.n1606 vss.n1605 3.011
R12638 vss.n1206 vss.n1205 3.011
R12639 vss.n1390 vss.n1389 3.011
R12640 vss.n1308 vss.n1307 3.011
R12641 vss.n376 vss.n375 3.011
R12642 vss.n261 vss.n260 3.011
R12643 vss.n278 vss.n277 3.011
R12644 vss.n52 vss.n51 3.011
R12645 vss.n77 vss.n76 3.011
R12646 vss.n972 vss.n971 3.011
R12647 vss.n102 vss.n101 3.011
R12648 vss.n127 vss.n126 3.011
R12649 vss.n846 vss.n845 3.011
R12650 vss.n752 vss.n751 3.011
R12651 vss.n758 vss.n757 3.011
R12652 vss.n403 vss.n402 3.011
R12653 vss.n409 vss.n408 3.011
R12654 vss.n534 vss.n533 3.011
R12655 vss.n486 vss.n485 3.011
R12656 vss.n34 vss.n33 3.011
R12657 vss.n701 vss.n700 3.011
R12658 vss.n1473 vss.n1471 2.635
R12659 vss.n1831 vss.n1827 2.635
R12660 vss.n1776 vss.n1772 2.635
R12661 vss.n1778 vss.n1776 2.635
R12662 vss.n1506 vss.n1504 2.635
R12663 vss.n1672 vss.n1668 2.635
R12664 vss.n1617 vss.n1613 2.635
R12665 vss.n1619 vss.n1617 2.635
R12666 vss.n276 vss.n275 2.635
R12667 vss.n950 vss.n949 2.635
R12668 vss.n821 vss.n820 2.635
R12669 vss.n471 vss.n470 2.635
R12670 vss.n638 vss.n637 2.635
R12671 vss.n42 vss.n41 2.635
R12672 vss.n675 vss.n671 2.635
R12673 vss.n1232 vss.n1230 2.527
R12674 vss.n1413 vss.n1411 2.527
R12675 vss.n1332 vss.n1330 2.527
R12676 vss.n331 vss.n329 2.527
R12677 vss.n300 vss.n298 2.527
R12678 vss.n1121 vss.n1120 2.356
R12679 vss.n1805 vss.n1804 2.258
R12680 vss.n1751 vss.n1750 2.258
R12681 vss.n1646 vss.n1645 2.258
R12682 vss.n1742 vss.n1741 2.258
R12683 vss.n1212 vss.n1211 2.258
R12684 vss.n1396 vss.n1395 2.258
R12685 vss.n1314 vss.n1313 2.258
R12686 vss.n1078 vss.n1077 2.258
R12687 vss.n314 vss.n313 2.258
R12688 vss.n283 vss.n282 2.258
R12689 vss.n250 vss.n249 2.258
R12690 vss.n188 vss.n187 2.258
R12691 vss.n56 vss.n55 2.258
R12692 vss.n81 vss.n80 2.258
R12693 vss.n976 vss.n975 2.258
R12694 vss.n106 vss.n105 2.258
R12695 vss.n131 vss.n130 2.258
R12696 vss.n836 vss.n835 2.258
R12697 vss.n763 vss.n762 2.258
R12698 vss.n769 vss.n768 2.258
R12699 vss.n411 vss.n410 2.258
R12700 vss.n417 vss.n416 2.258
R12701 vss.n524 vss.n523 2.258
R12702 vss.n490 vss.n489 2.258
R12703 vss.n23 vss.n22 2.258
R12704 vss.n691 vss.n690 2.258
R12705 vss.n710 vss.n709 2.258
R12706 vss.n686 vss.n685 2.24
R12707 vss.n159 vss.n158 2.219
R12708 vss.n1863 vss.n1862 1.965
R12709 vss.n1870 vss.n1869 1.965
R12710 vss.n1704 vss.n1703 1.965
R12711 vss.n1711 vss.n1710 1.965
R12712 vss.n1091 vss.n1090 1.965
R12713 vss.n195 vss.n194 1.965
R12714 vss.n783 vss.n782 1.965
R12715 vss.n433 vss.n432 1.965
R12716 vss.n1484 vss.n1482 1.882
R12717 vss.n1842 vss.n1838 1.882
R12718 vss.n1895 vss.n1891 1.882
R12719 vss.n1897 vss.n1895 1.882
R12720 vss.n1587 vss.n1585 1.882
R12721 vss.n1683 vss.n1679 1.882
R12722 vss.n1736 vss.n1732 1.882
R12723 vss.n1738 vss.n1736 1.882
R12724 vss.n1109 vss.n1108 1.882
R12725 vss.n220 vss.n219 1.882
R12726 vss.n806 vss.n802 1.882
R12727 vss.n456 vss.n452 1.882
R12728 vss.n675 vss.n674 1.882
R12729 vss.n1222 vss.n1221 1.821
R12730 vss.n1403 vss.n1402 1.821
R12731 vss.n1322 vss.n1321 1.821
R12732 vss.n321 vss.n320 1.821
R12733 vss.n287 vss.n286 1.821
R12734 vss.n720 vss.n716 1.665
R12735 vss.n666 vss.n665 1.603
R12736 vss.n1591 vss.n1590 1.601
R12737 vss.n144 vss.n143 1.601
R12738 vss.n505 vss.n504 1.601
R12739 vss.n164 vss.n163 1.572
R12740 vss.n738 vss.n172 1.572
R12741 vss.n171 vss.n170 1.572
R12742 vss.n1480 vss.n1479 1.519
R12743 vss.n1933 vss.n1490 1.514
R12744 vss.n1924 vss.n1595 1.514
R12745 vss.n1920 vss.n1747 1.514
R12746 vss.n1912 vss.n1754 1.512
R12747 vss.n680 vss.n679 1.505
R12748 vss.n825 vss.n824 1.484
R12749 vss.n959 vss.n151 1.484
R12750 vss.n513 vss.n512 1.484
R12751 vss.n647 vss.n474 1.484
R12752 vss.n999 vss.n98 1.484
R12753 vss.n964 vss.n123 1.484
R12754 vss.n1004 vss.n73 1.484
R12755 vss.n642 vss.n641 1.484
R12756 vss.n954 vss.n953 1.484
R12757 vss.n994 vss.n993 1.484
R12758 vss.n1318 vss.n1317 1.467
R12759 vss.n317 vss.n316 1.467
R12760 vss.n1218 vss.n1217 1.467
R12761 vss.n1399 vss.n1398 1.467
R12762 vss.n289 vss.n288 1.467
R12763 vss.n70 vss.n68 1.41
R12764 vss.n95 vss.n93 1.41
R12765 vss.n990 vss.n988 1.41
R12766 vss.n120 vss.n118 1.41
R12767 vss.n148 vss.n146 1.41
R12768 vss.n509 vss.n507 1.41
R12769 vss.n46 vss.n45 1.345
R12770 vss.n46 vss.n30 1.342
R12771 vss.n1055 vss.n1052 1.137
R12772 vss.n1055 vss.n1054 1.137
R12773 vss.n1055 vss.n1051 1.137
R12774 vss.n1957 vss.n1947 1.137
R12775 vss.n1957 vss.n1949 1.137
R12776 vss.n1957 vss.n1945 1.137
R12777 vss.n1957 vss.n1952 1.137
R12778 vss.n1957 vss.n1942 1.137
R12779 vss.n1957 vss.n1954 1.137
R12780 vss.n1957 vss.n1456 1.137
R12781 vss.n1957 vss.n1956 1.137
R12782 vss.n1957 vss.n1453 1.137
R12783 vss.n1957 vss.n1449 1.137
R12784 vss.n1957 vss.n2 1.137
R12785 vss.n1055 vss.n5 1.136
R12786 vss.n1933 vss.n1486 1.13
R12787 vss.n1924 vss.n1589 1.13
R12788 vss.n1920 vss.n1740 1.13
R12789 vss.n1912 vss.n1899 1.13
R12790 vss.n1853 vss.n1849 1.129
R12791 vss.n1882 vss.n1878 1.129
R12792 vss.n1694 vss.n1690 1.129
R12793 vss.n1723 vss.n1719 1.129
R12794 vss.n1084 vss.n1083 1.129
R12795 vss.n207 vss.n206 1.129
R12796 vss.n795 vss.n791 1.129
R12797 vss.n445 vss.n441 1.129
R12798 vss.n673 vss.n672 1.129
R12799 vss.n715 vss.n714 1.125
R12800 vss.n1790 vss.n1789 1.095
R12801 vss.n1517 vss.n1516 1.095
R12802 vss.n1630 vss.n1629 1.095
R12803 vss.n1156 vss.n1155 1.095
R12804 vss.n1357 vss.n1356 1.095
R12805 vss.n1275 vss.n1274 1.095
R12806 vss.n1265 vss.n1264 1.095
R12807 vss.n1173 vss.n1172 1.095
R12808 vss.n1250 vss.n1249 1.095
R12809 vss.n344 vss.n343 1.095
R12810 vss.n235 vss.n234 1.095
R12811 vss.n855 vss.n854 1.095
R12812 vss.n871 vss.n870 1.095
R12813 vss.n543 vss.n542 1.095
R12814 vss.n559 vss.n558 1.095
R12815 vss.n161 vss.n160 1.087
R12816 vss.n39 vss.n38 1.053
R12817 vss.n385 vss.n309 0.903
R12818 vss.n1421 vss.n1419 0.903
R12819 vss.n1137 vss.n1121 0.903
R12820 vss.n390 vss.n280 0.903
R12821 vss.n381 vss.n378 0.903
R12822 vss.n1048 vss.n1047 0.854
R12823 vss.n1439 vss.n1438 0.853
R12824 vss.n735 vss.n733 0.768
R12825 vss.n1791 vss.n1787 0.752
R12826 vss.n1518 vss.n1514 0.752
R12827 vss.n1631 vss.n1627 0.752
R12828 vss.n1157 vss.n1153 0.752
R12829 vss.n1358 vss.n1354 0.752
R12830 vss.n1276 vss.n1272 0.752
R12831 vss.n1266 vss.n1262 0.752
R12832 vss.n1174 vss.n1170 0.752
R12833 vss.n1251 vss.n1247 0.752
R12834 vss.n1111 vss.n1109 0.752
R12835 vss.n1086 vss.n1084 0.752
R12836 vss.n345 vss.n341 0.752
R12837 vss.n278 vss.n276 0.752
R12838 vss.n222 vss.n220 0.752
R12839 vss.n209 vss.n207 0.752
R12840 vss.n236 vss.n232 0.752
R12841 vss.n856 vss.n852 0.752
R12842 vss.n872 vss.n868 0.752
R12843 vss.n544 vss.n540 0.752
R12844 vss.n560 vss.n556 0.752
R12845 vss.n674 vss.n673 0.752
R12846 vss.n746 vss.n745 0.721
R12847 vss.n395 vss.n394 0.721
R12848 vss.n1342 vss.n1338 0.707
R12849 vss.n1241 vss.n1238 0.707
R12850 vss.n723 vss.n720 0.699
R12851 vss.n1429 vss.n1425 0.682
R12852 vss.n1244 vss.n1065 0.682
R12853 vss.n1922 vss.n1921 0.682
R12854 vss.n383 vss.n382 0.682
R12855 vss.n1002 vss.n1001 0.682
R12856 vss.n997 vss.n996 0.682
R12857 vss.n967 vss.n966 0.682
R12858 vss.n962 vss.n961 0.682
R12859 vss.n1242 vss.n1241 0.682
R12860 vss.n1031 vss.n1022 0.682
R12861 vss.n1040 vss.n16 0.682
R12862 vss.n40 vss.n39 0.637
R12863 vss.n1123 vss.n1122 0.621
R12864 vss.n1133 vss.n1130 0.614
R12865 vss.n309 vss.n281 0.593
R12866 vss.n318 vss.n317 0.573
R12867 vss.n1400 vss.n1399 0.573
R12868 vss.n1219 vss.n1218 0.572
R12869 vss.n1319 vss.n1318 0.572
R12870 vss.n1942 vss.n1941 0.568
R12871 vss.n290 vss.n289 0.559
R12872 vss.n1926 vss.n1925 0.534
R12873 comparator_top_0.VSS vss 0.511
R12874 vss.n1488 vss.n1487 0.461
R12875 vss.n1593 vss.n1592 0.461
R12876 vss.n1189 vss.n1188 0.461
R12877 vss.n1373 vss.n1372 0.461
R12878 vss.n1291 vss.n1290 0.461
R12879 vss.n359 vss.n358 0.461
R12880 vss.n54 vss.n53 0.461
R12881 vss.n79 vss.n78 0.461
R12882 vss.n974 vss.n973 0.461
R12883 vss.n104 vss.n103 0.461
R12884 vss.n129 vss.n128 0.461
R12885 vss.n887 vss.n886 0.461
R12886 vss.n834 vss.n833 0.461
R12887 vss.n575 vss.n574 0.461
R12888 vss.n522 vss.n521 0.461
R12889 vss.n488 vss.n487 0.461
R12890 vss.n21 vss.n20 0.461
R12891 vss.n708 vss.n707 0.461
R12892 vss.n1533 vss.n1532 0.46
R12893 vss.n1459 vss.n1458 0.43
R12894 vss.n1492 vss.n1491 0.43
R12895 vss.n1196 vss.n1195 0.43
R12896 vss.n1380 vss.n1379 0.43
R12897 vss.n1298 vss.n1297 0.43
R12898 vss.n366 vss.n365 0.43
R12899 vss.n50 vss.n49 0.43
R12900 vss.n75 vss.n74 0.43
R12901 vss.n970 vss.n969 0.43
R12902 vss.n100 vss.n99 0.43
R12903 vss.n125 vss.n124 0.43
R12904 vss.n894 vss.n893 0.43
R12905 vss.n844 vss.n843 0.43
R12906 vss.n582 vss.n581 0.43
R12907 vss.n532 vss.n531 0.43
R12908 vss.n484 vss.n483 0.43
R12909 vss.n32 vss.n31 0.43
R12910 vss.n699 vss.n698 0.43
R12911 vss.n1540 vss.n1539 0.429
R12912 vss.n1799 vss.n1797 0.418
R12913 vss.n244 vss.n242 0.418
R12914 vss.n1640 vss.n1638 0.418
R12915 vss.n1471 vss.n1470 0.398
R12916 vss.n1504 vss.n1503 0.398
R12917 vss.n901 vss.n900 0.398
R12918 vss.n589 vss.n588 0.398
R12919 vss.n1547 vss.n1546 0.398
R12920 vss.n1915 vss.n1914 0.384
R12921 vss.n1479 vss.n1478 0.377
R12922 vss.n1864 vss.n1860 0.376
R12923 vss.n1871 vss.n1867 0.376
R12924 vss.n1705 vss.n1701 0.376
R12925 vss.n1712 vss.n1708 0.376
R12926 vss.n1210 vss.n1208 0.376
R12927 vss.n1213 vss.n1212 0.376
R12928 vss.n1394 vss.n1392 0.376
R12929 vss.n1397 vss.n1396 0.376
R12930 vss.n1312 vss.n1310 0.376
R12931 vss.n1315 vss.n1314 0.376
R12932 vss.n1117 vss.n1115 0.376
R12933 vss.n1079 vss.n1078 0.376
R12934 vss.n1092 vss.n1089 0.376
R12935 vss.n312 vss.n310 0.376
R12936 vss.n315 vss.n314 0.376
R12937 vss.n306 vss.n304 0.376
R12938 vss.n284 vss.n283 0.376
R12939 vss.n186 vss.n184 0.376
R12940 vss.n189 vss.n188 0.376
R12941 vss.n196 vss.n192 0.376
R12942 vss.n784 vss.n780 0.376
R12943 vss.n434 vss.n431 0.376
R12944 vss.n1585 vss.n1584 0.366
R12945 vss.n908 vss.n907 0.366
R12946 vss.n596 vss.n595 0.366
R12947 vss.n1554 vss.n1553 0.366
R12948 vss.n937 vss.n936 0.366
R12949 vss.n625 vss.n624 0.366
R12950 vss.n1753 vss.n1752 0.337
R12951 vss.n1746 vss.n1743 0.337
R12952 vss.n1576 vss.n1575 0.334
R12953 vss.n915 vss.n914 0.334
R12954 vss.n603 vss.n602 0.334
R12955 vss.n1561 vss.n1560 0.333
R12956 vss.n930 vss.n929 0.333
R12957 vss.n618 vss.n617 0.333
R12958 vss.n388 vss.n387 0.324
R12959 vss.n645 vss.n644 0.324
R12960 vss.n516 vss.n515 0.324
R12961 vss.n957 vss.n956 0.324
R12962 vss.n828 vss.n827 0.324
R12963 vss.n353 vss.n351 0.314
R12964 vss.n1527 vss.n1525 0.314
R12965 comparator_top_0.comparator_bias_0.VSS vss.n1917 0.312
R12966 vss.n1490 vss.n1489 0.297
R12967 vss.n1595 vss.n1594 0.297
R12968 vss.n720 vss.n649 0.297
R12969 vss.n96 vss.n95 0.25
R12970 vss.n149 vss.n148 0.25
R12971 vss.n510 vss.n509 0.25
R12972 vss.n991 vss.n990 0.25
R12973 vss.n121 vss.n120 0.25
R12974 vss.n71 vss.n70 0.25
R12975 vss.n1424 vss.n1423 0.233
R12976 vss.n667 vss.n666 0.23
R12977 vss.n1181 vss.n1164 0.228
R12978 vss.n1181 vss.n1180 0.228
R12979 vss.n1283 vss.n1257 0.228
R12980 vss.n1283 vss.n1282 0.228
R12981 vss.n1365 vss.n1349 0.228
R12982 vss.n1365 vss.n1364 0.228
R12983 vss.n879 vss.n863 0.228
R12984 vss.n879 vss.n878 0.228
R12985 vss.n567 vss.n551 0.228
R12986 vss.n567 vss.n566 0.228
R12987 vss.n735 vss.n723 0.212
R12988 vss.n1367 vss.n1365 0.19
R12989 vss.n1285 vss.n1283 0.19
R12990 vss.n1183 vss.n1181 0.19
R12991 vss.n881 vss.n879 0.19
R12992 vss.n569 vss.n567 0.19
R12993 vss.n1872 vss.n1865 0.19
R12994 vss.n1570 vss.n1568 0.19
R12995 vss.n1713 vss.n1706 0.19
R12996 vss.n1175 vss.n1168 0.19
R12997 vss.n1277 vss.n1270 0.19
R12998 vss.n1270 vss.n1267 0.19
R12999 vss.n924 vss.n922 0.19
R13000 vss.n612 vss.n610 0.19
R13001 vss.n1801 vss.n1799 0.164
R13002 vss.n1642 vss.n1640 0.164
R13003 vss.n1369 vss.n1367 0.164
R13004 vss.n1287 vss.n1285 0.164
R13005 vss.n1185 vss.n1183 0.164
R13006 vss.n246 vss.n244 0.164
R13007 vss.n883 vss.n881 0.164
R13008 vss.n571 vss.n569 0.164
R13009 vss.n1797 vss.n1796 0.158
R13010 vss.n1525 vss.n1523 0.158
R13011 vss.n1638 vss.n1636 0.158
R13012 vss.n1164 vss.n1162 0.158
R13013 vss.n1180 vss.n1179 0.158
R13014 vss.n1257 vss.n1256 0.158
R13015 vss.n1282 vss.n1281 0.158
R13016 vss.n1349 vss.n1348 0.158
R13017 vss.n1364 vss.n1363 0.158
R13018 vss.n351 vss.n350 0.158
R13019 vss.n242 vss.n241 0.158
R13020 vss.n863 vss.n861 0.158
R13021 vss.n878 vss.n877 0.158
R13022 vss.n551 vss.n549 0.158
R13023 vss.n566 vss.n565 0.158
R13024 vss.n481 vss.n480 0.156
R13025 vss.n1443 vss.n1442 0.146
R13026 vss.n1812 vss.n1810 0.144
R13027 vss.n1823 vss.n1821 0.144
R13028 vss.n1834 vss.n1832 0.144
R13029 vss.n1845 vss.n1843 0.144
R13030 vss.n1856 vss.n1854 0.144
R13031 vss.n1883 vss.n1876 0.144
R13032 vss.n1536 vss.n1534 0.144
R13033 vss.n1543 vss.n1541 0.144
R13034 vss.n1550 vss.n1548 0.144
R13035 vss.n1557 vss.n1555 0.144
R13036 vss.n1564 vss.n1562 0.144
R13037 vss.n1577 vss.n1574 0.144
R13038 vss.n1653 vss.n1651 0.144
R13039 vss.n1664 vss.n1662 0.144
R13040 vss.n1675 vss.n1673 0.144
R13041 vss.n1686 vss.n1684 0.144
R13042 vss.n1697 vss.n1695 0.144
R13043 vss.n1724 vss.n1717 0.144
R13044 vss.n1376 vss.n1374 0.144
R13045 vss.n1383 vss.n1381 0.144
R13046 vss.n1294 vss.n1292 0.144
R13047 vss.n1301 vss.n1299 0.144
R13048 vss.n1192 vss.n1190 0.144
R13049 vss.n1199 vss.n1197 0.144
R13050 vss.n362 vss.n360 0.144
R13051 vss.n369 vss.n367 0.144
R13052 vss.n257 vss.n255 0.144
R13053 vss.n268 vss.n266 0.144
R13054 vss.n890 vss.n888 0.144
R13055 vss.n897 vss.n895 0.144
R13056 vss.n904 vss.n902 0.144
R13057 vss.n911 vss.n909 0.144
R13058 vss.n918 vss.n916 0.144
R13059 vss.n931 vss.n928 0.144
R13060 vss.n938 vss.n935 0.144
R13061 vss.n796 vss.n789 0.144
R13062 vss.n807 vss.n800 0.144
R13063 vss.n446 vss.n439 0.144
R13064 vss.n457 vss.n450 0.144
R13065 vss.n578 vss.n576 0.144
R13066 vss.n585 vss.n583 0.144
R13067 vss.n592 vss.n590 0.144
R13068 vss.n599 vss.n597 0.144
R13069 vss.n606 vss.n604 0.144
R13070 vss.n619 vss.n616 0.144
R13071 vss.n626 vss.n623 0.144
R13072 vss.n1529 vss.n1527 0.141
R13073 vss.n355 vss.n353 0.141
R13074 vss.n1204 vss.n1203 0.125
R13075 vss.n1388 vss.n1387 0.125
R13076 vss.n1306 vss.n1305 0.125
R13077 vss.n374 vss.n373 0.125
R13078 vss.n948 vss.n947 0.125
R13079 vss.n636 vss.n635 0.125
R13080 vss.n945 vss.n942 0.121
R13081 vss.n814 vss.n811 0.121
R13082 vss.n464 vss.n461 0.121
R13083 vss.n633 vss.n630 0.121
R13084 comparator_top_0.VSS vss.n1957 0.116
R13085 vss.n392 vss.n391 0.113
R13086 vss.n1135 vss.n1134 0.113
R13087 vss.n1888 vss.n1887 0.105
R13088 vss.n1582 vss.n1581 0.105
R13089 vss.n1729 vss.n1728 0.105
R13090 vss.n1230 vss.n1229 0.09
R13091 vss.n1411 vss.n1410 0.09
R13092 vss.n1330 vss.n1329 0.09
R13093 vss.n329 vss.n328 0.09
R13094 vss.n298 vss.n297 0.09
R13095 vss.n1129 vss.n1127 0.085
R13096 vss.n1130 vss.n1129 0.076
R13097 vss.n30 vss.n29 0.074
R13098 vss.n378 vss.n336 0.069
R13099 vss.n280 vss.n227 0.069
R13100 vss.n1121 vss.n1119 0.069
R13101 vss.n1419 vss.n1418 0.068
R13102 vss.n309 vss.n308 0.068
R13103 vss.n396 vss.n395 0.067
R13104 vss.n745 vss.n744 0.067
R13105 vss.n202 vss.n201 0.066
R13106 vss.n1098 vss.n1097 0.066
R13107 vss.n1918 comparator_top_0.comparator_bias_0.VSS 0.065
R13108 vss vss.n748 0.065
R13109 vss.n1130 vss.n1124 0.062
R13110 vss.n1338 vss.n1337 0.062
R13111 vss.n1238 vss.n1237 0.062
R13112 vss.n1464 vss.n1463 0.06
R13113 vss.n1497 vss.n1496 0.06
R13114 vss.n1598 vss.n1597 0.06
R13115 vss.n1765 vss.n1764 0.06
R13116 vss.n98 vss.n92 0.059
R13117 vss.n151 vss.n142 0.059
R13118 vss.n824 vss.n777 0.059
R13119 vss.n474 vss.n428 0.059
R13120 vss.n512 vss.n501 0.059
R13121 vss.n123 vss.n117 0.059
R13122 vss.n73 vss.n67 0.059
R13123 vss.n1104 vss.n1103 0.059
R13124 vss.n993 vss.n987 0.059
R13125 vss.n953 vss.n848 0.059
R13126 vss.n641 vss.n536 0.059
R13127 vss.n64 vss.n63 0.057
R13128 vss.n89 vss.n88 0.057
R13129 vss.n984 vss.n983 0.057
R13130 vss.n114 vss.n113 0.057
R13131 vss.n139 vss.n138 0.057
R13132 vss.n841 vss.n840 0.057
R13133 vss.n774 vss.n773 0.057
R13134 vss.n425 vss.n424 0.057
R13135 vss.n529 vss.n528 0.057
R13136 vss.n498 vss.n497 0.057
R13137 vss.n1233 vss.n1228 0.057
R13138 vss.n1468 vss.n1467 0.055
R13139 vss.n1769 vss.n1768 0.055
R13140 vss.n1501 vss.n1500 0.055
R13141 vss.n1610 vss.n1609 0.055
R13142 vss.n180 vss.n179 0.055
R13143 vss.n155 vss.n154 0.055
R13144 vss.n1127 vss.n1126 0.055
R13145 vss.n1221 vss.n1220 0.054
R13146 vss.n1402 vss.n1401 0.054
R13147 vss.n1321 vss.n1320 0.054
R13148 vss.n320 vss.n319 0.054
R13149 vss.n286 vss.n285 0.054
R13150 vss.n45 vss.n37 0.054
R13151 vss.n656 vss.n655 0.052
R13152 vss.n1477 vss.n1476 0.051
R13153 vss.n1476 vss.n1475 0.051
R13154 vss.n1782 vss.n1781 0.051
R13155 vss.n1781 vss.n1780 0.051
R13156 vss.n1510 vss.n1509 0.051
R13157 vss.n1509 vss.n1508 0.051
R13158 vss.n1623 vss.n1622 0.051
R13159 vss.n1622 vss.n1621 0.051
R13160 vss.n1007 vss.n1006 0.049
R13161 vss.n45 vss.n44 0.049
R13162 vss.n687 vss.n684 0.048
R13163 vss.n696 vss.n695 0.048
R13164 vss.n705 vss.n704 0.048
R13165 vss.n749 vss 0.048
R13166 vss.n1469 vss.n1468 0.047
R13167 vss.n1770 vss.n1769 0.047
R13168 vss.n1502 vss.n1501 0.047
R13169 vss.n1611 vss.n1610 0.047
R13170 vss.n1140 vss.n1139 0.047
R13171 vss.n1328 vss.n1327 0.045
R13172 vss.n63 vss.n62 0.045
R13173 vss.n88 vss.n87 0.045
R13174 vss.n983 vss.n982 0.045
R13175 vss.n113 vss.n112 0.045
R13176 vss.n138 vss.n137 0.045
R13177 vss.n840 vss.n839 0.045
R13178 vss.n773 vss.n772 0.045
R13179 vss.n424 vss.n423 0.045
R13180 vss.n528 vss.n527 0.045
R13181 vss.n497 vss.n496 0.045
R13182 vss.n296 vss.n295 0.045
R13183 vss.n327 vss.n326 0.045
R13184 vss.n215 vss.n214 0.045
R13185 vss.n1409 vss.n1408 0.045
R13186 vss.n1414 vss.n1409 0.044
R13187 vss.n1425 vss.n1345 0.044
R13188 vss.n332 vss.n327 0.044
R13189 vss.n301 vss.n296 0.044
R13190 vss.n223 vss.n215 0.044
R13191 vss.n1065 vss.n1064 0.044
R13192 vss.n1333 vss.n1328 0.044
R13193 vss.n993 vss.n992 0.043
R13194 vss.n953 vss.n952 0.043
R13195 vss.n641 vss.n640 0.043
R13196 vss.n1858 vss.n1856 0.043
R13197 vss.n1876 vss.n1874 0.043
R13198 vss.n1566 vss.n1564 0.043
R13199 vss.n1574 vss.n1572 0.043
R13200 vss.n1699 vss.n1697 0.043
R13201 vss.n1717 vss.n1715 0.043
R13202 vss.n1097 vss.n1095 0.043
R13203 vss.n201 vss.n199 0.043
R13204 vss.n920 vss.n918 0.043
R13205 vss.n928 vss.n926 0.043
R13206 vss.n789 vss.n787 0.043
R13207 vss.n439 vss.n437 0.043
R13208 vss.n608 vss.n606 0.043
R13209 vss.n616 vss.n614 0.043
R13210 vss.n98 vss.n97 0.043
R13211 vss.n151 vss.n150 0.043
R13212 vss.n824 vss.n823 0.043
R13213 vss.n474 vss.n473 0.043
R13214 vss.n512 vss.n511 0.043
R13215 vss.n73 vss.n72 0.043
R13216 vss.n123 vss.n122 0.043
R13217 vss.n1764 vss.n1763 0.043
R13218 vss.n1463 vss.n1462 0.042
R13219 vss.n1496 vss.n1495 0.042
R13220 vss.n1597 vss.n1596 0.042
R13221 vss.n1908 vss.n1907 0.042
R13222 vss.n1907 vss.n1906 0.042
R13223 vss.n1906 vss.n1905 0.042
R13224 vss.n1905 vss.n1904 0.042
R13225 vss.n1904 vss.n1903 0.042
R13226 vss.n1903 vss.n1902 0.042
R13227 vss.n1900 vss.n1457 0.042
R13228 vss.n1941 vss.n1457 0.042
R13229 vss.n1941 vss.n1940 0.042
R13230 vss.n1940 vss.n1939 0.042
R13231 vss.n1939 vss.n1938 0.042
R13232 vss.n1938 vss.n1937 0.042
R13233 vss.n1937 vss.n1936 0.042
R13234 vss.n1930 vss.n1929 0.042
R13235 vss.n479 vss.n478 0.042
R13236 vss.n478 vss.n477 0.042
R13237 vss.n477 vss.n476 0.042
R13238 vss.n476 vss.n475 0.042
R13239 vss.n475 vss.n16 0.042
R13240 vss.n16 vss.n15 0.042
R13241 vss.n15 vss.n14 0.042
R13242 vss.n14 vss.n13 0.042
R13243 vss.n13 vss.n12 0.042
R13244 vss.n12 vss.n11 0.042
R13245 vss.n1022 vss.n1021 0.042
R13246 vss.n1021 vss.n1020 0.042
R13247 vss.n1020 vss.n1019 0.042
R13248 vss.n1019 vss.n1018 0.042
R13249 vss.n1018 vss.n1017 0.042
R13250 vss.n1017 vss.n1016 0.042
R13251 vss.n1014 vss.n1013 0.042
R13252 vss.n1013 vss.n1012 0.042
R13253 vss.n1012 vss.n1011 0.042
R13254 vss.n1011 vss.n1010 0.042
R13255 vss.n1010 vss.n1009 0.042
R13256 vss.n1009 vss.n1008 0.042
R13257 vss.n1142 vss.n1141 0.042
R13258 vss.n1143 vss.n1142 0.042
R13259 vss.n1146 vss.n1145 0.042
R13260 vss.n1147 vss.n1146 0.042
R13261 vss.n1063 vss.n1062 0.042
R13262 vss.n1060 vss.n1059 0.042
R13263 vss.n1065 vss.n1063 0.041
R13264 vss.n676 vss.n670 0.041
R13265 vss.n1340 vss.n1339 0.041
R13266 vss.n291 vss.n290 0.041
R13267 vss.n1796 vss.n1794 0.04
R13268 vss.n1523 vss.n1521 0.04
R13269 vss.n1636 vss.n1634 0.04
R13270 vss.n1162 vss.n1160 0.04
R13271 vss.n1179 vss.n1177 0.04
R13272 vss.n1256 vss.n1254 0.04
R13273 vss.n1281 vss.n1279 0.04
R13274 vss.n1363 vss.n1361 0.04
R13275 vss.n350 vss.n348 0.04
R13276 vss.n241 vss.n239 0.04
R13277 vss.n861 vss.n859 0.04
R13278 vss.n877 vss.n875 0.04
R13279 vss.n549 vss.n547 0.04
R13280 vss.n565 vss.n563 0.04
R13281 vss.n1847 vss.n1845 0.038
R13282 vss.n1887 vss.n1885 0.038
R13283 vss.n1559 vss.n1557 0.038
R13284 vss.n1581 vss.n1579 0.038
R13285 vss.n1688 vss.n1686 0.038
R13286 vss.n1728 vss.n1726 0.038
R13287 vss.n913 vss.n911 0.038
R13288 vss.n935 vss.n933 0.038
R13289 vss.n800 vss.n798 0.038
R13290 vss.n450 vss.n448 0.038
R13291 vss.n601 vss.n599 0.038
R13292 vss.n623 vss.n621 0.038
R13293 vss.n480 vss.n479 0.037
R13294 vss.n1008 vss.n1007 0.037
R13295 vss.n1928 vss.n1927 0.036
R13296 vss.n1022 vss.n48 0.036
R13297 vss.n1425 vss.n1424 0.036
R13298 vss.n669 vss.n668 0.035
R13299 vss.n704 vss.n703 0.035
R13300 vss.n1145 vss.n1144 0.035
R13301 vss.n1061 vss.n1060 0.035
R13302 vss.n1141 vss.n1140 0.034
R13303 vss.n1016 vss.n1015 0.033
R13304 vss.n1228 vss.n1227 0.032
R13305 vss.n1836 vss.n1834 0.032
R13306 vss.n1552 vss.n1550 0.032
R13307 vss.n1677 vss.n1675 0.032
R13308 vss.n1931 vss.n1930 0.032
R13309 vss.n906 vss.n904 0.032
R13310 vss.n942 vss.n940 0.032
R13311 vss.n811 vss.n809 0.032
R13312 vss.n461 vss.n459 0.032
R13313 vss.n594 vss.n592 0.032
R13314 vss.n630 vss.n628 0.032
R13315 vss.n713 vss.n712 0.031
R13316 vss.n659 vss.n658 0.031
R13317 vss.n663 vss.n662 0.031
R13318 vss.n1910 vss.n1909 0.03
R13319 vss.n1902 vss.n1901 0.03
R13320 vss.n1112 vss.n1104 0.029
R13321 vss.n1223 vss.n1219 0.029
R13322 vss.n1323 vss.n1319 0.029
R13323 vss.n1810 vss.n1803 0.029
R13324 vss.n1534 vss.n1531 0.029
R13325 vss.n1651 vss.n1644 0.029
R13326 vss.n1909 vss.n1908 0.029
R13327 vss.n1927 vss.n1926 0.029
R13328 vss.n1374 vss.n1371 0.029
R13329 vss.n1292 vss.n1289 0.029
R13330 vss.n1190 vss.n1187 0.029
R13331 vss.n360 vss.n357 0.029
R13332 vss.n255 vss.n248 0.029
R13333 vss.n59 vss.n58 0.029
R13334 vss.n84 vss.n83 0.029
R13335 vss.n979 vss.n978 0.029
R13336 vss.n109 vss.n108 0.029
R13337 vss.n134 vss.n133 0.029
R13338 vss.n888 vss.n885 0.029
R13339 vss.n832 vss.n831 0.029
R13340 vss.n761 vss.n760 0.029
R13341 vss.n420 vss.n419 0.029
R13342 vss.n576 vss.n573 0.029
R13343 vss.n520 vss.n519 0.029
R13344 vss.n493 vss.n492 0.029
R13345 vss.n30 vss.n28 0.029
R13346 vss.n1099 vss.n1098 0.028
R13347 vss.n1404 vss.n1400 0.028
R13348 vss.n653 vss.n652 0.028
R13349 vss.n322 vss.n318 0.028
R13350 vss.n210 vss.n202 0.028
R13351 vss.n1825 vss.n1823 0.027
R13352 vss.n1545 vss.n1543 0.027
R13353 vss.n1666 vss.n1664 0.027
R13354 vss.n899 vss.n897 0.027
R13355 vss.n587 vss.n585 0.027
R13356 vss.n695 vss.n694 0.027
R13357 vss.n716 vss.n715 0.027
R13358 vss.n1148 vss.n1147 0.027
R13359 vss.n652 vss.n651 0.026
R13360 vss.n715 vss.n663 0.026
R13361 vss.n681 vss.n678 0.025
R13362 vss.n1821 vss.n1814 0.024
R13363 vss.n1541 vss.n1538 0.024
R13364 vss.n1662 vss.n1655 0.024
R13365 vss.n1381 vss.n1378 0.024
R13366 vss.n1385 vss.n1383 0.024
R13367 vss.n1299 vss.n1296 0.024
R13368 vss.n1303 vss.n1301 0.024
R13369 vss.n1197 vss.n1194 0.024
R13370 vss.n1201 vss.n1199 0.024
R13371 vss.n367 vss.n364 0.024
R13372 vss.n371 vss.n369 0.024
R13373 vss.n266 vss.n259 0.024
R13374 vss.n270 vss.n268 0.024
R13375 vss.n895 vss.n892 0.024
R13376 vss.n583 vss.n580 0.024
R13377 vss.n1338 vss.n1309 0.024
R13378 vss.n1238 vss.n1207 0.024
R13379 vss.n1481 vss.n1480 0.023
R13380 vss.n1889 vss.n1888 0.023
R13381 vss.n1583 vss.n1582 0.023
R13382 vss.n1730 vss.n1729 0.023
R13383 vss.n683 vss.n682 0.023
R13384 vss.n720 vss.n719 0.022
R13385 vss.n662 vss.n661 0.022
R13386 vss.n1814 vss.n1812 0.021
R13387 vss.n1538 vss.n1536 0.021
R13388 vss.n1655 vss.n1653 0.021
R13389 vss.n1417 vss.n1416 0.021
R13390 vss.n1406 vss.n1405 0.021
R13391 vss.n1378 vss.n1376 0.021
R13392 vss.n1386 vss.n1385 0.021
R13393 vss.n1336 vss.n1335 0.021
R13394 vss.n1325 vss.n1324 0.021
R13395 vss.n1296 vss.n1294 0.021
R13396 vss.n1304 vss.n1303 0.021
R13397 vss.n1194 vss.n1192 0.021
R13398 vss.n1202 vss.n1201 0.021
R13399 vss.n1236 vss.n1235 0.021
R13400 vss.n1225 vss.n1224 0.021
R13401 vss.n1118 vss.n1114 0.021
R13402 vss.n1101 vss.n1100 0.021
R13403 vss.n364 vss.n362 0.021
R13404 vss.n372 vss.n371 0.021
R13405 vss.n335 vss.n334 0.021
R13406 vss.n324 vss.n323 0.021
R13407 vss.n307 vss.n303 0.021
R13408 vss.n293 vss.n292 0.021
R13409 vss.n259 vss.n257 0.021
R13410 vss.n271 vss.n270 0.021
R13411 vss.n226 vss.n225 0.021
R13412 vss.n212 vss.n211 0.021
R13413 vss.n892 vss.n890 0.021
R13414 vss.n580 vss.n578 0.021
R13415 vss.n28 vss.n27 0.021
R13416 vss.n692 vss.n688 0.021
R13417 vss.n714 vss.n706 0.021
R13418 vss.n660 vss.n659 0.021
R13419 vss.n1056 vss.n1055 0.021
R13420 vss.n26 vss.n25 0.021
R13421 vss.n1936 vss.n1935 0.02
R13422 vss.n654 vss.n653 0.02
R13423 vss.n1474 vss.n1469 0.019
R13424 vss.n1832 vss.n1825 0.019
R13425 vss.n1779 vss.n1770 0.019
R13426 vss.n1548 vss.n1545 0.019
R13427 vss.n1507 vss.n1502 0.019
R13428 vss.n1673 vss.n1666 0.019
R13429 vss.n1620 vss.n1611 0.019
R13430 vss.n902 vss.n899 0.019
R13431 vss.n951 vss.n946 0.019
R13432 vss.n822 vss.n815 0.019
R13433 vss.n472 vss.n465 0.019
R13434 vss.n590 vss.n587 0.019
R13435 vss.n639 vss.n634 0.019
R13436 vss.n684 vss.n683 0.019
R13437 vss.n706 vss.n705 0.019
R13438 vss.n62 vss.n61 0.019
R13439 vss.n982 vss.n981 0.019
R13440 vss.n112 vss.n111 0.019
R13441 vss.n839 vss.n838 0.019
R13442 vss.n527 vss.n526 0.019
R13443 vss.n496 vss.n495 0.019
R13444 vss.n1899 vss.n1782 0.019
R13445 vss.n1589 vss.n1510 0.019
R13446 vss.n1740 vss.n1623 0.019
R13447 vss.n1486 vss.n1477 0.019
R13448 vss.n1419 vss.n1391 0.018
R13449 vss.n378 vss.n377 0.018
R13450 vss.n280 vss.n279 0.018
R13451 vss.n1391 vss.n1386 0.017
R13452 vss.n1309 vss.n1304 0.017
R13453 vss.n1207 vss.n1202 0.017
R13454 vss.n377 vss.n372 0.017
R13455 vss.n279 vss.n271 0.017
R13456 vss.n382 vss.n381 0.017
R13457 vss.n391 vss.n390 0.017
R13458 vss.n67 vss.n66 0.017
R13459 vss.n92 vss.n91 0.017
R13460 vss.n87 vss.n86 0.017
R13461 vss.n987 vss.n986 0.017
R13462 vss.n117 vss.n116 0.017
R13463 vss.n142 vss.n141 0.017
R13464 vss.n137 vss.n136 0.017
R13465 vss.n848 vss.n847 0.017
R13466 vss.n777 vss.n776 0.017
R13467 vss.n772 vss.n771 0.017
R13468 vss.n428 vss.n427 0.017
R13469 vss.n423 vss.n422 0.017
R13470 vss.n536 vss.n535 0.017
R13471 vss.n501 vss.n500 0.017
R13472 vss.n37 vss.n36 0.017
R13473 vss.n702 vss.n697 0.017
R13474 vss.n658 vss.n657 0.017
R13475 vss.n1134 vss.n1133 0.017
R13476 vss.n1421 vss.n1420 0.017
R13477 vss.n1803 vss.n1801 0.016
R13478 vss.n1531 vss.n1529 0.016
R13479 vss.n1644 vss.n1642 0.016
R13480 vss.n1925 vss.n1924 0.016
R13481 vss.n1921 vss.n1920 0.016
R13482 vss.n1371 vss.n1369 0.016
R13483 vss.n1289 vss.n1287 0.016
R13484 vss.n1187 vss.n1185 0.016
R13485 vss.n357 vss.n355 0.016
R13486 vss.n248 vss.n246 0.016
R13487 vss.n885 vss.n883 0.016
R13488 vss.n573 vss.n571 0.016
R13489 vss.n1465 vss.n1464 0.015
R13490 vss.n1766 vss.n1765 0.015
R13491 vss.n1498 vss.n1497 0.015
R13492 vss.n1607 vss.n1598 0.015
R13493 vss.n697 vss.n696 0.015
R13494 vss.n703 vss.n702 0.015
R13495 vss.n657 vss.n656 0.015
R13496 vss.n18 vss.n17 0.015
R13497 vss.n1342 vss.n1341 0.014
R13498 vss.n1475 vss.n1474 0.013
R13499 vss.n1843 vss.n1836 0.013
R13500 vss.n1780 vss.n1779 0.013
R13501 vss.n1555 vss.n1552 0.013
R13502 vss.n1508 vss.n1507 0.013
R13503 vss.n1684 vss.n1677 0.013
R13504 vss.n1621 vss.n1620 0.013
R13505 vss.n1947 vss.n1946 0.013
R13506 vss.n1949 vss.n1948 0.013
R13507 vss.n1945 vss.n1943 0.013
R13508 vss.n1945 vss.n1944 0.013
R13509 vss.n1952 vss.n1951 0.013
R13510 vss.n1954 vss.n1953 0.013
R13511 vss.n1456 vss.n1454 0.013
R13512 vss.n1456 vss.n1455 0.013
R13513 vss.n1453 vss.n1450 0.013
R13514 vss.n1415 vss.n1414 0.013
R13515 vss.n1334 vss.n1333 0.013
R13516 vss.n1234 vss.n1233 0.013
R13517 vss.n1113 vss.n1112 0.013
R13518 vss.n333 vss.n332 0.013
R13519 vss.n302 vss.n301 0.013
R13520 vss.n224 vss.n223 0.013
R13521 vss.n72 vss.n71 0.013
R13522 vss.n97 vss.n96 0.013
R13523 vss.n992 vss.n991 0.013
R13524 vss.n122 vss.n121 0.013
R13525 vss.n150 vss.n149 0.013
R13526 vss.n909 vss.n906 0.013
R13527 vss.n940 vss.n938 0.013
R13528 vss.n946 vss.n945 0.013
R13529 vss.n952 vss.n951 0.013
R13530 vss.n809 vss.n807 0.013
R13531 vss.n815 vss.n814 0.013
R13532 vss.n823 vss.n822 0.013
R13533 vss.n459 vss.n457 0.013
R13534 vss.n465 vss.n464 0.013
R13535 vss.n473 vss.n472 0.013
R13536 vss.n597 vss.n594 0.013
R13537 vss.n628 vss.n626 0.013
R13538 vss.n634 vss.n633 0.013
R13539 vss.n640 vss.n639 0.013
R13540 vss.n511 vss.n510 0.013
R13541 vss.n44 vss.n43 0.013
R13542 vss.n1045 vss.n1044 0.013
R13543 vss.n1044 vss.n1043 0.013
R13544 vss.n1043 vss.n1042 0.013
R13545 vss.n1042 vss.n1041 0.013
R13546 vss.n1041 vss.n1040 0.013
R13547 vss.n1040 vss.n1039 0.013
R13548 vss.n1039 vss.n1038 0.013
R13549 vss.n1038 vss.n1037 0.013
R13550 vss.n1037 vss.n1036 0.013
R13551 vss.n1036 vss.n1035 0.013
R13552 vss.n1035 vss.n1034 0.013
R13553 vss.n1032 vss.n1031 0.013
R13554 vss.n1031 vss.n1030 0.013
R13555 vss.n1030 vss.n1029 0.013
R13556 vss.n1029 vss.n1028 0.013
R13557 vss.n1028 vss.n1027 0.013
R13558 vss.n1027 vss.n1026 0.013
R13559 vss.n1026 vss.n1025 0.013
R13560 vss.n1054 vss.n1053 0.013
R13561 vss.n1051 vss.n1049 0.013
R13562 vss.n1051 vss.n1050 0.013
R13563 vss.n677 vss.n676 0.013
R13564 vss.n1071 vss.n1070 0.013
R13565 vss.n1072 vss.n1071 0.013
R13566 vss.n1075 vss.n1074 0.013
R13567 vss.n1076 vss.n1075 0.013
R13568 vss.n1242 vss.n1076 0.013
R13569 vss.n1243 vss.n1242 0.013
R13570 vss.n1244 vss.n1243 0.013
R13571 vss.n1438 vss.n1244 0.013
R13572 vss.n1438 vss.n1437 0.013
R13573 vss.n1435 vss.n1434 0.013
R13574 vss.n1434 vss.n1433 0.013
R13575 vss.n1433 vss.n1432 0.013
R13576 vss.n1430 vss.n1429 0.013
R13577 vss.n1901 vss.n1900 0.012
R13578 vss.n1046 vss.n1045 0.012
R13579 vss.n655 vss.n654 0.012
R13580 vss.n1919 vss.n1918 0.012
R13581 vss.n1923 vss.n1922 0.012
R13582 vss.n1935 vss.n1934 0.012
R13583 vss.n393 vss.n392 0.011
R13584 vss.n748 vss.n747 0.011
R13585 vss.n1132 vss.n1131 0.011
R13586 vss.n1452 vss.n1451 0.011
R13587 vss.n1407 vss.n1406 0.011
R13588 vss.n1326 vss.n1325 0.011
R13589 vss.n1226 vss.n1225 0.011
R13590 vss.n1102 vss.n1101 0.011
R13591 vss.n325 vss.n324 0.011
R13592 vss.n294 vss.n293 0.011
R13593 vss.n213 vss.n212 0.011
R13594 vss.n66 vss.n65 0.011
R13595 vss.n60 vss.n59 0.011
R13596 vss.n85 vss.n84 0.011
R13597 vss.n986 vss.n985 0.011
R13598 vss.n980 vss.n979 0.011
R13599 vss.n116 vss.n115 0.011
R13600 vss.n110 vss.n109 0.011
R13601 vss.n135 vss.n134 0.011
R13602 vss.n847 vss.n842 0.011
R13603 vss.n837 vss.n832 0.011
R13604 vss.n770 vss.n761 0.011
R13605 vss.n421 vss.n420 0.011
R13606 vss.n535 vss.n530 0.011
R13607 vss.n525 vss.n520 0.011
R13608 vss.n500 vss.n499 0.011
R13609 vss.n494 vss.n493 0.011
R13610 vss.n27 vss.n26 0.011
R13611 vss.n688 vss.n687 0.011
R13612 vss.n693 vss.n692 0.011
R13613 vss.n694 vss.n693 0.011
R13614 vss.n714 vss.n713 0.011
R13615 vss.n1070 vss.n1069 0.011
R13616 vss.n1074 vss.n1073 0.011
R13617 vss.n1436 vss.n1435 0.011
R13618 vss.n1429 vss.n1428 0.011
R13619 vss.n1932 vss.n1931 0.01
R13620 vss.n1034 vss.n1033 0.01
R13621 vss.n1025 vss.n1024 0.01
R13622 vss.n661 vss.n660 0.01
R13623 vss.n47 vss.n46 0.01
R13624 vss.n1345 vss.n1344 0.01
R13625 vss.n736 vss.n735 0.009
R13626 vss.n394 vss.n183 0.009
R13627 vss.n746 vss.n153 0.009
R13628 vss.n1466 vss.n1465 0.009
R13629 vss.n1485 vss.n1481 0.009
R13630 vss.n1898 vss.n1889 0.009
R13631 vss.n1588 vss.n1583 0.009
R13632 vss.n1739 vss.n1730 0.009
R13633 vss.n1416 vss.n1415 0.009
R13634 vss.n1405 vss.n1404 0.009
R13635 vss.n1335 vss.n1334 0.009
R13636 vss.n1324 vss.n1323 0.009
R13637 vss.n1235 vss.n1234 0.009
R13638 vss.n1224 vss.n1223 0.009
R13639 vss.n1114 vss.n1113 0.009
R13640 vss.n1100 vss.n1099 0.009
R13641 vss.n334 vss.n333 0.009
R13642 vss.n323 vss.n322 0.009
R13643 vss.n303 vss.n302 0.009
R13644 vss.n292 vss.n291 0.009
R13645 vss.n225 vss.n224 0.009
R13646 vss.n211 vss.n210 0.009
R13647 vss.n1015 vss.n1014 0.009
R13648 vss.n1431 vss.n1430 0.009
R13649 vss.n90 vss.n89 0.009
R13650 vss.n140 vss.n139 0.009
R13651 vss.n775 vss.n774 0.009
R13652 vss.n426 vss.n425 0.009
R13653 vss.n1768 vss.n1767 0.009
R13654 vss.n1500 vss.n1499 0.009
R13655 vss.n1609 vss.n1608 0.009
R13656 vss.n1911 vss.n1910 0.009
R13657 vss.n1912 vss.n1911 0.009
R13658 vss.n387 vss.n386 0.009
R13659 vss.n386 vss.n385 0.009
R13660 vss.n646 vss.n645 0.009
R13661 vss.n642 vss.n517 0.009
R13662 vss.n482 vss.n481 0.009
R13663 vss.n1004 vss.n1003 0.009
R13664 vss.n998 vss.n997 0.009
R13665 vss.n968 vss.n967 0.009
R13666 vss.n964 vss.n963 0.009
R13667 vss.n958 vss.n957 0.009
R13668 vss.n954 vss.n829 0.009
R13669 vss.n750 vss.n749 0.009
R13670 vss.n513 vss.n482 0.009
R13671 vss.n517 vss.n516 0.009
R13672 vss.n647 vss.n646 0.009
R13673 vss.n825 vss.n750 0.009
R13674 vss.n829 vss.n828 0.009
R13675 vss.n959 vss.n958 0.009
R13676 vss.n994 vss.n968 0.009
R13677 vss.n963 vss.n962 0.009
R13678 vss.n999 vss.n998 0.009
R13679 vss.n1003 vss.n1002 0.009
R13680 vss.n1139 vss.n1138 0.009
R13681 vss.n1241 vss.n1240 0.009
R13682 vss.n1343 vss.n1342 0.009
R13683 vss.n1138 vss.n1137 0.009
R13684 vss.n1344 vss.n1343 0.009
R13685 vss.n1240 vss.n1239 0.009
R13686 vss.n183 vss.n182 0.009
R13687 vss.n153 vss.n152 0.009
R13688 vss.n1914 vss.n1913 0.008
R13689 vss.n1913 vss.n1912 0.008
R13690 vss.n381 vss.n380 0.008
R13691 vss.n384 vss.n383 0.008
R13692 vss.n390 vss.n389 0.008
R13693 vss.n389 vss.n388 0.008
R13694 vss.n385 vss.n384 0.008
R13695 vss.n380 vss.n379 0.008
R13696 vss.n648 vss.n647 0.008
R13697 vss.n643 vss.n642 0.008
R13698 vss.n515 vss.n514 0.008
R13699 vss.n46 vss.n19 0.008
R13700 vss.n1005 vss.n1004 0.008
R13701 vss.n1000 vss.n999 0.008
R13702 vss.n996 vss.n995 0.008
R13703 vss.n965 vss.n964 0.008
R13704 vss.n960 vss.n959 0.008
R13705 vss.n955 vss.n954 0.008
R13706 vss.n827 vss.n826 0.008
R13707 vss.n644 vss.n643 0.008
R13708 vss.n649 vss.n648 0.008
R13709 vss.n956 vss.n955 0.008
R13710 vss.n961 vss.n960 0.008
R13711 vss.n966 vss.n965 0.008
R13712 vss.n826 vss.n825 0.008
R13713 vss.n995 vss.n994 0.008
R13714 vss.n1001 vss.n1000 0.008
R13715 vss.n514 vss.n513 0.008
R13716 vss.n19 vss.n18 0.008
R13717 vss.n1006 vss.n1005 0.008
R13718 vss.n1137 vss.n1136 0.008
R13719 vss.n1422 vss.n1421 0.008
R13720 vss.n1136 vss.n1135 0.008
R13721 vss.n1423 vss.n1422 0.008
R13722 vss.n1854 vss.n1847 0.008
R13723 vss.n1885 vss.n1883 0.008
R13724 vss.n1562 vss.n1559 0.008
R13725 vss.n1579 vss.n1577 0.008
R13726 vss.n1695 vss.n1688 0.008
R13727 vss.n1726 vss.n1724 0.008
R13728 vss.n916 vss.n913 0.008
R13729 vss.n933 vss.n931 0.008
R13730 vss.n798 vss.n796 0.008
R13731 vss.n448 vss.n446 0.008
R13732 vss.n604 vss.n601 0.008
R13733 vss.n621 vss.n619 0.008
R13734 vss.n1767 vss.n1766 0.008
R13735 vss.n1499 vss.n1498 0.008
R13736 vss.n1608 vss.n1607 0.008
R13737 vss.n1241 vss.n1149 0.008
R13738 vss.n1149 vss.n1148 0.008
R13739 vss.n1467 vss.n1466 0.008
R13740 vss.n670 vss.n669 0.007
R13741 vss.n682 vss.n681 0.007
R13742 vss.n1144 vss.n1143 0.007
R13743 vss.n1062 vss.n1061 0.007
R13744 vss.n36 vss.n35 0.007
R13745 vss.n1924 vss.n1923 0.006
R13746 vss.n1920 vss.n1919 0.006
R13747 vss.n1933 vss.n1932 0.006
R13748 vss.n1929 vss.n1928 0.006
R13749 vss.n48 vss.n47 0.006
R13750 vss.n1427 vss.n1426 0.006
R13751 vss.n776 vss.n775 0.006
R13752 vss.n141 vss.n140 0.006
R13753 vss.n427 vss.n426 0.006
R13754 vss.n91 vss.n90 0.006
R13755 vss.n394 vss.n393 0.006
R13756 vss.n747 vss.n746 0.006
R13757 vss.n1133 vss.n1132 0.006
R13758 vss.n1934 vss.n1933 0.005
R13759 vss.n1794 vss.n1792 0.005
R13760 vss.n1521 vss.n1519 0.005
R13761 vss.n1634 vss.n1632 0.005
R13762 vss.n1160 vss.n1158 0.005
R13763 vss.n1177 vss.n1175 0.005
R13764 vss.n1254 vss.n1252 0.005
R13765 vss.n1279 vss.n1277 0.005
R13766 vss.n1267 vss.n1260 0.005
R13767 vss.n1361 vss.n1359 0.005
R13768 vss.n348 vss.n346 0.005
R13769 vss.n239 vss.n237 0.005
R13770 vss.n859 vss.n857 0.005
R13771 vss.n875 vss.n873 0.005
R13772 vss.n547 vss.n545 0.005
R13773 vss.n563 vss.n561 0.005
R13774 vss.n678 vss.n677 0.005
R13775 vss.n651 vss.n650 0.005
R13776 vss.n727 vss.n725 0.005
R13777 vss.n739 vss.n738 0.004
R13778 vss.n1486 vss.n1485 0.004
R13779 vss.n1589 vss.n1588 0.004
R13780 vss.n1740 vss.n1739 0.004
R13781 vss.n1899 vss.n1898 0.004
R13782 vss.n1448 vss.n1447 0.004
R13783 vss.n1952 vss.n1950 0.004
R13784 vss.n1 vss.n0 0.004
R13785 vss.n168 vss.n167 0.004
R13786 vss.n741 vss.n740 0.004
R13787 vss.n177 vss.n176 0.004
R13788 vss.n399 vss.n398 0.004
R13789 vss.n725 vss.n724 0.004
R13790 vss.n730 vss.n729 0.004
R13791 vss.n1432 vss.n1431 0.004
R13792 vss.n43 vss.n40 0.004
R13793 vss.n738 vss.n400 0.004
R13794 vss.n731 vss.n730 0.004
R13795 vss.n178 vss.n177 0.004
R13796 vss.n738 vss.n169 0.003
R13797 vss.n65 vss.n64 0.003
R13798 vss.n86 vss.n85 0.003
R13799 vss.n985 vss.n984 0.003
R13800 vss.n115 vss.n114 0.003
R13801 vss.n136 vss.n135 0.003
R13802 vss.n842 vss.n841 0.003
R13803 vss.n771 vss.n770 0.003
R13804 vss.n422 vss.n421 0.003
R13805 vss.n530 vss.n529 0.003
R13806 vss.n499 vss.n498 0.003
R13807 vss.n1033 vss.n1032 0.003
R13808 vss.n1024 vss.n1023 0.003
R13809 vss.n668 vss.n667 0.003
R13810 vss.n1067 vss.n1066 0.003
R13811 vss.n5 vss.n4 0.002
R13812 vss.n1048 vss.n10 0.002
R13813 vss.n1865 vss.n1858 0.002
R13814 vss.n1874 vss.n1872 0.002
R13815 vss.n1568 vss.n1566 0.002
R13816 vss.n1572 vss.n1570 0.002
R13817 vss.n1706 vss.n1699 0.002
R13818 vss.n1715 vss.n1713 0.002
R13819 vss.n1956 vss.n1955 0.002
R13820 vss.n1453 vss.n1452 0.002
R13821 vss.n1095 vss.n1093 0.002
R13822 vss.n199 vss.n197 0.002
R13823 vss.n922 vss.n920 0.002
R13824 vss.n926 vss.n924 0.002
R13825 vss.n787 vss.n785 0.002
R13826 vss.n437 vss.n435 0.002
R13827 vss.n610 vss.n608 0.002
R13828 vss.n614 vss.n612 0.002
R13829 vss.n1073 vss.n1072 0.002
R13830 vss.n1437 vss.n1436 0.002
R13831 vss.n1428 vss.n1427 0.002
R13832 vss.n61 vss.n60 0.002
R13833 vss.n981 vss.n980 0.002
R13834 vss.n111 vss.n110 0.002
R13835 vss.n838 vss.n837 0.002
R13836 vss.n526 vss.n525 0.002
R13837 vss.n495 vss.n494 0.002
R13838 vss.n1446 vss.n1445 0.002
R13839 vss.n1957 vss.n1446 0.002
R13840 vss.n169 vss.n168 0.002
R13841 vss.n1068 vss.n1067 0.001
R13842 vss.n1069 vss.n1068 0.001
R13843 vss.n1449 vss.n1448 0.001
R13844 vss.n2 vss.n1 0.001
R13845 vss.n735 vss.n727 0.001
R13846 vss.n738 vss.n178 0.001
R13847 vss.n735 vss.n731 0.001
R13848 vss.n400 vss.n399 0.001
R13849 vss.n1418 vss.n1417 0.001
R13850 vss.n1408 vss.n1407 0.001
R13851 vss.n1337 vss.n1336 0.001
R13852 vss.n1327 vss.n1326 0.001
R13853 vss.n1237 vss.n1236 0.001
R13854 vss.n1227 vss.n1226 0.001
R13855 vss.n1119 vss.n1118 0.001
R13856 vss.n1103 vss.n1102 0.001
R13857 vss.n336 vss.n335 0.001
R13858 vss.n326 vss.n325 0.001
R13859 vss.n308 vss.n307 0.001
R13860 vss.n295 vss.n294 0.001
R13861 vss.n227 vss.n226 0.001
R13862 vss.n214 vss.n213 0.001
R13863 vss.n1047 vss.n1046 0.001
R13864 vss.n4 vss.n3 0.001
R13865 vss.n1341 vss.n1340 0.001
R13866 vss.n1440 vss.n1439 0.001
R13867 vss.n1439 vss.n1058 0.001
R13868 vss.n1055 vss.n1048 0.001
R13869 vss.n740 vss.n739 0.001
R13870 vss.n719 vss.n717 0.001
R13871 vss.n1442 vss.n1441 0.001
R13872 vss.n1057 vss.n1056 0.001
R13873 vss.n10 vss.n9 0.001
R13874 vss.n8 vss.n7 0.001
R13875 vss.n1441 vss.n1440 0.001
R13876 vss.n1058 vss.n1057 0.001
R13877 vss.n9 vss.n8 0.001
R13878 vss.n7 vss.n6 0.001
R13879 vss.n1445 vss.n1444 0.001
R13880 vss.n1444 vss.n1443 0.001
R13881 a_2151_4783.n51 a_2151_4783.t8 60.25
R13882 a_2151_4783.n72 a_2151_4783.t9 60.25
R13883 a_2151_4783.n94 a_2151_4783.t6 60.25
R13884 a_2151_4783.n39 a_2151_4783.t4 60.25
R13885 a_2151_4783.n5 a_2151_4783.n60 9.3
R13886 a_2151_4783.n7 a_2151_4783.n64 9.3
R13887 a_2151_4783.n8 a_2151_4783.n82 9.3
R13888 a_2151_4783.n10 a_2151_4783.n86 9.3
R13889 a_2151_4783.n11 a_2151_4783.n104 9.3
R13890 a_2151_4783.n12 a_2151_4783.n48 9.3
R13891 a_2151_4783.n12 a_2151_4783.n47 9.3
R13892 a_2151_4783.n12 a_2151_4783.n46 9.3
R13893 a_2151_4783.n46 a_2151_4783.n45 9.3
R13894 a_2151_4783.n11 a_2151_4783.n103 9.3
R13895 a_2151_4783.n11 a_2151_4783.n102 9.3
R13896 a_2151_4783.n102 a_2151_4783.n101 9.3
R13897 a_2151_4783.n10 a_2151_4783.n87 9.3
R13898 a_2151_4783.n10 a_2151_4783.n93 9.3
R13899 a_2151_4783.n93 a_2151_4783.n92 9.3
R13900 a_2151_4783.n8 a_2151_4783.n81 9.3
R13901 a_2151_4783.n8 a_2151_4783.n80 9.3
R13902 a_2151_4783.n80 a_2151_4783.n79 9.3
R13903 a_2151_4783.n7 a_2151_4783.n65 9.3
R13904 a_2151_4783.n7 a_2151_4783.n71 9.3
R13905 a_2151_4783.n71 a_2151_4783.n70 9.3
R13906 a_2151_4783.n5 a_2151_4783.n58 9.3
R13907 a_2151_4783.n58 a_2151_4783.n57 9.3
R13908 a_2151_4783.n5 a_2151_4783.n59 9.3
R13909 a_2151_4783.n0 a_2151_4783.n109 9.3
R13910 a_2151_4783.n95 a_2151_4783.n94 8.764
R13911 a_2151_4783.n73 a_2151_4783.n72 8.764
R13912 a_2151_4783.n44 a_2151_4783.n43 7.453
R13913 a_2151_4783.n100 a_2151_4783.n99 7.453
R13914 a_2151_4783.n91 a_2151_4783.n90 7.453
R13915 a_2151_4783.n78 a_2151_4783.n77 7.453
R13916 a_2151_4783.n69 a_2151_4783.n68 7.453
R13917 a_2151_4783.n56 a_2151_4783.n55 7.453
R13918 a_2151_4783.n40 a_2151_4783.n39 6.803
R13919 a_2151_4783.n52 a_2151_4783.n51 6.8
R13920 a_2151_4783.n111 a_2151_4783.n110 6.316
R13921 a_2151_4783.n42 a_2151_4783.n41 5.647
R13922 a_2151_4783.n98 a_2151_4783.n97 5.647
R13923 a_2151_4783.n89 a_2151_4783.n88 5.647
R13924 a_2151_4783.n76 a_2151_4783.n75 5.647
R13925 a_2151_4783.n67 a_2151_4783.n66 5.647
R13926 a_2151_4783.n54 a_2151_4783.n53 5.647
R13927 a_2151_4783.n112 a_2151_4783.t5 5.539
R13928 a_2151_4783.t7 a_2151_4783.n112 5.539
R13929 a_2151_4783.n0 a_2151_4783.n108 4.955
R13930 a_2151_4783.n62 a_2151_4783.n61 4.735
R13931 a_2151_4783.n50 a_2151_4783.n49 4.735
R13932 a_2151_4783.n106 a_2151_4783.n105 4.735
R13933 a_2151_4783.n9 a_2151_4783.n85 4.735
R13934 a_2151_4783.n84 a_2151_4783.n83 4.735
R13935 a_2151_4783.n6 a_2151_4783.n63 4.735
R13936 a_2151_4783.n1 a_2151_4783.n13 4.662
R13937 a_2151_4783.n96 a_2151_4783.n95 4.65
R13938 a_2151_4783.n74 a_2151_4783.n73 4.65
R13939 a_2151_4783.n4 a_2151_4783.n31 4.5
R13940 a_2151_4783.n4 a_2151_4783.n28 4.5
R13941 a_2151_4783.n2 a_2151_4783.n20 4.5
R13942 a_2151_4783.n3 a_2151_4783.n23 4.5
R13943 a_2151_4783.n0 a_2151_4783.n38 4.5
R13944 a_2151_4783.n1 a_2151_4783.n36 4.5
R13945 a_2151_4783.n1 a_2151_4783.n15 4.5
R13946 a_2151_4783.n28 a_2151_4783.n27 4.141
R13947 a_2151_4783.n23 a_2151_4783.n22 4.141
R13948 a_2151_4783.n15 a_2151_4783.n14 3.764
R13949 a_2151_4783.n5 a_2151_4783.n52 3.427
R13950 a_2151_4783.n12 a_2151_4783.n40 3.426
R13951 a_2151_4783.n38 a_2151_4783.n37 3.388
R13952 a_2151_4783.n32 a_2151_4783.t1 3.306
R13953 a_2151_4783.n32 a_2151_4783.t0 3.306
R13954 a_2151_4783.n16 a_2151_4783.t3 3.306
R13955 a_2151_4783.n16 a_2151_4783.t2 3.306
R13956 a_2151_4783.n36 a_2151_4783.n35 3.011
R13957 a_2151_4783.n30 a_2151_4783.n29 2.258
R13958 a_2151_4783.n19 a_2151_4783.n18 2.258
R13959 a_2151_4783.n111 a_2151_4783.n1 1.503
R13960 a_2151_4783.n17 a_2151_4783.n16 1.467
R13961 a_2151_4783.n45 a_2151_4783.n44 0.993
R13962 a_2151_4783.n101 a_2151_4783.n100 0.993
R13963 a_2151_4783.n92 a_2151_4783.n91 0.993
R13964 a_2151_4783.n79 a_2151_4783.n78 0.993
R13965 a_2151_4783.n70 a_2151_4783.n69 0.993
R13966 a_2151_4783.n57 a_2151_4783.n56 0.993
R13967 a_2151_4783.n34 a_2151_4783.n25 0.92
R13968 a_2151_4783.n46 a_2151_4783.n42 0.752
R13969 a_2151_4783.n102 a_2151_4783.n98 0.752
R13970 a_2151_4783.n93 a_2151_4783.n89 0.752
R13971 a_2151_4783.n80 a_2151_4783.n76 0.752
R13972 a_2151_4783.n71 a_2151_4783.n67 0.752
R13973 a_2151_4783.n58 a_2151_4783.n54 0.752
R13974 a_2151_4783.n13 a_2151_4783.n3 0.701
R13975 a_2151_4783.n13 a_2151_4783.n34 0.699
R13976 a_2151_4783.n3 a_2151_4783.n24 0.602
R13977 a_2151_4783.n25 a_2151_4783.n33 0.593
R13978 a_2151_4783.n4 a_2151_4783.n32 2.109
R13979 a_2151_4783.n2 a_2151_4783.n17 0.552
R13980 a_2151_4783.n6 a_2151_4783.n62 0.456
R13981 a_2151_4783.n9 a_2151_4783.n84 0.456
R13982 a_2151_4783.n112 a_2151_4783.n111 0.4
R13983 a_2151_4783.n28 a_2151_4783.n26 0.376
R13984 a_2151_4783.n31 a_2151_4783.n30 0.376
R13985 a_2151_4783.n23 a_2151_4783.n21 0.376
R13986 a_2151_4783.n20 a_2151_4783.n19 0.376
R13987 a_2151_4783.n0 a_2151_4783.n107 0.353
R13988 a_2151_4783.n1 a_2151_4783.n0 0.302
R13989 a_2151_4783.n3 a_2151_4783.n2 0.279
R13990 a_2151_4783.n107 a_2151_4783.n50 0.228
R13991 a_2151_4783.n107 a_2151_4783.n106 0.228
R13992 a_2151_4783.n50 a_2151_4783.n12 0.203
R13993 a_2151_4783.n106 a_2151_4783.n11 0.203
R13994 a_2151_4783.n10 a_2151_4783.n9 0.203
R13995 a_2151_4783.n84 a_2151_4783.n8 0.203
R13996 a_2151_4783.n7 a_2151_4783.n6 0.203
R13997 a_2151_4783.n62 a_2151_4783.n5 0.203
R13998 a_2151_4783.n25 a_2151_4783.n4 0.202
R13999 a_2151_4783.n11 a_2151_4783.n96 0.19
R14000 a_2151_4783.n96 a_2151_4783.n10 0.19
R14001 a_2151_4783.n8 a_2151_4783.n74 0.19
R14002 a_2151_4783.n74 a_2151_4783.n7 0.19
R14003 a_2551_4880.n76 a_2551_4880.t2 60.25
R14004 a_2551_4880.n53 a_2551_4880.t7 60.25
R14005 a_2551_4880.n30 a_2551_4880.t6 60.25
R14006 a_2551_4880.n90 a_2551_4880.t0 60.25
R14007 a_2551_4880.n140 a_2551_4880.n10 10.325
R14008 a_2551_4880.n140 a_2551_4880.n11 9.572
R14009 a_2551_4880.n7 a_2551_4880.n98 9.3
R14010 a_2551_4880.n100 a_2551_4880.n99 9.3
R14011 a_2551_4880.n7 a_2551_4880.n97 9.3
R14012 a_2551_4880.n97 a_2551_4880.n96 9.3
R14013 a_2551_4880.n64 a_2551_4880.n63 9.3
R14014 a_2551_4880.n1 a_2551_4880.n45 9.3
R14015 a_2551_4880.n40 a_2551_4880.n39 9.3
R14016 a_2551_4880.n0 a_2551_4880.n38 9.3
R14017 a_2551_4880.n0 a_2551_4880.n37 9.3
R14018 a_2551_4880.n37 a_2551_4880.n36 9.3
R14019 a_2551_4880.n2 a_2551_4880.n46 9.3
R14020 a_2551_4880.n2 a_2551_4880.n52 9.3
R14021 a_2551_4880.n52 a_2551_4880.n51 9.3
R14022 a_2551_4880.n3 a_2551_4880.n62 9.3
R14023 a_2551_4880.n3 a_2551_4880.n61 9.3
R14024 a_2551_4880.n61 a_2551_4880.n60 9.3
R14025 a_2551_4880.n4 a_2551_4880.n68 9.3
R14026 a_2551_4880.n5 a_2551_4880.n75 9.3
R14027 a_2551_4880.n75 a_2551_4880.n74 9.3
R14028 a_2551_4880.n5 a_2551_4880.n69 9.3
R14029 a_2551_4880.n6 a_2551_4880.n84 9.3
R14030 a_2551_4880.n84 a_2551_4880.n83 9.3
R14031 a_2551_4880.n87 a_2551_4880.n86 9.3
R14032 a_2551_4880.n6 a_2551_4880.n85 9.3
R14033 a_2551_4880.n112 a_2551_4880.n113 9.3
R14034 a_2551_4880.n110 a_2551_4880.n111 9.3
R14035 a_2551_4880.n108 a_2551_4880.n109 9.3
R14036 a_2551_4880.n106 a_2551_4880.n107 9.3
R14037 a_2551_4880.n105 a_2551_4880.n104 9.3
R14038 a_2551_4880.n54 a_2551_4880.n53 8.764
R14039 a_2551_4880.n77 a_2551_4880.n76 8.764
R14040 a_2551_4880.n35 a_2551_4880.n34 8.215
R14041 a_2551_4880.n50 a_2551_4880.n49 8.215
R14042 a_2551_4880.n59 a_2551_4880.n58 8.215
R14043 a_2551_4880.n95 a_2551_4880.n94 8.215
R14044 a_2551_4880.n73 a_2551_4880.n72 8.215
R14045 a_2551_4880.n82 a_2551_4880.n81 8.215
R14046 a_2551_4880.n140 a_2551_4880.n27 8.139
R14047 a_2551_4880.n140 a_2551_4880.n24 8.111
R14048 a_2551_4880.n140 a_2551_4880.n21 8.083
R14049 a_2551_4880.n140 a_2551_4880.n18 8.056
R14050 a_2551_4880.n133 a_2551_4880.n132 8.042
R14051 a_2551_4880.n140 a_2551_4880.n15 8.029
R14052 a_2551_4880.n140 a_2551_4880.n12 8.003
R14053 a_2551_4880.n31 a_2551_4880.n30 6.922
R14054 a_2551_4880.n91 a_2551_4880.n90 6.92
R14055 a_2551_4880.n33 a_2551_4880.n32 5.647
R14056 a_2551_4880.n48 a_2551_4880.n47 5.647
R14057 a_2551_4880.n57 a_2551_4880.n56 5.647
R14058 a_2551_4880.n93 a_2551_4880.n92 5.647
R14059 a_2551_4880.n71 a_2551_4880.n70 5.647
R14060 a_2551_4880.n80 a_2551_4880.n79 5.647
R14061 a_2551_4880.n122 a_2551_4880.n120 5.629
R14062 a_2551_4880.n127 a_2551_4880.t4 5.539
R14063 a_2551_4880.n127 a_2551_4880.t5 5.539
R14064 a_2551_4880.n101 a_2551_4880.n89 4.764
R14065 a_2551_4880.n67 a_2551_4880.n29 4.764
R14066 a_2551_4880.n88 a_2551_4880.n28 4.764
R14067 a_2551_4880.n42 a_2551_4880.n41 4.764
R14068 a_2551_4880.n44 a_2551_4880.n43 4.764
R14069 a_2551_4880.n66 a_2551_4880.n65 4.764
R14070 a_2551_4880.n55 a_2551_4880.n54 4.65
R14071 a_2551_4880.n78 a_2551_4880.n77 4.65
R14072 a_2551_4880.n9 a_2551_4880.n130 4.5
R14073 a_2551_4880.n8 a_2551_4880.n126 4.5
R14074 a_2551_4880.n135 a_2551_4880.n137 4.5
R14075 a_2551_4880.n134 a_2551_4880.n133 4.5
R14076 a_2551_4880.n117 a_2551_4880.n118 4.5
R14077 a_2551_4880.n114 a_2551_4880.n116 4.5
R14078 a_2551_4880.n14 a_2551_4880.n13 4.141
R14079 a_2551_4880.n130 a_2551_4880.n129 3.764
R14080 a_2551_4880.n7 a_2551_4880.n91 3.477
R14081 a_2551_4880.n0 a_2551_4880.n31 3.476
R14082 a_2551_4880.n126 a_2551_4880.n123 3.388
R14083 a_2551_4880.n17 a_2551_4880.n16 3.388
R14084 a_2551_4880.t3 a_2551_4880.n140 3.306
R14085 a_2551_4880.n140 a_2551_4880.t1 3.306
R14086 a_2551_4880.n126 a_2551_4880.n125 3.011
R14087 a_2551_4880.n130 a_2551_4880.n128 2.635
R14088 a_2551_4880.n20 a_2551_4880.n19 2.635
R14089 a_2551_4880.n137 a_2551_4880.n136 2.635
R14090 a_2551_4880.n116 a_2551_4880.n115 2.258
R14091 a_2551_4880.n9 a_2551_4880.n127 1.903
R14092 a_2551_4880.n23 a_2551_4880.n22 1.882
R14093 a_2551_4880.n140 a_2551_4880.n139 1.525
R14094 a_2551_4880.n26 a_2551_4880.n25 1.129
R14095 a_2551_4880.n36 a_2551_4880.n35 1.095
R14096 a_2551_4880.n51 a_2551_4880.n50 1.095
R14097 a_2551_4880.n60 a_2551_4880.n59 1.095
R14098 a_2551_4880.n96 a_2551_4880.n95 1.095
R14099 a_2551_4880.n74 a_2551_4880.n73 1.095
R14100 a_2551_4880.n83 a_2551_4880.n82 1.095
R14101 a_2551_4880.n139 a_2551_4880.n138 0.936
R14102 a_2551_4880.n37 a_2551_4880.n33 0.752
R14103 a_2551_4880.n52 a_2551_4880.n48 0.752
R14104 a_2551_4880.n61 a_2551_4880.n57 0.752
R14105 a_2551_4880.n97 a_2551_4880.n93 0.752
R14106 a_2551_4880.n75 a_2551_4880.n71 0.752
R14107 a_2551_4880.n84 a_2551_4880.n80 0.752
R14108 a_2551_4880.n15 a_2551_4880.n14 0.461
R14109 a_2551_4880.n67 a_2551_4880.n66 0.456
R14110 a_2551_4880.n44 a_2551_4880.n42 0.456
R14111 a_2551_4880.n18 a_2551_4880.n17 0.43
R14112 a_2551_4880.n21 a_2551_4880.n20 0.398
R14113 a_2551_4880.n24 a_2551_4880.n23 0.366
R14114 a_2551_4880.n27 a_2551_4880.n26 0.334
R14115 a_2551_4880.n119 a_2551_4880.n122 0.278
R14116 a_2551_4880.n102 a_2551_4880.n88 0.228
R14117 a_2551_4880.n102 a_2551_4880.n101 0.228
R14118 a_2551_4880.n103 a_2551_4880.n102 0.19
R14119 a_2551_4880.n55 a_2551_4880.n2 0.19
R14120 a_2551_4880.n3 a_2551_4880.n55 0.19
R14121 a_2551_4880.n78 a_2551_4880.n5 0.19
R14122 a_2551_4880.n6 a_2551_4880.n78 0.19
R14123 a_2551_4880.n110 a_2551_4880.n108 0.19
R14124 a_2551_4880.n106 a_2551_4880.n105 0.189
R14125 a_2551_4880.n108 a_2551_4880.n106 0.189
R14126 a_2551_4880.n112 a_2551_4880.n110 0.189
R14127 a_2551_4880.n114 a_2551_4880.n112 0.165
R14128 a_2551_4880.n105 a_2551_4880.n103 0.164
R14129 a_2551_4880.n120 a_2551_4880.n121 0.161
R14130 a_2551_4880.n42 a_2551_4880.n40 0.158
R14131 a_2551_4880.n1 a_2551_4880.n44 0.158
R14132 a_2551_4880.n66 a_2551_4880.n64 0.158
R14133 a_2551_4880.n4 a_2551_4880.n67 0.158
R14134 a_2551_4880.n88 a_2551_4880.n87 0.158
R14135 a_2551_4880.n101 a_2551_4880.n100 0.158
R14136 a_2551_4880.n123 a_2551_4880.n124 0.15
R14137 a_2551_4880.n9 a_2551_4880.n8 0.139
R14138 a_2551_4880.n8 a_2551_4880.n119 0.132
R14139 a_2551_4880.n100 a_2551_4880.n7 0.045
R14140 a_2551_4880.n87 a_2551_4880.n6 0.045
R14141 a_2551_4880.n5 a_2551_4880.n4 0.045
R14142 a_2551_4880.n64 a_2551_4880.n3 0.045
R14143 a_2551_4880.n2 a_2551_4880.n1 0.045
R14144 a_2551_4880.n40 a_2551_4880.n0 0.045
R14145 a_2551_4880.n134 a_2551_4880.n131 0.044
R14146 a_2551_4880.n131 a_2551_4880.n117 0.043
R14147 a_2551_4880.n117 a_2551_4880.n114 0.043
R14148 a_2551_4880.n135 a_2551_4880.n134 0.043
R14149 a_2551_4880.n138 a_2551_4880.n135 0.042
R14150 a_2551_4880.n131 a_2551_4880.n9 7.513
R14151 a_8881_1782.n109 a_8881_1782.t2 120.5
R14152 a_8881_1782.n21 a_8881_1782.t0 69.205
R14153 a_8881_1782.n59 a_8881_1782.t3 60.25
R14154 a_8881_1782.n46 a_8881_1782.n45 31.448
R14155 a_8881_1782.n24 a_8881_1782.n23 27.517
R14156 a_8881_1782.n7 a_8881_1782.n3 26.106
R14157 a_8881_1782.n35 a_8881_1782.n34 23.586
R14158 a_8881_1782.n13 a_8881_1782.n12 19.655
R14159 a_8881_1782.n3 a_8881_1782.n2 15.724
R14160 a_8881_1782.n14 a_8881_1782.n13 13.758
R14161 a_8881_1782.n36 a_8881_1782.n35 9.827
R14162 a_8881_1782.n86 a_8881_1782.n85 9.3
R14163 a_8881_1782.n69 a_8881_1782.n68 9.3
R14164 a_8881_1782.n123 a_8881_1782.n122 9.3
R14165 a_8881_1782.n104 a_8881_1782.n103 9.3
R14166 a_8881_1782.n50 a_8881_1782.n52 9.3
R14167 a_8881_1782.n15 a_8881_1782.n14 9.3
R14168 a_8881_1782.n37 a_8881_1782.n36 9.3
R14169 a_8881_1782.n28 a_8881_1782.n38 9.3
R14170 a_8881_1782.n26 a_8881_1782.n25 9.3
R14171 a_8881_1782.n39 a_8881_1782.n41 9.3
R14172 a_8881_1782.n48 a_8881_1782.n47 9.3
R14173 a_8881_1782.n1 a_8881_1782.n139 9.3
R14174 a_8881_1782.n131 a_8881_1782.n146 9.3
R14175 a_8881_1782.n1 a_8881_1782.n138 9.3
R14176 a_8881_1782.n0 a_8881_1782.n134 9.3
R14177 a_8881_1782.n131 a_8881_1782.n145 9.3
R14178 a_8881_1782.n60 a_8881_1782.n59 8.764
R14179 a_8881_1782.n110 a_8881_1782.n109 8.764
R14180 a_8881_1782.n67 a_8881_1782.n66 8.215
R14181 a_8881_1782.n84 a_8881_1782.n83 8.215
R14182 a_8881_1782.n102 a_8881_1782.n101 7.453
R14183 a_8881_1782.n121 a_8881_1782.n120 7.453
R14184 a_8881_1782.n25 a_8881_1782.n24 5.896
R14185 a_8881_1782.n150 a_8881_1782.n149 5.38
R14186 a_8881_1782.n8 a_8881_1782.n7 5.201
R14187 a_8881_1782.n56 a_8881_1782.n54 4.869
R14188 a_8881_1782.n89 a_8881_1782.n74 4.863
R14189 a_8881_1782.n92 a_8881_1782.n90 4.838
R14190 a_8881_1782.n126 a_8881_1782.n108 4.837
R14191 a_8881_1782.n111 a_8881_1782.n110 4.65
R14192 a_8881_1782.n0 a_8881_1782.n133 4.529
R14193 a_8881_1782.n30 a_8881_1782.n31 4.517
R14194 a_8881_1782.n33 a_8881_1782.n32 4.517
R14195 a_8881_1782.n55 a_8881_1782.n70 4.5
R14196 a_8881_1782.n57 a_8881_1782.n63 4.5
R14197 a_8881_1782.n77 a_8881_1782.n81 4.5
R14198 a_8881_1782.n82 a_8881_1782.n88 4.5
R14199 a_8881_1782.n91 a_8881_1782.n105 4.5
R14200 a_8881_1782.n93 a_8881_1782.n98 4.5
R14201 a_8881_1782.n114 a_8881_1782.n118 4.5
R14202 a_8881_1782.n119 a_8881_1782.n125 4.5
R14203 a_8881_1782.n8 a_8881_1782.n16 4.5
R14204 a_8881_1782.n42 a_8881_1782.n49 4.5
R14205 a_8881_1782.n29 a_8881_1782.n27 4.5
R14206 a_8881_1782.n94 a_8881_1782.n95 4.5
R14207 a_8881_1782.n113 a_8881_1782.n112 4.5
R14208 a_8881_1782.n1 a_8881_1782.n137 4.5
R14209 a_8881_1782.n130 a_8881_1782.n144 4.5
R14210 a_8881_1782.n58 a_8881_1782.n60 4.141
R14211 a_8881_1782.n76 a_8881_1782.n75 4.141
R14212 a_8881_1782.n49 a_8881_1782.n43 4.141
R14213 a_8881_1782.n88 a_8881_1782.n86 3.764
R14214 a_8881_1782.n125 a_8881_1782.n123 3.764
R14215 a_8881_1782.n16 a_8881_1782.n9 3.764
R14216 a_8881_1782.n11 a_8881_1782.n10 3.764
R14217 a_8881_1782.n70 a_8881_1782.n69 3.388
R14218 a_8881_1782.n105 a_8881_1782.n104 3.388
R14219 a_8881_1782.n6 a_8881_1782.n5 3.388
R14220 a_8881_1782.n130 a_8881_1782.n141 3.169
R14221 a_8881_1782.n70 a_8881_1782.n64 3.011
R14222 a_8881_1782.n81 a_8881_1782.n80 3.011
R14223 a_8881_1782.n105 a_8881_1782.n99 3.011
R14224 a_8881_1782.n98 a_8881_1782.n96 3.011
R14225 a_8881_1782.n5 a_8881_1782.n4 3.011
R14226 a_8881_1782.t1 a_8881_1782.n151 2.769
R14227 a_8881_1782.n63 a_8881_1782.n61 2.635
R14228 a_8881_1782.n88 a_8881_1782.n87 2.635
R14229 a_8881_1782.n118 a_8881_1782.n117 2.635
R14230 a_8881_1782.n125 a_8881_1782.n124 2.635
R14231 a_8881_1782.n16 a_8881_1782.n15 2.635
R14232 a_8881_1782.n15 a_8881_1782.n11 2.635
R14233 a_8881_1782.n53 a_8881_1782.n21 2.414
R14234 a_8881_1782.n107 a_8881_1782.n127 2.281
R14235 a_8881_1782.n49 a_8881_1782.n48 2.258
R14236 a_8881_1782.n52 a_8881_1782.n51 2.258
R14237 a_8881_1782.n47 a_8881_1782.n46 1.965
R14238 a_8881_1782.n30 a_8881_1782.n37 1.882
R14239 a_8881_1782.n37 a_8881_1782.n33 1.882
R14240 a_8881_1782.n151 a_8881_1782.n150 1.844
R14241 a_8881_1782.n81 a_8881_1782.n78 1.505
R14242 a_8881_1782.n118 a_8881_1782.n115 1.505
R14243 a_8881_1782.n117 a_8881_1782.n116 1.505
R14244 a_8881_1782.n27 a_8881_1782.n26 1.505
R14245 a_8881_1782.n41 a_8881_1782.n40 1.505
R14246 a_8881_1782.n151 a_8881_1782.n140 1.318
R14247 a_8881_1782.n151 a_8881_1782.n148 1.297
R14248 a_8881_1782.n18 a_8881_1782.n129 1.245
R14249 a_8881_1782.n107 a_8881_1782.n92 1.211
R14250 a_8881_1782.n71 a_8881_1782.n89 1.156
R14251 a_8881_1782.n73 a_8881_1782.n56 1.209
R14252 a_8881_1782.n106 a_8881_1782.n126 1.154
R14253 a_8881_1782.n63 a_8881_1782.n62 1.129
R14254 a_8881_1782.n80 a_8881_1782.n79 1.129
R14255 a_8881_1782.n98 a_8881_1782.n97 1.129
R14256 a_8881_1782.n26 a_8881_1782.n22 1.129
R14257 a_8881_1782.n68 a_8881_1782.n67 1.095
R14258 a_8881_1782.n85 a_8881_1782.n84 1.095
R14259 a_8881_1782.n1 a_8881_1782.n132 1.047
R14260 a_8881_1782.n147 a_8881_1782.n127 0.996
R14261 a_8881_1782.n17 a_8881_1782.n53 0.993
R14262 a_8881_1782.n103 a_8881_1782.n102 0.993
R14263 a_8881_1782.n122 a_8881_1782.n121 0.993
R14264 a_8881_1782.n72 a_8881_1782.n128 0.962
R14265 a_8881_1782.n69 a_8881_1782.n65 0.752
R14266 a_8881_1782.n104 a_8881_1782.n100 0.752
R14267 a_8881_1782.n137 a_8881_1782.n135 0.752
R14268 a_8881_1782.n140 a_8881_1782.n1 0.417
R14269 a_8881_1782.n148 a_8881_1782.n147 0.385
R14270 a_8881_1782.n48 a_8881_1782.n44 0.376
R14271 a_8881_1782.n144 a_8881_1782.n142 0.376
R14272 a_8881_1782.n7 a_8881_1782.n6 0.319
R14273 a_8881_1782.n135 a_8881_1782.n136 0.121
R14274 a_8881_1782.n142 a_8881_1782.n143 0.109
R14275 a_8881_1782.n147 a_8881_1782.n131 0.082
R14276 a_8881_1782.n53 a_8881_1782.n50 0.081
R14277 a_8881_1782.n107 a_8881_1782.n106 0.057
R14278 a_8881_1782.n42 a_8881_1782.n39 0.097
R14279 a_8881_1782.n126 a_8881_1782.n119 0.035
R14280 a_8881_1782.n131 a_8881_1782.n130 0.032
R14281 a_8881_1782.n20 a_8881_1782.n19 0.027
R14282 a_8881_1782.n128 a_8881_1782.n107 0.027
R14283 a_8881_1782.n129 a_8881_1782.n73 0.027
R14284 a_8881_1782.n20 a_8881_1782.n18 0.027
R14285 a_8881_1782.n73 a_8881_1782.n72 0.027
R14286 a_8881_1782.n113 a_8881_1782.n111 0.023
R14287 a_8881_1782.n77 a_8881_1782.n76 4.588
R14288 a_8881_1782.n114 a_8881_1782.n113 0.088
R14289 a_8881_1782.n93 a_8881_1782.n94 0.087
R14290 a_8881_1782.n57 a_8881_1782.n58 4.587
R14291 a_8881_1782.n20 a_8881_1782.n17 0.118
R14292 a_8881_1782.n28 a_8881_1782.n30 4.612
R14293 a_8881_1782.n73 a_8881_1782.n71 0.057
R14294 a_8881_1782.n82 a_8881_1782.n77 0.043
R14295 a_8881_1782.n119 a_8881_1782.n114 0.043
R14296 a_8881_1782.n91 a_8881_1782.n93 0.043
R14297 a_8881_1782.n55 a_8881_1782.n57 0.043
R14298 a_8881_1782.n92 a_8881_1782.n91 0.037
R14299 a_8881_1782.n89 a_8881_1782.n82 0.037
R14300 a_8881_1782.n56 a_8881_1782.n55 0.035
R14301 a_8881_1782.n50 a_8881_1782.n42 0.032
R14302 a_8881_1782.n39 a_8881_1782.n29 0.032
R14303 a_8881_1782.n29 a_8881_1782.n28 0.025
R14304 a_8881_1782.n20 a_8881_1782.n8 1.594
R14305 a_8881_1782.n1 a_8881_1782.n0 0.219
R14306 dvss.n2705 dvss.n2704 4919.86
R14307 dvss.n2639 dvss.n2638 4919.86
R14308 dvss.n2529 dvss.n2528 4919.86
R14309 dvss.n1378 dvss.n1377 4919.86
R14310 dvss.n2458 dvss.n1890 4919.86
R14311 dvss.n1996 dvss.n1995 4919.86
R14312 dvss.n2804 dvss.n659 4919.86
R14313 dvss.n765 dvss.n764 4919.86
R14314 dvss.n153 dvss.n152 4919.86
R14315 dvss.n2883 dvss.n2882 4919.86
R14316 dvss.n2705 dvss.n2698 4911.63
R14317 dvss.n2713 dvss.n2698 4911.63
R14318 dvss.n2714 dvss.n2713 4911.63
R14319 dvss.n2715 dvss.n2714 4911.63
R14320 dvss.n2715 dvss.n2690 4911.63
R14321 dvss.n2746 dvss.n2690 4911.63
R14322 dvss.n2639 dvss.n2632 4911.63
R14323 dvss.n2647 dvss.n2632 4911.63
R14324 dvss.n2648 dvss.n2647 4911.63
R14325 dvss.n2651 dvss.n2648 4911.63
R14326 dvss.n2651 dvss.n2650 4911.63
R14327 dvss.n2538 dvss.n2537 4911.63
R14328 dvss.n2537 dvss.n1271 4911.63
R14329 dvss.n2529 dvss.n1271 4911.63
R14330 dvss.n1327 dvss.n1326 4911.63
R14331 dvss.n1328 dvss.n1327 4911.63
R14332 dvss.n1328 dvss.n1300 4911.63
R14333 dvss.n1336 dvss.n1300 4911.63
R14334 dvss.n2469 dvss.n2468 4911.63
R14335 dvss.n2468 dvss.n2467 4911.63
R14336 dvss.n2467 dvss.n1890 4911.63
R14337 dvss.n1945 dvss.n1944 4911.63
R14338 dvss.n1946 dvss.n1945 4911.63
R14339 dvss.n1946 dvss.n1918 4911.63
R14340 dvss.n1954 dvss.n1918 4911.63
R14341 dvss.n2815 dvss.n2814 4911.63
R14342 dvss.n2814 dvss.n2813 4911.63
R14343 dvss.n2813 dvss.n659 4911.63
R14344 dvss.n714 dvss.n713 4911.63
R14345 dvss.n715 dvss.n714 4911.63
R14346 dvss.n715 dvss.n687 4911.63
R14347 dvss.n723 dvss.n687 4911.63
R14348 dvss.n102 dvss.n101 4911.63
R14349 dvss.n103 dvss.n102 4911.63
R14350 dvss.n103 dvss.n75 4911.63
R14351 dvss.n111 dvss.n75 4911.63
R14352 dvss.n2892 dvss.n43 4911.63
R14353 dvss.n2884 dvss.n43 4911.63
R14354 dvss.n2884 dvss.n2883 4911.63
R14355 dvss.n1337 dvss.n1336 4618.19
R14356 dvss.n1955 dvss.n1954 4618.19
R14357 dvss.n724 dvss.n723 4618.19
R14358 dvss.n112 dvss.n111 4618.19
R14359 dvss.n1377 dvss.n1281 4450.52
R14360 dvss.n1995 dvss.n1899 4450.52
R14361 dvss.n764 dvss.n668 4450.52
R14362 dvss.n152 dvss.n56 4450.52
R14363 dvss.n2577 dvss.n1233 3746.13
R14364 dvss.n2509 dvss.n2508 3746.13
R14365 dvss.n2853 dvss.n623 3746.13
R14366 dvss.n2926 dvss.n8 3746.13
R14367 dvss.t180 dvss.t178 3581.4
R14368 dvss.t174 dvss.t180 2984.5
R14369 dvss.n2539 dvss.n2538 2801.03
R14370 dvss.n2469 dvss.n1889 2801.03
R14371 dvss.n2815 dvss.n658 2801.03
R14372 dvss.n2893 dvss.n2892 2801.03
R14373 dvss.t119 dvss.t145 2244.48
R14374 dvss.n2747 dvss.n2746 1841.86
R14375 dvss.n2680 dvss.n2614 1665.19
R14376 dvss.n1326 dvss.n1306 1484.03
R14377 dvss.n1944 dvss.n1924 1484.03
R14378 dvss.n713 dvss.n693 1484.03
R14379 dvss.n101 dvss.n81 1484.03
R14380 dvss.n2650 dvss.n2649 1461.47
R14381 dvss.n1686 dvss.n1685 1308.2
R14382 dvss.n1679 dvss.n1675 1308.2
R14383 dvss.n2304 dvss.n2303 1308.2
R14384 dvss.n2297 dvss.n2293 1308.2
R14385 dvss.n1073 dvss.n1072 1308.2
R14386 dvss.n1066 dvss.n1062 1308.2
R14387 dvss.n461 dvss.n460 1308.2
R14388 dvss.n454 dvss.n450 1308.2
R14389 dvss.n1314 dvss.n1313 1295.7
R14390 dvss.n1932 dvss.n1931 1295.7
R14391 dvss.n701 dvss.n700 1295.7
R14392 dvss.n89 dvss.n88 1295.7
R14393 dvss.n2590 dvss.n2589 1260.9
R14394 dvss.n2519 dvss.n2518 1260.9
R14395 dvss.n2791 dvss.n2790 1260.9
R14396 dvss.n2866 dvss.n2865 1260.9
R14397 dvss.n2747 dvss.t147 1224.74
R14398 dvss.t4 dvss.n1227 1178.11
R14399 dvss.t57 dvss.n1842 1178.11
R14400 dvss.t153 dvss.n2775 1178.11
R14401 dvss.t165 dvss.n613 1178.11
R14402 dvss.t32 dvss.n1310 1156.39
R14403 dvss.t121 dvss.n1928 1156.39
R14404 dvss.t159 dvss.n697 1156.39
R14405 dvss.t112 dvss.n85 1156.39
R14406 dvss.n2664 dvss.n2663 1147.83
R14407 dvss.n2666 dvss.n2664 1147.83
R14408 dvss.n2554 dvss.n2553 1088.66
R14409 dvss.n2553 dvss.n2552 1088.66
R14410 dvss.n2485 dvss.n2484 1088.66
R14411 dvss.n2484 dvss.n1877 1088.66
R14412 dvss.n2831 dvss.n2830 1088.66
R14413 dvss.n2830 dvss.n646 1088.66
R14414 dvss.n2904 dvss.n2903 1088.66
R14415 dvss.n2903 dvss.n33 1088.66
R14416 dvss.n2663 dvss.t27 1076.09
R14417 dvss.n1687 dvss.n1549 1013.97
R14418 dvss.n1684 dvss.n1550 1013.97
R14419 dvss.n1678 dvss.n1677 1013.97
R14420 dvss.n1680 dvss.n1552 1013.97
R14421 dvss.n2305 dvss.n2167 1013.97
R14422 dvss.n2302 dvss.n2168 1013.97
R14423 dvss.n2296 dvss.n2295 1013.97
R14424 dvss.n2298 dvss.n2170 1013.97
R14425 dvss.n1074 dvss.n936 1013.97
R14426 dvss.n1071 dvss.n937 1013.97
R14427 dvss.n1065 dvss.n1064 1013.97
R14428 dvss.n1067 dvss.n939 1013.97
R14429 dvss.n462 dvss.n324 1013.97
R14430 dvss.n459 dvss.n325 1013.97
R14431 dvss.n453 dvss.n452 1013.97
R14432 dvss.n455 dvss.n327 1013.97
R14433 dvss.n2554 dvss.n1263 908.359
R14434 dvss.n2486 dvss.n2485 908.359
R14435 dvss.n2832 dvss.n2831 908.359
R14436 dvss.n2905 dvss.n2904 908.359
R14437 dvss.n2577 dvss.n2576 887.394
R14438 dvss.n2566 dvss.n1248 887.394
R14439 dvss.n2564 dvss.n1249 887.394
R14440 dvss.n1339 dvss.n1337 887.394
R14441 dvss.n1350 dvss.n1349 887.394
R14442 dvss.n1360 dvss.n1359 887.394
R14443 dvss.n1351 dvss.n1281 887.394
R14444 dvss.n2508 dvss.n1850 887.394
R14445 dvss.n2496 dvss.n1864 887.394
R14446 dvss.n2494 dvss.n1865 887.394
R14447 dvss.n1957 dvss.n1955 887.394
R14448 dvss.n1968 dvss.n1967 887.394
R14449 dvss.n1978 dvss.n1977 887.394
R14450 dvss.n1969 dvss.n1899 887.394
R14451 dvss.n2853 dvss.n2852 887.394
R14452 dvss.n2842 dvss.n633 887.394
R14453 dvss.n2840 dvss.n634 887.394
R14454 dvss.n726 dvss.n724 887.394
R14455 dvss.n737 dvss.n736 887.394
R14456 dvss.n747 dvss.n746 887.394
R14457 dvss.n738 dvss.n668 887.394
R14458 dvss.n114 dvss.n112 887.394
R14459 dvss.n125 dvss.n124 887.394
R14460 dvss.n135 dvss.n134 887.394
R14461 dvss.n126 dvss.n56 887.394
R14462 dvss.n2926 dvss.n2925 887.394
R14463 dvss.n2915 dvss.n20 887.394
R14464 dvss.n2913 dvss.n21 887.394
R14465 dvss.t47 dvss.n2575 841.176
R14466 dvss.n1863 dvss.t79 841.176
R14467 dvss.t16 dvss.n2851 841.176
R14468 dvss.t131 dvss.n2924 841.176
R14469 dvss.n2565 dvss.t41 822.689
R14470 dvss.n2495 dvss.t71 822.689
R14471 dvss.n2841 dvss.t10 822.689
R14472 dvss.n2914 dvss.t133 822.689
R14473 dvss.n1338 dvss.t103 794.957
R14474 dvss.n1956 dvss.t85 794.957
R14475 dvss.n725 dvss.t190 794.957
R14476 dvss.n113 dvss.t63 794.957
R14477 dvss.n2665 dvss.n2614 789.13
R14478 dvss.n1313 dvss.t163 782.822
R14479 dvss.n1931 dvss.t157 782.822
R14480 dvss.n700 dvss.t107 782.822
R14481 dvss.n88 dvss.t138 782.822
R14482 dvss.t101 dvss.n1358 757.983
R14483 dvss.t83 dvss.n1976 757.983
R14484 dvss.t188 dvss.n745 757.983
R14485 dvss.t59 dvss.n133 757.983
R14486 dvss.t174 dvss.n2665 753.26
R14487 dvss.n2589 dvss.t6 696.119
R14488 dvss.n2518 dvss.t55 696.119
R14489 dvss.n2790 dvss.t25 696.119
R14490 dvss.n2865 dvss.t167 696.119
R14491 dvss.n1358 dvss.t97 684.033
R14492 dvss.n1976 dvss.t87 684.033
R14493 dvss.n745 dvss.t186 684.033
R14494 dvss.n133 dvss.t69 684.033
R14495 dvss.n2552 dvss.t95 669.072
R14496 dvss.t91 dvss.n1877 669.072
R14497 dvss.t194 dvss.n646 669.072
R14498 dvss.t67 dvss.n33 669.072
R14499 dvss.n1589 dvss.n1568 668.499
R14500 dvss.n1593 dvss.n1570 668.499
R14501 dvss.n1650 dvss.n1604 668.499
R14502 dvss.n1655 dvss.n1654 668.499
R14503 dvss.n1662 dvss.n1557 668.499
R14504 dvss.n1660 dvss.n1560 668.499
R14505 dvss.n1709 dvss.n1529 668.499
R14506 dvss.n1669 dvss.n1532 668.499
R14507 dvss.n1475 dvss.n1470 668.499
R14508 dvss.n1736 dvss.n1472 668.499
R14509 dvss.n1818 dvss.n1389 668.499
R14510 dvss.n1799 dvss.n1386 668.499
R14511 dvss.n2207 dvss.n2186 668.499
R14512 dvss.n2211 dvss.n2188 668.499
R14513 dvss.n2268 dvss.n2222 668.499
R14514 dvss.n2273 dvss.n2272 668.499
R14515 dvss.n2280 dvss.n2175 668.499
R14516 dvss.n2278 dvss.n2178 668.499
R14517 dvss.n2327 dvss.n2147 668.499
R14518 dvss.n2287 dvss.n2150 668.499
R14519 dvss.n2093 dvss.n2088 668.499
R14520 dvss.n2354 dvss.n2090 668.499
R14521 dvss.n2436 dvss.n2007 668.499
R14522 dvss.n2417 dvss.n2004 668.499
R14523 dvss.n976 dvss.n955 668.499
R14524 dvss.n980 dvss.n957 668.499
R14525 dvss.n1037 dvss.n991 668.499
R14526 dvss.n1042 dvss.n1041 668.499
R14527 dvss.n1049 dvss.n944 668.499
R14528 dvss.n1047 dvss.n947 668.499
R14529 dvss.n1096 dvss.n916 668.499
R14530 dvss.n1056 dvss.n919 668.499
R14531 dvss.n862 dvss.n857 668.499
R14532 dvss.n1123 dvss.n859 668.499
R14533 dvss.n1205 dvss.n776 668.499
R14534 dvss.n1186 dvss.n773 668.499
R14535 dvss.n364 dvss.n343 668.499
R14536 dvss.n368 dvss.n345 668.499
R14537 dvss.n425 dvss.n379 668.499
R14538 dvss.n430 dvss.n429 668.499
R14539 dvss.n437 dvss.n332 668.499
R14540 dvss.n435 dvss.n335 668.499
R14541 dvss.n484 dvss.n304 668.499
R14542 dvss.n444 dvss.n307 668.499
R14543 dvss.n250 dvss.n245 668.499
R14544 dvss.n511 dvss.n247 668.499
R14545 dvss.n593 dvss.n164 668.499
R14546 dvss.n574 dvss.n161 668.499
R14547 dvss.t105 dvss.n1338 647.058
R14548 dvss.t93 dvss.n1956 647.058
R14549 dvss.t192 dvss.n725 647.058
R14550 dvss.t65 dvss.n113 647.058
R14551 dvss.n1439 dvss.n1432 623.66
R14552 dvss.n1781 dvss.n1392 623.66
R14553 dvss.n2057 dvss.n2050 623.66
R14554 dvss.n2399 dvss.n2010 623.66
R14555 dvss.n826 dvss.n819 623.66
R14556 dvss.n1168 dvss.n779 623.66
R14557 dvss.n214 dvss.n207 623.66
R14558 dvss.n556 dvss.n167 623.66
R14559 dvss.t43 dvss.n2565 619.327
R14560 dvss.t75 dvss.n2495 619.327
R14561 dvss.t12 dvss.n2841 619.327
R14562 dvss.t127 dvss.n2914 619.327
R14563 dvss.n2575 dvss.t45 600.84
R14564 dvss.t77 dvss.n1863 600.84
R14565 dvss.n2851 dvss.t14 600.84
R14566 dvss.n2924 dvss.t129 600.84
R14567 dvss.n0 dvss.t117 571.478
R14568 dvss.n2767 dvss.t39 571.478
R14569 dvss.t6 dvss.n2588 571.478
R14570 dvss.t55 dvss.n2517 571.478
R14571 dvss.t25 dvss.n2789 571.478
R14572 dvss.t167 dvss.n2864 571.478
R14573 dvss.t81 dvss.n1270 555.67
R14574 dvss.t155 dvss.n1888 555.67
R14575 dvss.t172 dvss.n657 555.67
R14576 dvss.n2894 dvss.t182 555.67
R14577 dvss.n1591 dvss.n1569 545.089
R14578 dvss.n1653 dvss.n1652 545.089
R14579 dvss.n1661 dvss.n1558 545.089
R14580 dvss.n1707 dvss.n1531 545.089
R14581 dvss.n1734 dvss.n1471 545.089
R14582 dvss.n1755 dvss.n1439 545.089
R14583 dvss.n1793 dvss.n1392 545.089
R14584 dvss.n1816 dvss.n1387 545.089
R14585 dvss.n2209 dvss.n2187 545.089
R14586 dvss.n2271 dvss.n2270 545.089
R14587 dvss.n2279 dvss.n2176 545.089
R14588 dvss.n2325 dvss.n2149 545.089
R14589 dvss.n2352 dvss.n2089 545.089
R14590 dvss.n2373 dvss.n2057 545.089
R14591 dvss.n2411 dvss.n2010 545.089
R14592 dvss.n2434 dvss.n2005 545.089
R14593 dvss.n978 dvss.n956 545.089
R14594 dvss.n1040 dvss.n1039 545.089
R14595 dvss.n1048 dvss.n945 545.089
R14596 dvss.n1094 dvss.n918 545.089
R14597 dvss.n1121 dvss.n858 545.089
R14598 dvss.n1142 dvss.n826 545.089
R14599 dvss.n1180 dvss.n779 545.089
R14600 dvss.n1203 dvss.n774 545.089
R14601 dvss.n366 dvss.n344 545.089
R14602 dvss.n428 dvss.n427 545.089
R14603 dvss.n436 dvss.n333 545.089
R14604 dvss.n482 dvss.n306 545.089
R14605 dvss.n509 dvss.n246 545.089
R14606 dvss.n530 dvss.n214 545.089
R14607 dvss.n568 dvss.n167 545.089
R14608 dvss.n591 dvss.n162 545.089
R14609 dvss.n2706 dvss.n2703 539.294
R14610 dvss.n2706 dvss.n2699 539.294
R14611 dvss.n2712 dvss.n2699 539.294
R14612 dvss.n2712 dvss.n2697 539.294
R14613 dvss.n2716 dvss.n2697 539.294
R14614 dvss.n2716 dvss.n2691 539.294
R14615 dvss.n2745 dvss.n2691 539.294
R14616 dvss.n2745 dvss.n2692 539.294
R14617 dvss.n2738 dvss.n2723 539.294
R14618 dvss.n2733 dvss.n2732 539.294
R14619 dvss.n2730 dvss.n2686 539.294
R14620 dvss.n2640 dvss.n2637 539.294
R14621 dvss.n2640 dvss.n2633 539.294
R14622 dvss.n2646 dvss.n2633 539.294
R14623 dvss.n2646 dvss.n2630 539.294
R14624 dvss.n2652 dvss.n2630 539.294
R14625 dvss.n2652 dvss.n2631 539.294
R14626 dvss.n2631 dvss.n2624 539.294
R14627 dvss.n2662 dvss.n2624 539.294
R14628 dvss.n2662 dvss.n2623 539.294
R14629 dvss.n2667 dvss.n2623 539.294
R14630 dvss.n2667 dvss.n2616 539.294
R14631 dvss.n2678 dvss.n2616 539.294
R14632 dvss.n2615 dvss.n2613 539.294
R14633 dvss.n2591 dvss.n1227 539.294
R14634 dvss.n2591 dvss.n1228 539.294
R14635 dvss.n2587 dvss.n1228 539.294
R14636 dvss.n2579 dvss.n2578 539.294
R14637 dvss.n2578 dvss.n1236 539.294
R14638 dvss.n2574 dvss.n1236 539.294
R14639 dvss.n2574 dvss.n1237 539.294
R14640 dvss.n2567 dvss.n1237 539.294
R14641 dvss.n2567 dvss.n1247 539.294
R14642 dvss.n2563 dvss.n1247 539.294
R14643 dvss.n2563 dvss.n1250 539.294
R14644 dvss.n1261 dvss.n1250 539.294
R14645 dvss.n2555 dvss.n1261 539.294
R14646 dvss.n2555 dvss.n1262 539.294
R14647 dvss.n2551 dvss.n1262 539.294
R14648 dvss.n2551 dvss.n1264 539.294
R14649 dvss.n2540 dvss.n1264 539.294
R14650 dvss.n2540 dvss.n1269 539.294
R14651 dvss.n2536 dvss.n1269 539.294
R14652 dvss.n2536 dvss.n1272 539.294
R14653 dvss.n2530 dvss.n1272 539.294
R14654 dvss.n2530 dvss.n1276 539.294
R14655 dvss.n1315 dvss.n1310 539.294
R14656 dvss.n1315 dvss.n1312 539.294
R14657 dvss.n1312 dvss.n1307 539.294
R14658 dvss.n1325 dvss.n1307 539.294
R14659 dvss.n1325 dvss.n1305 539.294
R14660 dvss.n1329 dvss.n1305 539.294
R14661 dvss.n1329 dvss.n1301 539.294
R14662 dvss.n1335 dvss.n1301 539.294
R14663 dvss.n1335 dvss.n1299 539.294
R14664 dvss.n1340 dvss.n1299 539.294
R14665 dvss.n1340 dvss.n1295 539.294
R14666 dvss.n1348 dvss.n1295 539.294
R14667 dvss.n1348 dvss.n1293 539.294
R14668 dvss.n1361 dvss.n1293 539.294
R14669 dvss.n1361 dvss.n1294 539.294
R14670 dvss.n1357 dvss.n1294 539.294
R14671 dvss.n1357 dvss.n1352 539.294
R14672 dvss.n1352 dvss.n1282 539.294
R14673 dvss.n1376 dvss.n1282 539.294
R14674 dvss.n1376 dvss.n1280 539.294
R14675 dvss.n2520 dvss.n1842 539.294
R14676 dvss.n2520 dvss.n1843 539.294
R14677 dvss.n2516 dvss.n1843 539.294
R14678 dvss.n2507 dvss.n1849 539.294
R14679 dvss.n2507 dvss.n1851 539.294
R14680 dvss.n1862 dvss.n1851 539.294
R14681 dvss.n1862 dvss.n1859 539.294
R14682 dvss.n2497 dvss.n1859 539.294
R14683 dvss.n2497 dvss.n1861 539.294
R14684 dvss.n2493 dvss.n1861 539.294
R14685 dvss.n2493 dvss.n1866 539.294
R14686 dvss.n2487 dvss.n1866 539.294
R14687 dvss.n2487 dvss.n1876 539.294
R14688 dvss.n2483 dvss.n1876 539.294
R14689 dvss.n2483 dvss.n1878 539.294
R14690 dvss.n1887 dvss.n1878 539.294
R14691 dvss.n1887 dvss.n1884 539.294
R14692 dvss.n2470 dvss.n1884 539.294
R14693 dvss.n2470 dvss.n1886 539.294
R14694 dvss.n2466 dvss.n1886 539.294
R14695 dvss.n2466 dvss.n1891 539.294
R14696 dvss.n2459 dvss.n1891 539.294
R14697 dvss.n1933 dvss.n1928 539.294
R14698 dvss.n1933 dvss.n1930 539.294
R14699 dvss.n1930 dvss.n1925 539.294
R14700 dvss.n1943 dvss.n1925 539.294
R14701 dvss.n1943 dvss.n1923 539.294
R14702 dvss.n1947 dvss.n1923 539.294
R14703 dvss.n1947 dvss.n1919 539.294
R14704 dvss.n1953 dvss.n1919 539.294
R14705 dvss.n1953 dvss.n1917 539.294
R14706 dvss.n1958 dvss.n1917 539.294
R14707 dvss.n1958 dvss.n1913 539.294
R14708 dvss.n1966 dvss.n1913 539.294
R14709 dvss.n1966 dvss.n1911 539.294
R14710 dvss.n1979 dvss.n1911 539.294
R14711 dvss.n1979 dvss.n1912 539.294
R14712 dvss.n1975 dvss.n1912 539.294
R14713 dvss.n1975 dvss.n1970 539.294
R14714 dvss.n1970 dvss.n1900 539.294
R14715 dvss.n1994 dvss.n1900 539.294
R14716 dvss.n1994 dvss.n1898 539.294
R14717 dvss.n2792 dvss.n2775 539.294
R14718 dvss.n2792 dvss.n2778 539.294
R14719 dvss.n2779 dvss.n2778 539.294
R14720 dvss.n2854 dvss.n620 539.294
R14721 dvss.n2854 dvss.n622 539.294
R14722 dvss.n2850 dvss.n622 539.294
R14723 dvss.n2850 dvss.n624 539.294
R14724 dvss.n2843 dvss.n624 539.294
R14725 dvss.n2843 dvss.n632 539.294
R14726 dvss.n2839 dvss.n632 539.294
R14727 dvss.n2839 dvss.n635 539.294
R14728 dvss.n2833 dvss.n635 539.294
R14729 dvss.n2833 dvss.n645 539.294
R14730 dvss.n2829 dvss.n645 539.294
R14731 dvss.n2829 dvss.n647 539.294
R14732 dvss.n656 dvss.n647 539.294
R14733 dvss.n656 dvss.n653 539.294
R14734 dvss.n2816 dvss.n653 539.294
R14735 dvss.n2816 dvss.n655 539.294
R14736 dvss.n2812 dvss.n655 539.294
R14737 dvss.n2812 dvss.n660 539.294
R14738 dvss.n2805 dvss.n660 539.294
R14739 dvss.n702 dvss.n697 539.294
R14740 dvss.n702 dvss.n699 539.294
R14741 dvss.n699 dvss.n694 539.294
R14742 dvss.n712 dvss.n694 539.294
R14743 dvss.n712 dvss.n692 539.294
R14744 dvss.n716 dvss.n692 539.294
R14745 dvss.n716 dvss.n688 539.294
R14746 dvss.n722 dvss.n688 539.294
R14747 dvss.n722 dvss.n686 539.294
R14748 dvss.n727 dvss.n686 539.294
R14749 dvss.n727 dvss.n682 539.294
R14750 dvss.n735 dvss.n682 539.294
R14751 dvss.n735 dvss.n680 539.294
R14752 dvss.n748 dvss.n680 539.294
R14753 dvss.n748 dvss.n681 539.294
R14754 dvss.n744 dvss.n681 539.294
R14755 dvss.n744 dvss.n739 539.294
R14756 dvss.n739 dvss.n669 539.294
R14757 dvss.n763 dvss.n669 539.294
R14758 dvss.n763 dvss.n667 539.294
R14759 dvss.n2867 dvss.n613 539.294
R14760 dvss.n2867 dvss.n614 539.294
R14761 dvss.n2863 dvss.n614 539.294
R14762 dvss.n90 dvss.n85 539.294
R14763 dvss.n90 dvss.n87 539.294
R14764 dvss.n87 dvss.n82 539.294
R14765 dvss.n100 dvss.n82 539.294
R14766 dvss.n100 dvss.n80 539.294
R14767 dvss.n104 dvss.n80 539.294
R14768 dvss.n104 dvss.n76 539.294
R14769 dvss.n110 dvss.n76 539.294
R14770 dvss.n110 dvss.n74 539.294
R14771 dvss.n115 dvss.n74 539.294
R14772 dvss.n115 dvss.n70 539.294
R14773 dvss.n123 dvss.n70 539.294
R14774 dvss.n123 dvss.n68 539.294
R14775 dvss.n136 dvss.n68 539.294
R14776 dvss.n136 dvss.n69 539.294
R14777 dvss.n132 dvss.n69 539.294
R14778 dvss.n132 dvss.n127 539.294
R14779 dvss.n127 dvss.n57 539.294
R14780 dvss.n151 dvss.n57 539.294
R14781 dvss.n151 dvss.n55 539.294
R14782 dvss.n2928 dvss.n2927 539.294
R14783 dvss.n2927 dvss.n9 539.294
R14784 dvss.n2923 dvss.n9 539.294
R14785 dvss.n2923 dvss.n10 539.294
R14786 dvss.n2916 dvss.n10 539.294
R14787 dvss.n2916 dvss.n19 539.294
R14788 dvss.n2912 dvss.n19 539.294
R14789 dvss.n2912 dvss.n22 539.294
R14790 dvss.n2906 dvss.n22 539.294
R14791 dvss.n2906 dvss.n32 539.294
R14792 dvss.n2902 dvss.n32 539.294
R14793 dvss.n2902 dvss.n34 539.294
R14794 dvss.n2895 dvss.n34 539.294
R14795 dvss.n2895 dvss.n42 539.294
R14796 dvss.n2891 dvss.n42 539.294
R14797 dvss.n2891 dvss.n44 539.294
R14798 dvss.n2885 dvss.n44 539.294
R14799 dvss.n2885 dvss.n50 539.294
R14800 dvss.n51 dvss.n50 539.294
R14801 dvss.n2539 dvss.t81 532.989
R14802 dvss.n1889 dvss.t155 532.989
R14803 dvss.n658 dvss.t172 532.989
R14804 dvss.t182 dvss.n2893 532.989
R14805 dvss.t163 dvss.n1306 512.883
R14806 dvss.t157 dvss.n1924 512.883
R14807 dvss.t107 dvss.n693 512.883
R14808 dvss.t138 dvss.n81 512.883
R14809 dvss.n2704 dvss.n2701 498.1
R14810 dvss.n2638 dvss.n2635 498.1
R14811 dvss.n2528 dvss.n2527 494.37
R14812 dvss.n1379 dvss.n1378 494.37
R14813 dvss.n2510 dvss.n2509 494.37
R14814 dvss.n1997 dvss.n1996 494.37
R14815 dvss.n623 dvss.n618 494.37
R14816 dvss.n766 dvss.n765 494.37
R14817 dvss.n154 dvss.n153 494.37
R14818 dvss.n2882 dvss.n2881 494.37
R14819 dvss.n2581 dvss.n1233 494.369
R14820 dvss.n2458 dvss.n2457 494.369
R14821 dvss.n2804 dvss.n2803 494.369
R14822 dvss.n8 dvss.n5 494.369
R14823 dvss.t49 dvss.n1249 489.915
R14824 dvss.t73 dvss.n1865 489.915
R14825 dvss.t8 dvss.n634 489.915
R14826 dvss.t125 dvss.n21 489.915
R14827 dvss.t99 dvss.n1350 462.184
R14828 dvss.t89 dvss.n1968 462.184
R14829 dvss.t184 dvss.n737 462.184
R14830 dvss.t61 dvss.n125 462.184
R14831 dvss.n1685 dvss.n1551 432.369
R14832 dvss.n1675 dvss.n1551 432.369
R14833 dvss.n2303 dvss.n2169 432.369
R14834 dvss.n2293 dvss.n2169 432.369
R14835 dvss.n1072 dvss.n938 432.369
R14836 dvss.n1062 dvss.n938 432.369
R14837 dvss.n460 dvss.n326 432.369
R14838 dvss.n450 dvss.n326 432.369
R14839 dvss.n1360 dvss.t99 425.21
R14840 dvss.n1978 dvss.t89 425.21
R14841 dvss.n747 dvss.t184 425.21
R14842 dvss.n135 dvss.t61 425.21
R14843 dvss.n1270 dvss.t95 419.587
R14844 dvss.n1888 dvss.t91 419.587
R14845 dvss.n657 dvss.t194 419.587
R14846 dvss.n2894 dvss.t67 419.587
R14847 dvss.n2789 dvss.n2788 403.934
R14848 dvss.n2588 dvss.n1229 403.934
R14849 dvss.n2517 dvss.n1844 403.934
R14850 dvss.n2864 dvss.n615 403.934
R14851 dvss.t176 dvss.t150 401.104
R14852 dvss.n1263 dvss.t49 397.478
R14853 dvss.n2486 dvss.t73 397.478
R14854 dvss.n2832 dvss.t8 397.478
R14855 dvss.n2905 dvss.t125 397.478
R14856 dvss.n2666 dvss.t174 394.565
R14857 dvss.n1684 dvss.n1552 394
R14858 dvss.n2302 dvss.n2170 394
R14859 dvss.n1071 dvss.n939 394
R14860 dvss.n459 dvss.n327 394
R14861 dvss.n1400 dvss.n1391 366.841
R14862 dvss.n1415 dvss.n1394 366.841
R14863 dvss.n1448 dvss.n1437 366.841
R14864 dvss.n1464 dvss.n1441 366.841
R14865 dvss.n2018 dvss.n2009 366.841
R14866 dvss.n2033 dvss.n2012 366.841
R14867 dvss.n2066 dvss.n2055 366.841
R14868 dvss.n2082 dvss.n2059 366.841
R14869 dvss.n787 dvss.n778 366.841
R14870 dvss.n802 dvss.n781 366.841
R14871 dvss.n835 dvss.n824 366.841
R14872 dvss.n851 dvss.n828 366.841
R14873 dvss.n175 dvss.n166 366.841
R14874 dvss.n190 dvss.n169 366.841
R14875 dvss.n223 dvss.n212 366.841
R14876 dvss.n239 dvss.n216 366.841
R14877 dvss.n1599 dvss.n1569 333.928
R14878 dvss.n1653 dvss.n1565 333.928
R14879 dvss.n1661 dvss.n1559 333.928
R14880 dvss.n1667 dvss.n1531 333.928
R14881 dvss.n1741 dvss.n1471 333.928
R14882 dvss.n1755 dvss.n1438 333.928
R14883 dvss.n1762 dvss.n1432 333.928
R14884 dvss.n1775 dvss.n1426 333.928
R14885 dvss.n1781 dvss.n1422 333.928
R14886 dvss.n1793 dvss.n1393 333.928
R14887 dvss.n1823 dvss.n1387 333.928
R14888 dvss.n2217 dvss.n2187 333.928
R14889 dvss.n2271 dvss.n2183 333.928
R14890 dvss.n2279 dvss.n2177 333.928
R14891 dvss.n2285 dvss.n2149 333.928
R14892 dvss.n2359 dvss.n2089 333.928
R14893 dvss.n2373 dvss.n2056 333.928
R14894 dvss.n2380 dvss.n2050 333.928
R14895 dvss.n2393 dvss.n2044 333.928
R14896 dvss.n2399 dvss.n2040 333.928
R14897 dvss.n2411 dvss.n2011 333.928
R14898 dvss.n2441 dvss.n2005 333.928
R14899 dvss.n986 dvss.n956 333.928
R14900 dvss.n1040 dvss.n952 333.928
R14901 dvss.n1048 dvss.n946 333.928
R14902 dvss.n1054 dvss.n918 333.928
R14903 dvss.n1128 dvss.n858 333.928
R14904 dvss.n1142 dvss.n825 333.928
R14905 dvss.n1149 dvss.n819 333.928
R14906 dvss.n1162 dvss.n813 333.928
R14907 dvss.n1168 dvss.n809 333.928
R14908 dvss.n1180 dvss.n780 333.928
R14909 dvss.n1210 dvss.n774 333.928
R14910 dvss.n374 dvss.n344 333.928
R14911 dvss.n428 dvss.n340 333.928
R14912 dvss.n436 dvss.n334 333.928
R14913 dvss.n442 dvss.n306 333.928
R14914 dvss.n516 dvss.n246 333.928
R14915 dvss.n530 dvss.n213 333.928
R14916 dvss.n537 dvss.n207 333.928
R14917 dvss.n550 dvss.n201 333.928
R14918 dvss.n556 dvss.n197 333.928
R14919 dvss.n568 dvss.n168 333.928
R14920 dvss.n598 dvss.n162 333.928
R14921 dvss.n1441 dvss.n1431 306.258
R14922 dvss.n1782 dvss.n1394 306.258
R14923 dvss.n1437 dvss.n1433 306.258
R14924 dvss.n1780 dvss.n1391 306.258
R14925 dvss.n2059 dvss.n2049 306.258
R14926 dvss.n2400 dvss.n2012 306.258
R14927 dvss.n2055 dvss.n2051 306.258
R14928 dvss.n2398 dvss.n2009 306.258
R14929 dvss.n828 dvss.n818 306.258
R14930 dvss.n1169 dvss.n781 306.258
R14931 dvss.n824 dvss.n820 306.258
R14932 dvss.n1167 dvss.n778 306.258
R14933 dvss.n216 dvss.n206 306.258
R14934 dvss.n557 dvss.n169 306.258
R14935 dvss.n212 dvss.n208 306.258
R14936 dvss.n555 dvss.n166 306.258
R14937 dvss.n1654 dvss.n1561 292.5
R14938 dvss.n1654 dvss.n1653 292.5
R14939 dvss.n1598 dvss.n1597 292.5
R14940 dvss.n1599 dvss.n1598 292.5
R14941 dvss.n1596 dvss.n1564 292.5
R14942 dvss.n1565 dvss.n1564 292.5
R14943 dvss.n1595 dvss.n1570 292.5
R14944 dvss.n1570 dvss.n1569 292.5
R14945 dvss.n1589 dvss.n1588 292.5
R14946 dvss.n1587 dvss.n1576 292.5
R14947 dvss.n1586 dvss.n1585 292.5
R14948 dvss.n1584 dvss.n1583 292.5
R14949 dvss.n1582 dvss.n1581 292.5
R14950 dvss.n1580 dvss.n1579 292.5
R14951 dvss.n1578 dvss.n1577 292.5
R14952 dvss.n1572 dvss.n1571 292.5
R14953 dvss.n1594 dvss.n1593 292.5
R14954 dvss.n1670 dvss.n1669 292.5
R14955 dvss.n1669 dvss.n1531 292.5
R14956 dvss.n1668 dvss.n1553 292.5
R14957 dvss.n1668 dvss.n1667 292.5
R14958 dvss.n1658 dvss.n1554 292.5
R14959 dvss.n1559 dvss.n1554 292.5
R14960 dvss.n1660 dvss.n1659 292.5
R14961 dvss.n1661 dvss.n1660 292.5
R14962 dvss.n1682 dvss.n1552 292.5
R14963 dvss.n1675 dvss.n1552 292.5
R14964 dvss.n1684 dvss.n1683 292.5
R14965 dvss.n1685 dvss.n1684 292.5
R14966 dvss.n1681 dvss.n1680 292.5
R14967 dvss.n1678 dvss.n1674 292.5
R14968 dvss.n1688 dvss.n1687 292.5
R14969 dvss.n1690 dvss.n1689 292.5
R14970 dvss.n1671 dvss.n1532 292.5
R14971 dvss.n1707 dvss.n1532 292.5
R14972 dvss.n1672 dvss.n1550 292.5
R14973 dvss.n1677 dvss.n1675 292.5
R14974 dvss.n1685 dvss.n1549 292.5
R14975 dvss.n1547 dvss.n1546 292.5
R14976 dvss.n1696 dvss.n1695 292.5
R14977 dvss.n1699 dvss.n1698 292.5
R14978 dvss.n1541 dvss.n1540 292.5
R14979 dvss.n1705 dvss.n1704 292.5
R14980 dvss.n1538 dvss.n1530 292.5
R14981 dvss.n1710 dvss.n1709 292.5
R14982 dvss.n1531 dvss.n1529 292.5
R14983 dvss.n1529 dvss.n1527 292.5
R14984 dvss.n1666 dvss.n1665 292.5
R14985 dvss.n1667 dvss.n1666 292.5
R14986 dvss.n1664 dvss.n1555 292.5
R14987 dvss.n1559 dvss.n1555 292.5
R14988 dvss.n1663 dvss.n1662 292.5
R14989 dvss.n1662 dvss.n1661 292.5
R14990 dvss.n1653 dvss.n1604 292.5
R14991 dvss.n1568 dvss.n1567 292.5
R14992 dvss.n1569 dvss.n1568 292.5
R14993 dvss.n1601 dvss.n1600 292.5
R14994 dvss.n1600 dvss.n1599 292.5
R14995 dvss.n1602 dvss.n1566 292.5
R14996 dvss.n1566 dvss.n1565 292.5
R14997 dvss.n1604 dvss.n1603 292.5
R14998 dvss.n1656 dvss.n1560 292.5
R14999 dvss.n1650 dvss.n1649 292.5
R15000 dvss.n1649 dvss.n1557 292.5
R15001 dvss.n1610 dvss.n1608 292.5
R15002 dvss.n1615 dvss.n1610 292.5
R15003 dvss.n1644 dvss.n1612 292.5
R15004 dvss.n1644 dvss.n1643 292.5
R15005 dvss.n1618 dvss.n1617 292.5
R15006 dvss.n1642 dvss.n1618 292.5
R15007 dvss.n1639 dvss.n1621 292.5
R15008 dvss.n1640 dvss.n1639 292.5
R15009 dvss.n1623 dvss.n1622 292.5
R15010 dvss.n1623 dvss.n1619 292.5
R15011 dvss.n1634 dvss.n1627 292.5
R15012 dvss.n1634 dvss.n1633 292.5
R15013 dvss.n1632 dvss.n1630 292.5
R15014 dvss.n1630 dvss.n1629 292.5
R15015 dvss.n1656 dvss.n1655 292.5
R15016 dvss.n1737 dvss.n1736 292.5
R15017 dvss.n1722 dvss.n1721 292.5
R15018 dvss.n1724 dvss.n1723 292.5
R15019 dvss.n1726 dvss.n1725 292.5
R15020 dvss.n1728 dvss.n1727 292.5
R15021 dvss.n1730 dvss.n1729 292.5
R15022 dvss.n1732 dvss.n1731 292.5
R15023 dvss.n1474 dvss.n1473 292.5
R15024 dvss.n1720 dvss.n1475 292.5
R15025 dvss.n1734 dvss.n1475 292.5
R15026 dvss.n1400 dvss.n1399 292.5
R15027 dvss.n1400 dvss.n1392 292.5
R15028 dvss.n1413 dvss.n1395 292.5
R15029 dvss.n1412 dvss.n1411 292.5
R15030 dvss.n1410 dvss.n1409 292.5
R15031 dvss.n1408 dvss.n1397 292.5
R15032 dvss.n1406 dvss.n1405 292.5
R15033 dvss.n1404 dvss.n1398 292.5
R15034 dvss.n1403 dvss.n1402 292.5
R15035 dvss.n1416 dvss.n1415 292.5
R15036 dvss.n1450 dvss.n1447 292.5
R15037 dvss.n1463 dvss.n1443 292.5
R15038 dvss.n1461 dvss.n1460 292.5
R15039 dvss.n1459 dvss.n1458 292.5
R15040 dvss.n1456 dvss.n1445 292.5
R15041 dvss.n1454 dvss.n1453 292.5
R15042 dvss.n1452 dvss.n1451 292.5
R15043 dvss.n1465 dvss.n1464 292.5
R15044 dvss.n1464 dvss.n1439 292.5
R15045 dvss.n1448 dvss.n1434 292.5
R15046 dvss.n1820 dvss.n1389 292.5
R15047 dvss.n1389 dvss.n1387 292.5
R15048 dvss.n1822 dvss.n1821 292.5
R15049 dvss.n1823 dvss.n1822 292.5
R15050 dvss.n1796 dvss.n1388 292.5
R15051 dvss.n1393 dvss.n1388 292.5
R15052 dvss.n1795 dvss.n1794 292.5
R15053 dvss.n1794 dvss.n1793 292.5
R15054 dvss.n1780 dvss.n1779 292.5
R15055 dvss.n1781 dvss.n1780 292.5
R15056 dvss.n1778 dvss.n1423 292.5
R15057 dvss.n1423 dvss.n1422 292.5
R15058 dvss.n1777 dvss.n1776 292.5
R15059 dvss.n1776 dvss.n1775 292.5
R15060 dvss.n1425 dvss.n1424 292.5
R15061 dvss.n1426 dvss.n1425 292.5
R15062 dvss.n1761 dvss.n1760 292.5
R15063 dvss.n1762 dvss.n1761 292.5
R15064 dvss.n1759 dvss.n1433 292.5
R15065 dvss.n1433 dvss.n1432 292.5
R15066 dvss.n1757 dvss.n1756 292.5
R15067 dvss.n1756 dvss.n1755 292.5
R15068 dvss.n1436 dvss.n1435 292.5
R15069 dvss.n1438 dvss.n1436 292.5
R15070 dvss.n1740 dvss.n1739 292.5
R15071 dvss.n1741 dvss.n1740 292.5
R15072 dvss.n1738 dvss.n1472 292.5
R15073 dvss.n1472 dvss.n1471 292.5
R15074 dvss.n1819 dvss.n1818 292.5
R15075 dvss.n1798 dvss.n1797 292.5
R15076 dvss.n1814 dvss.n1813 292.5
R15077 dvss.n1812 dvss.n1803 292.5
R15078 dvss.n1811 dvss.n1810 292.5
R15079 dvss.n1809 dvss.n1808 292.5
R15080 dvss.n1807 dvss.n1806 292.5
R15081 dvss.n1805 dvss.n1804 292.5
R15082 dvss.n1799 dvss.n1381 292.5
R15083 dvss.n2272 dvss.n2179 292.5
R15084 dvss.n2272 dvss.n2271 292.5
R15085 dvss.n2216 dvss.n2215 292.5
R15086 dvss.n2217 dvss.n2216 292.5
R15087 dvss.n2214 dvss.n2182 292.5
R15088 dvss.n2183 dvss.n2182 292.5
R15089 dvss.n2213 dvss.n2188 292.5
R15090 dvss.n2188 dvss.n2187 292.5
R15091 dvss.n2207 dvss.n2206 292.5
R15092 dvss.n2205 dvss.n2194 292.5
R15093 dvss.n2204 dvss.n2203 292.5
R15094 dvss.n2202 dvss.n2201 292.5
R15095 dvss.n2200 dvss.n2199 292.5
R15096 dvss.n2198 dvss.n2197 292.5
R15097 dvss.n2196 dvss.n2195 292.5
R15098 dvss.n2190 dvss.n2189 292.5
R15099 dvss.n2212 dvss.n2211 292.5
R15100 dvss.n2288 dvss.n2287 292.5
R15101 dvss.n2287 dvss.n2149 292.5
R15102 dvss.n2286 dvss.n2171 292.5
R15103 dvss.n2286 dvss.n2285 292.5
R15104 dvss.n2276 dvss.n2172 292.5
R15105 dvss.n2177 dvss.n2172 292.5
R15106 dvss.n2278 dvss.n2277 292.5
R15107 dvss.n2279 dvss.n2278 292.5
R15108 dvss.n2300 dvss.n2170 292.5
R15109 dvss.n2293 dvss.n2170 292.5
R15110 dvss.n2302 dvss.n2301 292.5
R15111 dvss.n2303 dvss.n2302 292.5
R15112 dvss.n2299 dvss.n2298 292.5
R15113 dvss.n2296 dvss.n2292 292.5
R15114 dvss.n2306 dvss.n2305 292.5
R15115 dvss.n2308 dvss.n2307 292.5
R15116 dvss.n2289 dvss.n2150 292.5
R15117 dvss.n2325 dvss.n2150 292.5
R15118 dvss.n2290 dvss.n2168 292.5
R15119 dvss.n2295 dvss.n2293 292.5
R15120 dvss.n2303 dvss.n2167 292.5
R15121 dvss.n2165 dvss.n2164 292.5
R15122 dvss.n2314 dvss.n2313 292.5
R15123 dvss.n2317 dvss.n2316 292.5
R15124 dvss.n2159 dvss.n2158 292.5
R15125 dvss.n2323 dvss.n2322 292.5
R15126 dvss.n2156 dvss.n2148 292.5
R15127 dvss.n2328 dvss.n2327 292.5
R15128 dvss.n2149 dvss.n2147 292.5
R15129 dvss.n2147 dvss.n2145 292.5
R15130 dvss.n2284 dvss.n2283 292.5
R15131 dvss.n2285 dvss.n2284 292.5
R15132 dvss.n2282 dvss.n2173 292.5
R15133 dvss.n2177 dvss.n2173 292.5
R15134 dvss.n2281 dvss.n2280 292.5
R15135 dvss.n2280 dvss.n2279 292.5
R15136 dvss.n2271 dvss.n2222 292.5
R15137 dvss.n2186 dvss.n2185 292.5
R15138 dvss.n2187 dvss.n2186 292.5
R15139 dvss.n2219 dvss.n2218 292.5
R15140 dvss.n2218 dvss.n2217 292.5
R15141 dvss.n2220 dvss.n2184 292.5
R15142 dvss.n2184 dvss.n2183 292.5
R15143 dvss.n2222 dvss.n2221 292.5
R15144 dvss.n2274 dvss.n2178 292.5
R15145 dvss.n2268 dvss.n2267 292.5
R15146 dvss.n2267 dvss.n2175 292.5
R15147 dvss.n2228 dvss.n2226 292.5
R15148 dvss.n2233 dvss.n2228 292.5
R15149 dvss.n2262 dvss.n2230 292.5
R15150 dvss.n2262 dvss.n2261 292.5
R15151 dvss.n2236 dvss.n2235 292.5
R15152 dvss.n2260 dvss.n2236 292.5
R15153 dvss.n2257 dvss.n2239 292.5
R15154 dvss.n2258 dvss.n2257 292.5
R15155 dvss.n2241 dvss.n2240 292.5
R15156 dvss.n2241 dvss.n2237 292.5
R15157 dvss.n2252 dvss.n2245 292.5
R15158 dvss.n2252 dvss.n2251 292.5
R15159 dvss.n2250 dvss.n2248 292.5
R15160 dvss.n2248 dvss.n2247 292.5
R15161 dvss.n2274 dvss.n2273 292.5
R15162 dvss.n2355 dvss.n2354 292.5
R15163 dvss.n2340 dvss.n2339 292.5
R15164 dvss.n2342 dvss.n2341 292.5
R15165 dvss.n2344 dvss.n2343 292.5
R15166 dvss.n2346 dvss.n2345 292.5
R15167 dvss.n2348 dvss.n2347 292.5
R15168 dvss.n2350 dvss.n2349 292.5
R15169 dvss.n2092 dvss.n2091 292.5
R15170 dvss.n2338 dvss.n2093 292.5
R15171 dvss.n2352 dvss.n2093 292.5
R15172 dvss.n2018 dvss.n2017 292.5
R15173 dvss.n2018 dvss.n2010 292.5
R15174 dvss.n2031 dvss.n2013 292.5
R15175 dvss.n2030 dvss.n2029 292.5
R15176 dvss.n2028 dvss.n2027 292.5
R15177 dvss.n2026 dvss.n2015 292.5
R15178 dvss.n2024 dvss.n2023 292.5
R15179 dvss.n2022 dvss.n2016 292.5
R15180 dvss.n2021 dvss.n2020 292.5
R15181 dvss.n2034 dvss.n2033 292.5
R15182 dvss.n2068 dvss.n2065 292.5
R15183 dvss.n2081 dvss.n2061 292.5
R15184 dvss.n2079 dvss.n2078 292.5
R15185 dvss.n2077 dvss.n2076 292.5
R15186 dvss.n2074 dvss.n2063 292.5
R15187 dvss.n2072 dvss.n2071 292.5
R15188 dvss.n2070 dvss.n2069 292.5
R15189 dvss.n2083 dvss.n2082 292.5
R15190 dvss.n2082 dvss.n2057 292.5
R15191 dvss.n2066 dvss.n2052 292.5
R15192 dvss.n2438 dvss.n2007 292.5
R15193 dvss.n2007 dvss.n2005 292.5
R15194 dvss.n2440 dvss.n2439 292.5
R15195 dvss.n2441 dvss.n2440 292.5
R15196 dvss.n2414 dvss.n2006 292.5
R15197 dvss.n2011 dvss.n2006 292.5
R15198 dvss.n2413 dvss.n2412 292.5
R15199 dvss.n2412 dvss.n2411 292.5
R15200 dvss.n2398 dvss.n2397 292.5
R15201 dvss.n2399 dvss.n2398 292.5
R15202 dvss.n2396 dvss.n2041 292.5
R15203 dvss.n2041 dvss.n2040 292.5
R15204 dvss.n2395 dvss.n2394 292.5
R15205 dvss.n2394 dvss.n2393 292.5
R15206 dvss.n2043 dvss.n2042 292.5
R15207 dvss.n2044 dvss.n2043 292.5
R15208 dvss.n2379 dvss.n2378 292.5
R15209 dvss.n2380 dvss.n2379 292.5
R15210 dvss.n2377 dvss.n2051 292.5
R15211 dvss.n2051 dvss.n2050 292.5
R15212 dvss.n2375 dvss.n2374 292.5
R15213 dvss.n2374 dvss.n2373 292.5
R15214 dvss.n2054 dvss.n2053 292.5
R15215 dvss.n2056 dvss.n2054 292.5
R15216 dvss.n2358 dvss.n2357 292.5
R15217 dvss.n2359 dvss.n2358 292.5
R15218 dvss.n2356 dvss.n2090 292.5
R15219 dvss.n2090 dvss.n2089 292.5
R15220 dvss.n2437 dvss.n2436 292.5
R15221 dvss.n2416 dvss.n2415 292.5
R15222 dvss.n2432 dvss.n2431 292.5
R15223 dvss.n2430 dvss.n2421 292.5
R15224 dvss.n2429 dvss.n2428 292.5
R15225 dvss.n2427 dvss.n2426 292.5
R15226 dvss.n2425 dvss.n2424 292.5
R15227 dvss.n2423 dvss.n2422 292.5
R15228 dvss.n2417 dvss.n1999 292.5
R15229 dvss.n1041 dvss.n948 292.5
R15230 dvss.n1041 dvss.n1040 292.5
R15231 dvss.n985 dvss.n984 292.5
R15232 dvss.n986 dvss.n985 292.5
R15233 dvss.n983 dvss.n951 292.5
R15234 dvss.n952 dvss.n951 292.5
R15235 dvss.n982 dvss.n957 292.5
R15236 dvss.n957 dvss.n956 292.5
R15237 dvss.n976 dvss.n975 292.5
R15238 dvss.n974 dvss.n963 292.5
R15239 dvss.n973 dvss.n972 292.5
R15240 dvss.n971 dvss.n970 292.5
R15241 dvss.n969 dvss.n968 292.5
R15242 dvss.n967 dvss.n966 292.5
R15243 dvss.n965 dvss.n964 292.5
R15244 dvss.n959 dvss.n958 292.5
R15245 dvss.n981 dvss.n980 292.5
R15246 dvss.n1057 dvss.n1056 292.5
R15247 dvss.n1056 dvss.n918 292.5
R15248 dvss.n1055 dvss.n940 292.5
R15249 dvss.n1055 dvss.n1054 292.5
R15250 dvss.n1045 dvss.n941 292.5
R15251 dvss.n946 dvss.n941 292.5
R15252 dvss.n1047 dvss.n1046 292.5
R15253 dvss.n1048 dvss.n1047 292.5
R15254 dvss.n1069 dvss.n939 292.5
R15255 dvss.n1062 dvss.n939 292.5
R15256 dvss.n1071 dvss.n1070 292.5
R15257 dvss.n1072 dvss.n1071 292.5
R15258 dvss.n1068 dvss.n1067 292.5
R15259 dvss.n1065 dvss.n1061 292.5
R15260 dvss.n1075 dvss.n1074 292.5
R15261 dvss.n1077 dvss.n1076 292.5
R15262 dvss.n1058 dvss.n919 292.5
R15263 dvss.n1094 dvss.n919 292.5
R15264 dvss.n1059 dvss.n937 292.5
R15265 dvss.n1064 dvss.n1062 292.5
R15266 dvss.n1072 dvss.n936 292.5
R15267 dvss.n934 dvss.n933 292.5
R15268 dvss.n1083 dvss.n1082 292.5
R15269 dvss.n1086 dvss.n1085 292.5
R15270 dvss.n928 dvss.n927 292.5
R15271 dvss.n1092 dvss.n1091 292.5
R15272 dvss.n925 dvss.n917 292.5
R15273 dvss.n1097 dvss.n1096 292.5
R15274 dvss.n918 dvss.n916 292.5
R15275 dvss.n916 dvss.n914 292.5
R15276 dvss.n1053 dvss.n1052 292.5
R15277 dvss.n1054 dvss.n1053 292.5
R15278 dvss.n1051 dvss.n942 292.5
R15279 dvss.n946 dvss.n942 292.5
R15280 dvss.n1050 dvss.n1049 292.5
R15281 dvss.n1049 dvss.n1048 292.5
R15282 dvss.n1040 dvss.n991 292.5
R15283 dvss.n955 dvss.n954 292.5
R15284 dvss.n956 dvss.n955 292.5
R15285 dvss.n988 dvss.n987 292.5
R15286 dvss.n987 dvss.n986 292.5
R15287 dvss.n989 dvss.n953 292.5
R15288 dvss.n953 dvss.n952 292.5
R15289 dvss.n991 dvss.n990 292.5
R15290 dvss.n1043 dvss.n947 292.5
R15291 dvss.n1037 dvss.n1036 292.5
R15292 dvss.n1036 dvss.n944 292.5
R15293 dvss.n997 dvss.n995 292.5
R15294 dvss.n1002 dvss.n997 292.5
R15295 dvss.n1031 dvss.n999 292.5
R15296 dvss.n1031 dvss.n1030 292.5
R15297 dvss.n1005 dvss.n1004 292.5
R15298 dvss.n1029 dvss.n1005 292.5
R15299 dvss.n1026 dvss.n1008 292.5
R15300 dvss.n1027 dvss.n1026 292.5
R15301 dvss.n1010 dvss.n1009 292.5
R15302 dvss.n1010 dvss.n1006 292.5
R15303 dvss.n1021 dvss.n1014 292.5
R15304 dvss.n1021 dvss.n1020 292.5
R15305 dvss.n1019 dvss.n1017 292.5
R15306 dvss.n1017 dvss.n1016 292.5
R15307 dvss.n1043 dvss.n1042 292.5
R15308 dvss.n1124 dvss.n1123 292.5
R15309 dvss.n1109 dvss.n1108 292.5
R15310 dvss.n1111 dvss.n1110 292.5
R15311 dvss.n1113 dvss.n1112 292.5
R15312 dvss.n1115 dvss.n1114 292.5
R15313 dvss.n1117 dvss.n1116 292.5
R15314 dvss.n1119 dvss.n1118 292.5
R15315 dvss.n861 dvss.n860 292.5
R15316 dvss.n1107 dvss.n862 292.5
R15317 dvss.n1121 dvss.n862 292.5
R15318 dvss.n787 dvss.n786 292.5
R15319 dvss.n787 dvss.n779 292.5
R15320 dvss.n800 dvss.n782 292.5
R15321 dvss.n799 dvss.n798 292.5
R15322 dvss.n797 dvss.n796 292.5
R15323 dvss.n795 dvss.n784 292.5
R15324 dvss.n793 dvss.n792 292.5
R15325 dvss.n791 dvss.n785 292.5
R15326 dvss.n790 dvss.n789 292.5
R15327 dvss.n803 dvss.n802 292.5
R15328 dvss.n837 dvss.n834 292.5
R15329 dvss.n850 dvss.n830 292.5
R15330 dvss.n848 dvss.n847 292.5
R15331 dvss.n846 dvss.n845 292.5
R15332 dvss.n843 dvss.n832 292.5
R15333 dvss.n841 dvss.n840 292.5
R15334 dvss.n839 dvss.n838 292.5
R15335 dvss.n852 dvss.n851 292.5
R15336 dvss.n851 dvss.n826 292.5
R15337 dvss.n835 dvss.n821 292.5
R15338 dvss.n1207 dvss.n776 292.5
R15339 dvss.n776 dvss.n774 292.5
R15340 dvss.n1209 dvss.n1208 292.5
R15341 dvss.n1210 dvss.n1209 292.5
R15342 dvss.n1183 dvss.n775 292.5
R15343 dvss.n780 dvss.n775 292.5
R15344 dvss.n1182 dvss.n1181 292.5
R15345 dvss.n1181 dvss.n1180 292.5
R15346 dvss.n1167 dvss.n1166 292.5
R15347 dvss.n1168 dvss.n1167 292.5
R15348 dvss.n1165 dvss.n810 292.5
R15349 dvss.n810 dvss.n809 292.5
R15350 dvss.n1164 dvss.n1163 292.5
R15351 dvss.n1163 dvss.n1162 292.5
R15352 dvss.n812 dvss.n811 292.5
R15353 dvss.n813 dvss.n812 292.5
R15354 dvss.n1148 dvss.n1147 292.5
R15355 dvss.n1149 dvss.n1148 292.5
R15356 dvss.n1146 dvss.n820 292.5
R15357 dvss.n820 dvss.n819 292.5
R15358 dvss.n1144 dvss.n1143 292.5
R15359 dvss.n1143 dvss.n1142 292.5
R15360 dvss.n823 dvss.n822 292.5
R15361 dvss.n825 dvss.n823 292.5
R15362 dvss.n1127 dvss.n1126 292.5
R15363 dvss.n1128 dvss.n1127 292.5
R15364 dvss.n1125 dvss.n859 292.5
R15365 dvss.n859 dvss.n858 292.5
R15366 dvss.n1206 dvss.n1205 292.5
R15367 dvss.n1185 dvss.n1184 292.5
R15368 dvss.n1201 dvss.n1200 292.5
R15369 dvss.n1199 dvss.n1190 292.5
R15370 dvss.n1198 dvss.n1197 292.5
R15371 dvss.n1196 dvss.n1195 292.5
R15372 dvss.n1194 dvss.n1193 292.5
R15373 dvss.n1192 dvss.n1191 292.5
R15374 dvss.n1186 dvss.n768 292.5
R15375 dvss.n429 dvss.n336 292.5
R15376 dvss.n429 dvss.n428 292.5
R15377 dvss.n373 dvss.n372 292.5
R15378 dvss.n374 dvss.n373 292.5
R15379 dvss.n371 dvss.n339 292.5
R15380 dvss.n340 dvss.n339 292.5
R15381 dvss.n370 dvss.n345 292.5
R15382 dvss.n345 dvss.n344 292.5
R15383 dvss.n364 dvss.n363 292.5
R15384 dvss.n362 dvss.n351 292.5
R15385 dvss.n361 dvss.n360 292.5
R15386 dvss.n359 dvss.n358 292.5
R15387 dvss.n357 dvss.n356 292.5
R15388 dvss.n355 dvss.n354 292.5
R15389 dvss.n353 dvss.n352 292.5
R15390 dvss.n347 dvss.n346 292.5
R15391 dvss.n369 dvss.n368 292.5
R15392 dvss.n445 dvss.n444 292.5
R15393 dvss.n444 dvss.n306 292.5
R15394 dvss.n443 dvss.n328 292.5
R15395 dvss.n443 dvss.n442 292.5
R15396 dvss.n433 dvss.n329 292.5
R15397 dvss.n334 dvss.n329 292.5
R15398 dvss.n435 dvss.n434 292.5
R15399 dvss.n436 dvss.n435 292.5
R15400 dvss.n457 dvss.n327 292.5
R15401 dvss.n450 dvss.n327 292.5
R15402 dvss.n459 dvss.n458 292.5
R15403 dvss.n460 dvss.n459 292.5
R15404 dvss.n456 dvss.n455 292.5
R15405 dvss.n453 dvss.n449 292.5
R15406 dvss.n463 dvss.n462 292.5
R15407 dvss.n465 dvss.n464 292.5
R15408 dvss.n446 dvss.n307 292.5
R15409 dvss.n482 dvss.n307 292.5
R15410 dvss.n447 dvss.n325 292.5
R15411 dvss.n452 dvss.n450 292.5
R15412 dvss.n460 dvss.n324 292.5
R15413 dvss.n322 dvss.n321 292.5
R15414 dvss.n471 dvss.n470 292.5
R15415 dvss.n474 dvss.n473 292.5
R15416 dvss.n316 dvss.n315 292.5
R15417 dvss.n480 dvss.n479 292.5
R15418 dvss.n313 dvss.n305 292.5
R15419 dvss.n485 dvss.n484 292.5
R15420 dvss.n306 dvss.n304 292.5
R15421 dvss.n304 dvss.n302 292.5
R15422 dvss.n441 dvss.n440 292.5
R15423 dvss.n442 dvss.n441 292.5
R15424 dvss.n439 dvss.n330 292.5
R15425 dvss.n334 dvss.n330 292.5
R15426 dvss.n438 dvss.n437 292.5
R15427 dvss.n437 dvss.n436 292.5
R15428 dvss.n428 dvss.n379 292.5
R15429 dvss.n343 dvss.n342 292.5
R15430 dvss.n344 dvss.n343 292.5
R15431 dvss.n376 dvss.n375 292.5
R15432 dvss.n375 dvss.n374 292.5
R15433 dvss.n377 dvss.n341 292.5
R15434 dvss.n341 dvss.n340 292.5
R15435 dvss.n379 dvss.n378 292.5
R15436 dvss.n431 dvss.n335 292.5
R15437 dvss.n425 dvss.n424 292.5
R15438 dvss.n424 dvss.n332 292.5
R15439 dvss.n385 dvss.n383 292.5
R15440 dvss.n390 dvss.n385 292.5
R15441 dvss.n419 dvss.n387 292.5
R15442 dvss.n419 dvss.n418 292.5
R15443 dvss.n393 dvss.n392 292.5
R15444 dvss.n417 dvss.n393 292.5
R15445 dvss.n414 dvss.n396 292.5
R15446 dvss.n415 dvss.n414 292.5
R15447 dvss.n398 dvss.n397 292.5
R15448 dvss.n398 dvss.n394 292.5
R15449 dvss.n409 dvss.n402 292.5
R15450 dvss.n409 dvss.n408 292.5
R15451 dvss.n407 dvss.n405 292.5
R15452 dvss.n405 dvss.n404 292.5
R15453 dvss.n431 dvss.n430 292.5
R15454 dvss.n512 dvss.n511 292.5
R15455 dvss.n497 dvss.n496 292.5
R15456 dvss.n499 dvss.n498 292.5
R15457 dvss.n501 dvss.n500 292.5
R15458 dvss.n503 dvss.n502 292.5
R15459 dvss.n505 dvss.n504 292.5
R15460 dvss.n507 dvss.n506 292.5
R15461 dvss.n249 dvss.n248 292.5
R15462 dvss.n495 dvss.n250 292.5
R15463 dvss.n509 dvss.n250 292.5
R15464 dvss.n175 dvss.n174 292.5
R15465 dvss.n175 dvss.n167 292.5
R15466 dvss.n188 dvss.n170 292.5
R15467 dvss.n187 dvss.n186 292.5
R15468 dvss.n185 dvss.n184 292.5
R15469 dvss.n183 dvss.n172 292.5
R15470 dvss.n181 dvss.n180 292.5
R15471 dvss.n179 dvss.n173 292.5
R15472 dvss.n178 dvss.n177 292.5
R15473 dvss.n191 dvss.n190 292.5
R15474 dvss.n225 dvss.n222 292.5
R15475 dvss.n238 dvss.n218 292.5
R15476 dvss.n236 dvss.n235 292.5
R15477 dvss.n234 dvss.n233 292.5
R15478 dvss.n231 dvss.n220 292.5
R15479 dvss.n229 dvss.n228 292.5
R15480 dvss.n227 dvss.n226 292.5
R15481 dvss.n240 dvss.n239 292.5
R15482 dvss.n239 dvss.n214 292.5
R15483 dvss.n223 dvss.n209 292.5
R15484 dvss.n595 dvss.n164 292.5
R15485 dvss.n164 dvss.n162 292.5
R15486 dvss.n597 dvss.n596 292.5
R15487 dvss.n598 dvss.n597 292.5
R15488 dvss.n571 dvss.n163 292.5
R15489 dvss.n168 dvss.n163 292.5
R15490 dvss.n570 dvss.n569 292.5
R15491 dvss.n569 dvss.n568 292.5
R15492 dvss.n555 dvss.n554 292.5
R15493 dvss.n556 dvss.n555 292.5
R15494 dvss.n553 dvss.n198 292.5
R15495 dvss.n198 dvss.n197 292.5
R15496 dvss.n552 dvss.n551 292.5
R15497 dvss.n551 dvss.n550 292.5
R15498 dvss.n200 dvss.n199 292.5
R15499 dvss.n201 dvss.n200 292.5
R15500 dvss.n536 dvss.n535 292.5
R15501 dvss.n537 dvss.n536 292.5
R15502 dvss.n534 dvss.n208 292.5
R15503 dvss.n208 dvss.n207 292.5
R15504 dvss.n532 dvss.n531 292.5
R15505 dvss.n531 dvss.n530 292.5
R15506 dvss.n211 dvss.n210 292.5
R15507 dvss.n213 dvss.n211 292.5
R15508 dvss.n515 dvss.n514 292.5
R15509 dvss.n516 dvss.n515 292.5
R15510 dvss.n513 dvss.n247 292.5
R15511 dvss.n247 dvss.n246 292.5
R15512 dvss.n594 dvss.n593 292.5
R15513 dvss.n573 dvss.n572 292.5
R15514 dvss.n589 dvss.n588 292.5
R15515 dvss.n587 dvss.n578 292.5
R15516 dvss.n586 dvss.n585 292.5
R15517 dvss.n584 dvss.n583 292.5
R15518 dvss.n582 dvss.n581 292.5
R15519 dvss.n580 dvss.n579 292.5
R15520 dvss.n574 dvss.n156 292.5
R15521 dvss.n1248 dvss.t45 286.554
R15522 dvss.n1864 dvss.t77 286.554
R15523 dvss.n633 dvss.t14 286.554
R15524 dvss.n20 dvss.t129 286.554
R15525 dvss.n1754 dvss.n1441 270.034
R15526 dvss.n1794 dvss.n1391 270.034
R15527 dvss.n1792 dvss.n1394 270.034
R15528 dvss.n1756 dvss.n1437 270.034
R15529 dvss.n2372 dvss.n2059 270.034
R15530 dvss.n2412 dvss.n2009 270.034
R15531 dvss.n2410 dvss.n2012 270.034
R15532 dvss.n2374 dvss.n2055 270.034
R15533 dvss.n1141 dvss.n828 270.034
R15534 dvss.n1181 dvss.n778 270.034
R15535 dvss.n1179 dvss.n781 270.034
R15536 dvss.n1143 dvss.n824 270.034
R15537 dvss.n529 dvss.n216 270.034
R15538 dvss.n569 dvss.n166 270.034
R15539 dvss.n567 dvss.n169 270.034
R15540 dvss.n531 dvss.n212 270.034
R15541 dvss.n2566 dvss.t43 268.067
R15542 dvss.n2496 dvss.t75 268.067
R15543 dvss.n2842 dvss.t12 268.067
R15544 dvss.n2915 dvss.t127 268.067
R15545 dvss.n1444 dvss.n1439 248.682
R15546 dvss.n1457 dvss.n1439 248.682
R15547 dvss.n1455 dvss.n1439 248.682
R15548 dvss.n2062 dvss.n2057 248.682
R15549 dvss.n2075 dvss.n2057 248.682
R15550 dvss.n2073 dvss.n2057 248.682
R15551 dvss.n831 dvss.n826 248.682
R15552 dvss.n844 dvss.n826 248.682
R15553 dvss.n842 dvss.n826 248.682
R15554 dvss.n219 dvss.n214 248.682
R15555 dvss.n232 dvss.n214 248.682
R15556 dvss.n230 dvss.n214 248.682
R15557 dvss.n1707 dvss.n1534 245.511
R15558 dvss.n1707 dvss.n1535 245.511
R15559 dvss.n1707 dvss.n1536 245.511
R15560 dvss.n1707 dvss.n1537 245.511
R15561 dvss.n1707 dvss.n1706 245.511
R15562 dvss.n1734 dvss.n1477 245.511
R15563 dvss.n1734 dvss.n1478 245.511
R15564 dvss.n1734 dvss.n1479 245.511
R15565 dvss.n1734 dvss.n1480 245.511
R15566 dvss.n1734 dvss.n1733 245.511
R15567 dvss.n2325 dvss.n2152 245.511
R15568 dvss.n2325 dvss.n2153 245.511
R15569 dvss.n2325 dvss.n2154 245.511
R15570 dvss.n2325 dvss.n2155 245.511
R15571 dvss.n2325 dvss.n2324 245.511
R15572 dvss.n2352 dvss.n2095 245.511
R15573 dvss.n2352 dvss.n2096 245.511
R15574 dvss.n2352 dvss.n2097 245.511
R15575 dvss.n2352 dvss.n2098 245.511
R15576 dvss.n2352 dvss.n2351 245.511
R15577 dvss.n1094 dvss.n921 245.511
R15578 dvss.n1094 dvss.n922 245.511
R15579 dvss.n1094 dvss.n923 245.511
R15580 dvss.n1094 dvss.n924 245.511
R15581 dvss.n1094 dvss.n1093 245.511
R15582 dvss.n1121 dvss.n864 245.511
R15583 dvss.n1121 dvss.n865 245.511
R15584 dvss.n1121 dvss.n866 245.511
R15585 dvss.n1121 dvss.n867 245.511
R15586 dvss.n1121 dvss.n1120 245.511
R15587 dvss.n482 dvss.n309 245.511
R15588 dvss.n482 dvss.n310 245.511
R15589 dvss.n482 dvss.n311 245.511
R15590 dvss.n482 dvss.n312 245.511
R15591 dvss.n482 dvss.n481 245.511
R15592 dvss.n509 dvss.n252 245.511
R15593 dvss.n509 dvss.n253 245.511
R15594 dvss.n509 dvss.n254 245.511
R15595 dvss.n509 dvss.n255 245.511
R15596 dvss.n509 dvss.n508 245.511
R15597 dvss.n2614 dvss.t176 241.6
R15598 dvss.n1339 dvss.t105 240.336
R15599 dvss.n1957 dvss.t93 240.336
R15600 dvss.n726 dvss.t192 240.336
R15601 dvss.n114 dvss.t65 240.336
R15602 dvss.n1585 dvss.n1584 223.931
R15603 dvss.n1581 dvss.n1580 223.931
R15604 dvss.n1577 dvss.n1572 223.931
R15605 dvss.n1600 dvss.n1568 223.931
R15606 dvss.n1600 dvss.n1566 223.931
R15607 dvss.n1604 dvss.n1566 223.931
R15608 dvss.n1617 dvss.n1612 223.931
R15609 dvss.n1622 dvss.n1621 223.931
R15610 dvss.n1629 dvss.n1627 223.931
R15611 dvss.n1598 dvss.n1570 223.931
R15612 dvss.n1598 dvss.n1564 223.931
R15613 dvss.n1654 dvss.n1564 223.931
R15614 dvss.n1643 dvss.n1642 223.931
R15615 dvss.n1640 dvss.n1619 223.931
R15616 dvss.n1633 dvss.n1632 223.931
R15617 dvss.n1662 dvss.n1555 223.931
R15618 dvss.n1666 dvss.n1555 223.931
R15619 dvss.n1666 dvss.n1529 223.931
R15620 dvss.n1689 dvss.n1532 223.931
R15621 dvss.n1660 dvss.n1554 223.931
R15622 dvss.n1668 dvss.n1554 223.931
R15623 dvss.n1669 dvss.n1668 223.931
R15624 dvss.n1742 dvss.n1470 223.931
R15625 dvss.n1742 dvss.n1440 223.931
R15626 dvss.n1754 dvss.n1440 223.931
R15627 dvss.n1721 dvss.n1475 223.931
R15628 dvss.n1794 dvss.n1388 223.931
R15629 dvss.n1822 dvss.n1388 223.931
R15630 dvss.n1822 dvss.n1389 223.931
R15631 dvss.n1814 dvss.n1803 223.931
R15632 dvss.n1810 dvss.n1809 223.931
R15633 dvss.n1806 dvss.n1805 223.931
R15634 dvss.n1792 dvss.n1385 223.931
R15635 dvss.n1824 dvss.n1385 223.931
R15636 dvss.n1824 dvss.n1386 223.931
R15637 dvss.n1763 dvss.n1431 223.931
R15638 dvss.n1763 dvss.n1427 223.931
R15639 dvss.n1774 dvss.n1427 223.931
R15640 dvss.n1774 dvss.n1421 223.931
R15641 dvss.n1782 dvss.n1421 223.931
R15642 dvss.n1761 dvss.n1433 223.931
R15643 dvss.n1761 dvss.n1425 223.931
R15644 dvss.n1776 dvss.n1425 223.931
R15645 dvss.n1776 dvss.n1423 223.931
R15646 dvss.n1780 dvss.n1423 223.931
R15647 dvss.n1740 dvss.n1472 223.931
R15648 dvss.n1740 dvss.n1436 223.931
R15649 dvss.n1756 dvss.n1436 223.931
R15650 dvss.n2203 dvss.n2202 223.931
R15651 dvss.n2199 dvss.n2198 223.931
R15652 dvss.n2195 dvss.n2190 223.931
R15653 dvss.n2218 dvss.n2186 223.931
R15654 dvss.n2218 dvss.n2184 223.931
R15655 dvss.n2222 dvss.n2184 223.931
R15656 dvss.n2235 dvss.n2230 223.931
R15657 dvss.n2240 dvss.n2239 223.931
R15658 dvss.n2247 dvss.n2245 223.931
R15659 dvss.n2216 dvss.n2188 223.931
R15660 dvss.n2216 dvss.n2182 223.931
R15661 dvss.n2272 dvss.n2182 223.931
R15662 dvss.n2261 dvss.n2260 223.931
R15663 dvss.n2258 dvss.n2237 223.931
R15664 dvss.n2251 dvss.n2250 223.931
R15665 dvss.n2280 dvss.n2173 223.931
R15666 dvss.n2284 dvss.n2173 223.931
R15667 dvss.n2284 dvss.n2147 223.931
R15668 dvss.n2307 dvss.n2150 223.931
R15669 dvss.n2278 dvss.n2172 223.931
R15670 dvss.n2286 dvss.n2172 223.931
R15671 dvss.n2287 dvss.n2286 223.931
R15672 dvss.n2360 dvss.n2088 223.931
R15673 dvss.n2360 dvss.n2058 223.931
R15674 dvss.n2372 dvss.n2058 223.931
R15675 dvss.n2339 dvss.n2093 223.931
R15676 dvss.n2412 dvss.n2006 223.931
R15677 dvss.n2440 dvss.n2006 223.931
R15678 dvss.n2440 dvss.n2007 223.931
R15679 dvss.n2432 dvss.n2421 223.931
R15680 dvss.n2428 dvss.n2427 223.931
R15681 dvss.n2424 dvss.n2423 223.931
R15682 dvss.n2410 dvss.n2003 223.931
R15683 dvss.n2442 dvss.n2003 223.931
R15684 dvss.n2442 dvss.n2004 223.931
R15685 dvss.n2381 dvss.n2049 223.931
R15686 dvss.n2381 dvss.n2045 223.931
R15687 dvss.n2392 dvss.n2045 223.931
R15688 dvss.n2392 dvss.n2039 223.931
R15689 dvss.n2400 dvss.n2039 223.931
R15690 dvss.n2379 dvss.n2051 223.931
R15691 dvss.n2379 dvss.n2043 223.931
R15692 dvss.n2394 dvss.n2043 223.931
R15693 dvss.n2394 dvss.n2041 223.931
R15694 dvss.n2398 dvss.n2041 223.931
R15695 dvss.n2358 dvss.n2090 223.931
R15696 dvss.n2358 dvss.n2054 223.931
R15697 dvss.n2374 dvss.n2054 223.931
R15698 dvss.n972 dvss.n971 223.931
R15699 dvss.n968 dvss.n967 223.931
R15700 dvss.n964 dvss.n959 223.931
R15701 dvss.n987 dvss.n955 223.931
R15702 dvss.n987 dvss.n953 223.931
R15703 dvss.n991 dvss.n953 223.931
R15704 dvss.n1004 dvss.n999 223.931
R15705 dvss.n1009 dvss.n1008 223.931
R15706 dvss.n1016 dvss.n1014 223.931
R15707 dvss.n985 dvss.n957 223.931
R15708 dvss.n985 dvss.n951 223.931
R15709 dvss.n1041 dvss.n951 223.931
R15710 dvss.n1030 dvss.n1029 223.931
R15711 dvss.n1027 dvss.n1006 223.931
R15712 dvss.n1020 dvss.n1019 223.931
R15713 dvss.n1049 dvss.n942 223.931
R15714 dvss.n1053 dvss.n942 223.931
R15715 dvss.n1053 dvss.n916 223.931
R15716 dvss.n1076 dvss.n919 223.931
R15717 dvss.n1047 dvss.n941 223.931
R15718 dvss.n1055 dvss.n941 223.931
R15719 dvss.n1056 dvss.n1055 223.931
R15720 dvss.n1129 dvss.n857 223.931
R15721 dvss.n1129 dvss.n827 223.931
R15722 dvss.n1141 dvss.n827 223.931
R15723 dvss.n1108 dvss.n862 223.931
R15724 dvss.n1181 dvss.n775 223.931
R15725 dvss.n1209 dvss.n775 223.931
R15726 dvss.n1209 dvss.n776 223.931
R15727 dvss.n1201 dvss.n1190 223.931
R15728 dvss.n1197 dvss.n1196 223.931
R15729 dvss.n1193 dvss.n1192 223.931
R15730 dvss.n1179 dvss.n772 223.931
R15731 dvss.n1211 dvss.n772 223.931
R15732 dvss.n1211 dvss.n773 223.931
R15733 dvss.n1150 dvss.n818 223.931
R15734 dvss.n1150 dvss.n814 223.931
R15735 dvss.n1161 dvss.n814 223.931
R15736 dvss.n1161 dvss.n808 223.931
R15737 dvss.n1169 dvss.n808 223.931
R15738 dvss.n1148 dvss.n820 223.931
R15739 dvss.n1148 dvss.n812 223.931
R15740 dvss.n1163 dvss.n812 223.931
R15741 dvss.n1163 dvss.n810 223.931
R15742 dvss.n1167 dvss.n810 223.931
R15743 dvss.n1127 dvss.n859 223.931
R15744 dvss.n1127 dvss.n823 223.931
R15745 dvss.n1143 dvss.n823 223.931
R15746 dvss.n360 dvss.n359 223.931
R15747 dvss.n356 dvss.n355 223.931
R15748 dvss.n352 dvss.n347 223.931
R15749 dvss.n375 dvss.n343 223.931
R15750 dvss.n375 dvss.n341 223.931
R15751 dvss.n379 dvss.n341 223.931
R15752 dvss.n392 dvss.n387 223.931
R15753 dvss.n397 dvss.n396 223.931
R15754 dvss.n404 dvss.n402 223.931
R15755 dvss.n373 dvss.n345 223.931
R15756 dvss.n373 dvss.n339 223.931
R15757 dvss.n429 dvss.n339 223.931
R15758 dvss.n418 dvss.n417 223.931
R15759 dvss.n415 dvss.n394 223.931
R15760 dvss.n408 dvss.n407 223.931
R15761 dvss.n437 dvss.n330 223.931
R15762 dvss.n441 dvss.n330 223.931
R15763 dvss.n441 dvss.n304 223.931
R15764 dvss.n464 dvss.n307 223.931
R15765 dvss.n435 dvss.n329 223.931
R15766 dvss.n443 dvss.n329 223.931
R15767 dvss.n444 dvss.n443 223.931
R15768 dvss.n517 dvss.n245 223.931
R15769 dvss.n517 dvss.n215 223.931
R15770 dvss.n529 dvss.n215 223.931
R15771 dvss.n496 dvss.n250 223.931
R15772 dvss.n569 dvss.n163 223.931
R15773 dvss.n597 dvss.n163 223.931
R15774 dvss.n597 dvss.n164 223.931
R15775 dvss.n589 dvss.n578 223.931
R15776 dvss.n585 dvss.n584 223.931
R15777 dvss.n581 dvss.n580 223.931
R15778 dvss.n567 dvss.n160 223.931
R15779 dvss.n599 dvss.n160 223.931
R15780 dvss.n599 dvss.n161 223.931
R15781 dvss.n538 dvss.n206 223.931
R15782 dvss.n538 dvss.n202 223.931
R15783 dvss.n549 dvss.n202 223.931
R15784 dvss.n549 dvss.n196 223.931
R15785 dvss.n557 dvss.n196 223.931
R15786 dvss.n536 dvss.n208 223.931
R15787 dvss.n536 dvss.n200 223.931
R15788 dvss.n551 dvss.n200 223.931
R15789 dvss.n551 dvss.n198 223.931
R15790 dvss.n555 dvss.n198 223.931
R15791 dvss.n515 dvss.n247 223.931
R15792 dvss.n515 dvss.n211 223.931
R15793 dvss.n531 dvss.n211 223.931
R15794 dvss.t20 dvss.n1426 220.982
R15795 dvss.n1775 dvss.t19 220.982
R15796 dvss.t136 dvss.n2044 220.982
R15797 dvss.n2393 dvss.t135 220.982
R15798 dvss.t24 dvss.n813 220.982
R15799 dvss.n1162 dvss.t114 220.982
R15800 dvss.t23 dvss.n201 220.982
R15801 dvss.n550 dvss.t137 220.982
R15802 dvss.n1402 dvss.n1400 206.158
R15803 dvss.n1406 dvss.n1398 206.158
R15804 dvss.n1409 dvss.n1408 206.158
R15805 dvss.n1413 dvss.n1412 206.158
R15806 dvss.n1451 dvss.n1450 206.158
R15807 dvss.n1464 dvss.n1463 206.158
R15808 dvss.n2020 dvss.n2018 206.158
R15809 dvss.n2024 dvss.n2016 206.158
R15810 dvss.n2027 dvss.n2026 206.158
R15811 dvss.n2031 dvss.n2030 206.158
R15812 dvss.n2069 dvss.n2068 206.158
R15813 dvss.n2082 dvss.n2081 206.158
R15814 dvss.n789 dvss.n787 206.158
R15815 dvss.n793 dvss.n785 206.158
R15816 dvss.n796 dvss.n795 206.158
R15817 dvss.n800 dvss.n799 206.158
R15818 dvss.n838 dvss.n837 206.158
R15819 dvss.n851 dvss.n850 206.158
R15820 dvss.n177 dvss.n175 206.158
R15821 dvss.n181 dvss.n173 206.158
R15822 dvss.n184 dvss.n183 206.158
R15823 dvss.n188 dvss.n187 206.158
R15824 dvss.n226 dvss.n225 206.158
R15825 dvss.n239 dvss.n238 206.158
R15826 dvss.n1351 dvss.t97 203.361
R15827 dvss.n1969 dvss.t87 203.361
R15828 dvss.n738 dvss.t186 203.361
R15829 dvss.n126 dvss.t69 203.361
R15830 dvss.t147 dvss.t119 187.113
R15831 dvss.n1521 dvss.n1508 185
R15832 dvss.n1523 dvss.n1522 185
R15833 dvss.n1500 dvss.n1487 185
R15834 dvss.n1502 dvss.n1501 185
R15835 dvss.n2139 dvss.n2126 185
R15836 dvss.n2141 dvss.n2140 185
R15837 dvss.n2118 dvss.n2105 185
R15838 dvss.n2120 dvss.n2119 185
R15839 dvss.n908 dvss.n895 185
R15840 dvss.n910 dvss.n909 185
R15841 dvss.n887 dvss.n874 185
R15842 dvss.n889 dvss.n888 185
R15843 dvss.n296 dvss.n283 185
R15844 dvss.n298 dvss.n297 185
R15845 dvss.n275 dvss.n262 185
R15846 dvss.n277 dvss.n276 185
R15847 dvss.n1599 dvss.t51 166.964
R15848 dvss.t51 dvss.n1565 166.964
R15849 dvss.n1559 dvss.t110 166.964
R15850 dvss.n1667 dvss.t110 166.964
R15851 dvss.n1741 dvss.t109 166.964
R15852 dvss.t109 dvss.n1438 166.964
R15853 dvss.n1393 dvss.t29 166.964
R15854 dvss.n1823 dvss.t29 166.964
R15855 dvss.n2217 dvss.t0 166.964
R15856 dvss.t0 dvss.n2183 166.964
R15857 dvss.n2177 dvss.t123 166.964
R15858 dvss.n2285 dvss.t123 166.964
R15859 dvss.n2359 dvss.t171 166.964
R15860 dvss.t171 dvss.n2056 166.964
R15861 dvss.n2011 dvss.t34 166.964
R15862 dvss.n2441 dvss.t34 166.964
R15863 dvss.n986 dvss.t35 166.964
R15864 dvss.t35 dvss.n952 166.964
R15865 dvss.n946 dvss.t161 166.964
R15866 dvss.n1054 dvss.t161 166.964
R15867 dvss.n1128 dvss.t140 166.964
R15868 dvss.t140 dvss.n825 166.964
R15869 dvss.n780 dvss.t18 166.964
R15870 dvss.n1210 dvss.t18 166.964
R15871 dvss.n374 dvss.t141 166.964
R15872 dvss.t141 dvss.n340 166.964
R15873 dvss.n334 dvss.t21 166.964
R15874 dvss.n442 dvss.t21 166.964
R15875 dvss.n516 dvss.t31 166.964
R15876 dvss.t31 dvss.n213 166.964
R15877 dvss.n168 dvss.t30 166.964
R15878 dvss.n598 dvss.t30 166.964
R15879 dvss.n1446 dvss.n1439 157.903
R15880 dvss.n2064 dvss.n2057 157.903
R15881 dvss.n833 dvss.n826 157.903
R15882 dvss.n221 dvss.n214 157.903
R15883 dvss.n1462 dvss.n1439 157.903
R15884 dvss.n2080 dvss.n2057 157.903
R15885 dvss.n849 dvss.n826 157.903
R15886 dvss.n237 dvss.n214 157.903
R15887 dvss.n1708 dvss.n1707 155.355
R15888 dvss.n2326 dvss.n2325 155.355
R15889 dvss.n1095 dvss.n1094 155.355
R15890 dvss.n483 dvss.n482 155.355
R15891 dvss.n1591 dvss.n1590 155.355
R15892 dvss.n1591 dvss.n1575 155.355
R15893 dvss.n1707 dvss.n1533 155.355
R15894 dvss.n1652 dvss.n1651 155.355
R15895 dvss.n1614 dvss.n1558 155.355
R15896 dvss.n1652 dvss.n1607 155.355
R15897 dvss.n1616 dvss.n1558 155.355
R15898 dvss.n1735 dvss.n1734 155.355
R15899 dvss.n1734 dvss.n1476 155.355
R15900 dvss.n1817 dvss.n1816 155.355
R15901 dvss.n1816 dvss.n1815 155.355
R15902 dvss.n2209 dvss.n2208 155.355
R15903 dvss.n2209 dvss.n2193 155.355
R15904 dvss.n2325 dvss.n2151 155.355
R15905 dvss.n2270 dvss.n2269 155.355
R15906 dvss.n2232 dvss.n2176 155.355
R15907 dvss.n2270 dvss.n2225 155.355
R15908 dvss.n2234 dvss.n2176 155.355
R15909 dvss.n2353 dvss.n2352 155.355
R15910 dvss.n2352 dvss.n2094 155.355
R15911 dvss.n2435 dvss.n2434 155.355
R15912 dvss.n2434 dvss.n2433 155.355
R15913 dvss.n978 dvss.n977 155.355
R15914 dvss.n978 dvss.n962 155.355
R15915 dvss.n1094 dvss.n920 155.355
R15916 dvss.n1039 dvss.n1038 155.355
R15917 dvss.n1001 dvss.n945 155.355
R15918 dvss.n1039 dvss.n994 155.355
R15919 dvss.n1003 dvss.n945 155.355
R15920 dvss.n1122 dvss.n1121 155.355
R15921 dvss.n1121 dvss.n863 155.355
R15922 dvss.n1204 dvss.n1203 155.355
R15923 dvss.n1203 dvss.n1202 155.355
R15924 dvss.n366 dvss.n365 155.355
R15925 dvss.n366 dvss.n350 155.355
R15926 dvss.n482 dvss.n308 155.355
R15927 dvss.n427 dvss.n426 155.355
R15928 dvss.n389 dvss.n333 155.355
R15929 dvss.n427 dvss.n382 155.355
R15930 dvss.n391 dvss.n333 155.355
R15931 dvss.n510 dvss.n509 155.355
R15932 dvss.n509 dvss.n251 155.355
R15933 dvss.n592 dvss.n591 155.355
R15934 dvss.n591 dvss.n590 155.355
R15935 dvss.n1314 dvss.t32 148.466
R15936 dvss.n1932 dvss.t121 148.466
R15937 dvss.n701 dvss.t159 148.466
R15938 dvss.n89 dvss.t112 148.466
R15939 dvss.n1359 dvss.t101 129.411
R15940 dvss.n1977 dvss.t83 129.411
R15941 dvss.n746 dvss.t188 129.411
R15942 dvss.n134 dvss.t59 129.411
R15943 dvss.n1516 dvss.t111 119.996
R15944 dvss.n1495 dvss.t52 119.996
R15945 dvss.n2134 dvss.t124 119.996
R15946 dvss.n2113 dvss.t1 119.996
R15947 dvss.n903 dvss.t162 119.996
R15948 dvss.n882 dvss.t36 119.996
R15949 dvss.n291 dvss.t22 119.996
R15950 dvss.n270 dvss.t142 119.996
R15951 dvss.n1708 dvss.n1530 118.937
R15952 dvss.n2326 dvss.n2148 118.937
R15953 dvss.n1095 dvss.n917 118.937
R15954 dvss.n483 dvss.n305 118.937
R15955 dvss.n1590 dvss.n1576 118.936
R15956 dvss.n1576 dvss.n1575 118.936
R15957 dvss.n1546 dvss.n1533 118.936
R15958 dvss.n1651 dvss.n1608 118.936
R15959 dvss.n1615 dvss.n1614 118.936
R15960 dvss.n1608 dvss.n1607 118.936
R15961 dvss.n1616 dvss.n1615 118.936
R15962 dvss.n1735 dvss.n1474 118.936
R15963 dvss.n1723 dvss.n1476 118.936
R15964 dvss.n1817 dvss.n1798 118.936
R15965 dvss.n1815 dvss.n1798 118.936
R15966 dvss.n2208 dvss.n2194 118.936
R15967 dvss.n2194 dvss.n2193 118.936
R15968 dvss.n2164 dvss.n2151 118.936
R15969 dvss.n2269 dvss.n2226 118.936
R15970 dvss.n2233 dvss.n2232 118.936
R15971 dvss.n2226 dvss.n2225 118.936
R15972 dvss.n2234 dvss.n2233 118.936
R15973 dvss.n2353 dvss.n2092 118.936
R15974 dvss.n2341 dvss.n2094 118.936
R15975 dvss.n2435 dvss.n2416 118.936
R15976 dvss.n2433 dvss.n2416 118.936
R15977 dvss.n977 dvss.n963 118.936
R15978 dvss.n963 dvss.n962 118.936
R15979 dvss.n933 dvss.n920 118.936
R15980 dvss.n1038 dvss.n995 118.936
R15981 dvss.n1002 dvss.n1001 118.936
R15982 dvss.n995 dvss.n994 118.936
R15983 dvss.n1003 dvss.n1002 118.936
R15984 dvss.n1122 dvss.n861 118.936
R15985 dvss.n1110 dvss.n863 118.936
R15986 dvss.n1204 dvss.n1185 118.936
R15987 dvss.n1202 dvss.n1185 118.936
R15988 dvss.n365 dvss.n351 118.936
R15989 dvss.n351 dvss.n350 118.936
R15990 dvss.n321 dvss.n308 118.936
R15991 dvss.n426 dvss.n383 118.936
R15992 dvss.n390 dvss.n389 118.936
R15993 dvss.n383 dvss.n382 118.936
R15994 dvss.n391 dvss.n390 118.936
R15995 dvss.n510 dvss.n249 118.936
R15996 dvss.n498 dvss.n251 118.936
R15997 dvss.n592 dvss.n573 118.936
R15998 dvss.n590 dvss.n573 118.936
R15999 dvss.n1680 dvss.n1679 117.718
R16000 dvss.n1687 dvss.n1686 117.718
R16001 dvss.n1677 dvss.n1676 117.718
R16002 dvss.n2298 dvss.n2297 117.718
R16003 dvss.n2305 dvss.n2304 117.718
R16004 dvss.n2295 dvss.n2294 117.718
R16005 dvss.n1067 dvss.n1066 117.718
R16006 dvss.n1074 dvss.n1073 117.718
R16007 dvss.n1064 dvss.n1063 117.718
R16008 dvss.n455 dvss.n454 117.718
R16009 dvss.n462 dvss.n461 117.718
R16010 dvss.n452 dvss.n451 117.718
R16011 dvss.n1686 dvss.n1550 117.718
R16012 dvss.n1676 dvss.n1549 117.718
R16013 dvss.n2304 dvss.n2168 117.718
R16014 dvss.n2294 dvss.n2167 117.718
R16015 dvss.n1073 dvss.n937 117.718
R16016 dvss.n1063 dvss.n936 117.718
R16017 dvss.n461 dvss.n325 117.718
R16018 dvss.n451 dvss.n324 117.718
R16019 dvss.n1679 dvss.n1678 117.718
R16020 dvss.n2297 dvss.n2296 117.718
R16021 dvss.n1066 dvss.n1065 117.718
R16022 dvss.n454 dvss.n453 117.718
R16023 dvss.n2721 dvss.t146 115.689
R16024 dvss.n2600 dvss.t116 114.244
R16025 dvss.n2757 dvss.t170 114.244
R16026 dvss.n1223 dvss.t5 114.244
R16027 dvss.n2523 dvss.t58 114.244
R16028 dvss.n2774 dvss.t154 114.244
R16029 dvss.n2870 dvss.t166 114.244
R16030 dvss.n2619 dvss.t179 113.738
R16031 dvss.n1762 dvss.t20 112.946
R16032 dvss.t19 dvss.n1422 112.946
R16033 dvss.n2380 dvss.t136 112.946
R16034 dvss.t135 dvss.n2040 112.946
R16035 dvss.n1149 dvss.t24 112.946
R16036 dvss.t114 dvss.n809 112.946
R16037 dvss.n537 dvss.t23 112.946
R16038 dvss.t137 dvss.n197 112.946
R16039 dvss.n1524 dvss.n1523 112.829
R16040 dvss.n1503 dvss.n1502 112.829
R16041 dvss.n2142 dvss.n2141 112.829
R16042 dvss.n2121 dvss.n2120 112.829
R16043 dvss.n911 dvss.n910 112.829
R16044 dvss.n890 dvss.n889 112.829
R16045 dvss.n299 dvss.n298 112.829
R16046 dvss.n278 dvss.n277 112.829
R16047 dvss.n1454 dvss.n1446 111.293
R16048 dvss.n2072 dvss.n2064 111.293
R16049 dvss.n841 dvss.n833 111.293
R16050 dvss.n229 dvss.n221 111.293
R16051 dvss.n1462 dvss.n1461 111.292
R16052 dvss.n2080 dvss.n2079 111.292
R16053 dvss.n849 dvss.n848 111.292
R16054 dvss.n237 dvss.n236 111.292
R16055 dvss.n1449 dvss.n1439 108.141
R16056 dvss.n2067 dvss.n2057 108.141
R16057 dvss.n836 dvss.n826 108.141
R16058 dvss.n224 dvss.n214 108.141
R16059 dvss.n1401 dvss.n1392 108.141
R16060 dvss.n1407 dvss.n1392 108.141
R16061 dvss.n1396 dvss.n1392 108.141
R16062 dvss.n1414 dvss.n1392 108.141
R16063 dvss.n2019 dvss.n2010 108.141
R16064 dvss.n2025 dvss.n2010 108.141
R16065 dvss.n2014 dvss.n2010 108.141
R16066 dvss.n2032 dvss.n2010 108.141
R16067 dvss.n788 dvss.n779 108.141
R16068 dvss.n794 dvss.n779 108.141
R16069 dvss.n783 dvss.n779 108.141
R16070 dvss.n801 dvss.n779 108.141
R16071 dvss.n176 dvss.n167 108.141
R16072 dvss.n182 dvss.n167 108.141
R16073 dvss.n171 dvss.n167 108.141
R16074 dvss.n189 dvss.n167 108.141
R16075 dvss.n2656 dvss.t28 108.037
R16076 dvss.n1631 dvss.n1558 105.765
R16077 dvss.n2249 dvss.n2176 105.765
R16078 dvss.n1018 dvss.n945 105.765
R16079 dvss.n406 dvss.n333 105.765
R16080 dvss.n1591 dvss.n1574 105.765
R16081 dvss.n1591 dvss.n1573 105.765
R16082 dvss.n1592 dvss.n1591 105.765
R16083 dvss.n1652 dvss.n1606 105.765
R16084 dvss.n1641 dvss.n1558 105.765
R16085 dvss.n1652 dvss.n1605 105.765
R16086 dvss.n1628 dvss.n1558 105.765
R16087 dvss.n1652 dvss.n1563 105.765
R16088 dvss.n1816 dvss.n1802 105.765
R16089 dvss.n1816 dvss.n1801 105.765
R16090 dvss.n1816 dvss.n1800 105.765
R16091 dvss.n2209 dvss.n2192 105.765
R16092 dvss.n2209 dvss.n2191 105.765
R16093 dvss.n2210 dvss.n2209 105.765
R16094 dvss.n2270 dvss.n2224 105.765
R16095 dvss.n2259 dvss.n2176 105.765
R16096 dvss.n2270 dvss.n2223 105.765
R16097 dvss.n2246 dvss.n2176 105.765
R16098 dvss.n2270 dvss.n2181 105.765
R16099 dvss.n2434 dvss.n2420 105.765
R16100 dvss.n2434 dvss.n2419 105.765
R16101 dvss.n2434 dvss.n2418 105.765
R16102 dvss.n978 dvss.n961 105.765
R16103 dvss.n978 dvss.n960 105.765
R16104 dvss.n979 dvss.n978 105.765
R16105 dvss.n1039 dvss.n993 105.765
R16106 dvss.n1028 dvss.n945 105.765
R16107 dvss.n1039 dvss.n992 105.765
R16108 dvss.n1015 dvss.n945 105.765
R16109 dvss.n1039 dvss.n950 105.765
R16110 dvss.n1203 dvss.n1189 105.765
R16111 dvss.n1203 dvss.n1188 105.765
R16112 dvss.n1203 dvss.n1187 105.765
R16113 dvss.n366 dvss.n349 105.765
R16114 dvss.n366 dvss.n348 105.765
R16115 dvss.n367 dvss.n366 105.765
R16116 dvss.n427 dvss.n381 105.765
R16117 dvss.n416 dvss.n333 105.765
R16118 dvss.n427 dvss.n380 105.765
R16119 dvss.n403 dvss.n333 105.765
R16120 dvss.n427 dvss.n338 105.765
R16121 dvss.n591 dvss.n577 105.765
R16122 dvss.n591 dvss.n576 105.765
R16123 dvss.n591 dvss.n575 105.765
R16124 dvss.n1519 dvss.n1518 104.172
R16125 dvss.n1498 dvss.n1497 104.172
R16126 dvss.n2137 dvss.n2136 104.172
R16127 dvss.n2116 dvss.n2115 104.172
R16128 dvss.n906 dvss.n905 104.172
R16129 dvss.n885 dvss.n884 104.172
R16130 dvss.n294 dvss.n293 104.172
R16131 dvss.n273 dvss.n272 104.172
R16132 dvss.n4 dvss.t118 101.037
R16133 dvss.n2772 dvss.t40 101.037
R16134 dvss.n1231 dvss.t7 101.037
R16135 dvss.n1846 dvss.t56 101.037
R16136 dvss.n2785 dvss.t26 101.037
R16137 dvss.n617 dvss.t168 101.037
R16138 dvss.n1706 dvss.n1705 93.979
R16139 dvss.n1540 dvss.n1537 93.979
R16140 dvss.n1698 dvss.n1536 93.979
R16141 dvss.n1695 dvss.n1535 93.979
R16142 dvss.n1546 dvss.n1534 93.979
R16143 dvss.n1695 dvss.n1534 93.979
R16144 dvss.n1698 dvss.n1535 93.979
R16145 dvss.n1540 dvss.n1536 93.979
R16146 dvss.n1705 dvss.n1537 93.979
R16147 dvss.n1706 dvss.n1530 93.979
R16148 dvss.n1733 dvss.n1732 93.979
R16149 dvss.n1729 dvss.n1480 93.979
R16150 dvss.n1727 dvss.n1479 93.979
R16151 dvss.n1725 dvss.n1478 93.979
R16152 dvss.n1723 dvss.n1477 93.979
R16153 dvss.n1732 dvss.n1480 93.979
R16154 dvss.n1729 dvss.n1479 93.979
R16155 dvss.n1727 dvss.n1478 93.979
R16156 dvss.n1725 dvss.n1477 93.979
R16157 dvss.n1733 dvss.n1474 93.979
R16158 dvss.n2324 dvss.n2323 93.979
R16159 dvss.n2158 dvss.n2155 93.979
R16160 dvss.n2316 dvss.n2154 93.979
R16161 dvss.n2313 dvss.n2153 93.979
R16162 dvss.n2164 dvss.n2152 93.979
R16163 dvss.n2313 dvss.n2152 93.979
R16164 dvss.n2316 dvss.n2153 93.979
R16165 dvss.n2158 dvss.n2154 93.979
R16166 dvss.n2323 dvss.n2155 93.979
R16167 dvss.n2324 dvss.n2148 93.979
R16168 dvss.n2351 dvss.n2350 93.979
R16169 dvss.n2347 dvss.n2098 93.979
R16170 dvss.n2345 dvss.n2097 93.979
R16171 dvss.n2343 dvss.n2096 93.979
R16172 dvss.n2341 dvss.n2095 93.979
R16173 dvss.n2350 dvss.n2098 93.979
R16174 dvss.n2347 dvss.n2097 93.979
R16175 dvss.n2345 dvss.n2096 93.979
R16176 dvss.n2343 dvss.n2095 93.979
R16177 dvss.n2351 dvss.n2092 93.979
R16178 dvss.n1093 dvss.n1092 93.979
R16179 dvss.n927 dvss.n924 93.979
R16180 dvss.n1085 dvss.n923 93.979
R16181 dvss.n1082 dvss.n922 93.979
R16182 dvss.n933 dvss.n921 93.979
R16183 dvss.n1082 dvss.n921 93.979
R16184 dvss.n1085 dvss.n922 93.979
R16185 dvss.n927 dvss.n923 93.979
R16186 dvss.n1092 dvss.n924 93.979
R16187 dvss.n1093 dvss.n917 93.979
R16188 dvss.n1120 dvss.n1119 93.979
R16189 dvss.n1116 dvss.n867 93.979
R16190 dvss.n1114 dvss.n866 93.979
R16191 dvss.n1112 dvss.n865 93.979
R16192 dvss.n1110 dvss.n864 93.979
R16193 dvss.n1119 dvss.n867 93.979
R16194 dvss.n1116 dvss.n866 93.979
R16195 dvss.n1114 dvss.n865 93.979
R16196 dvss.n1112 dvss.n864 93.979
R16197 dvss.n1120 dvss.n861 93.979
R16198 dvss.n481 dvss.n480 93.979
R16199 dvss.n315 dvss.n312 93.979
R16200 dvss.n473 dvss.n311 93.979
R16201 dvss.n470 dvss.n310 93.979
R16202 dvss.n321 dvss.n309 93.979
R16203 dvss.n470 dvss.n309 93.979
R16204 dvss.n473 dvss.n310 93.979
R16205 dvss.n315 dvss.n311 93.979
R16206 dvss.n480 dvss.n312 93.979
R16207 dvss.n481 dvss.n305 93.979
R16208 dvss.n508 dvss.n507 93.979
R16209 dvss.n504 dvss.n255 93.979
R16210 dvss.n502 dvss.n254 93.979
R16211 dvss.n500 dvss.n253 93.979
R16212 dvss.n498 dvss.n252 93.979
R16213 dvss.n507 dvss.n255 93.979
R16214 dvss.n504 dvss.n254 93.979
R16215 dvss.n502 dvss.n253 93.979
R16216 dvss.n500 dvss.n252 93.979
R16217 dvss.n508 dvss.n249 93.979
R16218 dvss.n1518 dvss.n1517 92.5
R16219 dvss.n1497 dvss.n1496 92.5
R16220 dvss.n2136 dvss.n2135 92.5
R16221 dvss.n2115 dvss.n2114 92.5
R16222 dvss.n905 dvss.n904 92.5
R16223 dvss.n884 dvss.n883 92.5
R16224 dvss.n293 dvss.n292 92.5
R16225 dvss.n272 dvss.n271 92.5
R16226 dvss.n1349 dvss.t103 92.436
R16227 dvss.n1967 dvss.t85 92.436
R16228 dvss.n736 dvss.t190 92.436
R16229 dvss.n124 dvss.t63 92.436
R16230 dvss.n2606 dvss.t115 91.94
R16231 dvss.n2758 dvss.t169 91.94
R16232 dvss.n2590 dvss.t4 91.94
R16233 dvss.n2519 dvss.t57 91.94
R16234 dvss.n2791 dvss.t153 91.94
R16235 dvss.n2866 dvss.t165 91.94
R16236 dvss.n2620 dvss.t175 91.196
R16237 dvss.n2619 dvss.t181 91.196
R16238 dvss.n1258 dvss.t50 90.702
R16239 dvss.n1873 dvss.t74 90.702
R16240 dvss.n642 dvss.t9 90.702
R16241 dvss.n29 dvss.t126 90.702
R16242 dvss.n1367 dvss.t98 90.701
R16243 dvss.n1985 dvss.t88 90.701
R16244 dvss.n754 dvss.t187 90.701
R16245 dvss.n142 dvss.t70 90.701
R16246 dvss.n1456 dvss.n1455 87.638
R16247 dvss.n1458 dvss.n1457 87.638
R16248 dvss.n1461 dvss.n1444 87.638
R16249 dvss.n1455 dvss.n1454 87.638
R16250 dvss.n1457 dvss.n1456 87.638
R16251 dvss.n1458 dvss.n1444 87.638
R16252 dvss.n2074 dvss.n2073 87.638
R16253 dvss.n2076 dvss.n2075 87.638
R16254 dvss.n2079 dvss.n2062 87.638
R16255 dvss.n2073 dvss.n2072 87.638
R16256 dvss.n2075 dvss.n2074 87.638
R16257 dvss.n2076 dvss.n2062 87.638
R16258 dvss.n843 dvss.n842 87.638
R16259 dvss.n845 dvss.n844 87.638
R16260 dvss.n848 dvss.n831 87.638
R16261 dvss.n842 dvss.n841 87.638
R16262 dvss.n844 dvss.n843 87.638
R16263 dvss.n845 dvss.n831 87.638
R16264 dvss.n231 dvss.n230 87.638
R16265 dvss.n233 dvss.n232 87.638
R16266 dvss.n236 dvss.n219 87.638
R16267 dvss.n230 dvss.n229 87.638
R16268 dvss.n232 dvss.n231 87.638
R16269 dvss.n233 dvss.n219 87.638
R16270 dvss.n1676 dvss.n1544 87.392
R16271 dvss.n2294 dvss.n2162 87.392
R16272 dvss.n1063 dvss.n931 87.392
R16273 dvss.n451 dvss.n319 87.392
R16274 dvss.n1631 dvss.n1560 80.972
R16275 dvss.n2249 dvss.n2178 80.972
R16276 dvss.n1018 dvss.n947 80.972
R16277 dvss.n406 dvss.n335 80.972
R16278 dvss.n1632 dvss.n1631 80.972
R16279 dvss.n2250 dvss.n2249 80.972
R16280 dvss.n1019 dvss.n1018 80.972
R16281 dvss.n407 dvss.n406 80.972
R16282 dvss.n1581 dvss.n1574 80.971
R16283 dvss.n1577 dvss.n1573 80.971
R16284 dvss.n1593 dvss.n1592 80.971
R16285 dvss.n1621 dvss.n1606 80.971
R16286 dvss.n1627 dvss.n1605 80.971
R16287 dvss.n1655 dvss.n1563 80.971
R16288 dvss.n1584 dvss.n1574 80.971
R16289 dvss.n1580 dvss.n1573 80.971
R16290 dvss.n1592 dvss.n1572 80.971
R16291 dvss.n1641 dvss.n1640 80.971
R16292 dvss.n1633 dvss.n1628 80.971
R16293 dvss.n1617 dvss.n1606 80.971
R16294 dvss.n1642 dvss.n1641 80.971
R16295 dvss.n1622 dvss.n1605 80.971
R16296 dvss.n1628 dvss.n1619 80.971
R16297 dvss.n1629 dvss.n1563 80.971
R16298 dvss.n1810 dvss.n1802 80.971
R16299 dvss.n1806 dvss.n1801 80.971
R16300 dvss.n1800 dvss.n1799 80.971
R16301 dvss.n1803 dvss.n1802 80.971
R16302 dvss.n1809 dvss.n1801 80.971
R16303 dvss.n1805 dvss.n1800 80.971
R16304 dvss.n2199 dvss.n2192 80.971
R16305 dvss.n2195 dvss.n2191 80.971
R16306 dvss.n2211 dvss.n2210 80.971
R16307 dvss.n2239 dvss.n2224 80.971
R16308 dvss.n2245 dvss.n2223 80.971
R16309 dvss.n2273 dvss.n2181 80.971
R16310 dvss.n2202 dvss.n2192 80.971
R16311 dvss.n2198 dvss.n2191 80.971
R16312 dvss.n2210 dvss.n2190 80.971
R16313 dvss.n2259 dvss.n2258 80.971
R16314 dvss.n2251 dvss.n2246 80.971
R16315 dvss.n2235 dvss.n2224 80.971
R16316 dvss.n2260 dvss.n2259 80.971
R16317 dvss.n2240 dvss.n2223 80.971
R16318 dvss.n2246 dvss.n2237 80.971
R16319 dvss.n2247 dvss.n2181 80.971
R16320 dvss.n2428 dvss.n2420 80.971
R16321 dvss.n2424 dvss.n2419 80.971
R16322 dvss.n2418 dvss.n2417 80.971
R16323 dvss.n2421 dvss.n2420 80.971
R16324 dvss.n2427 dvss.n2419 80.971
R16325 dvss.n2423 dvss.n2418 80.971
R16326 dvss.n968 dvss.n961 80.971
R16327 dvss.n964 dvss.n960 80.971
R16328 dvss.n980 dvss.n979 80.971
R16329 dvss.n1008 dvss.n993 80.971
R16330 dvss.n1014 dvss.n992 80.971
R16331 dvss.n1042 dvss.n950 80.971
R16332 dvss.n971 dvss.n961 80.971
R16333 dvss.n967 dvss.n960 80.971
R16334 dvss.n979 dvss.n959 80.971
R16335 dvss.n1028 dvss.n1027 80.971
R16336 dvss.n1020 dvss.n1015 80.971
R16337 dvss.n1004 dvss.n993 80.971
R16338 dvss.n1029 dvss.n1028 80.971
R16339 dvss.n1009 dvss.n992 80.971
R16340 dvss.n1015 dvss.n1006 80.971
R16341 dvss.n1016 dvss.n950 80.971
R16342 dvss.n1197 dvss.n1189 80.971
R16343 dvss.n1193 dvss.n1188 80.971
R16344 dvss.n1187 dvss.n1186 80.971
R16345 dvss.n1190 dvss.n1189 80.971
R16346 dvss.n1196 dvss.n1188 80.971
R16347 dvss.n1192 dvss.n1187 80.971
R16348 dvss.n356 dvss.n349 80.971
R16349 dvss.n352 dvss.n348 80.971
R16350 dvss.n368 dvss.n367 80.971
R16351 dvss.n396 dvss.n381 80.971
R16352 dvss.n402 dvss.n380 80.971
R16353 dvss.n430 dvss.n338 80.971
R16354 dvss.n359 dvss.n349 80.971
R16355 dvss.n355 dvss.n348 80.971
R16356 dvss.n367 dvss.n347 80.971
R16357 dvss.n416 dvss.n415 80.971
R16358 dvss.n408 dvss.n403 80.971
R16359 dvss.n392 dvss.n381 80.971
R16360 dvss.n417 dvss.n416 80.971
R16361 dvss.n397 dvss.n380 80.971
R16362 dvss.n403 dvss.n394 80.971
R16363 dvss.n404 dvss.n338 80.971
R16364 dvss.n585 dvss.n577 80.971
R16365 dvss.n581 dvss.n576 80.971
R16366 dvss.n575 dvss.n574 80.971
R16367 dvss.n578 dvss.n577 80.971
R16368 dvss.n584 dvss.n576 80.971
R16369 dvss.n580 dvss.n575 80.971
R16370 dvss.n1258 dvss.n1257 76.723
R16371 dvss.n1257 dvss.n1244 76.723
R16372 dvss.n1366 dvss.n1287 76.723
R16373 dvss.n1367 dvss.n1366 76.723
R16374 dvss.n2502 dvss.n1856 76.723
R16375 dvss.n1873 dvss.n1856 76.723
R16376 dvss.n1984 dvss.n1905 76.723
R16377 dvss.n1985 dvss.n1984 76.723
R16378 dvss.n642 dvss.n641 76.723
R16379 dvss.n641 dvss.n629 76.723
R16380 dvss.n753 dvss.n674 76.723
R16381 dvss.n754 dvss.n753 76.723
R16382 dvss.n141 dvss.n62 76.723
R16383 dvss.n142 dvss.n141 76.723
R16384 dvss.n29 dvss.n28 76.723
R16385 dvss.n28 dvss.n16 76.723
R16386 dvss.n1450 dvss.n1449 76.22
R16387 dvss.n2068 dvss.n2067 76.22
R16388 dvss.n837 dvss.n836 76.22
R16389 dvss.n225 dvss.n224 76.22
R16390 dvss.n1449 dvss.n1448 76.22
R16391 dvss.n2067 dvss.n2066 76.22
R16392 dvss.n836 dvss.n835 76.22
R16393 dvss.n224 dvss.n223 76.22
R16394 dvss.n1401 dvss.n1398 76.219
R16395 dvss.n1408 dvss.n1407 76.219
R16396 dvss.n1412 dvss.n1396 76.219
R16397 dvss.n1415 dvss.n1414 76.219
R16398 dvss.n1402 dvss.n1401 76.219
R16399 dvss.n1407 dvss.n1406 76.219
R16400 dvss.n1409 dvss.n1396 76.219
R16401 dvss.n1414 dvss.n1413 76.219
R16402 dvss.n2019 dvss.n2016 76.219
R16403 dvss.n2026 dvss.n2025 76.219
R16404 dvss.n2030 dvss.n2014 76.219
R16405 dvss.n2033 dvss.n2032 76.219
R16406 dvss.n2020 dvss.n2019 76.219
R16407 dvss.n2025 dvss.n2024 76.219
R16408 dvss.n2027 dvss.n2014 76.219
R16409 dvss.n2032 dvss.n2031 76.219
R16410 dvss.n788 dvss.n785 76.219
R16411 dvss.n795 dvss.n794 76.219
R16412 dvss.n799 dvss.n783 76.219
R16413 dvss.n802 dvss.n801 76.219
R16414 dvss.n789 dvss.n788 76.219
R16415 dvss.n794 dvss.n793 76.219
R16416 dvss.n796 dvss.n783 76.219
R16417 dvss.n801 dvss.n800 76.219
R16418 dvss.n176 dvss.n173 76.219
R16419 dvss.n183 dvss.n182 76.219
R16420 dvss.n187 dvss.n171 76.219
R16421 dvss.n190 dvss.n189 76.219
R16422 dvss.n177 dvss.n176 76.219
R16423 dvss.n182 dvss.n181 76.219
R16424 dvss.n184 dvss.n171 76.219
R16425 dvss.n189 dvss.n188 76.219
R16426 dvss.n2649 dvss.t27 71.739
R16427 dvss.n2546 dvss.n2544 69.321
R16428 dvss.n2477 dvss.n2475 69.321
R16429 dvss.n2823 dvss.n2821 69.321
R16430 dvss.n39 dvss.n38 69.321
R16431 dvss.n1518 dvss.t111 66.827
R16432 dvss.n1497 dvss.t52 66.827
R16433 dvss.n2136 dvss.t124 66.827
R16434 dvss.n2115 dvss.t1 66.827
R16435 dvss.n905 dvss.t162 66.827
R16436 dvss.n884 dvss.t36 66.827
R16437 dvss.n293 dvss.t22 66.827
R16438 dvss.n272 dvss.t142 66.827
R16439 dvss.t41 dvss.n2564 64.705
R16440 dvss.t71 dvss.n2494 64.705
R16441 dvss.t10 dvss.n2840 64.705
R16442 dvss.t133 dvss.n2913 64.705
R16443 dvss.n1709 dvss.n1708 59.469
R16444 dvss.n2327 dvss.n2326 59.469
R16445 dvss.n1096 dvss.n1095 59.469
R16446 dvss.n484 dvss.n483 59.469
R16447 dvss.n1590 dvss.n1589 59.468
R16448 dvss.n1585 dvss.n1575 59.468
R16449 dvss.n1651 dvss.n1650 59.468
R16450 dvss.n1612 dvss.n1607 59.468
R16451 dvss.n1614 dvss.n1557 59.468
R16452 dvss.n1643 dvss.n1616 59.468
R16453 dvss.n1689 dvss.n1533 59.468
R16454 dvss.n1736 dvss.n1735 59.468
R16455 dvss.n1721 dvss.n1476 59.468
R16456 dvss.n1818 dvss.n1817 59.468
R16457 dvss.n1815 dvss.n1814 59.468
R16458 dvss.n2208 dvss.n2207 59.468
R16459 dvss.n2203 dvss.n2193 59.468
R16460 dvss.n2269 dvss.n2268 59.468
R16461 dvss.n2230 dvss.n2225 59.468
R16462 dvss.n2232 dvss.n2175 59.468
R16463 dvss.n2261 dvss.n2234 59.468
R16464 dvss.n2307 dvss.n2151 59.468
R16465 dvss.n2354 dvss.n2353 59.468
R16466 dvss.n2339 dvss.n2094 59.468
R16467 dvss.n2436 dvss.n2435 59.468
R16468 dvss.n2433 dvss.n2432 59.468
R16469 dvss.n977 dvss.n976 59.468
R16470 dvss.n972 dvss.n962 59.468
R16471 dvss.n1038 dvss.n1037 59.468
R16472 dvss.n999 dvss.n994 59.468
R16473 dvss.n1001 dvss.n944 59.468
R16474 dvss.n1030 dvss.n1003 59.468
R16475 dvss.n1076 dvss.n920 59.468
R16476 dvss.n1123 dvss.n1122 59.468
R16477 dvss.n1108 dvss.n863 59.468
R16478 dvss.n1205 dvss.n1204 59.468
R16479 dvss.n1202 dvss.n1201 59.468
R16480 dvss.n365 dvss.n364 59.468
R16481 dvss.n360 dvss.n350 59.468
R16482 dvss.n426 dvss.n425 59.468
R16483 dvss.n387 dvss.n382 59.468
R16484 dvss.n389 dvss.n332 59.468
R16485 dvss.n418 dvss.n391 59.468
R16486 dvss.n464 dvss.n308 59.468
R16487 dvss.n511 dvss.n510 59.468
R16488 dvss.n496 dvss.n251 59.468
R16489 dvss.n593 dvss.n592 59.468
R16490 dvss.n590 dvss.n589 59.468
R16491 dvss.n2727 dvss.n2726 59.351
R16492 dvss.n2672 dvss.n2671 59.351
R16493 dvss.n1451 dvss.n1446 55.647
R16494 dvss.n2069 dvss.n2064 55.647
R16495 dvss.n838 dvss.n833 55.647
R16496 dvss.n226 dvss.n221 55.647
R16497 dvss.n1463 dvss.n1462 55.647
R16498 dvss.n2081 dvss.n2080 55.647
R16499 dvss.n850 dvss.n849 55.647
R16500 dvss.n238 dvss.n237 55.647
R16501 dvss.n1320 dvss.n1319 52.306
R16502 dvss.n1938 dvss.n1937 52.306
R16503 dvss.n707 dvss.n706 52.306
R16504 dvss.n95 dvss.n94 52.306
R16505 dvss.n2576 dvss.t47 46.218
R16506 dvss.t79 dvss.n1850 46.218
R16507 dvss.n2852 dvss.t16 46.218
R16508 dvss.n2925 dvss.t131 46.218
R16509 dvss.n1595 dvss.n1594 45.577
R16510 dvss.n1588 dvss.n1567 45.577
R16511 dvss.n2213 dvss.n2212 45.577
R16512 dvss.n2206 dvss.n2185 45.577
R16513 dvss.n982 dvss.n981 45.577
R16514 dvss.n975 dvss.n954 45.577
R16515 dvss.n370 dvss.n369 45.577
R16516 dvss.n363 dvss.n342 45.577
R16517 dvss.n2721 dvss.n2720 43.883
R16518 dvss.n1682 dvss.n1681 42.409
R16519 dvss.n2300 dvss.n2299 42.409
R16520 dvss.n1069 dvss.n1068 42.409
R16521 dvss.n457 dvss.n456 42.409
R16522 dvss.n1711 dvss.n1527 36.76
R16523 dvss.n2329 dvss.n2145 36.76
R16524 dvss.n1098 dvss.n914 36.76
R16525 dvss.n486 dvss.n302 36.76
R16526 dvss.n2707 dvss.n2702 36.141
R16527 dvss.n2707 dvss.n2700 36.141
R16528 dvss.n2711 dvss.n2700 36.141
R16529 dvss.n2711 dvss.n2696 36.141
R16530 dvss.n2717 dvss.n2696 36.141
R16531 dvss.n2717 dvss.n2693 36.141
R16532 dvss.n2744 dvss.n2693 36.141
R16533 dvss.n2744 dvss.n2694 36.141
R16534 dvss.n2740 dvss.n2694 36.141
R16535 dvss.n2740 dvss.n2739 36.141
R16536 dvss.n2739 dvss.n2724 36.141
R16537 dvss.n2734 dvss.n2724 36.141
R16538 dvss.n2734 dvss.n2731 36.141
R16539 dvss.n2731 dvss.n2685 36.141
R16540 dvss.n2749 dvss.n2685 36.141
R16541 dvss.n2641 dvss.n2636 36.141
R16542 dvss.n2641 dvss.n2634 36.141
R16543 dvss.n2645 dvss.n2634 36.141
R16544 dvss.n2645 dvss.n2628 36.141
R16545 dvss.n2653 dvss.n2628 36.141
R16546 dvss.n2653 dvss.n2629 36.141
R16547 dvss.n2629 dvss.n2625 36.141
R16548 dvss.n2661 dvss.n2625 36.141
R16549 dvss.n2661 dvss.n2622 36.141
R16550 dvss.n2668 dvss.n2622 36.141
R16551 dvss.n2668 dvss.n2617 36.141
R16552 dvss.n2677 dvss.n2617 36.141
R16553 dvss.n2677 dvss.n2618 36.141
R16554 dvss.n2618 dvss.n2612 36.141
R16555 dvss.n2682 dvss.n2612 36.141
R16556 dvss.n2592 dvss.n1225 36.141
R16557 dvss.n2592 dvss.n1226 36.141
R16558 dvss.n2586 dvss.n1226 36.141
R16559 dvss.n2586 dvss.n1229 36.141
R16560 dvss.n2581 dvss.n2580 36.141
R16561 dvss.n2580 dvss.n1234 36.141
R16562 dvss.n1238 dvss.n1234 36.141
R16563 dvss.n2573 dvss.n1238 36.141
R16564 dvss.n2573 dvss.n1239 36.141
R16565 dvss.n2568 dvss.n1239 36.141
R16566 dvss.n2568 dvss.n1246 36.141
R16567 dvss.n2562 dvss.n1246 36.141
R16568 dvss.n2562 dvss.n1251 36.141
R16569 dvss.n1254 dvss.n1251 36.141
R16570 dvss.n2556 dvss.n1254 36.141
R16571 dvss.n2556 dvss.n1260 36.141
R16572 dvss.n2550 dvss.n1260 36.141
R16573 dvss.n2550 dvss.n1265 36.141
R16574 dvss.n2541 dvss.n1265 36.141
R16575 dvss.n2541 dvss.n1268 36.141
R16576 dvss.n2535 dvss.n1268 36.141
R16577 dvss.n2535 dvss.n1273 36.141
R16578 dvss.n2531 dvss.n1273 36.141
R16579 dvss.n1316 dvss.n1311 36.141
R16580 dvss.n1311 dvss.n1308 36.141
R16581 dvss.n1324 dvss.n1308 36.141
R16582 dvss.n1324 dvss.n1304 36.141
R16583 dvss.n1330 dvss.n1304 36.141
R16584 dvss.n1330 dvss.n1302 36.141
R16585 dvss.n1334 dvss.n1302 36.141
R16586 dvss.n1334 dvss.n1298 36.141
R16587 dvss.n1341 dvss.n1298 36.141
R16588 dvss.n1341 dvss.n1296 36.141
R16589 dvss.n1347 dvss.n1296 36.141
R16590 dvss.n1347 dvss.n1291 36.141
R16591 dvss.n1362 dvss.n1291 36.141
R16592 dvss.n1362 dvss.n1292 36.141
R16593 dvss.n1356 dvss.n1292 36.141
R16594 dvss.n1356 dvss.n1353 36.141
R16595 dvss.n1353 dvss.n1283 36.141
R16596 dvss.n1375 dvss.n1283 36.141
R16597 dvss.n2521 dvss.n1839 36.141
R16598 dvss.n2521 dvss.n1841 36.141
R16599 dvss.n2515 dvss.n1841 36.141
R16600 dvss.n2515 dvss.n1844 36.141
R16601 dvss.n2510 dvss.n1848 36.141
R16602 dvss.n2506 dvss.n1848 36.141
R16603 dvss.n2506 dvss.n1852 36.141
R16604 dvss.n1858 dvss.n1852 36.141
R16605 dvss.n2499 dvss.n1858 36.141
R16606 dvss.n2499 dvss.n2498 36.141
R16607 dvss.n2498 dvss.n1860 36.141
R16608 dvss.n2492 dvss.n1860 36.141
R16609 dvss.n2492 dvss.n1867 36.141
R16610 dvss.n2488 dvss.n1867 36.141
R16611 dvss.n2488 dvss.n1875 36.141
R16612 dvss.n2482 dvss.n1875 36.141
R16613 dvss.n2482 dvss.n1879 36.141
R16614 dvss.n1883 dvss.n1879 36.141
R16615 dvss.n2472 dvss.n1883 36.141
R16616 dvss.n2472 dvss.n2471 36.141
R16617 dvss.n2471 dvss.n1885 36.141
R16618 dvss.n2465 dvss.n1885 36.141
R16619 dvss.n2465 dvss.n1892 36.141
R16620 dvss.n1934 dvss.n1929 36.141
R16621 dvss.n1929 dvss.n1926 36.141
R16622 dvss.n1942 dvss.n1926 36.141
R16623 dvss.n1942 dvss.n1922 36.141
R16624 dvss.n1948 dvss.n1922 36.141
R16625 dvss.n1948 dvss.n1920 36.141
R16626 dvss.n1952 dvss.n1920 36.141
R16627 dvss.n1952 dvss.n1916 36.141
R16628 dvss.n1959 dvss.n1916 36.141
R16629 dvss.n1959 dvss.n1914 36.141
R16630 dvss.n1965 dvss.n1914 36.141
R16631 dvss.n1965 dvss.n1909 36.141
R16632 dvss.n1980 dvss.n1909 36.141
R16633 dvss.n1980 dvss.n1910 36.141
R16634 dvss.n1974 dvss.n1910 36.141
R16635 dvss.n1974 dvss.n1971 36.141
R16636 dvss.n1971 dvss.n1901 36.141
R16637 dvss.n1993 dvss.n1901 36.141
R16638 dvss.n2794 dvss.n2793 36.141
R16639 dvss.n2793 dvss.n2776 36.141
R16640 dvss.n2780 dvss.n2776 36.141
R16641 dvss.n2788 dvss.n2780 36.141
R16642 dvss.n2856 dvss.n618 36.141
R16643 dvss.n2856 dvss.n2855 36.141
R16644 dvss.n2855 dvss.n621 36.141
R16645 dvss.n2849 dvss.n621 36.141
R16646 dvss.n2849 dvss.n625 36.141
R16647 dvss.n2844 dvss.n625 36.141
R16648 dvss.n2844 dvss.n631 36.141
R16649 dvss.n2838 dvss.n631 36.141
R16650 dvss.n2838 dvss.n636 36.141
R16651 dvss.n2834 dvss.n636 36.141
R16652 dvss.n2834 dvss.n644 36.141
R16653 dvss.n2828 dvss.n644 36.141
R16654 dvss.n2828 dvss.n648 36.141
R16655 dvss.n652 dvss.n648 36.141
R16656 dvss.n2818 dvss.n652 36.141
R16657 dvss.n2818 dvss.n2817 36.141
R16658 dvss.n2817 dvss.n654 36.141
R16659 dvss.n2811 dvss.n654 36.141
R16660 dvss.n2811 dvss.n661 36.141
R16661 dvss.n703 dvss.n698 36.141
R16662 dvss.n698 dvss.n695 36.141
R16663 dvss.n711 dvss.n695 36.141
R16664 dvss.n711 dvss.n691 36.141
R16665 dvss.n717 dvss.n691 36.141
R16666 dvss.n717 dvss.n689 36.141
R16667 dvss.n721 dvss.n689 36.141
R16668 dvss.n721 dvss.n685 36.141
R16669 dvss.n728 dvss.n685 36.141
R16670 dvss.n728 dvss.n683 36.141
R16671 dvss.n734 dvss.n683 36.141
R16672 dvss.n734 dvss.n678 36.141
R16673 dvss.n749 dvss.n678 36.141
R16674 dvss.n749 dvss.n679 36.141
R16675 dvss.n743 dvss.n679 36.141
R16676 dvss.n743 dvss.n740 36.141
R16677 dvss.n740 dvss.n670 36.141
R16678 dvss.n762 dvss.n670 36.141
R16679 dvss.n2868 dvss.n610 36.141
R16680 dvss.n2868 dvss.n612 36.141
R16681 dvss.n2862 dvss.n612 36.141
R16682 dvss.n2862 dvss.n615 36.141
R16683 dvss.n91 dvss.n86 36.141
R16684 dvss.n86 dvss.n83 36.141
R16685 dvss.n99 dvss.n83 36.141
R16686 dvss.n99 dvss.n79 36.141
R16687 dvss.n105 dvss.n79 36.141
R16688 dvss.n105 dvss.n77 36.141
R16689 dvss.n109 dvss.n77 36.141
R16690 dvss.n109 dvss.n73 36.141
R16691 dvss.n116 dvss.n73 36.141
R16692 dvss.n116 dvss.n71 36.141
R16693 dvss.n122 dvss.n71 36.141
R16694 dvss.n122 dvss.n66 36.141
R16695 dvss.n137 dvss.n66 36.141
R16696 dvss.n137 dvss.n67 36.141
R16697 dvss.n131 dvss.n67 36.141
R16698 dvss.n131 dvss.n128 36.141
R16699 dvss.n128 dvss.n58 36.141
R16700 dvss.n150 dvss.n58 36.141
R16701 dvss.n2929 dvss.n5 36.141
R16702 dvss.n2929 dvss.n7 36.141
R16703 dvss.n11 dvss.n7 36.141
R16704 dvss.n2922 dvss.n11 36.141
R16705 dvss.n2922 dvss.n12 36.141
R16706 dvss.n2917 dvss.n12 36.141
R16707 dvss.n2917 dvss.n18 36.141
R16708 dvss.n2911 dvss.n18 36.141
R16709 dvss.n2911 dvss.n23 36.141
R16710 dvss.n2907 dvss.n23 36.141
R16711 dvss.n2907 dvss.n31 36.141
R16712 dvss.n2901 dvss.n31 36.141
R16713 dvss.n2901 dvss.n35 36.141
R16714 dvss.n2896 dvss.n35 36.141
R16715 dvss.n2896 dvss.n41 36.141
R16716 dvss.n2890 dvss.n41 36.141
R16717 dvss.n2890 dvss.n45 36.141
R16718 dvss.n2886 dvss.n45 36.141
R16719 dvss.n2886 dvss.n49 36.141
R16720 dvss.n2531 dvss.n1275 35.388
R16721 dvss.n1657 dvss.n1561 35.388
R16722 dvss.n1659 dvss.n1657 35.388
R16723 dvss.n1673 dvss.n1670 35.388
R16724 dvss.n1663 dvss.n1556 35.388
R16725 dvss.n1603 dvss.n1556 35.388
R16726 dvss.n2461 dvss.n1892 35.388
R16727 dvss.n2275 dvss.n2179 35.388
R16728 dvss.n2277 dvss.n2275 35.388
R16729 dvss.n2291 dvss.n2288 35.388
R16730 dvss.n2281 dvss.n2174 35.388
R16731 dvss.n2221 dvss.n2174 35.388
R16732 dvss.n2807 dvss.n661 35.388
R16733 dvss.n1044 dvss.n948 35.388
R16734 dvss.n1046 dvss.n1044 35.388
R16735 dvss.n1060 dvss.n1057 35.388
R16736 dvss.n1050 dvss.n943 35.388
R16737 dvss.n990 dvss.n943 35.388
R16738 dvss.n432 dvss.n336 35.388
R16739 dvss.n434 dvss.n432 35.388
R16740 dvss.n448 dvss.n445 35.388
R16741 dvss.n438 dvss.n331 35.388
R16742 dvss.n378 dvss.n331 35.388
R16743 dvss.n2874 dvss.n49 35.388
R16744 dvss.n2726 dvss.t120 35.068
R16745 dvss.n2671 dvss.t151 35.068
R16746 dvss.n1375 dvss.n1284 35.011
R16747 dvss.n1993 dvss.n1902 35.011
R16748 dvss.n762 dvss.n671 35.011
R16749 dvss.n150 dvss.n59 35.011
R16750 dvss.n1399 dvss.n1390 34.133
R16751 dvss.n1758 dvss.n1434 34.133
R16752 dvss.n2017 dvss.n2008 34.133
R16753 dvss.n2376 dvss.n2052 34.133
R16754 dvss.n786 dvss.n777 34.133
R16755 dvss.n1145 dvss.n821 34.133
R16756 dvss.n174 dvss.n165 34.133
R16757 dvss.n533 dvss.n209 34.133
R16758 dvss.n1256 dvss.n1255 33.519
R16759 dvss.n1244 dvss.n1243 33.519
R16760 dvss.n1287 dvss.n1286 33.519
R16761 dvss.n1365 dvss.n1289 33.519
R16762 dvss.n2502 dvss.n1855 33.519
R16763 dvss.n1871 dvss.n1869 33.519
R16764 dvss.n1905 dvss.n1904 33.519
R16765 dvss.n1983 dvss.n1907 33.519
R16766 dvss.n640 dvss.n639 33.519
R16767 dvss.n629 dvss.n628 33.519
R16768 dvss.n674 dvss.n673 33.519
R16769 dvss.n752 dvss.n676 33.519
R16770 dvss.n62 dvss.n61 33.519
R16771 dvss.n140 dvss.n64 33.519
R16772 dvss.n27 dvss.n26 33.519
R16773 dvss.n16 dvss.n15 33.519
R16774 dvss.n2798 dvss.n2797 32.375
R16775 dvss.n1379 dvss.n1279 30.87
R16776 dvss.n1997 dvss.n1897 30.87
R16777 dvss.n766 dvss.n666 30.87
R16778 dvss.n154 dvss.n54 30.87
R16779 dvss.n2620 dvss.n2619 30.57
R16780 dvss.n2527 dvss.n1277 30.494
R16781 dvss.n2457 dvss.n1895 30.494
R16782 dvss.n2803 dvss.n664 30.494
R16783 dvss.n2881 dvss.n52 30.494
R16784 dvss.n1683 dvss.n1673 29.741
R16785 dvss.n2301 dvss.n2291 29.741
R16786 dvss.n1070 dvss.n1060 29.741
R16787 dvss.n458 dvss.n448 29.741
R16788 dvss.n1519 dvss.n1508 29.482
R16789 dvss.n1498 dvss.n1487 29.482
R16790 dvss.n2137 dvss.n2126 29.482
R16791 dvss.n2116 dvss.n2105 29.482
R16792 dvss.n906 dvss.n895 29.482
R16793 dvss.n885 dvss.n874 29.482
R16794 dvss.n294 dvss.n283 29.482
R16795 dvss.n273 dvss.n262 29.482
R16796 dvss.n1738 dvss.n1737 29.197
R16797 dvss.n1820 dvss.n1819 29.197
R16798 dvss.n2356 dvss.n2355 29.197
R16799 dvss.n2438 dvss.n2437 29.197
R16800 dvss.n1125 dvss.n1124 29.197
R16801 dvss.n1207 dvss.n1206 29.197
R16802 dvss.n513 dvss.n512 29.197
R16803 dvss.n595 dvss.n594 29.197
R16804 dvss.n1319 dvss.t164 28.12
R16805 dvss.n1937 dvss.t158 28.12
R16806 dvss.n706 dvss.t108 28.12
R16807 dvss.n94 dvss.t139 28.12
R16808 dvss.n2753 dvss 26.526
R16809 dvss.n1597 dvss.n1595 25.6
R16810 dvss.n1597 dvss.n1596 25.6
R16811 dvss.n1596 dvss.n1561 25.6
R16812 dvss.n1659 dvss.n1658 25.6
R16813 dvss.n1658 dvss.n1553 25.6
R16814 dvss.n1670 dvss.n1553 25.6
R16815 dvss.n1683 dvss.n1682 25.6
R16816 dvss.n1664 dvss.n1663 25.6
R16817 dvss.n1665 dvss.n1664 25.6
R16818 dvss.n1665 dvss.n1527 25.6
R16819 dvss.n1601 dvss.n1567 25.6
R16820 dvss.n1602 dvss.n1601 25.6
R16821 dvss.n1603 dvss.n1602 25.6
R16822 dvss.n2215 dvss.n2213 25.6
R16823 dvss.n2215 dvss.n2214 25.6
R16824 dvss.n2214 dvss.n2179 25.6
R16825 dvss.n2277 dvss.n2276 25.6
R16826 dvss.n2276 dvss.n2171 25.6
R16827 dvss.n2288 dvss.n2171 25.6
R16828 dvss.n2301 dvss.n2300 25.6
R16829 dvss.n2282 dvss.n2281 25.6
R16830 dvss.n2283 dvss.n2282 25.6
R16831 dvss.n2283 dvss.n2145 25.6
R16832 dvss.n2219 dvss.n2185 25.6
R16833 dvss.n2220 dvss.n2219 25.6
R16834 dvss.n2221 dvss.n2220 25.6
R16835 dvss.n984 dvss.n982 25.6
R16836 dvss.n984 dvss.n983 25.6
R16837 dvss.n983 dvss.n948 25.6
R16838 dvss.n1046 dvss.n1045 25.6
R16839 dvss.n1045 dvss.n940 25.6
R16840 dvss.n1057 dvss.n940 25.6
R16841 dvss.n1070 dvss.n1069 25.6
R16842 dvss.n1051 dvss.n1050 25.6
R16843 dvss.n1052 dvss.n1051 25.6
R16844 dvss.n1052 dvss.n914 25.6
R16845 dvss.n988 dvss.n954 25.6
R16846 dvss.n989 dvss.n988 25.6
R16847 dvss.n990 dvss.n989 25.6
R16848 dvss.n372 dvss.n370 25.6
R16849 dvss.n372 dvss.n371 25.6
R16850 dvss.n371 dvss.n336 25.6
R16851 dvss.n434 dvss.n433 25.6
R16852 dvss.n433 dvss.n328 25.6
R16853 dvss.n445 dvss.n328 25.6
R16854 dvss.n458 dvss.n457 25.6
R16855 dvss.n439 dvss.n438 25.6
R16856 dvss.n440 dvss.n439 25.6
R16857 dvss.n440 dvss.n302 25.6
R16858 dvss.n376 dvss.n342 25.6
R16859 dvss.n377 dvss.n376 25.6
R16860 dvss.n378 dvss.n377 25.6
R16861 dvss.n1403 dvss.n1399 22.317
R16862 dvss.n1404 dvss.n1403 22.317
R16863 dvss.n1405 dvss.n1404 22.317
R16864 dvss.n1405 dvss.n1397 22.317
R16865 dvss.n1410 dvss.n1397 22.317
R16866 dvss.n1411 dvss.n1410 22.317
R16867 dvss.n1411 dvss.n1395 22.317
R16868 dvss.n1416 dvss.n1395 22.317
R16869 dvss.n1447 dvss.n1434 22.317
R16870 dvss.n1452 dvss.n1447 22.317
R16871 dvss.n1453 dvss.n1452 22.317
R16872 dvss.n1453 dvss.n1445 22.317
R16873 dvss.n1459 dvss.n1445 22.317
R16874 dvss.n1460 dvss.n1459 22.317
R16875 dvss.n1460 dvss.n1443 22.317
R16876 dvss.n1465 dvss.n1443 22.317
R16877 dvss.n2021 dvss.n2017 22.317
R16878 dvss.n2022 dvss.n2021 22.317
R16879 dvss.n2023 dvss.n2022 22.317
R16880 dvss.n2023 dvss.n2015 22.317
R16881 dvss.n2028 dvss.n2015 22.317
R16882 dvss.n2029 dvss.n2028 22.317
R16883 dvss.n2029 dvss.n2013 22.317
R16884 dvss.n2034 dvss.n2013 22.317
R16885 dvss.n2065 dvss.n2052 22.317
R16886 dvss.n2070 dvss.n2065 22.317
R16887 dvss.n2071 dvss.n2070 22.317
R16888 dvss.n2071 dvss.n2063 22.317
R16889 dvss.n2077 dvss.n2063 22.317
R16890 dvss.n2078 dvss.n2077 22.317
R16891 dvss.n2078 dvss.n2061 22.317
R16892 dvss.n2083 dvss.n2061 22.317
R16893 dvss.n790 dvss.n786 22.317
R16894 dvss.n791 dvss.n790 22.317
R16895 dvss.n792 dvss.n791 22.317
R16896 dvss.n792 dvss.n784 22.317
R16897 dvss.n797 dvss.n784 22.317
R16898 dvss.n798 dvss.n797 22.317
R16899 dvss.n798 dvss.n782 22.317
R16900 dvss.n803 dvss.n782 22.317
R16901 dvss.n834 dvss.n821 22.317
R16902 dvss.n839 dvss.n834 22.317
R16903 dvss.n840 dvss.n839 22.317
R16904 dvss.n840 dvss.n832 22.317
R16905 dvss.n846 dvss.n832 22.317
R16906 dvss.n847 dvss.n846 22.317
R16907 dvss.n847 dvss.n830 22.317
R16908 dvss.n852 dvss.n830 22.317
R16909 dvss.n178 dvss.n174 22.317
R16910 dvss.n179 dvss.n178 22.317
R16911 dvss.n180 dvss.n179 22.317
R16912 dvss.n180 dvss.n172 22.317
R16913 dvss.n185 dvss.n172 22.317
R16914 dvss.n186 dvss.n185 22.317
R16915 dvss.n186 dvss.n170 22.317
R16916 dvss.n191 dvss.n170 22.317
R16917 dvss.n222 dvss.n209 22.317
R16918 dvss.n227 dvss.n222 22.317
R16919 dvss.n228 dvss.n227 22.317
R16920 dvss.n228 dvss.n220 22.317
R16921 dvss.n234 dvss.n220 22.317
R16922 dvss.n235 dvss.n234 22.317
R16923 dvss.n235 dvss.n218 22.317
R16924 dvss.n240 dvss.n218 22.317
R16925 dvss.n2726 dvss.t152 22.237
R16926 dvss.n2671 dvss.t177 22.237
R16927 dvss.n2720 dvss.t148 21.28
R16928 dvss.n2720 dvss.t149 21.28
R16929 dvss.n1319 dvss.t33 21.28
R16930 dvss.n1937 dvss.t122 21.28
R16931 dvss.n706 dvss.t160 21.28
R16932 dvss.n94 dvss.t113 21.28
R16933 dvss.n1417 dvss.n1416 20.348
R16934 dvss.n1466 dvss.n1465 20.348
R16935 dvss.n2035 dvss.n2034 20.348
R16936 dvss.n2084 dvss.n2083 20.348
R16937 dvss.n804 dvss.n803 20.348
R16938 dvss.n853 dvss.n852 20.348
R16939 dvss.n192 dvss.n191 20.348
R16940 dvss.n241 dvss.n240 20.348
R16941 dvss.n2544 dvss.t96 20
R16942 dvss.n2544 dvss.t82 20
R16943 dvss.n2475 dvss.t92 20
R16944 dvss.n2475 dvss.t156 20
R16945 dvss.n2821 dvss.t195 20
R16946 dvss.n2821 dvss.t173 20
R16947 dvss.n38 dvss.t68 20
R16948 dvss.n38 dvss.t183 20
R16949 dvss.n2749 dvss.n2748 18.009
R16950 dvss.n2682 dvss.n2681 18.009
R16951 dvss.n2547 dvss.n2543 17.171
R16952 dvss.n2548 dvss.n2547 17.171
R16953 dvss.n2478 dvss.n2474 17.171
R16954 dvss.n2479 dvss.n2478 17.171
R16955 dvss.n2824 dvss.n2820 17.171
R16956 dvss.n2825 dvss.n2824 17.171
R16957 dvss.n46 dvss.n37 17.171
R16958 dvss.n2898 dvss.n37 17.171
R16959 dvss.n1779 dvss.n1390 17.021
R16960 dvss.n2397 dvss.n2008 17.021
R16961 dvss.n1166 dvss.n777 17.021
R16962 dvss.n554 dvss.n165 17.021
R16963 dvss.n1759 dvss.n1758 16.885
R16964 dvss.n2377 dvss.n2376 16.885
R16965 dvss.n1146 dvss.n1145 16.885
R16966 dvss.n534 dvss.n533 16.885
R16967 dvss.n1758 dvss.n1757 15.523
R16968 dvss.n2376 dvss.n2375 15.523
R16969 dvss.n1145 dvss.n1144 15.523
R16970 dvss.n533 dvss.n532 15.523
R16971 dvss.n1517 dvss.n1516 15.463
R16972 dvss.n1496 dvss.n1495 15.463
R16973 dvss.n2135 dvss.n2134 15.463
R16974 dvss.n2114 dvss.n2113 15.463
R16975 dvss.n904 dvss.n903 15.463
R16976 dvss.n883 dvss.n882 15.463
R16977 dvss.n292 dvss.n291 15.463
R16978 dvss.n271 dvss.n270 15.463
R16979 dvss.n1795 dvss.n1390 15.387
R16980 dvss.n2413 dvss.n2008 15.387
R16981 dvss.n1182 dvss.n777 15.387
R16982 dvss.n570 dvss.n165 15.387
R16983 dvss.n2781 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 15
R16984 dvss.n2621 dvss.n2620 14.454
R16985 dvss.n2722 dvss.n2721 14.428
R16986 dvss.n1522 dvss.n1509 13.552
R16987 dvss.n1517 dvss.n1513 13.552
R16988 dvss.n1501 dvss.n1488 13.552
R16989 dvss.n1496 dvss.n1492 13.552
R16990 dvss.n2140 dvss.n2127 13.552
R16991 dvss.n2135 dvss.n2131 13.552
R16992 dvss.n2119 dvss.n2106 13.552
R16993 dvss.n2114 dvss.n2110 13.552
R16994 dvss.n909 dvss.n896 13.552
R16995 dvss.n904 dvss.n900 13.552
R16996 dvss.n888 dvss.n875 13.552
R16997 dvss.n883 dvss.n879 13.552
R16998 dvss.n297 dvss.n284 13.552
R16999 dvss.n292 dvss.n288 13.552
R17000 dvss.n276 dvss.n263 13.552
R17001 dvss.n271 dvss.n267 13.552
R17002 dvss.n1317 dvss.n1310 12.897
R17003 dvss.n1935 dvss.n1928 12.897
R17004 dvss.n704 dvss.n697 12.897
R17005 dvss.n92 dvss.n85 12.897
R17006 dvss.n1829 dvss.n1381 11.008
R17007 dvss.n2447 dvss.n1999 11.008
R17008 dvss.n1216 dvss.n768 11.008
R17009 dvss.n604 dvss.n156 11.008
R17010 dvss.n1243 dvss.t48 10.64
R17011 dvss.n1243 dvss.t46 10.64
R17012 dvss.n1255 dvss.t44 10.64
R17013 dvss.n1255 dvss.t42 10.64
R17014 dvss.n1286 dvss.t106 10.64
R17015 dvss.n1286 dvss.t104 10.64
R17016 dvss.n1289 dvss.t100 10.64
R17017 dvss.n1289 dvss.t102 10.64
R17018 dvss.n1855 dvss.t80 10.64
R17019 dvss.n1855 dvss.t78 10.64
R17020 dvss.n1869 dvss.t76 10.64
R17021 dvss.n1869 dvss.t72 10.64
R17022 dvss.n1904 dvss.t94 10.64
R17023 dvss.n1904 dvss.t86 10.64
R17024 dvss.n1907 dvss.t90 10.64
R17025 dvss.n1907 dvss.t84 10.64
R17026 dvss.n628 dvss.t17 10.64
R17027 dvss.n628 dvss.t15 10.64
R17028 dvss.n639 dvss.t13 10.64
R17029 dvss.n639 dvss.t11 10.64
R17030 dvss.n673 dvss.t193 10.64
R17031 dvss.n673 dvss.t191 10.64
R17032 dvss.n676 dvss.t185 10.64
R17033 dvss.n676 dvss.t189 10.64
R17034 dvss.n61 dvss.t66 10.64
R17035 dvss.n61 dvss.t64 10.64
R17036 dvss.n64 dvss.t62 10.64
R17037 dvss.n64 dvss.t60 10.64
R17038 dvss.n15 dvss.t132 10.64
R17039 dvss.n15 dvss.t130 10.64
R17040 dvss.n26 dvss.t128 10.64
R17041 dvss.n26 dvss.t134 10.64
R17042 dvss.n1674 dvss.n1548 10.424
R17043 dvss.n2292 dvss.n2166 10.424
R17044 dvss.n1061 dvss.n935 10.424
R17045 dvss.n449 dvss.n323 10.424
R17046 dvss.n1720 dvss.n1719 9.4
R17047 dvss.n2338 dvss.n2337 9.4
R17048 dvss.n1107 dvss.n1106 9.4
R17049 dvss.n495 dvss.n494 9.4
R17050 dvss.n1372 dvss.n1371 9.3
R17051 dvss.n1373 dvss.n1284 9.3
R17052 dvss.n1507 dvss.n1506 9.3
R17053 dvss.n1514 dvss.n1510 9.3
R17054 dvss.n1515 dvss.n1513 9.3
R17055 dvss.n1520 dvss.n1512 9.3
R17056 dvss.n1520 dvss.n1519 9.3
R17057 dvss.n1511 dvss.n1509 9.3
R17058 dvss.n1525 dvss.n1524 9.3
R17059 dvss.n1486 dvss.n1485 9.3
R17060 dvss.n1493 dvss.n1489 9.3
R17061 dvss.n1494 dvss.n1492 9.3
R17062 dvss.n1499 dvss.n1491 9.3
R17063 dvss.n1499 dvss.n1498 9.3
R17064 dvss.n1490 dvss.n1488 9.3
R17065 dvss.n1504 dvss.n1503 9.3
R17066 dvss.n1482 dvss.n1468 9.3
R17067 dvss.n1743 dvss.n1469 9.3
R17068 dvss.n1744 dvss.n1467 9.3
R17069 dvss.n1746 dvss.n1745 9.3
R17070 dvss.n1747 dvss.n1442 9.3
R17071 dvss.n1753 dvss.n1752 9.3
R17072 dvss.n1751 dvss.n1750 9.3
R17073 dvss.n1765 dvss.n1429 9.3
R17074 dvss.n1767 dvss.n1766 9.3
R17075 dvss.n1768 dvss.n1428 9.3
R17076 dvss.n1769 dvss.n1420 9.3
R17077 dvss.n1783 dvss.n1419 9.3
R17078 dvss.n1785 dvss.n1784 9.3
R17079 dvss.n1791 dvss.n1790 9.3
R17080 dvss.n1789 dvss.n1418 9.3
R17081 dvss.n1788 dvss.n1787 9.3
R17082 dvss.n1786 dvss.n1384 9.3
R17083 dvss.n1825 dvss.n1383 9.3
R17084 dvss.n1827 dvss.n1826 9.3
R17085 dvss.n1990 dvss.n1989 9.3
R17086 dvss.n1991 dvss.n1902 9.3
R17087 dvss.n2125 dvss.n2124 9.3
R17088 dvss.n2132 dvss.n2128 9.3
R17089 dvss.n2133 dvss.n2131 9.3
R17090 dvss.n2138 dvss.n2130 9.3
R17091 dvss.n2138 dvss.n2137 9.3
R17092 dvss.n2129 dvss.n2127 9.3
R17093 dvss.n2143 dvss.n2142 9.3
R17094 dvss.n2104 dvss.n2103 9.3
R17095 dvss.n2111 dvss.n2107 9.3
R17096 dvss.n2112 dvss.n2110 9.3
R17097 dvss.n2117 dvss.n2109 9.3
R17098 dvss.n2117 dvss.n2116 9.3
R17099 dvss.n2108 dvss.n2106 9.3
R17100 dvss.n2122 dvss.n2121 9.3
R17101 dvss.n2100 dvss.n2086 9.3
R17102 dvss.n2361 dvss.n2087 9.3
R17103 dvss.n2362 dvss.n2085 9.3
R17104 dvss.n2364 dvss.n2363 9.3
R17105 dvss.n2365 dvss.n2060 9.3
R17106 dvss.n2371 dvss.n2370 9.3
R17107 dvss.n2369 dvss.n2368 9.3
R17108 dvss.n2383 dvss.n2047 9.3
R17109 dvss.n2385 dvss.n2384 9.3
R17110 dvss.n2386 dvss.n2046 9.3
R17111 dvss.n2387 dvss.n2038 9.3
R17112 dvss.n2401 dvss.n2037 9.3
R17113 dvss.n2403 dvss.n2402 9.3
R17114 dvss.n2409 dvss.n2408 9.3
R17115 dvss.n2407 dvss.n2036 9.3
R17116 dvss.n2406 dvss.n2405 9.3
R17117 dvss.n2404 dvss.n2002 9.3
R17118 dvss.n2443 dvss.n2001 9.3
R17119 dvss.n2445 dvss.n2444 9.3
R17120 dvss.n2462 dvss.n2461 9.3
R17121 dvss.n2460 dvss.n1894 9.3
R17122 dvss.n1275 dvss.n1274 9.3
R17123 dvss.n1836 dvss.n1835 9.3
R17124 dvss.n759 dvss.n758 9.3
R17125 dvss.n760 dvss.n671 9.3
R17126 dvss.n894 dvss.n893 9.3
R17127 dvss.n901 dvss.n897 9.3
R17128 dvss.n902 dvss.n900 9.3
R17129 dvss.n907 dvss.n899 9.3
R17130 dvss.n907 dvss.n906 9.3
R17131 dvss.n898 dvss.n896 9.3
R17132 dvss.n912 dvss.n911 9.3
R17133 dvss.n873 dvss.n872 9.3
R17134 dvss.n880 dvss.n876 9.3
R17135 dvss.n881 dvss.n879 9.3
R17136 dvss.n886 dvss.n878 9.3
R17137 dvss.n886 dvss.n885 9.3
R17138 dvss.n877 dvss.n875 9.3
R17139 dvss.n891 dvss.n890 9.3
R17140 dvss.n869 dvss.n855 9.3
R17141 dvss.n1130 dvss.n856 9.3
R17142 dvss.n1131 dvss.n854 9.3
R17143 dvss.n1133 dvss.n1132 9.3
R17144 dvss.n1134 dvss.n829 9.3
R17145 dvss.n1140 dvss.n1139 9.3
R17146 dvss.n1138 dvss.n1137 9.3
R17147 dvss.n1152 dvss.n816 9.3
R17148 dvss.n1154 dvss.n1153 9.3
R17149 dvss.n1155 dvss.n815 9.3
R17150 dvss.n1156 dvss.n807 9.3
R17151 dvss.n1170 dvss.n806 9.3
R17152 dvss.n1172 dvss.n1171 9.3
R17153 dvss.n1178 dvss.n1177 9.3
R17154 dvss.n1176 dvss.n805 9.3
R17155 dvss.n1175 dvss.n1174 9.3
R17156 dvss.n1173 dvss.n771 9.3
R17157 dvss.n1212 dvss.n770 9.3
R17158 dvss.n1214 dvss.n1213 9.3
R17159 dvss.n147 dvss.n146 9.3
R17160 dvss.n148 dvss.n59 9.3
R17161 dvss.n282 dvss.n281 9.3
R17162 dvss.n289 dvss.n285 9.3
R17163 dvss.n290 dvss.n288 9.3
R17164 dvss.n295 dvss.n287 9.3
R17165 dvss.n295 dvss.n294 9.3
R17166 dvss.n286 dvss.n284 9.3
R17167 dvss.n300 dvss.n299 9.3
R17168 dvss.n261 dvss.n260 9.3
R17169 dvss.n268 dvss.n264 9.3
R17170 dvss.n269 dvss.n267 9.3
R17171 dvss.n274 dvss.n266 9.3
R17172 dvss.n274 dvss.n273 9.3
R17173 dvss.n265 dvss.n263 9.3
R17174 dvss.n279 dvss.n278 9.3
R17175 dvss.n257 dvss.n243 9.3
R17176 dvss.n518 dvss.n244 9.3
R17177 dvss.n519 dvss.n242 9.3
R17178 dvss.n521 dvss.n520 9.3
R17179 dvss.n522 dvss.n217 9.3
R17180 dvss.n528 dvss.n527 9.3
R17181 dvss.n526 dvss.n525 9.3
R17182 dvss.n540 dvss.n204 9.3
R17183 dvss.n542 dvss.n541 9.3
R17184 dvss.n543 dvss.n203 9.3
R17185 dvss.n544 dvss.n195 9.3
R17186 dvss.n558 dvss.n194 9.3
R17187 dvss.n560 dvss.n559 9.3
R17188 dvss.n566 dvss.n565 9.3
R17189 dvss.n564 dvss.n193 9.3
R17190 dvss.n563 dvss.n562 9.3
R17191 dvss.n561 dvss.n159 9.3
R17192 dvss.n600 dvss.n158 9.3
R17193 dvss.n602 dvss.n601 9.3
R17194 dvss.n2874 dvss.n2873 9.3
R17195 dvss.n2876 dvss.n2875 9.3
R17196 dvss.n2808 dvss.n2807 9.3
R17197 dvss.n2806 dvss.n663 9.3
R17198 dvss.n1739 dvss.n1738 9.259
R17199 dvss.n1739 dvss.n1435 9.259
R17200 dvss.n1757 dvss.n1435 9.259
R17201 dvss.n1760 dvss.n1759 9.259
R17202 dvss.n1760 dvss.n1424 9.259
R17203 dvss.n1777 dvss.n1424 9.259
R17204 dvss.n1778 dvss.n1777 9.259
R17205 dvss.n1779 dvss.n1778 9.259
R17206 dvss.n1796 dvss.n1795 9.259
R17207 dvss.n1821 dvss.n1796 9.259
R17208 dvss.n1821 dvss.n1820 9.259
R17209 dvss.n2357 dvss.n2356 9.259
R17210 dvss.n2357 dvss.n2053 9.259
R17211 dvss.n2375 dvss.n2053 9.259
R17212 dvss.n2378 dvss.n2377 9.259
R17213 dvss.n2378 dvss.n2042 9.259
R17214 dvss.n2395 dvss.n2042 9.259
R17215 dvss.n2396 dvss.n2395 9.259
R17216 dvss.n2397 dvss.n2396 9.259
R17217 dvss.n2414 dvss.n2413 9.259
R17218 dvss.n2439 dvss.n2414 9.259
R17219 dvss.n2439 dvss.n2438 9.259
R17220 dvss.n1126 dvss.n1125 9.259
R17221 dvss.n1126 dvss.n822 9.259
R17222 dvss.n1144 dvss.n822 9.259
R17223 dvss.n1147 dvss.n1146 9.259
R17224 dvss.n1147 dvss.n811 9.259
R17225 dvss.n1164 dvss.n811 9.259
R17226 dvss.n1165 dvss.n1164 9.259
R17227 dvss.n1166 dvss.n1165 9.259
R17228 dvss.n1183 dvss.n1182 9.259
R17229 dvss.n1208 dvss.n1183 9.259
R17230 dvss.n1208 dvss.n1207 9.259
R17231 dvss.n514 dvss.n513 9.259
R17232 dvss.n514 dvss.n210 9.259
R17233 dvss.n532 dvss.n210 9.259
R17234 dvss.n535 dvss.n534 9.259
R17235 dvss.n535 dvss.n199 9.259
R17236 dvss.n552 dvss.n199 9.259
R17237 dvss.n553 dvss.n552 9.259
R17238 dvss.n554 dvss.n553 9.259
R17239 dvss.n571 dvss.n570 9.259
R17240 dvss.n596 dvss.n571 9.259
R17241 dvss.n596 dvss.n595 9.259
R17242 dvss.n2745 dvss.n2744 9.154
R17243 dvss.n2746 dvss.n2745 9.154
R17244 dvss.n2693 dvss.n2691 9.154
R17245 dvss.n2691 dvss.n2690 9.154
R17246 dvss.n2717 dvss.n2716 9.154
R17247 dvss.n2716 dvss.n2715 9.154
R17248 dvss.n2697 dvss.n2696 9.154
R17249 dvss.n2714 dvss.n2697 9.154
R17250 dvss.n2712 dvss.n2711 9.154
R17251 dvss.n2713 dvss.n2712 9.154
R17252 dvss.n2700 dvss.n2699 9.154
R17253 dvss.n2699 dvss.n2698 9.154
R17254 dvss.n2707 dvss.n2706 9.154
R17255 dvss.n2706 dvss.n2705 9.154
R17256 dvss.n2703 dvss.n2702 9.154
R17257 dvss.n2694 dvss.n2692 9.154
R17258 dvss.n2686 dvss.n2685 9.154
R17259 dvss.n2731 dvss.n2730 9.154
R17260 dvss.n2734 dvss.n2733 9.154
R17261 dvss.n2732 dvss.n2724 9.154
R17262 dvss.n2739 dvss.n2738 9.154
R17263 dvss.n2740 dvss.n2723 9.154
R17264 dvss.n2637 dvss.n2636 9.154
R17265 dvss.n2641 dvss.n2640 9.154
R17266 dvss.n2640 dvss.n2639 9.154
R17267 dvss.n2634 dvss.n2633 9.154
R17268 dvss.n2633 dvss.n2632 9.154
R17269 dvss.n2646 dvss.n2645 9.154
R17270 dvss.n2647 dvss.n2646 9.154
R17271 dvss.n2630 dvss.n2628 9.154
R17272 dvss.n2648 dvss.n2630 9.154
R17273 dvss.n2653 dvss.n2652 9.154
R17274 dvss.n2652 dvss.n2651 9.154
R17275 dvss.n2631 dvss.n2629 9.154
R17276 dvss.n2650 dvss.n2631 9.154
R17277 dvss.n2625 dvss.n2624 9.154
R17278 dvss.n2649 dvss.n2624 9.154
R17279 dvss.n2662 dvss.n2661 9.154
R17280 dvss.n2663 dvss.n2662 9.154
R17281 dvss.n2623 dvss.n2622 9.154
R17282 dvss.n2664 dvss.n2623 9.154
R17283 dvss.n2668 dvss.n2667 9.154
R17284 dvss.n2667 dvss.n2666 9.154
R17285 dvss.n2617 dvss.n2616 9.154
R17286 dvss.n2665 dvss.n2616 9.154
R17287 dvss.n2678 dvss.n2677 9.154
R17288 dvss.n2618 dvss.n2615 9.154
R17289 dvss.n2613 dvss.n2612 9.154
R17290 dvss.n2598 dvss.n2597 9.154
R17291 dvss.n2755 dvss.n2754 9.154
R17292 dvss.n1227 dvss.n1225 9.154
R17293 dvss.n1316 dvss.n1315 9.154
R17294 dvss.n1315 dvss.n1314 9.154
R17295 dvss.n1312 dvss.n1311 9.154
R17296 dvss.n1313 dvss.n1312 9.154
R17297 dvss.n1308 dvss.n1307 9.154
R17298 dvss.n1307 dvss.n1306 9.154
R17299 dvss.n1325 dvss.n1324 9.154
R17300 dvss.n1326 dvss.n1325 9.154
R17301 dvss.n1305 dvss.n1304 9.154
R17302 dvss.n1327 dvss.n1305 9.154
R17303 dvss.n1330 dvss.n1329 9.154
R17304 dvss.n1329 dvss.n1328 9.154
R17305 dvss.n1302 dvss.n1301 9.154
R17306 dvss.n1301 dvss.n1300 9.154
R17307 dvss.n1335 dvss.n1334 9.154
R17308 dvss.n1336 dvss.n1335 9.154
R17309 dvss.n1299 dvss.n1298 9.154
R17310 dvss.n1337 dvss.n1299 9.154
R17311 dvss.n1341 dvss.n1340 9.154
R17312 dvss.n1340 dvss.n1339 9.154
R17313 dvss.n1296 dvss.n1295 9.154
R17314 dvss.n1338 dvss.n1295 9.154
R17315 dvss.n1348 dvss.n1347 9.154
R17316 dvss.n1349 dvss.n1348 9.154
R17317 dvss.n1293 dvss.n1291 9.154
R17318 dvss.n1350 dvss.n1293 9.154
R17319 dvss.n1362 dvss.n1361 9.154
R17320 dvss.n1361 dvss.n1360 9.154
R17321 dvss.n1294 dvss.n1292 9.154
R17322 dvss.n1359 dvss.n1294 9.154
R17323 dvss.n1357 dvss.n1356 9.154
R17324 dvss.n1358 dvss.n1357 9.154
R17325 dvss.n1353 dvss.n1352 9.154
R17326 dvss.n1352 dvss.n1351 9.154
R17327 dvss.n1283 dvss.n1282 9.154
R17328 dvss.n1282 dvss.n1281 9.154
R17329 dvss.n1376 dvss.n1375 9.154
R17330 dvss.n1377 dvss.n1376 9.154
R17331 dvss.n1371 dvss.n1280 9.154
R17332 dvss.n1842 dvss.n1839 9.154
R17333 dvss.n1934 dvss.n1933 9.154
R17334 dvss.n1933 dvss.n1932 9.154
R17335 dvss.n1930 dvss.n1929 9.154
R17336 dvss.n1931 dvss.n1930 9.154
R17337 dvss.n1926 dvss.n1925 9.154
R17338 dvss.n1925 dvss.n1924 9.154
R17339 dvss.n1943 dvss.n1942 9.154
R17340 dvss.n1944 dvss.n1943 9.154
R17341 dvss.n1923 dvss.n1922 9.154
R17342 dvss.n1945 dvss.n1923 9.154
R17343 dvss.n1948 dvss.n1947 9.154
R17344 dvss.n1947 dvss.n1946 9.154
R17345 dvss.n1920 dvss.n1919 9.154
R17346 dvss.n1919 dvss.n1918 9.154
R17347 dvss.n1953 dvss.n1952 9.154
R17348 dvss.n1954 dvss.n1953 9.154
R17349 dvss.n1917 dvss.n1916 9.154
R17350 dvss.n1955 dvss.n1917 9.154
R17351 dvss.n1959 dvss.n1958 9.154
R17352 dvss.n1958 dvss.n1957 9.154
R17353 dvss.n1914 dvss.n1913 9.154
R17354 dvss.n1956 dvss.n1913 9.154
R17355 dvss.n1966 dvss.n1965 9.154
R17356 dvss.n1967 dvss.n1966 9.154
R17357 dvss.n1911 dvss.n1909 9.154
R17358 dvss.n1968 dvss.n1911 9.154
R17359 dvss.n1980 dvss.n1979 9.154
R17360 dvss.n1979 dvss.n1978 9.154
R17361 dvss.n1912 dvss.n1910 9.154
R17362 dvss.n1977 dvss.n1912 9.154
R17363 dvss.n1975 dvss.n1974 9.154
R17364 dvss.n1976 dvss.n1975 9.154
R17365 dvss.n1971 dvss.n1970 9.154
R17366 dvss.n1970 dvss.n1969 9.154
R17367 dvss.n1901 dvss.n1900 9.154
R17368 dvss.n1900 dvss.n1899 9.154
R17369 dvss.n1994 dvss.n1993 9.154
R17370 dvss.n1995 dvss.n1994 9.154
R17371 dvss.n1989 dvss.n1898 9.154
R17372 dvss.n1849 dvss.n1848 9.154
R17373 dvss.n2507 dvss.n2506 9.154
R17374 dvss.n2508 dvss.n2507 9.154
R17375 dvss.n1852 dvss.n1851 9.154
R17376 dvss.n1851 dvss.n1850 9.154
R17377 dvss.n1862 dvss.n1858 9.154
R17378 dvss.n1863 dvss.n1862 9.154
R17379 dvss.n2499 dvss.n1859 9.154
R17380 dvss.n1864 dvss.n1859 9.154
R17381 dvss.n2498 dvss.n2497 9.154
R17382 dvss.n2497 dvss.n2496 9.154
R17383 dvss.n1861 dvss.n1860 9.154
R17384 dvss.n2495 dvss.n1861 9.154
R17385 dvss.n2493 dvss.n2492 9.154
R17386 dvss.n2494 dvss.n2493 9.154
R17387 dvss.n1867 dvss.n1866 9.154
R17388 dvss.n1866 dvss.n1865 9.154
R17389 dvss.n2488 dvss.n2487 9.154
R17390 dvss.n2487 dvss.n2486 9.154
R17391 dvss.n1876 dvss.n1875 9.154
R17392 dvss.n2485 dvss.n1876 9.154
R17393 dvss.n2483 dvss.n2482 9.154
R17394 dvss.n2484 dvss.n2483 9.154
R17395 dvss.n1879 dvss.n1878 9.154
R17396 dvss.n1878 dvss.n1877 9.154
R17397 dvss.n1887 dvss.n1883 9.154
R17398 dvss.n1888 dvss.n1887 9.154
R17399 dvss.n2472 dvss.n1884 9.154
R17400 dvss.n1889 dvss.n1884 9.154
R17401 dvss.n2471 dvss.n2470 9.154
R17402 dvss.n2470 dvss.n2469 9.154
R17403 dvss.n1886 dvss.n1885 9.154
R17404 dvss.n2468 dvss.n1886 9.154
R17405 dvss.n2466 dvss.n2465 9.154
R17406 dvss.n2467 dvss.n2466 9.154
R17407 dvss.n1892 dvss.n1891 9.154
R17408 dvss.n1891 dvss.n1890 9.154
R17409 dvss.n2460 dvss.n2459 9.154
R17410 dvss.n2521 dvss.n2520 9.154
R17411 dvss.n2520 dvss.n2519 9.154
R17412 dvss.n1843 dvss.n1841 9.154
R17413 dvss.n2518 dvss.n1843 9.154
R17414 dvss.n2516 dvss.n2515 9.154
R17415 dvss.n1835 dvss.n1276 9.154
R17416 dvss.n2531 dvss.n2530 9.154
R17417 dvss.n2530 dvss.n2529 9.154
R17418 dvss.n1273 dvss.n1272 9.154
R17419 dvss.n1272 dvss.n1271 9.154
R17420 dvss.n2536 dvss.n2535 9.154
R17421 dvss.n2537 dvss.n2536 9.154
R17422 dvss.n1269 dvss.n1268 9.154
R17423 dvss.n2538 dvss.n1269 9.154
R17424 dvss.n2541 dvss.n2540 9.154
R17425 dvss.n2540 dvss.n2539 9.154
R17426 dvss.n1265 dvss.n1264 9.154
R17427 dvss.n1270 dvss.n1264 9.154
R17428 dvss.n2551 dvss.n2550 9.154
R17429 dvss.n2552 dvss.n2551 9.154
R17430 dvss.n1262 dvss.n1260 9.154
R17431 dvss.n2553 dvss.n1262 9.154
R17432 dvss.n2556 dvss.n2555 9.154
R17433 dvss.n2555 dvss.n2554 9.154
R17434 dvss.n1261 dvss.n1254 9.154
R17435 dvss.n1263 dvss.n1261 9.154
R17436 dvss.n1251 dvss.n1250 9.154
R17437 dvss.n1250 dvss.n1249 9.154
R17438 dvss.n2563 dvss.n2562 9.154
R17439 dvss.n2564 dvss.n2563 9.154
R17440 dvss.n1247 dvss.n1246 9.154
R17441 dvss.n2565 dvss.n1247 9.154
R17442 dvss.n2568 dvss.n2567 9.154
R17443 dvss.n2567 dvss.n2566 9.154
R17444 dvss.n1239 dvss.n1237 9.154
R17445 dvss.n1248 dvss.n1237 9.154
R17446 dvss.n2574 dvss.n2573 9.154
R17447 dvss.n2575 dvss.n2574 9.154
R17448 dvss.n1238 dvss.n1236 9.154
R17449 dvss.n2576 dvss.n1236 9.154
R17450 dvss.n2578 dvss.n1234 9.154
R17451 dvss.n2578 dvss.n2577 9.154
R17452 dvss.n2580 dvss.n2579 9.154
R17453 dvss.n2780 dvss.n2779 9.154
R17454 dvss.n2778 dvss.n2776 9.154
R17455 dvss.n2790 dvss.n2778 9.154
R17456 dvss.n2793 dvss.n2792 9.154
R17457 dvss.n2792 dvss.n2791 9.154
R17458 dvss.n2794 dvss.n2775 9.154
R17459 dvss.n2592 dvss.n2591 9.154
R17460 dvss.n2591 dvss.n2590 9.154
R17461 dvss.n1228 dvss.n1226 9.154
R17462 dvss.n2589 dvss.n1228 9.154
R17463 dvss.n2587 dvss.n2586 9.154
R17464 dvss.n703 dvss.n702 9.154
R17465 dvss.n702 dvss.n701 9.154
R17466 dvss.n699 dvss.n698 9.154
R17467 dvss.n700 dvss.n699 9.154
R17468 dvss.n695 dvss.n694 9.154
R17469 dvss.n694 dvss.n693 9.154
R17470 dvss.n712 dvss.n711 9.154
R17471 dvss.n713 dvss.n712 9.154
R17472 dvss.n692 dvss.n691 9.154
R17473 dvss.n714 dvss.n692 9.154
R17474 dvss.n717 dvss.n716 9.154
R17475 dvss.n716 dvss.n715 9.154
R17476 dvss.n689 dvss.n688 9.154
R17477 dvss.n688 dvss.n687 9.154
R17478 dvss.n722 dvss.n721 9.154
R17479 dvss.n723 dvss.n722 9.154
R17480 dvss.n686 dvss.n685 9.154
R17481 dvss.n724 dvss.n686 9.154
R17482 dvss.n728 dvss.n727 9.154
R17483 dvss.n727 dvss.n726 9.154
R17484 dvss.n683 dvss.n682 9.154
R17485 dvss.n725 dvss.n682 9.154
R17486 dvss.n735 dvss.n734 9.154
R17487 dvss.n736 dvss.n735 9.154
R17488 dvss.n680 dvss.n678 9.154
R17489 dvss.n737 dvss.n680 9.154
R17490 dvss.n749 dvss.n748 9.154
R17491 dvss.n748 dvss.n747 9.154
R17492 dvss.n681 dvss.n679 9.154
R17493 dvss.n746 dvss.n681 9.154
R17494 dvss.n744 dvss.n743 9.154
R17495 dvss.n745 dvss.n744 9.154
R17496 dvss.n740 dvss.n739 9.154
R17497 dvss.n739 dvss.n738 9.154
R17498 dvss.n670 dvss.n669 9.154
R17499 dvss.n669 dvss.n668 9.154
R17500 dvss.n763 dvss.n762 9.154
R17501 dvss.n764 dvss.n763 9.154
R17502 dvss.n758 dvss.n667 9.154
R17503 dvss.n613 dvss.n610 9.154
R17504 dvss.n91 dvss.n90 9.154
R17505 dvss.n90 dvss.n89 9.154
R17506 dvss.n87 dvss.n86 9.154
R17507 dvss.n88 dvss.n87 9.154
R17508 dvss.n83 dvss.n82 9.154
R17509 dvss.n82 dvss.n81 9.154
R17510 dvss.n100 dvss.n99 9.154
R17511 dvss.n101 dvss.n100 9.154
R17512 dvss.n80 dvss.n79 9.154
R17513 dvss.n102 dvss.n80 9.154
R17514 dvss.n105 dvss.n104 9.154
R17515 dvss.n104 dvss.n103 9.154
R17516 dvss.n77 dvss.n76 9.154
R17517 dvss.n76 dvss.n75 9.154
R17518 dvss.n110 dvss.n109 9.154
R17519 dvss.n111 dvss.n110 9.154
R17520 dvss.n74 dvss.n73 9.154
R17521 dvss.n112 dvss.n74 9.154
R17522 dvss.n116 dvss.n115 9.154
R17523 dvss.n115 dvss.n114 9.154
R17524 dvss.n71 dvss.n70 9.154
R17525 dvss.n113 dvss.n70 9.154
R17526 dvss.n123 dvss.n122 9.154
R17527 dvss.n124 dvss.n123 9.154
R17528 dvss.n68 dvss.n66 9.154
R17529 dvss.n125 dvss.n68 9.154
R17530 dvss.n137 dvss.n136 9.154
R17531 dvss.n136 dvss.n135 9.154
R17532 dvss.n69 dvss.n67 9.154
R17533 dvss.n134 dvss.n69 9.154
R17534 dvss.n132 dvss.n131 9.154
R17535 dvss.n133 dvss.n132 9.154
R17536 dvss.n128 dvss.n127 9.154
R17537 dvss.n127 dvss.n126 9.154
R17538 dvss.n58 dvss.n57 9.154
R17539 dvss.n57 dvss.n56 9.154
R17540 dvss.n151 dvss.n150 9.154
R17541 dvss.n152 dvss.n151 9.154
R17542 dvss.n146 dvss.n55 9.154
R17543 dvss.n2886 dvss.n2885 9.154
R17544 dvss.n2885 dvss.n2884 9.154
R17545 dvss.n45 dvss.n44 9.154
R17546 dvss.n44 dvss.n43 9.154
R17547 dvss.n2891 dvss.n2890 9.154
R17548 dvss.n2892 dvss.n2891 9.154
R17549 dvss.n42 dvss.n41 9.154
R17550 dvss.n2893 dvss.n42 9.154
R17551 dvss.n2896 dvss.n2895 9.154
R17552 dvss.n2895 dvss.n2894 9.154
R17553 dvss.n35 dvss.n34 9.154
R17554 dvss.n34 dvss.n33 9.154
R17555 dvss.n2902 dvss.n2901 9.154
R17556 dvss.n2903 dvss.n2902 9.154
R17557 dvss.n32 dvss.n31 9.154
R17558 dvss.n2904 dvss.n32 9.154
R17559 dvss.n2907 dvss.n2906 9.154
R17560 dvss.n2906 dvss.n2905 9.154
R17561 dvss.n23 dvss.n22 9.154
R17562 dvss.n22 dvss.n21 9.154
R17563 dvss.n2912 dvss.n2911 9.154
R17564 dvss.n2913 dvss.n2912 9.154
R17565 dvss.n19 dvss.n18 9.154
R17566 dvss.n2914 dvss.n19 9.154
R17567 dvss.n2917 dvss.n2916 9.154
R17568 dvss.n2916 dvss.n2915 9.154
R17569 dvss.n12 dvss.n10 9.154
R17570 dvss.n20 dvss.n10 9.154
R17571 dvss.n2923 dvss.n2922 9.154
R17572 dvss.n2924 dvss.n2923 9.154
R17573 dvss.n11 dvss.n9 9.154
R17574 dvss.n2925 dvss.n9 9.154
R17575 dvss.n2927 dvss.n7 9.154
R17576 dvss.n2927 dvss.n2926 9.154
R17577 dvss.n2929 dvss.n2928 9.154
R17578 dvss.n2875 dvss.n51 9.154
R17579 dvss.n50 dvss.n49 9.154
R17580 dvss.n2883 dvss.n50 9.154
R17581 dvss.n2868 dvss.n2867 9.154
R17582 dvss.n2867 dvss.n2866 9.154
R17583 dvss.n614 dvss.n612 9.154
R17584 dvss.n2865 dvss.n614 9.154
R17585 dvss.n2863 dvss.n2862 9.154
R17586 dvss.n2856 dvss.n620 9.154
R17587 dvss.n2855 dvss.n2854 9.154
R17588 dvss.n2854 dvss.n2853 9.154
R17589 dvss.n622 dvss.n621 9.154
R17590 dvss.n2852 dvss.n622 9.154
R17591 dvss.n2850 dvss.n2849 9.154
R17592 dvss.n2851 dvss.n2850 9.154
R17593 dvss.n625 dvss.n624 9.154
R17594 dvss.n633 dvss.n624 9.154
R17595 dvss.n2844 dvss.n2843 9.154
R17596 dvss.n2843 dvss.n2842 9.154
R17597 dvss.n632 dvss.n631 9.154
R17598 dvss.n2841 dvss.n632 9.154
R17599 dvss.n2839 dvss.n2838 9.154
R17600 dvss.n2840 dvss.n2839 9.154
R17601 dvss.n636 dvss.n635 9.154
R17602 dvss.n635 dvss.n634 9.154
R17603 dvss.n2834 dvss.n2833 9.154
R17604 dvss.n2833 dvss.n2832 9.154
R17605 dvss.n645 dvss.n644 9.154
R17606 dvss.n2831 dvss.n645 9.154
R17607 dvss.n2829 dvss.n2828 9.154
R17608 dvss.n2830 dvss.n2829 9.154
R17609 dvss.n648 dvss.n647 9.154
R17610 dvss.n647 dvss.n646 9.154
R17611 dvss.n656 dvss.n652 9.154
R17612 dvss.n657 dvss.n656 9.154
R17613 dvss.n2818 dvss.n653 9.154
R17614 dvss.n658 dvss.n653 9.154
R17615 dvss.n2817 dvss.n2816 9.154
R17616 dvss.n2816 dvss.n2815 9.154
R17617 dvss.n655 dvss.n654 9.154
R17618 dvss.n2814 dvss.n655 9.154
R17619 dvss.n2812 dvss.n2811 9.154
R17620 dvss.n2813 dvss.n2812 9.154
R17621 dvss.n661 dvss.n660 9.154
R17622 dvss.n660 dvss.n659 9.154
R17623 dvss.n2806 dvss.n2805 9.154
R17624 dvss.n2760 dvss.n2759 9.154
R17625 dvss.n2759 dvss.n2758 9.154
R17626 dvss.n2764 dvss.n2763 9.154
R17627 dvss.n2763 dvss.n2762 9.154
R17628 dvss.n2769 dvss.n2768 9.154
R17629 dvss.n2608 dvss.n2607 9.154
R17630 dvss.n2607 dvss.n2606 9.154
R17631 dvss.n2604 dvss.n2603 9.154
R17632 dvss.n2603 dvss.n2602 9.154
R17633 dvss.n2 dvss.n1 9.154
R17634 dvss.n1387 dvss.n1386 9.013
R17635 dvss.n1824 dvss.n1823 9.013
R17636 dvss.n1393 dvss.n1385 9.013
R17637 dvss.n1793 dvss.n1792 9.013
R17638 dvss.n1782 dvss.n1781 9.013
R17639 dvss.n1422 dvss.n1421 9.013
R17640 dvss.n1775 dvss.n1774 9.013
R17641 dvss.n1427 dvss.n1426 9.013
R17642 dvss.n1763 dvss.n1762 9.013
R17643 dvss.n1432 dvss.n1431 9.013
R17644 dvss.n1755 dvss.n1754 9.013
R17645 dvss.n1440 dvss.n1438 9.013
R17646 dvss.n1742 dvss.n1741 9.013
R17647 dvss.n1471 dvss.n1470 9.013
R17648 dvss.n2005 dvss.n2004 9.013
R17649 dvss.n2442 dvss.n2441 9.013
R17650 dvss.n2011 dvss.n2003 9.013
R17651 dvss.n2411 dvss.n2410 9.013
R17652 dvss.n2400 dvss.n2399 9.013
R17653 dvss.n2040 dvss.n2039 9.013
R17654 dvss.n2393 dvss.n2392 9.013
R17655 dvss.n2045 dvss.n2044 9.013
R17656 dvss.n2381 dvss.n2380 9.013
R17657 dvss.n2050 dvss.n2049 9.013
R17658 dvss.n2373 dvss.n2372 9.013
R17659 dvss.n2058 dvss.n2056 9.013
R17660 dvss.n2360 dvss.n2359 9.013
R17661 dvss.n2089 dvss.n2088 9.013
R17662 dvss.n774 dvss.n773 9.013
R17663 dvss.n1211 dvss.n1210 9.013
R17664 dvss.n780 dvss.n772 9.013
R17665 dvss.n1180 dvss.n1179 9.013
R17666 dvss.n1169 dvss.n1168 9.013
R17667 dvss.n809 dvss.n808 9.013
R17668 dvss.n1162 dvss.n1161 9.013
R17669 dvss.n814 dvss.n813 9.013
R17670 dvss.n1150 dvss.n1149 9.013
R17671 dvss.n819 dvss.n818 9.013
R17672 dvss.n1142 dvss.n1141 9.013
R17673 dvss.n827 dvss.n825 9.013
R17674 dvss.n1129 dvss.n1128 9.013
R17675 dvss.n858 dvss.n857 9.013
R17676 dvss.n162 dvss.n161 9.013
R17677 dvss.n599 dvss.n598 9.013
R17678 dvss.n168 dvss.n160 9.013
R17679 dvss.n568 dvss.n567 9.013
R17680 dvss.n557 dvss.n556 9.013
R17681 dvss.n197 dvss.n196 9.013
R17682 dvss.n550 dvss.n549 9.013
R17683 dvss.n202 dvss.n201 9.013
R17684 dvss.n538 dvss.n537 9.013
R17685 dvss.n207 dvss.n206 9.013
R17686 dvss.n530 dvss.n529 9.013
R17687 dvss.n215 dvss.n213 9.013
R17688 dvss.n517 dvss.n516 9.013
R17689 dvss.n246 dvss.n245 9.013
R17690 dvss.n1483 dvss.n1470 9.013
R17691 dvss.n1743 dvss.n1742 9.013
R17692 dvss.n1745 dvss.n1440 9.013
R17693 dvss.n1754 dvss.n1753 9.013
R17694 dvss.n1749 dvss.n1431 9.013
R17695 dvss.n1764 dvss.n1763 9.013
R17696 dvss.n1766 dvss.n1427 9.013
R17697 dvss.n1774 dvss.n1773 9.013
R17698 dvss.n1770 dvss.n1421 9.013
R17699 dvss.n1783 dvss.n1782 9.013
R17700 dvss.n1792 dvss.n1791 9.013
R17701 dvss.n1787 dvss.n1385 9.013
R17702 dvss.n1825 dvss.n1824 9.013
R17703 dvss.n1386 dvss.n1382 9.013
R17704 dvss.n2101 dvss.n2088 9.013
R17705 dvss.n2361 dvss.n2360 9.013
R17706 dvss.n2363 dvss.n2058 9.013
R17707 dvss.n2372 dvss.n2371 9.013
R17708 dvss.n2367 dvss.n2049 9.013
R17709 dvss.n2382 dvss.n2381 9.013
R17710 dvss.n2384 dvss.n2045 9.013
R17711 dvss.n2392 dvss.n2391 9.013
R17712 dvss.n2388 dvss.n2039 9.013
R17713 dvss.n2401 dvss.n2400 9.013
R17714 dvss.n2410 dvss.n2409 9.013
R17715 dvss.n2405 dvss.n2003 9.013
R17716 dvss.n2443 dvss.n2442 9.013
R17717 dvss.n2004 dvss.n2000 9.013
R17718 dvss.n870 dvss.n857 9.013
R17719 dvss.n1130 dvss.n1129 9.013
R17720 dvss.n1132 dvss.n827 9.013
R17721 dvss.n1141 dvss.n1140 9.013
R17722 dvss.n1136 dvss.n818 9.013
R17723 dvss.n1151 dvss.n1150 9.013
R17724 dvss.n1153 dvss.n814 9.013
R17725 dvss.n1161 dvss.n1160 9.013
R17726 dvss.n1157 dvss.n808 9.013
R17727 dvss.n1170 dvss.n1169 9.013
R17728 dvss.n1179 dvss.n1178 9.013
R17729 dvss.n1174 dvss.n772 9.013
R17730 dvss.n1212 dvss.n1211 9.013
R17731 dvss.n773 dvss.n769 9.013
R17732 dvss.n258 dvss.n245 9.013
R17733 dvss.n518 dvss.n517 9.013
R17734 dvss.n520 dvss.n215 9.013
R17735 dvss.n529 dvss.n528 9.013
R17736 dvss.n524 dvss.n206 9.013
R17737 dvss.n539 dvss.n538 9.013
R17738 dvss.n541 dvss.n202 9.013
R17739 dvss.n549 dvss.n548 9.013
R17740 dvss.n545 dvss.n196 9.013
R17741 dvss.n558 dvss.n557 9.013
R17742 dvss.n567 dvss.n566 9.013
R17743 dvss.n562 dvss.n160 9.013
R17744 dvss.n600 dvss.n599 9.013
R17745 dvss.n161 dvss.n157 9.013
R17746 dvss.n1681 dvss.n1674 8.973
R17747 dvss.n2299 dvss.n2292 8.973
R17748 dvss.n1068 dvss.n1061 8.973
R17749 dvss.n456 dvss.n449 8.973
R17750 dvss.n2679 dvss.n2678 8.855
R17751 dvss.n2723 dvss.n2689 8.854
R17752 dvss.n2732 dvss.n2688 8.854
R17753 dvss.n2730 dvss.n2687 8.854
R17754 dvss.n2692 dvss.n2689 8.854
R17755 dvss.n2748 dvss.n2686 8.854
R17756 dvss.n2733 dvss.n2687 8.854
R17757 dvss.n2738 dvss.n2688 8.854
R17758 dvss.n2681 dvss.n2613 8.854
R17759 dvss.n2679 dvss.n2615 8.854
R17760 dvss.n1657 dvss.n1656 8.151
R17761 dvss.n2275 dvss.n2274 8.151
R17762 dvss.n1044 dvss.n1043 8.151
R17763 dvss.n432 dvss.n431 8.151
R17764 dvss.n1737 dvss.n1473 7.568
R17765 dvss.n1731 dvss.n1473 7.568
R17766 dvss.n1731 dvss.n1730 7.568
R17767 dvss.n1730 dvss.n1728 7.568
R17768 dvss.n1728 dvss.n1726 7.568
R17769 dvss.n1726 dvss.n1724 7.568
R17770 dvss.n1724 dvss.n1722 7.568
R17771 dvss.n1722 dvss.n1720 7.568
R17772 dvss.n1819 dvss.n1797 7.568
R17773 dvss.n1813 dvss.n1797 7.568
R17774 dvss.n1813 dvss.n1812 7.568
R17775 dvss.n1812 dvss.n1811 7.568
R17776 dvss.n1811 dvss.n1808 7.568
R17777 dvss.n1808 dvss.n1807 7.568
R17778 dvss.n1807 dvss.n1804 7.568
R17779 dvss.n1804 dvss.n1381 7.568
R17780 dvss.n2355 dvss.n2091 7.568
R17781 dvss.n2349 dvss.n2091 7.568
R17782 dvss.n2349 dvss.n2348 7.568
R17783 dvss.n2348 dvss.n2346 7.568
R17784 dvss.n2346 dvss.n2344 7.568
R17785 dvss.n2344 dvss.n2342 7.568
R17786 dvss.n2342 dvss.n2340 7.568
R17787 dvss.n2340 dvss.n2338 7.568
R17788 dvss.n2437 dvss.n2415 7.568
R17789 dvss.n2431 dvss.n2415 7.568
R17790 dvss.n2431 dvss.n2430 7.568
R17791 dvss.n2430 dvss.n2429 7.568
R17792 dvss.n2429 dvss.n2426 7.568
R17793 dvss.n2426 dvss.n2425 7.568
R17794 dvss.n2425 dvss.n2422 7.568
R17795 dvss.n2422 dvss.n1999 7.568
R17796 dvss.n1124 dvss.n860 7.568
R17797 dvss.n1118 dvss.n860 7.568
R17798 dvss.n1118 dvss.n1117 7.568
R17799 dvss.n1117 dvss.n1115 7.568
R17800 dvss.n1115 dvss.n1113 7.568
R17801 dvss.n1113 dvss.n1111 7.568
R17802 dvss.n1111 dvss.n1109 7.568
R17803 dvss.n1109 dvss.n1107 7.568
R17804 dvss.n1206 dvss.n1184 7.568
R17805 dvss.n1200 dvss.n1184 7.568
R17806 dvss.n1200 dvss.n1199 7.568
R17807 dvss.n1199 dvss.n1198 7.568
R17808 dvss.n1198 dvss.n1195 7.568
R17809 dvss.n1195 dvss.n1194 7.568
R17810 dvss.n1194 dvss.n1191 7.568
R17811 dvss.n1191 dvss.n768 7.568
R17812 dvss.n512 dvss.n248 7.568
R17813 dvss.n506 dvss.n248 7.568
R17814 dvss.n506 dvss.n505 7.568
R17815 dvss.n505 dvss.n503 7.568
R17816 dvss.n503 dvss.n501 7.568
R17817 dvss.n501 dvss.n499 7.568
R17818 dvss.n499 dvss.n497 7.568
R17819 dvss.n497 dvss.n495 7.568
R17820 dvss.n594 dvss.n572 7.568
R17821 dvss.n588 dvss.n572 7.568
R17822 dvss.n588 dvss.n587 7.568
R17823 dvss.n587 dvss.n586 7.568
R17824 dvss.n586 dvss.n583 7.568
R17825 dvss.n583 dvss.n582 7.568
R17826 dvss.n582 dvss.n579 7.568
R17827 dvss.n579 dvss.n156 7.568
R17828 dvss.n1673 dvss.n1672 6.467
R17829 dvss.n2291 dvss.n2290 6.467
R17830 dvss.n1060 dvss.n1059 6.467
R17831 dvss.n448 dvss.n447 6.467
R17832 dvss.n1588 dvss.n1587 5.726
R17833 dvss.n1587 dvss.n1586 5.726
R17834 dvss.n1586 dvss.n1583 5.726
R17835 dvss.n1583 dvss.n1582 5.726
R17836 dvss.n1582 dvss.n1579 5.726
R17837 dvss.n1579 dvss.n1578 5.726
R17838 dvss.n1578 dvss.n1571 5.726
R17839 dvss.n1594 dvss.n1571 5.726
R17840 dvss.n2206 dvss.n2205 5.726
R17841 dvss.n2205 dvss.n2204 5.726
R17842 dvss.n2204 dvss.n2201 5.726
R17843 dvss.n2201 dvss.n2200 5.726
R17844 dvss.n2200 dvss.n2197 5.726
R17845 dvss.n2197 dvss.n2196 5.726
R17846 dvss.n2196 dvss.n2189 5.726
R17847 dvss.n2212 dvss.n2189 5.726
R17848 dvss.n975 dvss.n974 5.726
R17849 dvss.n974 dvss.n973 5.726
R17850 dvss.n973 dvss.n970 5.726
R17851 dvss.n970 dvss.n969 5.726
R17852 dvss.n969 dvss.n966 5.726
R17853 dvss.n966 dvss.n965 5.726
R17854 dvss.n965 dvss.n958 5.726
R17855 dvss.n981 dvss.n958 5.726
R17856 dvss.n363 dvss.n362 5.726
R17857 dvss.n362 dvss.n361 5.726
R17858 dvss.n361 dvss.n358 5.726
R17859 dvss.n358 dvss.n357 5.726
R17860 dvss.n357 dvss.n354 5.726
R17861 dvss.n354 dvss.n353 5.726
R17862 dvss.n353 dvss.n346 5.726
R17863 dvss.n369 dvss.n346 5.726
R17864 dvss.n1835 dvss.n1277 5.647
R17865 dvss.n1521 dvss.n1520 5.647
R17866 dvss.n1520 dvss.n1510 5.647
R17867 dvss.n1500 dvss.n1499 5.647
R17868 dvss.n1499 dvss.n1489 5.647
R17869 dvss.n2460 dvss.n1895 5.647
R17870 dvss.n2139 dvss.n2138 5.647
R17871 dvss.n2138 dvss.n2128 5.647
R17872 dvss.n2118 dvss.n2117 5.647
R17873 dvss.n2117 dvss.n2107 5.647
R17874 dvss.n2806 dvss.n664 5.647
R17875 dvss.n908 dvss.n907 5.647
R17876 dvss.n907 dvss.n897 5.647
R17877 dvss.n887 dvss.n886 5.647
R17878 dvss.n886 dvss.n876 5.647
R17879 dvss.n296 dvss.n295 5.647
R17880 dvss.n295 dvss.n285 5.647
R17881 dvss.n275 dvss.n274 5.647
R17882 dvss.n274 dvss.n264 5.647
R17883 dvss.n2875 dvss.n52 5.647
R17884 dvss.n1750 dvss.n1749 5.579
R17885 dvss.n1784 dvss.n1783 5.579
R17886 dvss.n2368 dvss.n2367 5.579
R17887 dvss.n2402 dvss.n2401 5.579
R17888 dvss.n1137 dvss.n1136 5.579
R17889 dvss.n1171 dvss.n1170 5.579
R17890 dvss.n525 dvss.n524 5.579
R17891 dvss.n559 dvss.n558 5.579
R17892 dvss.n1753 dvss.n1466 5.345
R17893 dvss.n2371 dvss.n2084 5.345
R17894 dvss.n1140 dvss.n853 5.345
R17895 dvss.n528 dvss.n241 5.345
R17896 dvss.n1791 dvss.n1417 5.298
R17897 dvss.n2409 dvss.n2035 5.298
R17898 dvss.n1178 dvss.n804 5.298
R17899 dvss.n566 dvss.n192 5.298
R17900 dvss.n1371 dvss.n1279 5.27
R17901 dvss.n1989 dvss.n1897 5.27
R17902 dvss.n758 dvss.n666 5.27
R17903 dvss.n146 dvss.n54 5.27
R17904 dvss.n1524 dvss.n1507 4.894
R17905 dvss.n1503 dvss.n1486 4.894
R17906 dvss.n2142 dvss.n2125 4.894
R17907 dvss.n2121 dvss.n2104 4.894
R17908 dvss.n911 dvss.n894 4.894
R17909 dvss.n890 dvss.n873 4.894
R17910 dvss.n299 dvss.n282 4.894
R17911 dvss.n278 dvss.n261 4.894
R17912 dvss.n1692 dvss.n1545 4.742
R17913 dvss.n1625 dvss.n1562 4.742
R17914 dvss.n2310 dvss.n2163 4.742
R17915 dvss.n2243 dvss.n2180 4.742
R17916 dvss.n1079 dvss.n932 4.742
R17917 dvss.n1012 dvss.n949 4.742
R17918 dvss.n467 dvss.n320 4.742
R17919 dvss.n400 dvss.n337 4.742
R17920 dvss.n2750 dvss.n2749 4.65
R17921 dvss.n2728 dvss.n2727 4.65
R17922 dvss.n2727 dvss.n2725 4.65
R17923 dvss.n2744 dvss.n2743 4.65
R17924 dvss.n2719 dvss.n2693 4.65
R17925 dvss.n2718 dvss.n2717 4.65
R17926 dvss.n2696 dvss.n2695 4.65
R17927 dvss.n2711 dvss.n2710 4.65
R17928 dvss.n2709 dvss.n2700 4.65
R17929 dvss.n2708 dvss.n2707 4.65
R17930 dvss.n2742 dvss.n2694 4.65
R17931 dvss.n2685 dvss.n2684 4.65
R17932 dvss.n2731 dvss.n2729 4.65
R17933 dvss.n2735 dvss.n2734 4.65
R17934 dvss.n2736 dvss.n2724 4.65
R17935 dvss.n2739 dvss.n2737 4.65
R17936 dvss.n2741 dvss.n2740 4.65
R17937 dvss.n2656 dvss.n2655 4.65
R17938 dvss.n2657 dvss.n2656 4.65
R17939 dvss.n2675 dvss.n2672 4.65
R17940 dvss.n2673 dvss.n2672 4.65
R17941 dvss.n2642 dvss.n2641 4.65
R17942 dvss.n2643 dvss.n2634 4.65
R17943 dvss.n2645 dvss.n2644 4.65
R17944 dvss.n2628 dvss.n2627 4.65
R17945 dvss.n2654 dvss.n2653 4.65
R17946 dvss.n2629 dvss.n2626 4.65
R17947 dvss.n2658 dvss.n2625 4.65
R17948 dvss.n2661 dvss.n2660 4.65
R17949 dvss.n2659 dvss.n2622 4.65
R17950 dvss.n2669 dvss.n2668 4.65
R17951 dvss.n2670 dvss.n2617 4.65
R17952 dvss.n2677 dvss.n2676 4.65
R17953 dvss.n2674 dvss.n2618 4.65
R17954 dvss.n2612 dvss.n2611 4.65
R17955 dvss.n2683 dvss.n2682 4.65
R17956 dvss.n1365 dvss.n1288 4.65
R17957 dvss.n1365 dvss.n1364 4.65
R17958 dvss.n1345 dvss.n1287 4.65
R17959 dvss.n1343 dvss.n1287 4.65
R17960 dvss.n1321 dvss.n1320 4.65
R17961 dvss.n1320 dvss.n1318 4.65
R17962 dvss.n1311 dvss.n1309 4.65
R17963 dvss.n1322 dvss.n1308 4.65
R17964 dvss.n1324 dvss.n1323 4.65
R17965 dvss.n1304 dvss.n1303 4.65
R17966 dvss.n1331 dvss.n1330 4.65
R17967 dvss.n1332 dvss.n1302 4.65
R17968 dvss.n1334 dvss.n1333 4.65
R17969 dvss.n1298 dvss.n1297 4.65
R17970 dvss.n1342 dvss.n1341 4.65
R17971 dvss.n1344 dvss.n1296 4.65
R17972 dvss.n1347 dvss.n1346 4.65
R17973 dvss.n1291 dvss.n1290 4.65
R17974 dvss.n1363 dvss.n1362 4.65
R17975 dvss.n1354 dvss.n1292 4.65
R17976 dvss.n1356 dvss.n1355 4.65
R17977 dvss.n1353 dvss.n1285 4.65
R17978 dvss.n1369 dvss.n1283 4.65
R17979 dvss.n1375 dvss.n1374 4.65
R17980 dvss.n1692 dvss.n1691 4.65
R17981 dvss.n1712 dvss.n1711 4.65
R17982 dvss.n1694 dvss.n1693 4.65
R17983 dvss.n1697 dvss.n1543 4.65
R17984 dvss.n1701 dvss.n1700 4.65
R17985 dvss.n1703 dvss.n1702 4.65
R17986 dvss.n1542 dvss.n1539 4.65
R17987 dvss.n1528 dvss.n1526 4.65
R17988 dvss.n1609 dvss.n1505 4.65
R17989 dvss.n1636 dvss.n1635 4.65
R17990 dvss.n1638 dvss.n1637 4.65
R17991 dvss.n1624 dvss.n1620 4.65
R17992 dvss.n1613 dvss.n1611 4.65
R17993 dvss.n1646 dvss.n1645 4.65
R17994 dvss.n1648 dvss.n1647 4.65
R17995 dvss.n1626 dvss.n1625 4.65
R17996 dvss.n1983 dvss.n1906 4.65
R17997 dvss.n1983 dvss.n1982 4.65
R17998 dvss.n1963 dvss.n1905 4.65
R17999 dvss.n1961 dvss.n1905 4.65
R18000 dvss.n1939 dvss.n1938 4.65
R18001 dvss.n1938 dvss.n1936 4.65
R18002 dvss.n1929 dvss.n1927 4.65
R18003 dvss.n1940 dvss.n1926 4.65
R18004 dvss.n1942 dvss.n1941 4.65
R18005 dvss.n1922 dvss.n1921 4.65
R18006 dvss.n1949 dvss.n1948 4.65
R18007 dvss.n1950 dvss.n1920 4.65
R18008 dvss.n1952 dvss.n1951 4.65
R18009 dvss.n1916 dvss.n1915 4.65
R18010 dvss.n1960 dvss.n1959 4.65
R18011 dvss.n1962 dvss.n1914 4.65
R18012 dvss.n1965 dvss.n1964 4.65
R18013 dvss.n1909 dvss.n1908 4.65
R18014 dvss.n1981 dvss.n1980 4.65
R18015 dvss.n1972 dvss.n1910 4.65
R18016 dvss.n1974 dvss.n1973 4.65
R18017 dvss.n1971 dvss.n1903 4.65
R18018 dvss.n1987 dvss.n1901 4.65
R18019 dvss.n1993 dvss.n1992 4.65
R18020 dvss.n2310 dvss.n2309 4.65
R18021 dvss.n2330 dvss.n2329 4.65
R18022 dvss.n2312 dvss.n2311 4.65
R18023 dvss.n2315 dvss.n2161 4.65
R18024 dvss.n2319 dvss.n2318 4.65
R18025 dvss.n2321 dvss.n2320 4.65
R18026 dvss.n2160 dvss.n2157 4.65
R18027 dvss.n2146 dvss.n2144 4.65
R18028 dvss.n2227 dvss.n2123 4.65
R18029 dvss.n2254 dvss.n2253 4.65
R18030 dvss.n2256 dvss.n2255 4.65
R18031 dvss.n2242 dvss.n2238 4.65
R18032 dvss.n2231 dvss.n2229 4.65
R18033 dvss.n2264 dvss.n2263 4.65
R18034 dvss.n2266 dvss.n2265 4.65
R18035 dvss.n2244 dvss.n2243 4.65
R18036 dvss.n2477 dvss.n2476 4.65
R18037 dvss.n2502 dvss.n2501 4.65
R18038 dvss.n1871 dvss.n1870 4.65
R18039 dvss.n1872 dvss.n1871 4.65
R18040 dvss.n2503 dvss.n2502 4.65
R18041 dvss.n1853 dvss.n1848 4.65
R18042 dvss.n2506 dvss.n2505 4.65
R18043 dvss.n2504 dvss.n1852 4.65
R18044 dvss.n1858 dvss.n1854 4.65
R18045 dvss.n2500 dvss.n2499 4.65
R18046 dvss.n2498 dvss.n1857 4.65
R18047 dvss.n1868 dvss.n1860 4.65
R18048 dvss.n2492 dvss.n2491 4.65
R18049 dvss.n2490 dvss.n1867 4.65
R18050 dvss.n2489 dvss.n2488 4.65
R18051 dvss.n1880 dvss.n1875 4.65
R18052 dvss.n2482 dvss.n2481 4.65
R18053 dvss.n2480 dvss.n1879 4.65
R18054 dvss.n1883 dvss.n1881 4.65
R18055 dvss.n2473 dvss.n2472 4.65
R18056 dvss.n2471 dvss.n1882 4.65
R18057 dvss.n1893 dvss.n1885 4.65
R18058 dvss.n2465 dvss.n2464 4.65
R18059 dvss.n2463 dvss.n1892 4.65
R18060 dvss.n2511 dvss.n2510 4.65
R18061 dvss.n2524 dvss.n1839 4.65
R18062 dvss.n2522 dvss.n2521 4.65
R18063 dvss.n1841 dvss.n1840 4.65
R18064 dvss.n2515 dvss.n2514 4.65
R18065 dvss.n2513 dvss.n1844 4.65
R18066 dvss.n1846 dvss.n1845 4.65
R18067 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vss1p8 dvss.n1846 4.65
R18068 dvss.n2512 dvss.n1846 4.65
R18069 dvss.n2571 dvss.n1244 4.65
R18070 dvss.n2546 dvss.n2545 4.65
R18071 dvss.n2532 dvss.n2531 4.65
R18072 dvss.n2533 dvss.n1273 4.65
R18073 dvss.n2535 dvss.n2534 4.65
R18074 dvss.n1268 dvss.n1267 4.65
R18075 dvss.n2542 dvss.n2541 4.65
R18076 dvss.n1266 dvss.n1265 4.65
R18077 dvss.n2550 dvss.n2549 4.65
R18078 dvss.n1260 dvss.n1259 4.65
R18079 dvss.n2557 dvss.n2556 4.65
R18080 dvss.n2559 dvss.n1254 4.65
R18081 dvss.n2560 dvss.n1251 4.65
R18082 dvss.n2562 dvss.n2561 4.65
R18083 dvss.n1252 dvss.n1246 4.65
R18084 dvss.n2569 dvss.n2568 4.65
R18085 dvss.n2570 dvss.n1239 4.65
R18086 dvss.n2573 dvss.n2572 4.65
R18087 dvss.n1241 dvss.n1238 4.65
R18088 dvss.n1240 dvss.n1234 4.65
R18089 dvss.n2580 dvss.n1235 4.65
R18090 dvss.n1256 dvss.n1245 4.65
R18091 dvss.n1256 dvss.n1253 4.65
R18092 dvss.n1244 dvss.n1242 4.65
R18093 dvss.n2582 dvss.n2581 4.65
R18094 dvss.n2788 dvss.n2787 4.65
R18095 dvss.n2783 dvss.n2780 4.65
R18096 dvss.n2781 dvss.n2776 4.65
R18097 dvss.n2793 dvss.n2777 4.65
R18098 dvss.n2795 dvss.n2794 4.65
R18099 dvss.n2786 dvss.n2785 4.65
R18100 dvss.n2785 dvss.n2784 4.65
R18101 dvss.n2785 dvss.n2782 4.65
R18102 dvss.n1225 dvss.n1222 4.65
R18103 dvss.n2593 dvss.n2592 4.65
R18104 dvss.n1226 dvss.n1224 4.65
R18105 dvss.n2586 dvss.n2585 4.65
R18106 dvss.n2584 dvss.n1229 4.65
R18107 dvss.n1231 dvss.n1230 4.65
R18108 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vss1p8 dvss.n1231 4.65
R18109 dvss.n2583 dvss.n1231 4.65
R18110 dvss.n752 dvss.n675 4.65
R18111 dvss.n752 dvss.n751 4.65
R18112 dvss.n732 dvss.n674 4.65
R18113 dvss.n730 dvss.n674 4.65
R18114 dvss.n708 dvss.n707 4.65
R18115 dvss.n707 dvss.n705 4.65
R18116 dvss.n698 dvss.n696 4.65
R18117 dvss.n709 dvss.n695 4.65
R18118 dvss.n711 dvss.n710 4.65
R18119 dvss.n691 dvss.n690 4.65
R18120 dvss.n718 dvss.n717 4.65
R18121 dvss.n719 dvss.n689 4.65
R18122 dvss.n721 dvss.n720 4.65
R18123 dvss.n685 dvss.n684 4.65
R18124 dvss.n729 dvss.n728 4.65
R18125 dvss.n731 dvss.n683 4.65
R18126 dvss.n734 dvss.n733 4.65
R18127 dvss.n678 dvss.n677 4.65
R18128 dvss.n750 dvss.n749 4.65
R18129 dvss.n741 dvss.n679 4.65
R18130 dvss.n743 dvss.n742 4.65
R18131 dvss.n740 dvss.n672 4.65
R18132 dvss.n756 dvss.n670 4.65
R18133 dvss.n762 dvss.n761 4.65
R18134 dvss.n1079 dvss.n1078 4.65
R18135 dvss.n1099 dvss.n1098 4.65
R18136 dvss.n1081 dvss.n1080 4.65
R18137 dvss.n1084 dvss.n930 4.65
R18138 dvss.n1088 dvss.n1087 4.65
R18139 dvss.n1090 dvss.n1089 4.65
R18140 dvss.n929 dvss.n926 4.65
R18141 dvss.n915 dvss.n913 4.65
R18142 dvss.n996 dvss.n892 4.65
R18143 dvss.n1023 dvss.n1022 4.65
R18144 dvss.n1025 dvss.n1024 4.65
R18145 dvss.n1011 dvss.n1007 4.65
R18146 dvss.n1000 dvss.n998 4.65
R18147 dvss.n1033 dvss.n1032 4.65
R18148 dvss.n1035 dvss.n1034 4.65
R18149 dvss.n1013 dvss.n1012 4.65
R18150 dvss.n140 dvss.n63 4.65
R18151 dvss.n140 dvss.n139 4.65
R18152 dvss.n120 dvss.n62 4.65
R18153 dvss.n118 dvss.n62 4.65
R18154 dvss.n96 dvss.n95 4.65
R18155 dvss.n95 dvss.n93 4.65
R18156 dvss.n86 dvss.n84 4.65
R18157 dvss.n97 dvss.n83 4.65
R18158 dvss.n99 dvss.n98 4.65
R18159 dvss.n79 dvss.n78 4.65
R18160 dvss.n106 dvss.n105 4.65
R18161 dvss.n107 dvss.n77 4.65
R18162 dvss.n109 dvss.n108 4.65
R18163 dvss.n73 dvss.n72 4.65
R18164 dvss.n117 dvss.n116 4.65
R18165 dvss.n119 dvss.n71 4.65
R18166 dvss.n122 dvss.n121 4.65
R18167 dvss.n66 dvss.n65 4.65
R18168 dvss.n138 dvss.n137 4.65
R18169 dvss.n129 dvss.n67 4.65
R18170 dvss.n131 dvss.n130 4.65
R18171 dvss.n128 dvss.n60 4.65
R18172 dvss.n144 dvss.n58 4.65
R18173 dvss.n150 dvss.n149 4.65
R18174 dvss.n467 dvss.n466 4.65
R18175 dvss.n487 dvss.n486 4.65
R18176 dvss.n469 dvss.n468 4.65
R18177 dvss.n472 dvss.n318 4.65
R18178 dvss.n476 dvss.n475 4.65
R18179 dvss.n478 dvss.n477 4.65
R18180 dvss.n317 dvss.n314 4.65
R18181 dvss.n303 dvss.n301 4.65
R18182 dvss.n384 dvss.n280 4.65
R18183 dvss.n411 dvss.n410 4.65
R18184 dvss.n413 dvss.n412 4.65
R18185 dvss.n399 dvss.n395 4.65
R18186 dvss.n388 dvss.n386 4.65
R18187 dvss.n421 dvss.n420 4.65
R18188 dvss.n423 dvss.n422 4.65
R18189 dvss.n401 dvss.n400 4.65
R18190 dvss.n2932 dvss.n5 4.65
R18191 dvss.n16 dvss.n14 4.65
R18192 dvss.n2920 dvss.n16 4.65
R18193 dvss.n27 dvss.n17 4.65
R18194 dvss.n27 dvss.n25 4.65
R18195 dvss.n40 dvss.n39 4.65
R18196 dvss.n2887 dvss.n2886 4.65
R18197 dvss.n2888 dvss.n45 4.65
R18198 dvss.n2890 dvss.n2889 4.65
R18199 dvss.n47 dvss.n41 4.65
R18200 dvss.n2897 dvss.n2896 4.65
R18201 dvss.n2899 dvss.n35 4.65
R18202 dvss.n2901 dvss.n2900 4.65
R18203 dvss.n36 dvss.n31 4.65
R18204 dvss.n2908 dvss.n2907 4.65
R18205 dvss.n2909 dvss.n23 4.65
R18206 dvss.n2911 dvss.n2910 4.65
R18207 dvss.n24 dvss.n18 4.65
R18208 dvss.n2918 dvss.n2917 4.65
R18209 dvss.n2919 dvss.n12 4.65
R18210 dvss.n2922 dvss.n2921 4.65
R18211 dvss.n13 dvss.n11 4.65
R18212 dvss.n7 dvss.n6 4.65
R18213 dvss.n2930 dvss.n2929 4.65
R18214 dvss.n2872 dvss.n49 4.65
R18215 dvss.n2871 dvss.n610 4.65
R18216 dvss.n2869 dvss.n2868 4.65
R18217 dvss.n612 dvss.n611 4.65
R18218 dvss.n2862 dvss.n2861 4.65
R18219 dvss.n2860 dvss.n615 4.65
R18220 dvss.n617 dvss.n616 4.65
R18221 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vss1p8 dvss.n617 4.65
R18222 dvss.n2859 dvss.n617 4.65
R18223 dvss.n2823 dvss.n2822 4.65
R18224 dvss.n629 dvss.n627 4.65
R18225 dvss.n2847 dvss.n629 4.65
R18226 dvss.n640 dvss.n630 4.65
R18227 dvss.n640 dvss.n638 4.65
R18228 dvss.n2858 dvss.n618 4.65
R18229 dvss.n2857 dvss.n2856 4.65
R18230 dvss.n2855 dvss.n619 4.65
R18231 dvss.n626 dvss.n621 4.65
R18232 dvss.n2849 dvss.n2848 4.65
R18233 dvss.n2846 dvss.n625 4.65
R18234 dvss.n2845 dvss.n2844 4.65
R18235 dvss.n637 dvss.n631 4.65
R18236 dvss.n2838 dvss.n2837 4.65
R18237 dvss.n2836 dvss.n636 4.65
R18238 dvss.n2835 dvss.n2834 4.65
R18239 dvss.n649 dvss.n644 4.65
R18240 dvss.n2828 dvss.n2827 4.65
R18241 dvss.n2826 dvss.n648 4.65
R18242 dvss.n652 dvss.n650 4.65
R18243 dvss.n2819 dvss.n2818 4.65
R18244 dvss.n2817 dvss.n651 4.65
R18245 dvss.n662 dvss.n654 4.65
R18246 dvss.n2811 dvss.n2810 4.65
R18247 dvss.n2809 dvss.n661 4.65
R18248 dvss.n2756 dvss.n2755 4.65
R18249 dvss.n2761 dvss.n2760 4.65
R18250 dvss.n2765 dvss.n2764 4.65
R18251 dvss.n2770 dvss.n2769 4.65
R18252 dvss.n2596 dvss.n2595 4.65
R18253 dvss.n2772 dvss.n2771 4.65
R18254 dvss.n2773 dvss.n2772 4.65
R18255 dvss.n2599 dvss.n2598 4.65
R18256 dvss.n2609 dvss.n2608 4.65
R18257 dvss.n2605 dvss.n2604 4.65
R18258 dvss.n3 dvss.n2 4.65
R18259 dvss.n2935 dvss.n2934 4.65
R18260 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vss1p8 dvss.n4 4.65
R18261 dvss.n2933 dvss.n4 4.65
R18262 dvss.n1718 dvss.n1717 4.5
R18263 dvss.n1370 dvss.n1279 4.5
R18264 dvss.n1833 dvss.n1832 4.5
R18265 dvss.n2336 dvss.n2335 4.5
R18266 dvss.n1988 dvss.n1897 4.5
R18267 dvss.n2451 dvss.n2450 4.5
R18268 dvss.n2453 dvss.n1895 4.5
R18269 dvss.n1837 dvss.n1277 4.5
R18270 dvss.n1105 dvss.n1104 4.5
R18271 dvss.n757 dvss.n666 4.5
R18272 dvss.n1220 dvss.n1219 4.5
R18273 dvss.n493 dvss.n492 4.5
R18274 dvss.n145 dvss.n54 4.5
R18275 dvss.n608 dvss.n607 4.5
R18276 dvss.n2877 dvss.n52 4.5
R18277 dvss.n2799 dvss.n664 4.5
R18278 dvss.n1649 dvss.n1609 4.311
R18279 dvss.n2267 dvss.n2227 4.311
R18280 dvss.n1036 dvss.n996 4.311
R18281 dvss.n424 dvss.n384 4.311
R18282 dvss.n1648 dvss.n1610 4.042
R18283 dvss.n2266 dvss.n2228 4.042
R18284 dvss.n1035 dvss.n997 4.042
R18285 dvss.n423 dvss.n385 4.042
R18286 dvss.n1523 dvss.n1508 3.931
R18287 dvss.n1502 dvss.n1487 3.931
R18288 dvss.n2141 dvss.n2126 3.931
R18289 dvss.n2120 dvss.n2105 3.931
R18290 dvss.n910 dvss.n895 3.931
R18291 dvss.n889 dvss.n874 3.931
R18292 dvss.n298 dvss.n283 3.931
R18293 dvss.n277 dvss.n262 3.931
R18294 dvss.n1609 dvss.n1556 3.84
R18295 dvss.n2227 dvss.n2174 3.84
R18296 dvss.n996 dvss.n943 3.84
R18297 dvss.n384 dvss.n331 3.84
R18298 dvss.n1645 dvss.n1644 3.772
R18299 dvss.n2263 dvss.n2262 3.772
R18300 dvss.n1032 dvss.n1031 3.772
R18301 dvss.n420 dvss.n419 3.772
R18302 dvss.n2702 dvss.n2701 3.695
R18303 dvss.n2636 dvss.n2635 3.695
R18304 dvss.n1317 dvss.n1316 3.694
R18305 dvss.n1935 dvss.n1934 3.694
R18306 dvss.n704 dvss.n703 3.694
R18307 dvss.n92 dvss.n91 3.694
R18308 dvss.n1257 dvss.n1256 3.688
R18309 dvss.n1366 dvss.n1365 3.688
R18310 dvss.n1871 dvss.n1856 3.688
R18311 dvss.n1984 dvss.n1983 3.688
R18312 dvss.n641 dvss.n640 3.688
R18313 dvss.n753 dvss.n752 3.688
R18314 dvss.n141 dvss.n140 3.688
R18315 dvss.n28 dvss.n27 3.688
R18316 dvss.n1618 dvss.n1613 3.503
R18317 dvss.n2236 dvss.n2231 3.503
R18318 dvss.n1005 dvss.n1000 3.503
R18319 dvss.n393 dvss.n388 3.503
R18320 dvss.n1639 dvss.n1620 3.233
R18321 dvss.n2257 dvss.n2238 3.233
R18322 dvss.n1026 dvss.n1007 3.233
R18323 dvss.n414 dvss.n395 3.233
R18324 dvss.n1716 dvss.n1715 3.2
R18325 dvss.n2334 dvss.n2333 3.2
R18326 dvss.n1103 dvss.n1102 3.2
R18327 dvss.n491 dvss.n490 3.2
R18328 dvss.n1380 dvss.n1379 3.033
R18329 dvss.n1998 dvss.n1997 3.033
R18330 dvss.n2457 dvss.n2456 3.033
R18331 dvss.n2527 dvss.n2526 3.033
R18332 dvss.n767 dvss.n766 3.033
R18333 dvss.n155 dvss.n154 3.033
R18334 dvss.n2881 dvss.n2880 3.033
R18335 dvss.n2803 dvss.n2802 3.033
R18336 dvss.n1484 dvss.n1483 2.98
R18337 dvss.n2102 dvss.n2101 2.98
R18338 dvss.n871 dvss.n870 2.98
R18339 dvss.n259 dvss.n258 2.98
R18340 dvss.n1638 dvss.n1623 2.964
R18341 dvss.n2256 dvss.n2241 2.964
R18342 dvss.n1025 dvss.n1010 2.964
R18343 dvss.n413 dvss.n398 2.964
R18344 dvss.n2547 dvss.n2546 2.844
R18345 dvss.n2478 dvss.n2477 2.844
R18346 dvss.n2824 dvss.n2823 2.844
R18347 dvss.n39 dvss.n37 2.844
R18348 dvss.n2796 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 2.782
R18349 dvss.n1635 dvss.n1634 2.694
R18350 dvss.n2253 dvss.n2252 2.694
R18351 dvss.n1022 dvss.n1021 2.694
R18352 dvss.n410 dvss.n409 2.694
R18353 dvss.n1691 dvss.n1690 2.56
R18354 dvss.n2309 dvss.n2308 2.56
R18355 dvss.n1078 dvss.n1077 2.56
R18356 dvss.n466 dvss.n465 2.56
R18357 dvss.n1630 dvss.n1626 2.425
R18358 dvss.n1630 dvss.n1562 2.425
R18359 dvss.n2248 dvss.n2244 2.425
R18360 dvss.n2248 dvss.n2180 2.425
R18361 dvss.n1017 dvss.n1013 2.425
R18362 dvss.n1017 dvss.n949 2.425
R18363 dvss.n405 dvss.n401 2.425
R18364 dvss.n405 dvss.n337 2.425
R18365 dvss.n2789 dvss.n2779 2.413
R18366 dvss.n2517 dvss.n2516 2.413
R18367 dvss.n2588 dvss.n2587 2.413
R18368 dvss.n2864 dvss.n2863 2.413
R18369 dvss.n2768 dvss.n2767 2.413
R18370 dvss.n1 dvss.n0 2.413
R18371 dvss.n2798 dvss.n1222 2.387
R18372 dvss.n2558 dvss.n1258 2.316
R18373 dvss.n30 dvss.n29 2.315
R18374 dvss.n643 dvss.n642 2.315
R18375 dvss.n1368 dvss.n1367 2.314
R18376 dvss.n1986 dvss.n1985 2.314
R18377 dvss.n1874 dvss.n1873 2.314
R18378 dvss.n755 dvss.n754 2.314
R18379 dvss.n143 dvss.n142 2.314
R18380 dvss.n1671 dvss.n1545 2.29
R18381 dvss.n2289 dvss.n2163 2.29
R18382 dvss.n1058 dvss.n932 2.29
R18383 dvss.n446 dvss.n320 2.29
R18384 dvss.n2879 dvss.n2878 2.273
R18385 dvss.n2525 dvss.n1838 2.273
R18386 dvss.n2801 dvss.n2800 2.273
R18387 dvss.n2455 dvss.n2454 2.273
R18388 dvss.n1831 dvss.n1830 2.247
R18389 dvss.n2449 dvss.n2448 2.247
R18390 dvss.n1218 dvss.n1217 2.247
R18391 dvss.n606 dvss.n605 2.247
R18392 dvss.n1771 dvss.n1770 2.176
R18393 dvss.n2389 dvss.n2388 2.176
R18394 dvss.n1158 dvss.n1157 2.176
R18395 dvss.n546 dvss.n545 2.176
R18396 dvss.n1634 dvss.n1626 2.155
R18397 dvss.n1656 dvss.n1562 2.155
R18398 dvss.n2252 dvss.n2244 2.155
R18399 dvss.n2274 dvss.n2180 2.155
R18400 dvss.n1021 dvss.n1013 2.155
R18401 dvss.n1043 dvss.n949 2.155
R18402 dvss.n409 dvss.n401 2.155
R18403 dvss.n431 dvss.n337 2.155
R18404 dvss.n2756 dvss.n2753 2.009
R18405 dvss dvss.n2752 1.972
R18406 dvss.n2796 dvss.n2795 1.935
R18407 dvss.n1635 dvss.n1623 1.886
R18408 dvss.n2253 dvss.n2241 1.886
R18409 dvss.n1022 dvss.n1010 1.886
R18410 dvss.n410 dvss.n398 1.886
R18411 dvss.n1690 dvss.n1688 1.684
R18412 dvss.n1672 dvss.n1671 1.684
R18413 dvss.n2308 dvss.n2306 1.684
R18414 dvss.n2290 dvss.n2289 1.684
R18415 dvss.n1077 dvss.n1075 1.684
R18416 dvss.n1059 dvss.n1058 1.684
R18417 dvss.n465 dvss.n463 1.684
R18418 dvss.n447 dvss.n446 1.684
R18419 dvss.n1711 dvss.n1710 1.646
R18420 dvss.n2329 dvss.n2328 1.646
R18421 dvss.n1098 dvss.n1097 1.646
R18422 dvss.n486 dvss.n485 1.646
R18423 dvss.n1639 dvss.n1638 1.616
R18424 dvss.n2257 dvss.n2256 1.616
R18425 dvss.n1026 dvss.n1025 1.616
R18426 dvss.n414 dvss.n413 1.616
R18427 dvss.n1483 dvss.n1468 1.594
R18428 dvss.n1743 dvss.n1468 1.594
R18429 dvss.n1744 dvss.n1743 1.594
R18430 dvss.n1745 dvss.n1744 1.594
R18431 dvss.n1745 dvss.n1442 1.594
R18432 dvss.n1753 dvss.n1442 1.594
R18433 dvss.n1765 dvss.n1764 1.594
R18434 dvss.n1766 dvss.n1765 1.594
R18435 dvss.n1766 dvss.n1428 1.594
R18436 dvss.n1773 dvss.n1428 1.594
R18437 dvss.n1770 dvss.n1420 1.594
R18438 dvss.n1783 dvss.n1420 1.594
R18439 dvss.n1791 dvss.n1418 1.594
R18440 dvss.n1787 dvss.n1418 1.594
R18441 dvss.n1787 dvss.n1384 1.594
R18442 dvss.n1825 dvss.n1384 1.594
R18443 dvss.n1826 dvss.n1825 1.594
R18444 dvss.n1826 dvss.n1382 1.594
R18445 dvss.n2101 dvss.n2086 1.594
R18446 dvss.n2361 dvss.n2086 1.594
R18447 dvss.n2362 dvss.n2361 1.594
R18448 dvss.n2363 dvss.n2362 1.594
R18449 dvss.n2363 dvss.n2060 1.594
R18450 dvss.n2371 dvss.n2060 1.594
R18451 dvss.n2383 dvss.n2382 1.594
R18452 dvss.n2384 dvss.n2383 1.594
R18453 dvss.n2384 dvss.n2046 1.594
R18454 dvss.n2391 dvss.n2046 1.594
R18455 dvss.n2388 dvss.n2038 1.594
R18456 dvss.n2401 dvss.n2038 1.594
R18457 dvss.n2409 dvss.n2036 1.594
R18458 dvss.n2405 dvss.n2036 1.594
R18459 dvss.n2405 dvss.n2002 1.594
R18460 dvss.n2443 dvss.n2002 1.594
R18461 dvss.n2444 dvss.n2443 1.594
R18462 dvss.n2444 dvss.n2000 1.594
R18463 dvss.n870 dvss.n855 1.594
R18464 dvss.n1130 dvss.n855 1.594
R18465 dvss.n1131 dvss.n1130 1.594
R18466 dvss.n1132 dvss.n1131 1.594
R18467 dvss.n1132 dvss.n829 1.594
R18468 dvss.n1140 dvss.n829 1.594
R18469 dvss.n1152 dvss.n1151 1.594
R18470 dvss.n1153 dvss.n1152 1.594
R18471 dvss.n1153 dvss.n815 1.594
R18472 dvss.n1160 dvss.n815 1.594
R18473 dvss.n1157 dvss.n807 1.594
R18474 dvss.n1170 dvss.n807 1.594
R18475 dvss.n1178 dvss.n805 1.594
R18476 dvss.n1174 dvss.n805 1.594
R18477 dvss.n1174 dvss.n771 1.594
R18478 dvss.n1212 dvss.n771 1.594
R18479 dvss.n1213 dvss.n1212 1.594
R18480 dvss.n1213 dvss.n769 1.594
R18481 dvss.n258 dvss.n243 1.594
R18482 dvss.n518 dvss.n243 1.594
R18483 dvss.n519 dvss.n518 1.594
R18484 dvss.n520 dvss.n519 1.594
R18485 dvss.n520 dvss.n217 1.594
R18486 dvss.n528 dvss.n217 1.594
R18487 dvss.n540 dvss.n539 1.594
R18488 dvss.n541 dvss.n540 1.594
R18489 dvss.n541 dvss.n203 1.594
R18490 dvss.n548 dvss.n203 1.594
R18491 dvss.n545 dvss.n195 1.594
R18492 dvss.n558 dvss.n195 1.594
R18493 dvss.n566 dvss.n193 1.594
R18494 dvss.n562 dvss.n193 1.594
R18495 dvss.n562 dvss.n159 1.594
R18496 dvss.n600 dvss.n159 1.594
R18497 dvss.n601 dvss.n600 1.594
R18498 dvss.n601 dvss.n157 1.594
R18499 dvss.n1749 dvss.n1748 1.583
R18500 dvss.n2367 dvss.n2366 1.583
R18501 dvss.n1136 dvss.n1135 1.583
R18502 dvss.n524 dvss.n523 1.583
R18503 dvss.n1538 dvss.n1528 1.546
R18504 dvss.n2156 dvss.n2146 1.546
R18505 dvss.n925 dvss.n915 1.546
R18506 dvss.n313 dvss.n303 1.546
R18507 dvss.n1509 dvss.n1507 1.505
R18508 dvss.n1488 dvss.n1486 1.505
R18509 dvss.n2127 dvss.n2125 1.505
R18510 dvss.n2106 dvss.n2104 1.505
R18511 dvss.n896 dvss.n894 1.505
R18512 dvss.n875 dvss.n873 1.505
R18513 dvss.n284 dvss.n282 1.505
R18514 dvss.n263 dvss.n261 1.505
R18515 dvss.n1516 dvss.n1515 1.45
R18516 dvss.n1495 dvss.n1494 1.45
R18517 dvss.n2134 dvss.n2133 1.45
R18518 dvss.n2113 dvss.n2112 1.45
R18519 dvss.n903 dvss.n902 1.45
R18520 dvss.n882 dvss.n881 1.45
R18521 dvss.n291 dvss.n290 1.45
R18522 dvss.n270 dvss.n269 1.45
R18523 dvss.n1704 dvss.n1539 1.447
R18524 dvss.n2322 dvss.n2157 1.447
R18525 dvss.n1091 dvss.n926 1.447
R18526 dvss.n479 dvss.n314 1.447
R18527 dvss.n2751 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VNB 1.391
R18528 dvss.n2751 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VNB 1.389
R18529 dvss.n1703 dvss.n1541 1.347
R18530 dvss.n1620 dvss.n1618 1.347
R18531 dvss.n2321 dvss.n2159 1.347
R18532 dvss.n2238 dvss.n2236 1.347
R18533 dvss.n1090 dvss.n928 1.347
R18534 dvss.n1007 dvss.n1005 1.347
R18535 dvss.n478 dvss.n316 1.347
R18536 dvss.n395 dvss.n393 1.347
R18537 dvss.n1847 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 1.25
R18538 dvss.n1700 dvss.n1699 1.247
R18539 dvss.n2318 dvss.n2317 1.247
R18540 dvss.n1087 dvss.n1086 1.247
R18541 dvss.n475 dvss.n474 1.247
R18542 dvss.n2931 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 1.153
R18543 dvss.n1697 dvss.n1696 1.147
R18544 dvss.n2315 dvss.n2314 1.147
R18545 dvss.n1084 dvss.n1083 1.147
R18546 dvss.n472 dvss.n471 1.147
R18547 dvss.n1232 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 1.133
R18548 dvss.n1371 dvss.n1284 1.129
R18549 dvss.n1989 dvss.n1902 1.129
R18550 dvss.n758 dvss.n671 1.129
R18551 dvss.n146 dvss.n59 1.129
R18552 dvss.n1764 dvss.n1430 1.113
R18553 dvss.n2382 dvss.n2048 1.113
R18554 dvss.n1151 dvss.n817 1.113
R18555 dvss.n539 dvss.n205 1.113
R18556 dvss.n1834 dvss.n1833 1.106
R18557 dvss.n2452 dvss.n2451 1.106
R18558 dvss.n1221 dvss.n1220 1.106
R18559 dvss.n609 dvss.n608 1.106
R18560 dvss.n1691 dvss.n1548 1.077
R18561 dvss.n1644 dvss.n1613 1.077
R18562 dvss.n2309 dvss.n2166 1.077
R18563 dvss.n2262 dvss.n2231 1.077
R18564 dvss.n1078 dvss.n935 1.077
R18565 dvss.n1031 dvss.n1000 1.077
R18566 dvss.n466 dvss.n323 1.077
R18567 dvss.n419 dvss.n388 1.077
R18568 dvss.n1694 dvss.n1544 0.973
R18569 dvss.n2312 dvss.n2162 0.973
R18570 dvss.n1081 dvss.n931 0.973
R18571 dvss.n469 dvss.n319 0.973
R18572 dvss.n1378 dvss.n1280 0.903
R18573 dvss.n1996 dvss.n1898 0.903
R18574 dvss.n2509 dvss.n1849 0.903
R18575 dvss.n2528 dvss.n1276 0.903
R18576 dvss.n765 dvss.n667 0.903
R18577 dvss.n153 dvss.n55 0.903
R18578 dvss.n2882 dvss.n51 0.903
R18579 dvss.n623 dvss.n620 0.903
R18580 dvss.n2704 dvss.n2703 0.903
R18581 dvss.n2638 dvss.n2637 0.903
R18582 dvss.n2459 dvss.n2458 0.903
R18583 dvss.n2579 dvss.n1233 0.903
R18584 dvss.n2928 dvss.n8 0.903
R18585 dvss.n2805 dvss.n2804 0.903
R18586 dvss.n1645 dvss.n1610 0.808
R18587 dvss.n2263 dvss.n2228 0.808
R18588 dvss.n1032 dvss.n997 0.808
R18589 dvss.n420 dvss.n385 0.808
R18590 dvss.n1835 dvss.n1275 0.752
R18591 dvss.n1522 dvss.n1521 0.752
R18592 dvss.n1513 dvss.n1510 0.752
R18593 dvss.n1501 dvss.n1500 0.752
R18594 dvss.n1492 dvss.n1489 0.752
R18595 dvss.n2461 dvss.n2460 0.752
R18596 dvss.n2140 dvss.n2139 0.752
R18597 dvss.n2131 dvss.n2128 0.752
R18598 dvss.n2119 dvss.n2118 0.752
R18599 dvss.n2110 dvss.n2107 0.752
R18600 dvss.n2807 dvss.n2806 0.752
R18601 dvss.n909 dvss.n908 0.752
R18602 dvss.n900 dvss.n897 0.752
R18603 dvss.n888 dvss.n887 0.752
R18604 dvss.n879 dvss.n876 0.752
R18605 dvss.n297 dvss.n296 0.752
R18606 dvss.n288 dvss.n285 0.752
R18607 dvss.n276 dvss.n275 0.752
R18608 dvss.n267 dvss.n264 0.752
R18609 dvss.n2875 dvss.n2874 0.752
R18610 dvss.n1696 dvss.n1694 0.648
R18611 dvss.n2314 dvss.n2312 0.648
R18612 dvss.n1083 dvss.n1081 0.648
R18613 dvss.n471 dvss.n469 0.648
R18614 dvss.n1688 dvss.n1545 0.606
R18615 dvss.n2306 dvss.n2163 0.606
R18616 dvss.n1075 dvss.n932 0.606
R18617 dvss.n463 dvss.n320 0.606
R18618 dvss.n1699 dvss.n1697 0.548
R18619 dvss.n2317 dvss.n2315 0.548
R18620 dvss.n1086 dvss.n1084 0.548
R18621 dvss.n474 dvss.n472 0.548
R18622 dvss.n1649 dvss.n1648 0.538
R18623 dvss.n2267 dvss.n2266 0.538
R18624 dvss.n1036 dvss.n1035 0.538
R18625 dvss.n424 dvss.n423 0.538
R18626 dvss.n2708 dvss.n2701 0.525
R18627 dvss.n2642 dvss.n2635 0.525
R18628 dvss.n1318 dvss.n1317 0.501
R18629 dvss.n1936 dvss.n1935 0.501
R18630 dvss.n705 dvss.n704 0.501
R18631 dvss.n93 dvss.n92 0.501
R18632 dvss.n1700 dvss.n1541 0.449
R18633 dvss.n2318 dvss.n2159 0.449
R18634 dvss.n1087 dvss.n928 0.449
R18635 dvss.n475 dvss.n316 0.449
R18636 dvss.n1704 dvss.n1703 0.349
R18637 dvss.n1548 dvss.n1547 0.349
R18638 dvss.n2322 dvss.n2321 0.349
R18639 dvss.n2166 dvss.n2165 0.349
R18640 dvss.n1091 dvss.n1090 0.349
R18641 dvss.n935 dvss.n934 0.349
R18642 dvss.n479 dvss.n478 0.349
R18643 dvss.n323 dvss.n322 0.349
R18644 dvss.n1713 dvss.n1525 0.336
R18645 dvss.n1715 dvss.n1504 0.336
R18646 dvss.n2331 dvss.n2143 0.336
R18647 dvss.n2333 dvss.n2122 0.336
R18648 dvss.n1100 dvss.n912 0.336
R18649 dvss.n1102 dvss.n891 0.336
R18650 dvss.n488 dvss.n300 0.336
R18651 dvss.n490 dvss.n279 0.336
R18652 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB dvss.n2798 0.315
R18653 dvss.n2752 comparator_top_0.DVSS 0.299
R18654 dvss.n1784 dvss.n1417 0.281
R18655 dvss.n2402 dvss.n2035 0.281
R18656 dvss.n1171 dvss.n804 0.281
R18657 dvss.n559 dvss.n192 0.281
R18658 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.vss3p3 dvss.n1829 0.27
R18659 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.vss3p3 dvss.n2447 0.27
R18660 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.vss3p3 dvss.n1216 0.27
R18661 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.vss3p3 dvss.n604 0.27
R18662 dvss.n2753 dvss.n2610 0.256
R18663 dvss.n1539 dvss.n1538 0.249
R18664 dvss.n2157 dvss.n2156 0.249
R18665 dvss.n926 dvss.n925 0.249
R18666 dvss.n314 dvss.n313 0.249
R18667 dvss.n1750 dvss.n1466 0.234
R18668 dvss.n2368 dvss.n2084 0.234
R18669 dvss.n1137 dvss.n853 0.234
R18670 dvss.n525 dvss.n241 0.234
R18671 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB EF_AMUX21m_1.vss 0.224
R18672 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB EF_AMUX21m_2.vss 0.22
R18673 dvss.n2797 dvss.n2594 0.213
R18674 dvss.n2797 dvss.n2796 0.21
R18675 dvss.n1713 dvss.n1712 0.197
R18676 dvss.n2331 dvss.n2330 0.197
R18677 dvss.n1100 dvss.n1099 0.197
R18678 dvss.n488 dvss.n487 0.197
R18679 dvss.n1715 dvss.n1714 0.196
R18680 dvss.n2333 dvss.n2332 0.196
R18681 dvss.n1102 dvss.n1101 0.196
R18682 dvss.n490 dvss.n489 0.196
R18683 dvss.n48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 0.186
R18684 dvss.n2751 comparator_top_0.DVSS 0.177
R18685 dvss.n2680 dvss.n2679 0.151
R18686 dvss.n2748 dvss.n2747 0.151
R18687 dvss.n2747 dvss.n2687 0.151
R18688 dvss.n2747 dvss.n2688 0.151
R18689 dvss.n2747 dvss.n2689 0.151
R18690 dvss.n2681 dvss.n2680 0.151
R18691 dvss.n1710 dvss.n1528 0.149
R18692 dvss.n2328 dvss.n2146 0.149
R18693 dvss.n1097 dvss.n915 0.149
R18694 dvss.n485 dvss.n303 0.149
R18695 dvss.n1832 EF_AMUX21m_1.array_1ls_1tgm_0.vss 0.146
R18696 dvss.n2450 EF_AMUX21m_1.array_1ls_1tgm_1.vss 0.146
R18697 dvss.n1219 EF_AMUX21m_2.array_1ls_1tgm_1.vss 0.146
R18698 dvss.n607 EF_AMUX21m_2.array_1ls_1tgm_0.vss 0.146
R18699 EF_AMUX21m_1.vss dvss.n2524 0.145
R18700 EF_AMUX21m_2.vss dvss.n2871 0.142
R18701 dvss.n1773 dvss.n1772 0.138
R18702 dvss.n2391 dvss.n2390 0.138
R18703 dvss.n1160 dvss.n1159 0.138
R18704 dvss.n548 dvss.n547 0.138
R18705 EF_AMUX21m_1.array_1ls_1tgm_0.vss EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.vss3p3 0.137
R18706 EF_AMUX21m_1.array_1ls_1tgm_1.vss EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.vss3p3 0.137
R18707 EF_AMUX21m_2.array_1ls_1tgm_1.vss EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.vss3p3 0.137
R18708 EF_AMUX21m_2.array_1ls_1tgm_0.vss EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.vss3p3 0.137
R18709 dvss.n2752 dvss.n2751 0.126
R18710 dvss.n1828 dvss.n1382 0.093
R18711 dvss.n2446 dvss.n2000 0.093
R18712 dvss.n1215 dvss.n769 0.093
R18713 dvss.n603 dvss.n157 0.093
R18714 dvss.n1712 dvss.n1526 0.092
R18715 dvss.n1542 dvss.n1526 0.092
R18716 dvss.n1702 dvss.n1542 0.092
R18717 dvss.n1702 dvss.n1701 0.092
R18718 dvss.n1701 dvss.n1543 0.092
R18719 dvss.n1693 dvss.n1543 0.092
R18720 dvss.n1693 dvss.n1692 0.092
R18721 dvss.n1647 dvss.n1505 0.092
R18722 dvss.n1647 dvss.n1646 0.092
R18723 dvss.n1646 dvss.n1611 0.092
R18724 dvss.n1624 dvss.n1611 0.092
R18725 dvss.n1637 dvss.n1624 0.092
R18726 dvss.n1637 dvss.n1636 0.092
R18727 dvss.n1636 dvss.n1625 0.092
R18728 dvss.n2330 dvss.n2144 0.092
R18729 dvss.n2160 dvss.n2144 0.092
R18730 dvss.n2320 dvss.n2160 0.092
R18731 dvss.n2320 dvss.n2319 0.092
R18732 dvss.n2319 dvss.n2161 0.092
R18733 dvss.n2311 dvss.n2161 0.092
R18734 dvss.n2311 dvss.n2310 0.092
R18735 dvss.n2265 dvss.n2123 0.092
R18736 dvss.n2265 dvss.n2264 0.092
R18737 dvss.n2264 dvss.n2229 0.092
R18738 dvss.n2242 dvss.n2229 0.092
R18739 dvss.n2255 dvss.n2242 0.092
R18740 dvss.n2255 dvss.n2254 0.092
R18741 dvss.n2254 dvss.n2243 0.092
R18742 dvss.n1099 dvss.n913 0.092
R18743 dvss.n929 dvss.n913 0.092
R18744 dvss.n1089 dvss.n929 0.092
R18745 dvss.n1089 dvss.n1088 0.092
R18746 dvss.n1088 dvss.n930 0.092
R18747 dvss.n1080 dvss.n930 0.092
R18748 dvss.n1080 dvss.n1079 0.092
R18749 dvss.n1034 dvss.n892 0.092
R18750 dvss.n1034 dvss.n1033 0.092
R18751 dvss.n1033 dvss.n998 0.092
R18752 dvss.n1011 dvss.n998 0.092
R18753 dvss.n1024 dvss.n1011 0.092
R18754 dvss.n1024 dvss.n1023 0.092
R18755 dvss.n1023 dvss.n1012 0.092
R18756 dvss.n487 dvss.n301 0.092
R18757 dvss.n317 dvss.n301 0.092
R18758 dvss.n477 dvss.n317 0.092
R18759 dvss.n477 dvss.n476 0.092
R18760 dvss.n476 dvss.n318 0.092
R18761 dvss.n468 dvss.n318 0.092
R18762 dvss.n468 dvss.n467 0.092
R18763 dvss.n422 dvss.n280 0.092
R18764 dvss.n422 dvss.n421 0.092
R18765 dvss.n421 dvss.n386 0.092
R18766 dvss.n399 dvss.n386 0.092
R18767 dvss.n412 dvss.n399 0.092
R18768 dvss.n412 dvss.n411 0.092
R18769 dvss.n411 dvss.n400 0.092
R18770 dvss.n1714 dvss.n1713 0.086
R18771 dvss.n2332 dvss.n2331 0.086
R18772 dvss.n1101 dvss.n1100 0.086
R18773 dvss.n489 dvss.n488 0.086
R18774 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND dvss.n2511 0.084
R18775 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND dvss.n2858 0.083
R18776 dvss.n1751 dvss.n1748 0.081
R18777 dvss.n2369 dvss.n2366 0.081
R18778 dvss.n1138 dvss.n1135 0.081
R18779 dvss.n526 dvss.n523 0.081
R18780 dvss.n1512 dvss.n1511 0.078
R18781 dvss.n1491 dvss.n1490 0.078
R18782 dvss.n2130 dvss.n2129 0.078
R18783 dvss.n2109 dvss.n2108 0.078
R18784 dvss.n899 dvss.n898 0.078
R18785 dvss.n878 dvss.n877 0.078
R18786 dvss.n287 dvss.n286 0.078
R18787 dvss.n266 dvss.n265 0.078
R18788 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND dvss.n2932 0.078
R18789 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND dvss.n2582 0.077
R18790 dvss.n1547 dvss.n1544 0.074
R18791 dvss.n2165 dvss.n2162 0.074
R18792 dvss.n934 dvss.n931 0.074
R18793 dvss.n322 dvss.n319 0.074
R18794 dvss.n2781 dvss.n2777 0.073
R18795 dvss.n2765 dvss.n2761 0.071
R18796 dvss.n1752 dvss.n1751 0.063
R18797 dvss.n1785 dvss.n1419 0.063
R18798 dvss.n1790 dvss.n1785 0.063
R18799 dvss.n2370 dvss.n2369 0.063
R18800 dvss.n2403 dvss.n2037 0.063
R18801 dvss.n2408 dvss.n2403 0.063
R18802 dvss.n2777 dvss.n2774 0.063
R18803 dvss.n1139 dvss.n1138 0.063
R18804 dvss.n1172 dvss.n806 0.063
R18805 dvss.n1177 dvss.n1172 0.063
R18806 dvss.n527 dvss.n526 0.063
R18807 dvss.n560 dvss.n194 0.063
R18808 dvss.n565 dvss.n560 0.063
R18809 dvss.n2505 dvss.n1853 0.061
R18810 dvss.n2505 dvss.n2504 0.061
R18811 dvss.n2500 dvss.n1857 0.061
R18812 dvss.n2491 dvss.n2490 0.061
R18813 dvss.n2481 dvss.n1880 0.061
R18814 dvss.n2481 dvss.n2480 0.061
R18815 dvss.n2473 dvss.n1882 0.061
R18816 dvss.n1893 dvss.n1882 0.061
R18817 dvss.n2464 dvss.n2463 0.061
R18818 dvss.n2761 dvss.n2757 0.061
R18819 dvss.n1323 dvss.n1322 0.06
R18820 dvss.n1323 dvss.n1303 0.06
R18821 dvss.n1331 dvss.n1303 0.06
R18822 dvss.n1332 dvss.n1331 0.06
R18823 dvss.n1333 dvss.n1332 0.06
R18824 dvss.n1333 dvss.n1297 0.06
R18825 dvss.n1342 dvss.n1297 0.06
R18826 dvss.n1346 dvss.n1290 0.06
R18827 dvss.n1355 dvss.n1354 0.06
R18828 dvss.n1355 dvss.n1285 0.06
R18829 dvss.n1374 dvss.n1369 0.06
R18830 dvss.n1941 dvss.n1940 0.06
R18831 dvss.n1941 dvss.n1921 0.06
R18832 dvss.n1949 dvss.n1921 0.06
R18833 dvss.n1950 dvss.n1949 0.06
R18834 dvss.n1951 dvss.n1950 0.06
R18835 dvss.n1951 dvss.n1915 0.06
R18836 dvss.n1960 dvss.n1915 0.06
R18837 dvss.n1964 dvss.n1908 0.06
R18838 dvss.n1973 dvss.n1972 0.06
R18839 dvss.n1973 dvss.n1903 0.06
R18840 dvss.n1992 dvss.n1987 0.06
R18841 dvss.n2490 dvss.n2489 0.06
R18842 dvss.n710 dvss.n709 0.06
R18843 dvss.n710 dvss.n690 0.06
R18844 dvss.n718 dvss.n690 0.06
R18845 dvss.n719 dvss.n718 0.06
R18846 dvss.n720 dvss.n719 0.06
R18847 dvss.n720 dvss.n684 0.06
R18848 dvss.n729 dvss.n684 0.06
R18849 dvss.n733 dvss.n677 0.06
R18850 dvss.n742 dvss.n741 0.06
R18851 dvss.n742 dvss.n672 0.06
R18852 dvss.n761 dvss.n756 0.06
R18853 dvss.n98 dvss.n97 0.06
R18854 dvss.n98 dvss.n78 0.06
R18855 dvss.n106 dvss.n78 0.06
R18856 dvss.n107 dvss.n106 0.06
R18857 dvss.n108 dvss.n107 0.06
R18858 dvss.n108 dvss.n72 0.06
R18859 dvss.n117 dvss.n72 0.06
R18860 dvss.n121 dvss.n65 0.06
R18861 dvss.n130 dvss.n129 0.06
R18862 dvss.n130 dvss.n60 0.06
R18863 dvss.n149 dvss.n144 0.06
R18864 dvss.n2463 dvss.n2462 0.059
R18865 dvss.n1364 dvss.n1290 0.058
R18866 dvss.n1374 dvss.n1373 0.058
R18867 dvss.n1982 dvss.n1908 0.058
R18868 dvss.n1992 dvss.n1991 0.058
R18869 dvss.n751 dvss.n677 0.058
R18870 dvss.n761 dvss.n760 0.058
R18871 dvss.n139 dvss.n65 0.058
R18872 dvss.n149 dvss.n148 0.058
R18873 dvss.n2858 dvss.n2857 0.057
R18874 dvss.n2857 dvss.n619 0.057
R18875 dvss.n626 dvss.n619 0.057
R18876 dvss.n2846 dvss.n2845 0.057
R18877 dvss.n2837 dvss.n2836 0.057
R18878 dvss.n2836 dvss.n2835 0.057
R18879 dvss.n2827 dvss.n649 0.057
R18880 dvss.n2827 dvss.n2826 0.057
R18881 dvss.n2819 dvss.n651 0.057
R18882 dvss.n662 dvss.n651 0.057
R18883 dvss.n2810 dvss.n2809 0.057
R18884 dvss.n1322 dvss.n1321 0.056
R18885 dvss.n1940 dvss.n1939 0.056
R18886 dvss.n709 dvss.n708 0.056
R18887 dvss.n97 dvss.n96 0.056
R18888 dvss.n2930 dvss.n6 0.056
R18889 dvss.n13 dvss.n6 0.056
R18890 dvss.n2919 dvss.n2918 0.056
R18891 dvss.n2910 dvss.n2909 0.056
R18892 dvss.n2900 dvss.n36 0.056
R18893 dvss.n2900 dvss.n2899 0.056
R18894 dvss.n2889 dvss.n47 0.056
R18895 dvss.n2889 dvss.n2888 0.056
R18896 dvss.n2809 dvss.n2808 0.056
R18897 dvss.n1240 dvss.n1235 0.055
R18898 dvss.n1241 dvss.n1240 0.055
R18899 dvss.n2570 dvss.n2569 0.055
R18900 dvss.n2561 dvss.n2560 0.055
R18901 dvss.n2557 dvss.n1259 0.055
R18902 dvss.n2549 dvss.n1259 0.055
R18903 dvss.n2542 dvss.n1267 0.055
R18904 dvss.n2534 dvss.n1267 0.055
R18905 dvss.n2533 dvss.n2532 0.055
R18906 dvss.n2909 dvss.n2908 0.055
R18907 dvss.n1717 dvss.n1481 0.054
R18908 dvss.n2335 dvss.n2099 0.054
R18909 dvss.n2560 dvss.n2559 0.054
R18910 dvss.n2532 dvss.n1274 0.054
R18911 dvss.n1104 dvss.n868 0.054
R18912 dvss.n492 dvss.n256 0.054
R18913 dvss.n2873 dvss.n2872 0.054
R18914 dvss.n1484 dvss.n1482 0.052
R18915 dvss.n2102 dvss.n2100 0.052
R18916 dvss.n871 dvss.n869 0.052
R18917 dvss.n259 dvss.n257 0.052
R18918 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vss1p8 dvss.n1893 0.047
R18919 dvss.n2501 dvss.n2500 0.046
R18920 dvss.n2709 dvss.n2708 0.045
R18921 dvss.n2710 dvss.n2709 0.045
R18922 dvss.n2710 dvss.n2695 0.045
R18923 dvss.n2718 dvss.n2695 0.045
R18924 dvss.n2719 dvss.n2718 0.045
R18925 dvss.n2743 dvss.n2719 0.045
R18926 dvss.n2743 dvss.n2742 0.045
R18927 dvss.n2742 dvss.n2741 0.045
R18928 dvss.n2737 dvss.n2736 0.045
R18929 dvss.n2736 dvss.n2735 0.045
R18930 dvss.n2750 dvss.n2684 0.045
R18931 dvss.n2643 dvss.n2642 0.045
R18932 dvss.n2644 dvss.n2643 0.045
R18933 dvss.n2644 dvss.n2627 0.045
R18934 dvss.n2654 dvss.n2627 0.045
R18935 dvss.n2660 dvss.n2658 0.045
R18936 dvss.n2660 dvss.n2659 0.045
R18937 dvss.n2670 dvss.n2669 0.045
R18938 dvss.n2676 dvss.n2670 0.045
R18939 dvss.n2683 dvss.n2611 0.045
R18940 dvss.n1853 dvss.n1847 0.045
R18941 dvss.n1870 dvss.n1857 0.045
R18942 dvss.n2476 dvss.n2474 0.045
R18943 dvss.n2872 dvss.n48 0.044
R18944 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vss1p8 dvss.n662 0.044
R18945 dvss.n1771 dvss.n1769 0.043
R18946 dvss.n2389 dvss.n2387 0.043
R18947 dvss.n1158 dvss.n1156 0.043
R18948 dvss.n546 dvss.n544 0.043
R18949 dvss.n2782 dvss.n2781 0.043
R18950 dvss.n2888 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vss1p8 0.043
R18951 dvss.n2847 dvss.n2846 0.043
R18952 dvss.n2822 dvss.n2820 0.043
R18953 dvss.n1343 dvss.n1342 0.042
R18954 dvss.n1363 dvss.n1288 0.042
R18955 dvss.n1961 dvss.n1960 0.042
R18956 dvss.n1981 dvss.n1906 0.042
R18957 dvss.n2479 dvss.n1881 0.042
R18958 dvss.n2571 dvss.n2570 0.042
R18959 dvss.n2534 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vss1p8 0.042
R18960 dvss.n730 dvss.n729 0.042
R18961 dvss.n750 dvss.n675 0.042
R18962 dvss.n118 dvss.n117 0.042
R18963 dvss.n138 dvss.n63 0.042
R18964 dvss.n2931 dvss.n2930 0.042
R18965 dvss.n2920 dvss.n2919 0.042
R18966 dvss.n46 dvss.n40 0.042
R18967 dvss.n2845 dvss.n630 0.042
R18968 dvss.n2771 dvss.n2765 0.042
R18969 dvss.n2655 dvss.n2654 0.041
R18970 dvss.n1318 dvss.n1309 0.041
R18971 dvss.n1936 dvss.n1927 0.041
R18972 dvss.n1235 dvss.n1232 0.041
R18973 dvss.n2545 dvss.n2543 0.041
R18974 dvss.n2784 EF_AMUX21m_1.invm_0.vss3p3 0.041
R18975 dvss.n705 dvss.n696 0.041
R18976 dvss.n93 dvss.n84 0.041
R18977 dvss.n2918 dvss.n17 0.041
R18978 dvss.n2569 dvss.n1245 0.04
R18979 dvss.n2766 EF_AMUX21m_2.invm_0.vss3p3 0.04
R18980 dvss.n2825 dvss.n650 0.039
R18981 dvss.n2548 dvss.n1266 0.038
R18982 dvss.n2898 dvss.n2897 0.038
R18983 dvss.n1880 dvss.n1874 0.038
R18984 dvss.n649 dvss.n643 0.037
R18985 dvss.n2454 dvss.n2453 0.037
R18986 dvss.n36 dvss.n30 0.036
R18987 dvss.n1370 dvss.n1278 0.035
R18988 dvss.n1988 dvss.n1896 0.035
R18989 dvss.n757 dvss.n665 0.035
R18990 dvss.n145 dvss.n53 0.035
R18991 dvss.n1368 dvss.n1285 0.035
R18992 dvss.n1986 dvss.n1903 0.035
R18993 dvss.n755 dvss.n672 0.035
R18994 dvss.n143 dvss.n60 0.035
R18995 dvss.n2558 dvss.n2557 0.035
R18996 dvss.n1838 dvss.n1837 0.034
R18997 dvss.n2800 dvss.n2799 0.034
R18998 dvss.n2878 dvss.n2877 0.033
R18999 dvss.n1346 dvss.n1345 0.032
R19000 dvss.n1964 dvss.n1963 0.032
R19001 dvss.n733 dvss.n732 0.032
R19002 dvss.n121 dvss.n120 0.032
R19003 dvss.n2503 dvss.n1854 0.031
R19004 dvss.n2491 dvss.n1872 0.031
R19005 dvss.n1430 dvss.n1429 0.031
R19006 dvss.n2048 dvss.n2047 0.031
R19007 dvss.n817 dvss.n816 0.031
R19008 dvss.n205 dvss.n204 0.031
R19009 dvss.n2735 dvss.n2725 0.029
R19010 dvss.n2657 dvss.n2626 0.029
R19011 dvss.n2676 dvss.n2675 0.029
R19012 dvss.n2504 dvss.n2503 0.029
R19013 dvss.n1872 dvss.n1868 0.029
R19014 dvss.n2783 dvss.n2782 0.029
R19015 dvss.n2786 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 0.029
R19016 dvss.n2848 dvss.n627 0.029
R19017 dvss.n2837 dvss.n638 0.029
R19018 dvss.n2771 dvss.n2770 0.029
R19019 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND dvss.n2773 0.029
R19020 dvss.n1717 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.vss 0.028
R19021 dvss.n2335 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.vss 0.028
R19022 dvss.n2572 dvss.n1242 0.028
R19023 dvss.n2561 dvss.n1253 0.028
R19024 dvss.n1104 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.vss 0.028
R19025 dvss.n492 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.vss 0.028
R19026 dvss.n2921 dvss.n14 0.028
R19027 dvss.n2910 dvss.n25 0.028
R19028 dvss.n627 dvss.n626 0.028
R19029 dvss.n638 dvss.n637 0.028
R19030 dvss.n2728 dvss.n2684 0.027
R19031 dvss.n2673 dvss.n2611 0.027
R19032 dvss.n1345 dvss.n1344 0.027
R19033 dvss.n1963 dvss.n1962 0.027
R19034 dvss.n1242 dvss.n1241 0.027
R19035 dvss.n1253 dvss.n1252 0.027
R19036 dvss.n732 dvss.n731 0.027
R19037 dvss.n120 dvss.n119 0.027
R19038 dvss.n14 dvss.n13 0.027
R19039 dvss.n25 dvss.n24 0.027
R19040 dvss.n2741 dvss.n2722 0.027
R19041 dvss.n2784 dvss.n2783 0.025
R19042 dvss.n1369 dvss.n1368 0.025
R19043 dvss.n1987 dvss.n1986 0.025
R19044 dvss.n756 dvss.n755 0.025
R19045 dvss.n144 dvss.n143 0.025
R19046 dvss.n2659 dvss.n2621 0.024
R19047 dvss.n2522 dvss.n1840 0.024
R19048 dvss.n2869 dvss.n611 0.024
R19049 dvss.n2770 dvss.n2766 0.024
R19050 dvss.n2593 dvss.n1224 0.023
R19051 dvss.n2609 dvss.n2605 0.023
R19052 dvss.n1830 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VGND 0.023
R19053 dvss.n2448 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VGND 0.023
R19054 dvss.n1217 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VGND 0.023
R19055 dvss.n605 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VGND 0.023
R19056 dvss.n2489 dvss.n1874 0.023
R19057 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VNB dvss.n2750 0.022
R19058 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.VNB dvss.n2683 0.022
R19059 dvss.n1514 dvss.n1512 0.022
R19060 dvss.n1493 dvss.n1491 0.022
R19061 dvss.n2132 dvss.n2130 0.022
R19062 dvss.n2111 dvss.n2109 0.022
R19063 dvss.n901 dvss.n899 0.022
R19064 dvss.n880 dvss.n878 0.022
R19065 dvss.n289 dvss.n287 0.022
R19066 dvss.n268 dvss.n266 0.022
R19067 dvss.n2455 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 0.022
R19068 dvss.n2835 dvss.n643 0.022
R19069 dvss.n2669 dvss.n2621 0.021
R19070 dvss.n2908 dvss.n30 0.021
R19071 dvss.n2559 dvss.n2558 0.021
R19072 dvss.n2801 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 0.021
R19073 dvss.n2525 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 0.02
R19074 dvss.n2879 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.VNB 0.02
R19075 dvss.n2523 dvss.n2522 0.02
R19076 dvss.n2870 dvss.n2869 0.02
R19077 dvss.n1828 dvss.n1827 0.019
R19078 dvss.n2446 dvss.n2445 0.019
R19079 dvss.n1215 dvss.n1214 0.019
R19080 dvss.n603 dvss.n602 0.019
R19081 dvss.n1772 dvss.n1768 0.019
R19082 dvss.n2390 dvss.n2386 0.019
R19083 dvss.n1159 dvss.n1155 0.019
R19084 dvss.n547 dvss.n543 0.019
R19085 dvss.n1525 dvss.n1506 0.019
R19086 dvss.n1504 dvss.n1485 0.019
R19087 dvss.n2143 dvss.n2124 0.019
R19088 dvss.n2122 dvss.n2103 0.019
R19089 dvss.n2480 dvss.n2479 0.019
R19090 dvss.n912 dvss.n893 0.019
R19091 dvss.n891 dvss.n872 0.019
R19092 dvss.n300 dvss.n281 0.019
R19093 dvss.n279 dvss.n260 0.019
R19094 dvss.n1831 dvss.n1278 0.018
R19095 dvss.n2449 dvss.n1896 0.018
R19096 dvss.n1218 dvss.n665 0.018
R19097 dvss.n606 dvss.n53 0.018
R19098 dvss.n1482 dvss.n1469 0.018
R19099 dvss.n1469 dvss.n1467 0.018
R19100 dvss.n1746 dvss.n1467 0.018
R19101 dvss.n1747 dvss.n1746 0.018
R19102 dvss.n1752 dvss.n1747 0.018
R19103 dvss.n1767 dvss.n1429 0.018
R19104 dvss.n1768 dvss.n1767 0.018
R19105 dvss.n1769 dvss.n1419 0.018
R19106 dvss.n1790 dvss.n1789 0.018
R19107 dvss.n1789 dvss.n1788 0.018
R19108 dvss.n1788 dvss.n1786 0.018
R19109 dvss.n1786 dvss.n1383 0.018
R19110 dvss.n1827 dvss.n1383 0.018
R19111 dvss.n2100 dvss.n2087 0.018
R19112 dvss.n2087 dvss.n2085 0.018
R19113 dvss.n2364 dvss.n2085 0.018
R19114 dvss.n2365 dvss.n2364 0.018
R19115 dvss.n2370 dvss.n2365 0.018
R19116 dvss.n2385 dvss.n2047 0.018
R19117 dvss.n2386 dvss.n2385 0.018
R19118 dvss.n2387 dvss.n2037 0.018
R19119 dvss.n2408 dvss.n2407 0.018
R19120 dvss.n2407 dvss.n2406 0.018
R19121 dvss.n2406 dvss.n2404 0.018
R19122 dvss.n2404 dvss.n2001 0.018
R19123 dvss.n2445 dvss.n2001 0.018
R19124 dvss.n869 dvss.n856 0.018
R19125 dvss.n856 dvss.n854 0.018
R19126 dvss.n1133 dvss.n854 0.018
R19127 dvss.n1134 dvss.n1133 0.018
R19128 dvss.n1139 dvss.n1134 0.018
R19129 dvss.n1154 dvss.n816 0.018
R19130 dvss.n1155 dvss.n1154 0.018
R19131 dvss.n1156 dvss.n806 0.018
R19132 dvss.n1177 dvss.n1176 0.018
R19133 dvss.n1176 dvss.n1175 0.018
R19134 dvss.n1175 dvss.n1173 0.018
R19135 dvss.n1173 dvss.n770 0.018
R19136 dvss.n1214 dvss.n770 0.018
R19137 dvss.n257 dvss.n244 0.018
R19138 dvss.n244 dvss.n242 0.018
R19139 dvss.n521 dvss.n242 0.018
R19140 dvss.n522 dvss.n521 0.018
R19141 dvss.n527 dvss.n522 0.018
R19142 dvss.n542 dvss.n204 0.018
R19143 dvss.n543 dvss.n542 0.018
R19144 dvss.n544 dvss.n194 0.018
R19145 dvss.n565 dvss.n564 0.018
R19146 dvss.n564 dvss.n563 0.018
R19147 dvss.n563 dvss.n561 0.018
R19148 dvss.n561 dvss.n158 0.018
R19149 dvss.n602 dvss.n158 0.018
R19150 dvss.n2826 dvss.n2825 0.018
R19151 dvss.n2729 dvss.n2728 0.017
R19152 dvss.n2674 dvss.n2673 0.017
R19153 dvss.n1344 dvss.n1343 0.017
R19154 dvss.n1354 dvss.n1288 0.017
R19155 dvss.n1833 dvss.n1380 0.017
R19156 dvss.n1832 dvss.n1831 0.017
R19157 dvss.n1962 dvss.n1961 0.017
R19158 dvss.n1972 dvss.n1906 0.017
R19159 dvss.n2451 dvss.n1998 0.017
R19160 dvss.n2450 dvss.n2449 0.017
R19161 dvss.n2549 dvss.n2548 0.017
R19162 dvss.n731 dvss.n730 0.017
R19163 dvss.n741 dvss.n675 0.017
R19164 dvss.n1220 dvss.n767 0.017
R19165 dvss.n1219 dvss.n1218 0.017
R19166 dvss.n119 dvss.n118 0.017
R19167 dvss.n129 dvss.n63 0.017
R19168 dvss.n608 dvss.n155 0.017
R19169 dvss.n607 dvss.n606 0.017
R19170 dvss.n2899 dvss.n2898 0.017
R19171 dvss.n2737 dvss.n2722 0.017
R19172 dvss.n1829 dvss.n1828 0.017
R19173 dvss.n2447 dvss.n2446 0.017
R19174 dvss.n1216 dvss.n1215 0.017
R19175 dvss.n604 dvss.n603 0.017
R19176 dvss.n1718 dvss.n1484 0.017
R19177 dvss.n2336 dvss.n2102 0.017
R19178 dvss.n1105 dvss.n871 0.017
R19179 dvss.n493 dvss.n259 0.017
R19180 dvss.n2675 dvss.n2674 0.016
R19181 dvss.n2729 dvss.n2725 0.015
R19182 dvss.n2658 dvss.n2657 0.015
R19183 dvss.n1870 dvss.n1868 0.015
R19184 dvss.n2456 dvss.n2452 0.015
R19185 dvss.n637 dvss.n630 0.015
R19186 dvss.n2802 dvss.n1221 0.015
R19187 dvss.n2501 dvss.n1854 0.014
R19188 dvss.n2464 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vss1p8 0.014
R19189 dvss.n2511 dvss.n1847 0.014
R19190 dvss.n1845 dvss.n1840 0.014
R19191 dvss.n1252 dvss.n1245 0.014
R19192 dvss.n2526 dvss.n1834 0.014
R19193 dvss.n24 dvss.n17 0.014
R19194 dvss.n2880 dvss.n609 0.014
R19195 dvss.n616 dvss.n611 0.014
R19196 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vss1p8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.vss3p3 0.013
R19197 dvss.n2572 dvss.n2571 0.013
R19198 dvss.n2582 dvss.n1232 0.013
R19199 dvss.n2594 dvss.n1223 0.013
R19200 dvss.n1230 dvss.n1224 0.013
R19201 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vss1p8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.vss3p3 0.013
R19202 dvss.n2932 dvss.n2931 0.013
R19203 dvss.n2921 dvss.n2920 0.013
R19204 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vss1p8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.vss3p3 0.013
R19205 dvss.n2848 dvss.n2847 0.013
R19206 dvss.n2810 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vss1p8 0.013
R19207 dvss.n2610 dvss.n2600 0.013
R19208 dvss.n2605 dvss.n2601 0.013
R19209 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vss1p8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.vss3p3 0.013
R19210 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vss1p8 dvss.n2533 0.012
R19211 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vss1p8 dvss.n2887 0.012
R19212 dvss.n1772 dvss.n1771 0.011
R19213 dvss.n2390 dvss.n2389 0.011
R19214 dvss.n1159 dvss.n1158 0.011
R19215 dvss.n547 dvss.n546 0.011
R19216 dvss.n2474 dvss.n2473 0.011
R19217 dvss.n1719 dvss.n1481 0.011
R19218 dvss.n2337 dvss.n2099 0.011
R19219 dvss.n1106 dvss.n868 0.011
R19220 dvss.n494 dvss.n256 0.011
R19221 dvss.n2543 dvss.n2542 0.01
R19222 dvss.n47 dvss.n46 0.01
R19223 dvss.n2887 dvss.n48 0.01
R19224 dvss.n2820 dvss.n2819 0.01
R19225 dvss.n2453 dvss.n1894 0.009
R19226 dvss.n2514 dvss.n1845 0.009
R19227 dvss.n2512 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 0.009
R19228 dvss.n2795 dvss.n2774 0.009
R19229 dvss.n2585 dvss.n1230 0.009
R19230 dvss.n2583 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 0.009
R19231 dvss.n2861 dvss.n616 0.009
R19232 dvss.n2859 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 0.009
R19233 dvss.n2799 dvss.n663 0.009
R19234 dvss.n2757 dvss.n2756 0.009
R19235 dvss.n2601 dvss.n3 0.009
R19236 dvss.n2933 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.VGND 0.009
R19237 dvss.n1372 dvss.n1370 0.008
R19238 dvss.n1990 dvss.n1988 0.008
R19239 dvss.n1837 dvss.n1836 0.008
R19240 dvss.n759 dvss.n757 0.008
R19241 dvss.n147 dvss.n145 0.008
R19242 dvss.n2877 dvss.n2876 0.008
R19243 dvss.n1830 dvss.n1380 0.008
R19244 dvss.n2448 dvss.n1998 0.008
R19245 dvss.n2456 dvss.n2455 0.008
R19246 dvss.n1217 dvss.n767 0.008
R19247 dvss.n605 dvss.n155 0.008
R19248 dvss.n2802 dvss.n2801 0.008
R19249 dvss.n2526 dvss.n2525 0.007
R19250 dvss.n2880 dvss.n2879 0.007
R19251 dvss.n2514 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vss1p8 0.007
R19252 dvss.n2585 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vss1p8 0.007
R19253 dvss.n2861 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vss1p8 0.007
R19254 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vss1p8 dvss.n3 0.007
R19255 dvss.n1748 dvss.n1430 0.007
R19256 dvss.n2366 dvss.n2048 0.007
R19257 dvss.n1135 dvss.n817 0.007
R19258 dvss.n523 dvss.n205 0.007
R19259 dvss.n2787 EF_AMUX21m_1.invm_0.vss3p3 0.006
R19260 dvss.n2787 dvss.n2786 0.006
R19261 dvss.n2594 dvss.n2593 0.006
R19262 dvss.n2773 dvss.n2596 0.006
R19263 dvss.n2610 dvss.n2609 0.006
R19264 dvss.n1511 dvss.n1506 0.005
R19265 dvss.n1714 dvss.n1505 0.005
R19266 dvss.n1490 dvss.n1485 0.005
R19267 dvss.n2129 dvss.n2124 0.005
R19268 dvss.n2332 dvss.n2123 0.005
R19269 dvss.n2108 dvss.n2103 0.005
R19270 dvss.n898 dvss.n893 0.005
R19271 dvss.n1101 dvss.n892 0.005
R19272 dvss.n877 dvss.n872 0.005
R19273 dvss.n286 dvss.n281 0.005
R19274 dvss.n489 dvss.n280 0.005
R19275 dvss.n265 dvss.n260 0.005
R19276 EF_AMUX21m_2.invm_0.vss3p3 dvss.n2596 0.005
R19277 dvss.n2655 dvss.n2626 0.004
R19278 dvss.n1321 dvss.n1309 0.004
R19279 dvss.n1939 dvss.n1927 0.004
R19280 dvss.n708 dvss.n696 0.004
R19281 dvss.n96 dvss.n84 0.004
R19282 dvss.n2476 dvss.n1881 0.003
R19283 dvss.n2524 dvss.n2523 0.003
R19284 dvss.n2545 dvss.n1266 0.003
R19285 dvss.n1223 dvss.n1222 0.003
R19286 dvss.n2897 dvss.n40 0.003
R19287 dvss.n2871 dvss.n2870 0.003
R19288 dvss.n2822 dvss.n650 0.003
R19289 dvss.n2600 dvss.n2599 0.003
R19290 dvss.n1718 dvss.n1716 0.003
R19291 dvss.n2336 dvss.n2334 0.003
R19292 dvss.n1105 dvss.n1103 0.003
R19293 dvss.n493 dvss.n491 0.003
R19294 dvss.n1364 dvss.n1363 0.002
R19295 dvss.n1515 dvss.n1514 0.002
R19296 dvss.n1494 dvss.n1493 0.002
R19297 dvss.n1982 dvss.n1981 0.002
R19298 dvss.n2133 dvss.n2132 0.002
R19299 dvss.n2112 dvss.n2111 0.002
R19300 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.vss3p3 dvss.n2513 0.002
R19301 dvss.n2513 dvss.n2512 0.002
R19302 dvss.n2584 dvss.n2583 0.002
R19303 dvss.n751 dvss.n750 0.002
R19304 dvss.n902 dvss.n901 0.002
R19305 dvss.n881 dvss.n880 0.002
R19306 dvss.n139 dvss.n138 0.002
R19307 dvss.n290 dvss.n289 0.002
R19308 dvss.n269 dvss.n268 0.002
R19309 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.vss3p3 dvss.n2860 0.002
R19310 dvss.n2860 dvss.n2859 0.002
R19311 dvss.n2935 dvss.n2933 0.002
R19312 dvss.n1719 dvss.n1718 0.001
R19313 dvss.n2337 dvss.n2336 0.001
R19314 dvss.n1106 dvss.n1105 0.001
R19315 dvss.n494 dvss.n493 0.001
R19316 dvss.n1373 dvss.n1372 0.001
R19317 dvss.n1991 dvss.n1990 0.001
R19318 dvss.n2462 dvss.n1894 0.001
R19319 dvss.n1836 dvss.n1274 0.001
R19320 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.vss3p3 dvss.n2584 0.001
R19321 dvss.n760 dvss.n759 0.001
R19322 dvss.n148 dvss.n147 0.001
R19323 dvss.n2876 dvss.n2873 0.001
R19324 dvss.n2808 dvss.n663 0.001
R19325 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.vss3p3 dvss.n2935 0.001
R19326 dvss.n2454 dvss.n2452 0.001
R19327 dvss.n1838 dvss.n1834 0.001
R19328 dvss.n2800 dvss.n1221 0.001
R19329 dvss.n2878 dvss.n609 0.001
R19330 dvss.n1833 dvss.n1278 0.001
R19331 dvss.n2451 dvss.n1896 0.001
R19332 dvss.n1220 dvss.n665 0.001
R19333 dvss.n608 dvss.n53 0.001
R19334 dvss.n1716 dvss.n1481 0.001
R19335 dvss.n2334 dvss.n2099 0.001
R19336 dvss.n1103 dvss.n868 0.001
R19337 dvss.n491 dvss.n256 0.001
R19338 a_570_n5724.n2 a_570_n5724.t0 333.409
R19339 a_570_n5724.n1 a_570_n5724.n0 177.236
R19340 a_570_n5724.t5 a_570_n5724.n7 153.872
R19341 a_570_n5724.n1 a_570_n5724.t8 139.997
R19342 a_570_n5724.n0 a_570_n5724.t7 124.47
R19343 a_570_n5724.n5 a_570_n5724.n4 104.473
R19344 a_570_n5724.n0 a_570_n5724.t6 88.32
R19345 a_570_n5724.n2 a_570_n5724.n1 65.236
R19346 a_570_n5724.n6 a_570_n5724.n5 60.509
R19347 a_570_n5724.n5 a_570_n5724.n3 43.964
R19348 a_570_n5724.n6 a_570_n5724.n2 22.109
R19349 a_570_n5724.n7 a_570_n5724.n6 20.908
R19350 a_570_n5724.n3 a_570_n5724.t2 10.64
R19351 a_570_n5724.n3 a_570_n5724.t4 10.64
R19352 a_570_n5724.n4 a_570_n5724.t1 10.64
R19353 a_570_n5724.n4 a_570_n5724.t3 10.64
R19354 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 136.803
R19355 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 136.324
R19356 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 119.998
R19357 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 93.901
R19358 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 93.303
R19359 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 93.083
R19360 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n4 92.5
R19361 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 92.462
R19362 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 69.227
R19363 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 29.482
R19364 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 27.695
R19365 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 27.695
R19366 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 15.462
R19367 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n16 9.3
R19368 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n8 9.3
R19369 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n7 9.3
R19370 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 9.3
R19371 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 9.3
R19372 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n15 9.3
R19373 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n17 9.3
R19374 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 9.02
R19375 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 9.02
R19376 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n34 8.282
R19377 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n21 8.282
R19378 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 5.647
R19379 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 5.316
R19380 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n42 4.141
R19381 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n28 4.141
R19382 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 4.067
R19383 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n11 3.931
R19384 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n40 3.764
R19385 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n33 3.764
R19386 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n24 3.764
R19387 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n19 3.764
R19388 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n36 3.388
R19389 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n22 3.388
R19390 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 3.072
R19391 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 3.072
R19392 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 3.07
R19393 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 3.043
R19394 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 3.033
R19395 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 3.033
R19396 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 3.033
R19397 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n39 2.635
R19398 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n20 2.635
R19399 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 2.362
R19400 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 2.273
R19401 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 2.258
R19402 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 2.258
R19403 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 1.806
R19404 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n30 1.613
R19405 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 1.455
R19406 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 1.192
R19407 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n9 0.752
R19408 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 0.719
R19409 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 0.224
R19410 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 0.175
R19411 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 2.362
R19412 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 1.142
R19413 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 0.994
R19414 b1.n59 b1.n58 185
R19415 b1.n57 b1.n50 185
R19416 b1.n17 b1.n8 185
R19417 b1.n16 b1.n15 185
R19418 b1.n62 b1.t5 120.035
R19419 b1.t6 b1.n7 120.035
R19420 b1.n52 b1.n50 112.829
R19421 b1.n15 b1.n14 112.829
R19422 b1.n61 b1.n60 104.172
R19423 b1.n20 b1.n19 104.172
R19424 b1.n61 b1.n49 92.5
R19425 b1.n21 b1.n20 92.5
R19426 b1.t5 b1.n61 66.827
R19427 b1.n20 b1.t6 66.827
R19428 b1.n76 b1.t2 35.203
R19429 b1.n73 b1.t3 34.056
R19430 b1.n60 b1.n59 29.482
R19431 b1.n19 b1.n8 29.482
R19432 b1.n71 b1.t7 27.695
R19433 b1.n71 b1.t4 27.695
R19434 b1.n38 b1.n37 19.093
R19435 b1.n62 b1.n49 15.455
R19436 b1.n21 b1.n7 15.455
R19437 b1.n57 b1.n56 13.552
R19438 b1.n16 b1.n11 13.552
R19439 b1.n72 b1.n71 9.676
R19440 b1.n34 b1.n27 9.305
R19441 b1.n52 b1.n51 9.304
R19442 b1.n14 b1.n13 9.304
R19443 b1.n33 b1.n32 9.3
R19444 b1.n39 b1.n38 9.3
R19445 b1.n64 b1.n63 9.3
R19446 b1.n48 b1.n45 9.3
R19447 b1.n60 b1.n48 9.3
R19448 b1.n56 b1.n55 9.3
R19449 b1.n65 b1.n47 9.3
R19450 b1.n22 b1.n6 9.3
R19451 b1.n18 b1.n4 9.3
R19452 b1.n19 b1.n18 9.3
R19453 b1.n11 b1.n10 9.3
R19454 b1.n24 b1.n23 9.3
R19455 b1.n64 b1.n49 9.035
R19456 b1.n22 b1.n21 9.035
R19457 b1.n36 b1.n34 8.493
R19458 b1.n36 b1.t1 8.265
R19459 b1.n36 b1.t0 8.265
R19460 b1.n37 b1.n36 7.977
R19461 b1.n35 b1.n33 7.266
R19462 b1.n36 b1.n35 6.152
R19463 b1.n58 b1.n48 5.647
R19464 b1.n18 b1.n17 5.647
R19465 b1.n34 b1.n28 4.894
R19466 b1.n53 b1.n52 4.894
R19467 b1.n14 b1.n12 4.894
R19468 b1.n66 b1.n48 4.517
R19469 b1.n65 b1.n64 4.517
R19470 b1.n18 b1.n5 4.517
R19471 b1.n23 b1.n22 4.517
R19472 b1.n75 b1.n74 4.5
R19473 b1.n74 b1.n72 4.5
R19474 b1.n44 b1.n2 4.5
R19475 b1.n42 b1.n2 4.5
R19476 b1.n44 b1.n43 4.5
R19477 b1.n43 b1.n42 4.5
R19478 b1.n67 b1.n46 4.5
R19479 b1.n68 b1.n1 4.5
R19480 b1.n46 b1.n1 4.5
R19481 b1.n68 b1.n67 4.5
R19482 b1.n41 b1.n25 4.5
R19483 b1.n40 b1.n29 4.5
R19484 b1.n41 b1.n40 4.5
R19485 b1.n29 b1.n25 4.5
R19486 b1.n31 b1.n26 4.5
R19487 b1.n59 b1.n50 3.931
R19488 b1.n15 b1.n8 3.931
R19489 b1.n12 b1.n2 3.033
R19490 b1.n43 b1.n5 3.033
R19491 b1.n53 b1.n1 3.033
R19492 b1.n67 b1.n66 3.033
R19493 b1.n40 b1.n28 3.033
R19494 b1.n73 b1.n70 2.27
R19495 b1.n13 b1.n3 2.252
R19496 b1.n51 b1.n0 2.252
R19497 b1.n27 b1.n26 2.251
R19498 b1.n30 b1.n26 2.244
R19499 b1.n66 b1.n65 1.882
R19500 b1.n23 b1.n5 1.882
R19501 b1.n38 b1.n28 1.505
R19502 b1.n56 b1.n53 1.505
R19503 b1.n12 b1.n11 1.505
R19504 b1.n9 b1.n3 1.492
R19505 b1.n54 b1.n0 1.492
R19506 b1.n63 b1.n62 1.491
R19507 b1.n7 b1.n6 1.49
R19508 b1.n58 b1.n57 0.752
R19509 b1.n17 b1.n16 0.752
R19510 b1.n37 b1.n33 0.521
R19511 EF_AMUX21m_2.a EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.in0 0.456
R19512 b1.n77 b1.n76 0.297
R19513 b1 EF_AMUX21m_2.array_1ls_1tgm_1.in0 0.239
R19514 b1.n42 b1.n41 0.238
R19515 EF_AMUX21m_2.array_1ls_1tgm_1.in0 b1 0.213
R19516 b1.n77 b1.n69 0.195
R19517 b1 b1.n77 0.185
R19518 b1.n76 b1.n75 0.149
R19519 b1.n68 b1.n44 0.124
R19520 b1.n35 b1.n25 0.057
R19521 b1.n55 b1.n54 0.038
R19522 b1.n10 b1.n9 0.037
R19523 b1.n39 b1.n30 0.03
R19524 b1.n75 b1.n70 0.027
R19525 b1.n32 b1.n30 0.025
R19526 b1.n54 b1.n45 0.019
R19527 b1.n9 b1.n4 0.019
R19528 b1.n44 b1.n3 0.016
R19529 b1.n29 b1.n26 0.015
R19530 b1.n67 b1.n45 0.012
R19531 b1.n63 b1.n47 0.012
R19532 b1.n43 b1.n4 0.012
R19533 b1.n24 b1.n6 0.012
R19534 b1.n31 b1.n25 0.011
R19535 b1.n51 b1.n1 0.01
R19536 b1.n13 b1.n2 0.01
R19537 EF_AMUX21m_2.a b1 0.01
R19538 b1.n69 b1.n0 0.009
R19539 b1.n40 b1.n27 0.009
R19540 b1.n67 b1.n47 0.005
R19541 b1.n43 b1.n24 0.005
R19542 b1.n40 b1.n39 0.004
R19543 b1.n55 b1.n1 0.004
R19544 b1.n10 b1.n2 0.004
R19545 b1.n46 b1.n0 0.004
R19546 b1.n69 b1.n68 0.004
R19547 b1.n72 b1.n70 0.003
R19548 b1.n32 b1.n31 0.003
R19549 b1.n41 b1.n26 0.002
R19550 b1.n74 b1.n73 0.001
R19551 b1.n42 b1.n3 0.001
R19552 a_2221_8623.n123 a_2221_8623.t9 60.25
R19553 a_2221_8623.n101 a_2221_8623.t6 60.25
R19554 a_2221_8623.n87 a_2221_8623.t8 60.25
R19555 a_2221_8623.n65 a_2221_8623.t7 60.25
R19556 a_2221_8623.n2 a_2221_8623.n28 9.3
R19557 a_2221_8623.n2 a_2221_8623.n26 9.3
R19558 a_2221_8623.n6 a_2221_8623.n109 9.3
R19559 a_2221_8623.n6 a_2221_8623.n110 9.3
R19560 a_2221_8623.n6 a_2221_8623.n108 9.3
R19561 a_2221_8623.n108 a_2221_8623.n107 9.3
R19562 a_2221_8623.n7 a_2221_8623.n116 9.3
R19563 a_2221_8623.n8 a_2221_8623.n133 9.3
R19564 a_2221_8623.n7 a_2221_8623.n122 9.3
R19565 a_2221_8623.n122 a_2221_8623.n121 9.3
R19566 a_2221_8623.n7 a_2221_8623.n115 9.3
R19567 a_2221_8623.n8 a_2221_8623.n131 9.3
R19568 a_2221_8623.n131 a_2221_8623.n130 9.3
R19569 a_2221_8623.n8 a_2221_8623.n132 9.3
R19570 a_2221_8623.n5 a_2221_8623.n73 9.3
R19571 a_2221_8623.n5 a_2221_8623.n74 9.3
R19572 a_2221_8623.n5 a_2221_8623.n72 9.3
R19573 a_2221_8623.n72 a_2221_8623.n71 9.3
R19574 a_2221_8623.n4 a_2221_8623.n80 9.3
R19575 a_2221_8623.n4 a_2221_8623.n86 9.3
R19576 a_2221_8623.n86 a_2221_8623.n85 9.3
R19577 a_2221_8623.n4 a_2221_8623.n79 9.3
R19578 a_2221_8623.n3 a_2221_8623.n95 9.3
R19579 a_2221_8623.n95 a_2221_8623.n94 9.3
R19580 a_2221_8623.n3 a_2221_8623.n97 9.3
R19581 a_2221_8623.n3 a_2221_8623.n96 9.3
R19582 a_2221_8623.n9 a_2221_8623.n64 9.3
R19583 a_2221_8623.n10 a_2221_8623.n59 9.3
R19584 a_2221_8623.n157 a_2221_8623.n154 9.3
R19585 a_2221_8623.n157 a_2221_8623.n155 9.3
R19586 a_2221_8623.n124 a_2221_8623.n123 8.764
R19587 a_2221_8623.n88 a_2221_8623.n87 8.764
R19588 a_2221_8623.n129 a_2221_8623.n128 7.453
R19589 a_2221_8623.n120 a_2221_8623.n119 7.453
R19590 a_2221_8623.n106 a_2221_8623.n105 7.453
R19591 a_2221_8623.n84 a_2221_8623.n83 7.453
R19592 a_2221_8623.n93 a_2221_8623.n92 7.453
R19593 a_2221_8623.n70 a_2221_8623.n69 7.453
R19594 a_2221_8623.n102 a_2221_8623.n101 6.8
R19595 a_2221_8623.n66 a_2221_8623.n65 6.8
R19596 a_2221_8623.n127 a_2221_8623.n126 5.647
R19597 a_2221_8623.n118 a_2221_8623.n117 5.647
R19598 a_2221_8623.n104 a_2221_8623.n103 5.647
R19599 a_2221_8623.n82 a_2221_8623.n81 5.647
R19600 a_2221_8623.n91 a_2221_8623.n90 5.647
R19601 a_2221_8623.n68 a_2221_8623.n67 5.647
R19602 a_2221_8623.n13 a_2221_8623.t4 5.539
R19603 a_2221_8623.n13 a_2221_8623.t3 5.539
R19604 a_2221_8623.t5 a_2221_8623.n157 5.539
R19605 a_2221_8623.n157 a_2221_8623.t2 5.539
R19606 a_2221_8623.n114 a_2221_8623.n113 4.735
R19607 a_2221_8623.n78 a_2221_8623.n77 4.735
R19608 a_2221_8623.n112 a_2221_8623.n111 4.735
R19609 a_2221_8623.n76 a_2221_8623.n75 4.735
R19610 a_2221_8623.n125 a_2221_8623.n124 4.65
R19611 a_2221_8623.n89 a_2221_8623.n88 4.65
R19612 a_2221_8623.n32 a_2221_8623.n31 4.517
R19613 a_2221_8623.n62 a_2221_8623.n61 4.517
R19614 a_2221_8623.n52 a_2221_8623.n51 4.517
R19615 a_2221_8623.n2 a_2221_8623.n25 4.5
R19616 a_2221_8623.n0 a_2221_8623.n30 4.5
R19617 a_2221_8623.n1 a_2221_8623.n22 4.5
R19618 a_2221_8623.n1 a_2221_8623.n17 4.5
R19619 a_2221_8623.n9 a_2221_8623.n57 4.5
R19620 a_2221_8623.n10 a_2221_8623.n62 4.5
R19621 a_2221_8623.n145 a_2221_8623.n150 4.5
R19622 a_2221_8623.n44 a_2221_8623.n43 4.5
R19623 a_2221_8623.n49 a_2221_8623.n48 4.5
R19624 a_2221_8623.n38 a_2221_8623.n36 4.5
R19625 a_2221_8623.n157 a_2221_8623.n156 4.357
R19626 a_2221_8623.n135 a_2221_8623.n137 4.244
R19627 a_2221_8623.n98 a_2221_8623.n100 4.244
R19628 a_2221_8623.n57 a_2221_8623.n56 3.764
R19629 a_2221_8623.n6 a_2221_8623.n102 3.427
R19630 a_2221_8623.n5 a_2221_8623.n66 3.427
R19631 a_2221_8623.n22 a_2221_8623.n18 3.388
R19632 a_2221_8623.n43 a_2221_8623.n40 3.388
R19633 a_2221_8623.n28 a_2221_8623.n27 3.384
R19634 a_2221_8623.n153 a_2221_8623.n152 3.384
R19635 a_2221_8623.n140 a_2221_8623.t1 3.306
R19636 a_2221_8623.n140 a_2221_8623.t0 3.306
R19637 a_2221_8623.n150 a_2221_8623.n148 3.28
R19638 a_2221_8623.n142 a_2221_8623.n141 3.158
R19639 a_2221_8623.n1 a_2221_8623.n32 3.033
R19640 a_2221_8623.n50 a_2221_8623.n52 3.033
R19641 a_2221_8623.n150 a_2221_8623.n149 3.011
R19642 a_2221_8623.n57 a_2221_8623.n55 2.635
R19643 a_2221_8623.n59 a_2221_8623.n58 2.616
R19644 a_2221_8623.n2 a_2221_8623.n23 2.577
R19645 a_2221_8623.n21 a_2221_8623.n20 2.258
R19646 a_2221_8623.n42 a_2221_8623.n41 2.258
R19647 a_2221_8623.n64 a_2221_8623.n63 2.246
R19648 a_2221_8623.n17 a_2221_8623.n15 2.223
R19649 a_2221_8623.n48 a_2221_8623.n46 2.223
R19650 a_2221_8623.n157 a_2221_8623.n45 1.985
R19651 a_2221_8623.n62 a_2221_8623.n60 1.882
R19652 a_2221_8623.n14 a_2221_8623.n13 1.717
R19653 a_2221_8623.n142 a_2221_8623.n140 1.615
R19654 a_2221_8623.n151 a_2221_8623.n139 1.514
R19655 a_2221_8623.n139 a_2221_8623.n9 1.513
R19656 a_2221_8623.n25 a_2221_8623.n24 1.505
R19657 a_2221_8623.n154 a_2221_8623.n153 1.505
R19658 a_2221_8623.n37 a_2221_8623.n39 1.505
R19659 a_2221_8623.n144 a_2221_8623.n143 1.129
R19660 a_2221_8623.n12 a_2221_8623.n138 3.286
R19661 a_2221_8623.n130 a_2221_8623.n129 0.993
R19662 a_2221_8623.n121 a_2221_8623.n120 0.993
R19663 a_2221_8623.n107 a_2221_8623.n106 0.993
R19664 a_2221_8623.n85 a_2221_8623.n84 0.993
R19665 a_2221_8623.n94 a_2221_8623.n93 0.993
R19666 a_2221_8623.n71 a_2221_8623.n70 0.993
R19667 a_2221_8623.n11 a_2221_8623.n53 0.829
R19668 a_2221_8623.n30 a_2221_8623.n29 0.752
R19669 a_2221_8623.n131 a_2221_8623.n127 0.752
R19670 a_2221_8623.n122 a_2221_8623.n118 0.752
R19671 a_2221_8623.n108 a_2221_8623.n104 0.752
R19672 a_2221_8623.n86 a_2221_8623.n82 0.752
R19673 a_2221_8623.n95 a_2221_8623.n91 0.752
R19674 a_2221_8623.n72 a_2221_8623.n68 0.752
R19675 a_2221_8623.n36 a_2221_8623.n35 0.752
R19676 a_2221_8623.n34 a_2221_8623.n33 0.754
R19677 a_2221_8623.n137 a_2221_8623.n136 0.709
R19678 a_2221_8623.n100 a_2221_8623.n99 0.709
R19679 a_2221_8623.n11 a_2221_8623.n34 0.678
R19680 a_2221_8623.n114 a_2221_8623.n112 0.456
R19681 a_2221_8623.n78 a_2221_8623.n76 0.456
R19682 a_2221_8623.n22 a_2221_8623.n21 0.376
R19683 a_2221_8623.n20 a_2221_8623.n19 0.376
R19684 a_2221_8623.n147 a_2221_8623.n146 0.376
R19685 a_2221_8623.n43 a_2221_8623.n42 0.376
R19686 a_2221_8623.n33 a_2221_8623.n14 0.224
R19687 a_2221_8623.n151 a_2221_8623.n142 0.223
R19688 a_2221_8623.n8 a_2221_8623.n125 0.19
R19689 a_2221_8623.n125 a_2221_8623.n7 0.19
R19690 a_2221_8623.n89 a_2221_8623.n4 0.19
R19691 a_2221_8623.n3 a_2221_8623.n89 0.19
R19692 a_2221_8623.n138 a_2221_8623.n98 0.158
R19693 a_2221_8623.n138 a_2221_8623.n135 0.158
R19694 a_2221_8623.n148 a_2221_8623.n147 0.09
R19695 a_2221_8623.n151 a_2221_8623.n145 0.085
R19696 a_2221_8623.n53 a_2221_8623.n50 0.05
R19697 a_2221_8623.n53 a_2221_8623.n44 0.039
R19698 a_2221_8623.n15 a_2221_8623.n16 0.03
R19699 a_2221_8623.n46 a_2221_8623.n47 0.03
R19700 a_2221_8623.n145 a_2221_8623.n144 4.543
R19701 a_2221_8623.n44 a_2221_8623.n38 0.042
R19702 a_2221_8623.n139 a_2221_8623.n12 0.903
R19703 a_2221_8623.n49 a_2221_8623.n45 0.011
R19704 a_2221_8623.n50 a_2221_8623.n49 0.043
R19705 a_2221_8623.n11 a_2221_8623.n12 1.082
R19706 a_2221_8623.n135 a_2221_8623.n134 0.039
R19707 a_2221_8623.n9 a_2221_8623.n54 2.769
R19708 a_2221_8623.n38 a_2221_8623.n37 4.629
R19709 a_2221_8623.n7 a_2221_8623.n114 0.203
R19710 a_2221_8623.n112 a_2221_8623.n6 0.203
R19711 a_2221_8623.n76 a_2221_8623.n5 0.203
R19712 a_2221_8623.n4 a_2221_8623.n78 0.203
R19713 a_2221_8623.n98 a_2221_8623.n3 0.173
R19714 a_2221_8623.n0 a_2221_8623.n2 0.166
R19715 a_2221_8623.n9 a_2221_8623.n10 0.162
R19716 a_2221_8623.n134 a_2221_8623.n8 0.136
R19717 a_2221_8623.n1 a_2221_8623.n0 0.132
R19718 a_2221_8623.n33 a_2221_8623.n1 0.103
R19719 comparator_top_0.comparator_0.VBP.n54 comparator_top_0.comparator_0.VBP.t3 116.84
R19720 comparator_top_0.comparator_0.VBP.n81 comparator_top_0.comparator_0.VBP.t2 60.25
R19721 comparator_top_0.comparator_0.VBP.n13 comparator_top_0.comparator_0.VBP.t4 60.25
R19722 comparator_top_0.comparator_0.VBP.n25 comparator_top_0.comparator_0.VBP.t5 60.25
R19723 comparator_top_0.comparator_0.VBP.n58 comparator_top_0.comparator_0.VBP.n57 52.689
R19724 comparator_top_0.comparator_0.VBP.n66 comparator_top_0.comparator_0.VBP.n65 46.103
R19725 comparator_top_0.comparator_0.VBP.n114 comparator_top_0.comparator_0.VBP.n113 39.517
R19726 comparator_top_0.comparator_0.VBP.n106 comparator_top_0.comparator_0.VBP.n105 32.931
R19727 comparator_top_0.comparator_0.VBP.n97 comparator_top_0.comparator_0.VBP.n96 29.637
R19728 comparator_top_0.comparator_0.VBP.n96 comparator_top_0.comparator_0.VBP.n95 26.344
R19729 comparator_top_0.comparator_0.VBP.n107 comparator_top_0.comparator_0.VBP.n106 23.051
R19730 comparator_top_0.comparator_0.VBP.n115 comparator_top_0.comparator_0.VBP.n114 16.465
R19731 comparator_top_0.comparator_0.VBP.n67 comparator_top_0.comparator_0.VBP.n66 9.879
R19732 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n61 9.3
R19733 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n69 9.3
R19734 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n68 9.3
R19735 comparator_top_0.comparator_0.VBP.n68 comparator_top_0.comparator_0.VBP.n67 9.3
R19736 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n62 9.3
R19737 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n60 9.3
R19738 comparator_top_0.comparator_0.VBP.n60 comparator_top_0.comparator_0.VBP.n59 9.3
R19739 comparator_top_0.comparator_0.VBP.n8 comparator_top_0.comparator_0.VBP.n101 9.3
R19740 comparator_top_0.comparator_0.VBP.n108 comparator_top_0.comparator_0.VBP.n107 9.3
R19741 comparator_top_0.comparator_0.VBP.n116 comparator_top_0.comparator_0.VBP.n115 9.3
R19742 comparator_top_0.comparator_0.VBP.n8 comparator_top_0.comparator_0.VBP.n98 9.3
R19743 comparator_top_0.comparator_0.VBP.n98 comparator_top_0.comparator_0.VBP.n97 9.3
R19744 comparator_top_0.comparator_0.VBP.n90 comparator_top_0.comparator_0.VBP.n89 9.3
R19745 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n84 9.3
R19746 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n73 9.3
R19747 comparator_top_0.comparator_0.VBP.n79 comparator_top_0.comparator_0.VBP.n78 9.3
R19748 comparator_top_0.comparator_0.VBP.n4 comparator_top_0.comparator_0.VBP.n22 9.3
R19749 comparator_top_0.comparator_0.VBP.n4 comparator_top_0.comparator_0.VBP.n20 9.3
R19750 comparator_top_0.comparator_0.VBP.n20 comparator_top_0.comparator_0.VBP.n19 9.3
R19751 comparator_top_0.comparator_0.VBP.n4 comparator_top_0.comparator_0.VBP.n21 9.3
R19752 comparator_top_0.comparator_0.VBP.n5 comparator_top_0.comparator_0.VBP.n32 9.3
R19753 comparator_top_0.comparator_0.VBP.n32 comparator_top_0.comparator_0.VBP.n31 9.3
R19754 comparator_top_0.comparator_0.VBP.n5 comparator_top_0.comparator_0.VBP.n34 9.3
R19755 comparator_top_0.comparator_0.VBP.n5 comparator_top_0.comparator_0.VBP.n33 9.3
R19756 comparator_top_0.comparator_0.VBP.n6 comparator_top_0.comparator_0.VBP.n43 9.3
R19757 comparator_top_0.comparator_0.VBP.n6 comparator_top_0.comparator_0.VBP.n38 9.3
R19758 comparator_top_0.comparator_0.VBP.n82 comparator_top_0.comparator_0.VBP.n81 8.764
R19759 comparator_top_0.comparator_0.VBP.n77 comparator_top_0.comparator_0.VBP.n76 7.453
R19760 comparator_top_0.comparator_0.VBP.n88 comparator_top_0.comparator_0.VBP.n87 7.453
R19761 comparator_top_0.comparator_0.VBP.n18 comparator_top_0.comparator_0.VBP.n17 7.453
R19762 comparator_top_0.comparator_0.VBP.n30 comparator_top_0.comparator_0.VBP.n29 7.453
R19763 comparator_top_0.comparator_0.VBP.n14 comparator_top_0.comparator_0.VBP.n13 6.8
R19764 comparator_top_0.comparator_0.VBP.n26 comparator_top_0.comparator_0.VBP.n25 6.8
R19765 comparator_top_0.comparator_0.VBP.n56 comparator_top_0.comparator_0.VBP.n55 6.023
R19766 comparator_top_0.comparator_0.VBP.n2 comparator_top_0.comparator_0.VBP.n118 6
R19767 comparator_top_0.comparator_0.VBP.n2 comparator_top_0.comparator_0.VBP.n111 6
R19768 comparator_top_0.comparator_0.VBP.n75 comparator_top_0.comparator_0.VBP.n74 5.647
R19769 comparator_top_0.comparator_0.VBP.n86 comparator_top_0.comparator_0.VBP.n85 5.647
R19770 comparator_top_0.comparator_0.VBP.n16 comparator_top_0.comparator_0.VBP.n15 5.647
R19771 comparator_top_0.comparator_0.VBP.n28 comparator_top_0.comparator_0.VBP.n27 5.647
R19772 comparator_top_0.comparator_0.VBP.n64 comparator_top_0.comparator_0.VBP.n63 5.27
R19773 comparator_top_0.comparator_0.VBP.n10 comparator_top_0.comparator_0.VBP.n94 5.25
R19774 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n72 4.88
R19775 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n83 4.878
R19776 comparator_top_0.comparator_0.VBP.n1 comparator_top_0.comparator_0.VBP.n9 4.543
R19777 comparator_top_0.comparator_0.VBP.n41 comparator_top_0.comparator_0.VBP.n40 4.517
R19778 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n80 4.5
R19779 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n91 4.5
R19780 comparator_top_0.comparator_0.VBP.n8 comparator_top_0.comparator_0.VBP.n103 4.5
R19781 comparator_top_0.comparator_0.VBP.n10 comparator_top_0.comparator_0.VBP.n93 4.5
R19782 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n71 4.5
R19783 comparator_top_0.comparator_0.VBP.n6 comparator_top_0.comparator_0.VBP.n41 4.5
R19784 comparator_top_0.comparator_0.VBP.n6 comparator_top_0.comparator_0.VBP.n46 4.5
R19785 comparator_top_0.comparator_0.VBP.n1 comparator_top_0.comparator_0.VBP.n51 4.5
R19786 comparator_top_0.comparator_0.VBP.n4 comparator_top_0.comparator_0.VBP.n12 4.244
R19787 comparator_top_0.comparator_0.VBP.n5 comparator_top_0.comparator_0.VBP.n24 4.244
R19788 comparator_top_0.comparator_0.VBP.n3 comparator_top_0.comparator_0.VBP.n54 4.235
R19789 comparator_top_0.comparator_0.VBP.n118 comparator_top_0.comparator_0.VBP.n112 4.141
R19790 comparator_top_0.comparator_0.VBP.n46 comparator_top_0.comparator_0.VBP.n45 3.764
R19791 comparator_top_0.comparator_0.VBP.n5 comparator_top_0.comparator_0.VBP.n26 3.428
R19792 comparator_top_0.comparator_0.VBP.n4 comparator_top_0.comparator_0.VBP.n14 3.427
R19793 comparator_top_0.comparator_0.VBP.n111 comparator_top_0.comparator_0.VBP.n104 3.388
R19794 comparator_top_0.comparator_0.VBP.n52 comparator_top_0.comparator_0.VBP.t1 3.306
R19795 comparator_top_0.comparator_0.VBP.n52 comparator_top_0.comparator_0.VBP.t0 3.306
R19796 comparator_top_0.comparator_0.VBP.n59 comparator_top_0.comparator_0.VBP.n58 3.293
R19797 comparator_top_0.comparator_0.VBP.n51 comparator_top_0.comparator_0.VBP.n49 3.746
R19798 comparator_top_0.comparator_0.VBP comparator_top_0.comparator_0.VBP.n120 3.264
R19799 comparator_top_0.comparator_0.VBP.n1 comparator_top_0.comparator_0.VBP.n53 3.158
R19800 comparator_top_0.comparator_0.VBP.n0 comparator_top_0.comparator_0.VBP.n82 3.033
R19801 comparator_top_0.comparator_0.VBP.n100 comparator_top_0.comparator_0.VBP.n99 3.011
R19802 comparator_top_0.comparator_0.VBP.n51 comparator_top_0.comparator_0.VBP.n50 3.011
R19803 comparator_top_0.comparator_0.VBP.n6 comparator_top_0.comparator_0.VBP.n36 2.769
R19804 comparator_top_0.comparator_0.VBP.n46 comparator_top_0.comparator_0.VBP.n44 2.635
R19805 comparator_top_0.comparator_0.VBP.n38 comparator_top_0.comparator_0.VBP.n37 2.616
R19806 comparator_top_0.comparator_0.VBP.n110 comparator_top_0.comparator_0.VBP.n109 2.258
R19807 comparator_top_0.comparator_0.VBP.n43 comparator_top_0.comparator_0.VBP.n42 2.246
R19808 comparator_top_0.comparator_0.VBP.n117 comparator_top_0.comparator_0.VBP.n116 1.882
R19809 comparator_top_0.comparator_0.VBP.n101 comparator_top_0.comparator_0.VBP.n100 1.882
R19810 comparator_top_0.comparator_0.VBP.n41 comparator_top_0.comparator_0.VBP.n39 1.882
R19811 comparator_top_0.comparator_0.VBP.n7 comparator_top_0.comparator_0.VBP.n0 1.841
R19812 comparator_top_0.comparator_0.VBP.n47 comparator_top_0.comparator_0.VBP.n1 1.822
R19813 comparator_top_0.comparator_0.VBP.n35 comparator_top_0.comparator_0.VBP.n5 1.754
R19814 comparator_top_0.comparator_0.VBP.n2 comparator_top_0.comparator_0.VBP.n3 1.743
R19815 comparator_top_0.comparator_0.VBP.n47 comparator_top_0.comparator_0.VBP.n6 1.675
R19816 comparator_top_0.comparator_0.VBP.n1 comparator_top_0.comparator_0.VBP.n52 1.615
R19817 comparator_top_0.comparator_0.VBP.n2 comparator_top_0.comparator_0.VBP.n8 1.604
R19818 comparator_top_0.comparator_0.VBP.n2 comparator_top_0.comparator_0.VBP.n10 1.549
R19819 comparator_top_0.comparator_0.VBP.n93 comparator_top_0.comparator_0.VBP.n92 1.505
R19820 comparator_top_0.comparator_0.VBP comparator_top_0.comparator_0.VBP.n35 1.314
R19821 comparator_top_0.comparator_0.VBP.n68 comparator_top_0.comparator_0.VBP.n64 1.129
R19822 comparator_top_0.comparator_0.VBP.n9 comparator_top_0.comparator_0.VBP.n48 1.129
R19823 comparator_top_0.comparator_0.VBP.n120 comparator_top_0.comparator_0.VBP.n47 1.042
R19824 comparator_top_0.comparator_0.VBP.n78 comparator_top_0.comparator_0.VBP.n77 0.993
R19825 comparator_top_0.comparator_0.VBP.n89 comparator_top_0.comparator_0.VBP.n88 0.993
R19826 comparator_top_0.comparator_0.VBP.n19 comparator_top_0.comparator_0.VBP.n18 0.993
R19827 comparator_top_0.comparator_0.VBP.n31 comparator_top_0.comparator_0.VBP.n30 0.993
R19828 comparator_top_0.comparator_0.VBP.n119 comparator_top_0.comparator_0.VBP.n2 0.79
R19829 comparator_top_0.comparator_0.VBP.n71 comparator_top_0.comparator_0.VBP.n70 0.752
R19830 comparator_top_0.comparator_0.VBP.n103 comparator_top_0.comparator_0.VBP.n102 0.752
R19831 comparator_top_0.comparator_0.VBP.n80 comparator_top_0.comparator_0.VBP.n79 0.752
R19832 comparator_top_0.comparator_0.VBP.n79 comparator_top_0.comparator_0.VBP.n75 0.752
R19833 comparator_top_0.comparator_0.VBP.n90 comparator_top_0.comparator_0.VBP.n86 0.752
R19834 comparator_top_0.comparator_0.VBP.n91 comparator_top_0.comparator_0.VBP.n90 0.752
R19835 comparator_top_0.comparator_0.VBP.n20 comparator_top_0.comparator_0.VBP.n16 0.752
R19836 comparator_top_0.comparator_0.VBP.n32 comparator_top_0.comparator_0.VBP.n28 0.752
R19837 comparator_top_0.comparator_0.VBP.n2 comparator_top_0.comparator_0.VBP.n7 0.735
R19838 comparator_top_0.comparator_0.VBP.n12 comparator_top_0.comparator_0.VBP.n11 0.709
R19839 comparator_top_0.comparator_0.VBP.n24 comparator_top_0.comparator_0.VBP.n23 0.709
R19840 comparator_top_0.comparator_0.VBP.n5 comparator_top_0.comparator_0.VBP.n4 0.664
R19841 comparator_top_0.comparator_0.VBP.n120 comparator_top_0.comparator_0.VBP.n119 0.575
R19842 comparator_top_0.comparator_0.VBP.n7 comparator_top_0.comparator_bias_0.VBP 0.536
R19843 comparator_top_0.comparator_0.VBP.n60 comparator_top_0.comparator_0.VBP.n56 0.376
R19844 comparator_top_0.comparator_0.VBP.n118 comparator_top_0.comparator_0.VBP.n117 0.376
R19845 comparator_top_0.comparator_0.VBP.n111 comparator_top_0.comparator_0.VBP.n110 0.376
R19846 comparator_top_0.comparator_0.VBP.n109 comparator_top_0.comparator_0.VBP.n108 0.376
R19847 a_2093_3714.n46 a_2093_3714.n45 6.316
R19848 a_2093_3714.n9 a_2093_3714.n40 6.125
R19849 a_2093_3714.n3 a_2093_3714.n18 6.124
R19850 a_2093_3714.n5 a_2093_3714.n24 6.124
R19851 a_2093_3714.n16 a_2093_3714.t4 5.539
R19852 a_2093_3714.n16 a_2093_3714.t10 5.539
R19853 a_2093_3714.n22 a_2093_3714.t11 5.539
R19854 a_2093_3714.n22 a_2093_3714.t9 5.539
R19855 a_2093_3714.n28 a_2093_3714.t8 5.539
R19856 a_2093_3714.n28 a_2093_3714.t3 5.539
R19857 a_2093_3714.n33 a_2093_3714.t2 5.539
R19858 a_2093_3714.n33 a_2093_3714.t1 5.539
R19859 a_2093_3714.n35 a_2093_3714.t6 5.539
R19860 a_2093_3714.n35 a_2093_3714.t7 5.539
R19861 a_2093_3714.n50 a_2093_3714.t0 5.539
R19862 a_2093_3714.t5 a_2093_3714.n50 5.539
R19863 a_2093_3714.n48 a_2093_3714.n47 5.268
R19864 a_2093_3714.n6 a_2093_3714.n32 4.5
R19865 a_2093_3714.n8 a_2093_3714.n39 4.5
R19866 a_2093_3714.n4 a_2093_3714.n21 4.5
R19867 a_2093_3714.n7 a_2093_3714.n27 4.5
R19868 a_2093_3714.n2 a_2093_3714.n15 4.5
R19869 a_2093_3714.n1 a_2093_3714.n44 4.5
R19870 a_2093_3714.n1 a_2093_3714.n42 4.5
R19871 a_2093_3714.n50 a_2093_3714.n49 4.273
R19872 a_2093_3714.n15 a_2093_3714.n13 3.764
R19873 a_2093_3714.n21 a_2093_3714.n19 3.764
R19874 a_2093_3714.n27 a_2093_3714.n25 3.764
R19875 a_2093_3714.n32 a_2093_3714.n30 3.764
R19876 a_2093_3714.n39 a_2093_3714.n37 3.764
R19877 a_2093_3714.n44 a_2093_3714.n43 3.764
R19878 a_2093_3714.n42 a_2093_3714.n41 3.011
R19879 a_2093_3714.n15 a_2093_3714.n14 2.635
R19880 a_2093_3714.n21 a_2093_3714.n20 2.635
R19881 a_2093_3714.n27 a_2093_3714.n26 2.635
R19882 a_2093_3714.n32 a_2093_3714.n31 2.635
R19883 a_2093_3714.n39 a_2093_3714.n38 2.635
R19884 a_2093_3714.n11 a_2093_3714.n3 2.201
R19885 a_2093_3714.n0 a_2093_3714.n9 2.183
R19886 a_2093_3714.n49 a_2093_3714.n48 1.896
R19887 a_2093_3714.n1 a_2093_3714.n0 1.56
R19888 a_2093_3714.n11 a_2093_3714.n5 1.484
R19889 a_2093_3714.n10 a_2093_3714.n6 1.738
R19890 a_2093_3714.n12 a_2093_3714.n7 1.737
R19891 a_2093_3714.n46 a_2093_3714.n1 1.641
R19892 a_2093_3714.n7 a_2093_3714.n29 1.463
R19893 a_2093_3714.n8 a_2093_3714.n36 1.463
R19894 a_2093_3714.n2 a_2093_3714.n17 1.463
R19895 a_2093_3714.n4 a_2093_3714.n23 1.463
R19896 a_2093_3714.n6 a_2093_3714.n34 1.463
R19897 a_2093_3714.n0 a_2093_3714.n10 0.752
R19898 a_2093_3714.n10 a_2093_3714.n12 0.717
R19899 a_2093_3714.n12 a_2093_3714.n11 0.7
R19900 a_2093_3714.n29 a_2093_3714.n28 0.4
R19901 a_2093_3714.n36 a_2093_3714.n35 0.4
R19902 a_2093_3714.n17 a_2093_3714.n16 0.4
R19903 a_2093_3714.n23 a_2093_3714.n22 0.4
R19904 a_2093_3714.n34 a_2093_3714.n33 0.4
R19905 a_2093_3714.n50 a_2093_3714.n46 0.4
R19906 a_2093_3714.n3 a_2093_3714.n2 0.254
R19907 a_2093_3714.n5 a_2093_3714.n4 0.254
R19908 a_2093_3714.n9 a_2093_3714.n8 0.253
R19909 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 136.803
R19910 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 136.324
R19911 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 119.998
R19912 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 93.901
R19913 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 93.303
R19914 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 93.083
R19915 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n4 92.5
R19916 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 92.462
R19917 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 69.227
R19918 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 29.482
R19919 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 27.695
R19920 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 27.695
R19921 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n5 15.462
R19922 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n16 9.3
R19923 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n8 9.3
R19924 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n7 9.3
R19925 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 9.3
R19926 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n13 9.3
R19927 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n15 9.3
R19928 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n17 9.3
R19929 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n43 9.02
R19930 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n26 9.02
R19931 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n34 8.282
R19932 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n21 8.282
R19933 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 5.647
R19934 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 5.316
R19935 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n42 4.141
R19936 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n28 4.141
R19937 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 4.067
R19938 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n11 3.931
R19939 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n40 3.764
R19940 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n33 3.764
R19941 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n24 3.764
R19942 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n19 3.764
R19943 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n36 3.388
R19944 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n22 3.388
R19945 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 3.072
R19946 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n37 3.072
R19947 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n35 3.07
R19948 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 3.043
R19949 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 3.033
R19950 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n25 3.033
R19951 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n23 3.033
R19952 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n39 2.635
R19953 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n20 2.635
R19954 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n38 2.362
R19955 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n46 2.273
R19956 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n44 2.258
R19957 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n27 2.258
R19958 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 1.806
R19959 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n30 1.613
R19960 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n6 1.455
R19961 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n3 1.192
R19962 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n9 0.752
R19963 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 0.719
R19964 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 0.224
R19965 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n48 0.175
R19966 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n2 2.362
R19967 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n1 1.142
R19968 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.n0 0.994
R19969 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 120.008
R19970 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 92.941
R19971 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n4 92.5
R19972 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 92.462
R19973 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 73.192
R19974 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 72.162
R19975 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 29.482
R19976 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 27.695
R19977 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 27.695
R19978 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 15.46
R19979 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 9.3
R19980 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 9.3
R19981 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 9.02
R19982 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 9.019
R19983 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n26 8.282
R19984 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n16 8.282
R19985 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 5.647
R19986 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 5.32
R19987 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 5.318
R19988 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n31 4.141
R19989 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n23 4.141
R19990 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n19 4.141
R19991 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 4.033
R19992 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n9 3.931
R19993 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n33 3.764
R19994 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n14 3.764
R19995 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 3.202
R19996 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 3.071
R19997 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 3.044
R19998 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 3.033
R19999 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 3.033
R20000 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 3.033
R20001 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n27 3.011
R20002 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n17 3.011
R20003 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n34 2.635
R20004 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n15 2.635
R20005 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 2.27
R20006 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 2.258
R20007 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 2.258
R20008 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 1.509
R20009 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n7 0.752
R20010 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 2.478
R20011 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 1.148
R20012 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 1.04
R20013 a_2151_594.n7 a_2151_594.t4 60.25
R20014 a_2151_594.n64 a_2151_594.t6 60.25
R20015 a_2151_594.n21 a_2151_594.t9 60.25
R20016 a_2151_594.n42 a_2151_594.t8 60.25
R20017 a_2151_594.n4 a_2151_594.n73 9.3
R20018 a_2151_594.n3 a_2151_594.n57 9.3
R20019 a_2151_594.n2 a_2151_594.n51 9.3
R20020 a_2151_594.n1 a_2151_594.n35 9.3
R20021 a_2151_594.n1 a_2151_594.n34 9.3
R20022 a_2151_594.n2 a_2151_594.n52 9.3
R20023 a_2151_594.n2 a_2151_594.n50 9.3
R20024 a_2151_594.n50 a_2151_594.n49 9.3
R20025 a_2151_594.n1 a_2151_594.n41 9.3
R20026 a_2151_594.n41 a_2151_594.n40 9.3
R20027 a_2151_594.n0 a_2151_594.n29 9.3
R20028 a_2151_594.n0 a_2151_594.n30 9.3
R20029 a_2151_594.n0 a_2151_594.n28 9.3
R20030 a_2151_594.n28 a_2151_594.n27 9.3
R20031 a_2151_594.n4 a_2151_594.n74 9.3
R20032 a_2151_594.n4 a_2151_594.n72 9.3
R20033 a_2151_594.n72 a_2151_594.n71 9.3
R20034 a_2151_594.n3 a_2151_594.n63 9.3
R20035 a_2151_594.n63 a_2151_594.n62 9.3
R20036 a_2151_594.n3 a_2151_594.n56 9.3
R20037 a_2151_594.n5 a_2151_594.n14 9.3
R20038 a_2151_594.n14 a_2151_594.n13 9.3
R20039 a_2151_594.n5 a_2151_594.n16 9.3
R20040 a_2151_594.n5 a_2151_594.n15 9.3
R20041 a_2151_594.n43 a_2151_594.n42 8.764
R20042 a_2151_594.n65 a_2151_594.n64 8.764
R20043 a_2151_594.n26 a_2151_594.n25 8.215
R20044 a_2151_594.n48 a_2151_594.n47 8.215
R20045 a_2151_594.n39 a_2151_594.n38 8.215
R20046 a_2151_594.n70 a_2151_594.n69 8.215
R20047 a_2151_594.n61 a_2151_594.n60 8.215
R20048 a_2151_594.n12 a_2151_594.n11 8.215
R20049 a_2151_594.n22 a_2151_594.n21 6.92
R20050 a_2151_594.n8 a_2151_594.n7 6.919
R20051 a_2151_594.n24 a_2151_594.n23 5.647
R20052 a_2151_594.n46 a_2151_594.n45 5.647
R20053 a_2151_594.n37 a_2151_594.n36 5.647
R20054 a_2151_594.n68 a_2151_594.n67 5.647
R20055 a_2151_594.n59 a_2151_594.n58 5.647
R20056 a_2151_594.n10 a_2151_594.n9 5.647
R20057 a_2151_594.n97 a_2151_594.t2 5.539
R20058 a_2151_594.n97 a_2151_594.t1 5.539
R20059 a_2151_594.n115 a_2151_594.t0 5.539
R20060 a_2151_594.t3 a_2151_594.n115 5.539
R20061 a_2151_594.n78 a_2151_594.n77 5.274
R20062 a_2151_594.n31 a_2151_594.n20 4.764
R20063 a_2151_594.n53 a_2151_594.n19 4.764
R20064 a_2151_594.n75 a_2151_594.n18 4.764
R20065 a_2151_594.n55 a_2151_594.n54 4.764
R20066 a_2151_594.n17 a_2151_594.n6 4.764
R20067 a_2151_594.n33 a_2151_594.n32 4.764
R20068 a_2151_594.n44 a_2151_594.n43 4.65
R20069 a_2151_594.n66 a_2151_594.n65 4.65
R20070 a_2151_594.n104 a_2151_594.n103 4.517
R20071 a_2151_594.n109 a_2151_594.n108 4.517
R20072 a_2151_594.n79 a_2151_594.n90 6
R20073 a_2151_594.n80 a_2151_594.n82 4.5
R20074 a_2151_594.n96 a_2151_594.n101 4.5
R20075 a_2151_594.n92 a_2151_594.n112 4.5
R20076 a_2151_594.n5 a_2151_594.n8 3.478
R20077 a_2151_594.n0 a_2151_594.n22 3.477
R20078 a_2151_594.n90 a_2151_594.n89 3.381
R20079 a_2151_594.n95 a_2151_594.t5 3.306
R20080 a_2151_594.n95 a_2151_594.t7 3.306
R20081 a_2151_594.n84 a_2151_594.n95 3.206
R20082 a_2151_594.n102 a_2151_594.n104 3.033
R20083 a_2151_594.n93 a_2151_594.n109 3.033
R20084 a_2151_594.n115 a_2151_594.n91 2.851
R20085 a_2151_594.n94 a_2151_594.n84 2.628
R20086 a_2151_594.n100 a_2151_594.n99 2.258
R20087 a_2151_594.n111 a_2151_594.n110 2.258
R20088 a_2151_594.n90 a_2151_594.n88 1.882
R20089 a_2151_594.n115 a_2151_594.n114 1.642
R20090 a_2151_594.n98 a_2151_594.n97 1.642
R20091 a_2151_594.n94 a_2151_594.n106 1.619
R20092 a_2151_594.n83 a_2151_594.n86 6
R20093 a_2151_594.n86 a_2151_594.n85 1.129
R20094 a_2151_594.n27 a_2151_594.n26 1.095
R20095 a_2151_594.n49 a_2151_594.n48 1.095
R20096 a_2151_594.n40 a_2151_594.n39 1.095
R20097 a_2151_594.n71 a_2151_594.n70 1.095
R20098 a_2151_594.n62 a_2151_594.n61 1.095
R20099 a_2151_594.n13 a_2151_594.n12 1.095
R20100 a_2151_594.n101 a_2151_594.n100 0.752
R20101 a_2151_594.n28 a_2151_594.n24 0.752
R20102 a_2151_594.n50 a_2151_594.n46 0.752
R20103 a_2151_594.n41 a_2151_594.n37 0.752
R20104 a_2151_594.n72 a_2151_594.n68 0.752
R20105 a_2151_594.n63 a_2151_594.n59 0.752
R20106 a_2151_594.n14 a_2151_594.n10 0.752
R20107 a_2151_594.n88 a_2151_594.n87 0.752
R20108 a_2151_594.n112 a_2151_594.n111 0.752
R20109 a_2151_594.n107 a_2151_594.n94 0.6
R20110 a_2151_594.n106 a_2151_594.n105 0.56
R20111 a_2151_594.n114 a_2151_594.n113 0.46
R20112 a_2151_594.n55 a_2151_594.n53 0.456
R20113 a_2151_594.n33 a_2151_594.n31 0.456
R20114 a_2151_594.n82 a_2151_594.n81 0.376
R20115 a_2151_594.n76 a_2151_594.n17 0.228
R20116 a_2151_594.n76 a_2151_594.n75 0.228
R20117 a_2151_594.n78 a_2151_594.n76 0.19
R20118 a_2151_594.n4 a_2151_594.n66 0.19
R20119 a_2151_594.n66 a_2151_594.n3 0.19
R20120 a_2151_594.n2 a_2151_594.n44 0.19
R20121 a_2151_594.n44 a_2151_594.n1 0.19
R20122 a_2151_594.n83 a_2151_594.n84 0.093
R20123 a_2151_594.n102 a_2151_594.n96 0.132
R20124 a_2151_594.n92 a_2151_594.n93 0.131
R20125 a_2151_594.n79 a_2151_594.n83 0.074
R20126 a_2151_594.n80 a_2151_594.n78 0.121
R20127 a_2151_594.n106 a_2151_594.n102 0.07
R20128 a_2151_594.n93 a_2151_594.n107 0.051
R20129 a_2151_594.n113 a_2151_594.n92 0.09
R20130 a_2151_594.n96 a_2151_594.n98 0.551
R20131 a_2151_594.n80 a_2151_594.n79 1.538
R20132 a_2151_594.n17 a_2151_594.n5 0.203
R20133 a_2151_594.n75 a_2151_594.n4 0.203
R20134 a_2151_594.n3 a_2151_594.n55 0.203
R20135 a_2151_594.n53 a_2151_594.n2 0.203
R20136 a_2151_594.n1 a_2151_594.n33 0.203
R20137 a_2151_594.n31 a_2151_594.n0 0.203
R20138 a_2551_620.n27 a_2551_620.t6 60.25
R20139 a_2551_620.n48 a_2551_620.t7 60.25
R20140 a_2551_620.n70 a_2551_620.t4 60.25
R20141 a_2551_620.n82 a_2551_620.t2 60.25
R20142 a_2551_620.n1 a_2551_620.n90 9.3
R20143 a_2551_620.n1 a_2551_620.n91 9.3
R20144 a_2551_620.n1 a_2551_620.n89 9.3
R20145 a_2551_620.n89 a_2551_620.n88 9.3
R20146 a_2551_620.n2 a_2551_620.n79 9.3
R20147 a_2551_620.n3 a_2551_620.n63 9.3
R20148 a_2551_620.n3 a_2551_620.n62 9.3
R20149 a_2551_620.n3 a_2551_620.n69 9.3
R20150 a_2551_620.n69 a_2551_620.n68 9.3
R20151 a_2551_620.n2 a_2551_620.n78 9.3
R20152 a_2551_620.n78 a_2551_620.n77 9.3
R20153 a_2551_620.n2 a_2551_620.n80 9.3
R20154 a_2551_620.n4 a_2551_620.n57 9.3
R20155 a_2551_620.n5 a_2551_620.n41 9.3
R20156 a_2551_620.n5 a_2551_620.n40 9.3
R20157 a_2551_620.n5 a_2551_620.n47 9.3
R20158 a_2551_620.n47 a_2551_620.n46 9.3
R20159 a_2551_620.n4 a_2551_620.n56 9.3
R20160 a_2551_620.n56 a_2551_620.n55 9.3
R20161 a_2551_620.n4 a_2551_620.n58 9.3
R20162 a_2551_620.n6 a_2551_620.n35 9.3
R20163 a_2551_620.n6 a_2551_620.n34 9.3
R20164 a_2551_620.n34 a_2551_620.n33 9.3
R20165 a_2551_620.n6 a_2551_620.n36 9.3
R20166 a_2551_620.n7 a_2551_620.n98 9.3
R20167 a_2551_620.n7 a_2551_620.n97 9.3
R20168 a_2551_620.n100 a_2551_620.n99 9.3
R20169 a_2551_620.n102 a_2551_620.n101 9.3
R20170 a_2551_620.n104 a_2551_620.n103 9.3
R20171 a_2551_620.n0 a_2551_620.n105 9.3
R20172 a_2551_620.n125 a_2551_620.n112 9.908
R20173 a_2551_620.n125 a_2551_620.n113 11.038
R20174 a_2551_620.n125 a_2551_620.n124 8.891
R20175 a_2551_620.n125 a_2551_620.n121 8.88
R20176 a_2551_620.n125 a_2551_620.n118 8.869
R20177 a_2551_620.n125 a_2551_620.n115 8.858
R20178 a_2551_620.n71 a_2551_620.n70 8.764
R20179 a_2551_620.n49 a_2551_620.n48 8.764
R20180 a_2551_620.n32 a_2551_620.n31 7.453
R20181 a_2551_620.n45 a_2551_620.n44 7.453
R20182 a_2551_620.n54 a_2551_620.n53 7.453
R20183 a_2551_620.n67 a_2551_620.n66 7.453
R20184 a_2551_620.n76 a_2551_620.n75 7.453
R20185 a_2551_620.n87 a_2551_620.n86 7.453
R20186 a_2551_620.n20 a_2551_620.n19 7.451
R20187 a_2551_620.n28 a_2551_620.n27 6.8
R20188 a_2551_620.n83 a_2551_620.n82 6.8
R20189 a_2551_620.n0 a_2551_620.n11 6.291
R20190 a_2551_620.n30 a_2551_620.n29 5.647
R20191 a_2551_620.n43 a_2551_620.n42 5.647
R20192 a_2551_620.n52 a_2551_620.n51 5.647
R20193 a_2551_620.n65 a_2551_620.n64 5.647
R20194 a_2551_620.n74 a_2551_620.n73 5.647
R20195 a_2551_620.n85 a_2551_620.n84 5.647
R20196 a_2551_620.n125 a_2551_620.t5 5.539
R20197 a_2551_620.t3 a_2551_620.n125 5.539
R20198 a_2551_620.n96 a_2551_620.n95 4.955
R20199 a_2551_620.n37 a_2551_620.n26 4.735
R20200 a_2551_620.n59 a_2551_620.n25 4.735
R20201 a_2551_620.n81 a_2551_620.n24 4.735
R20202 a_2551_620.n39 a_2551_620.n38 4.735
R20203 a_2551_620.n61 a_2551_620.n60 4.735
R20204 a_2551_620.n93 a_2551_620.n92 4.735
R20205 a_2551_620.n72 a_2551_620.n71 4.65
R20206 a_2551_620.n50 a_2551_620.n49 4.65
R20207 a_2551_620.n8 a_2551_620.n21 4.5
R20208 a_2551_620.n9 a_2551_620.n20 4.5
R20209 a_2551_620.n8 a_2551_620.n108 4.5
R20210 a_2551_620.n0 a_2551_620.n23 4.5
R20211 a_2551_620.n9 a_2551_620.n110 4.5
R20212 a_2551_620.n6 a_2551_620.n28 3.427
R20213 a_2551_620.n1 a_2551_620.n83 3.427
R20214 a_2551_620.n110 a_2551_620.n109 3.388
R20215 a_2551_620.n117 a_2551_620.n116 3.388
R20216 a_2551_620.n17 a_2551_620.n16 3.381
R20217 a_2551_620.n106 a_2551_620.t1 3.306
R20218 a_2551_620.n106 a_2551_620.t0 3.306
R20219 a_2551_620.n11 a_2551_620.n106 3.206
R20220 a_2551_620.n20 a_2551_620.n18 2.635
R20221 a_2551_620.n120 a_2551_620.n119 2.635
R20222 a_2551_620.n17 a_2551_620.n15 1.882
R20223 a_2551_620.n23 a_2551_620.n22 1.882
R20224 a_2551_620.n123 a_2551_620.n122 1.882
R20225 a_2551_620.n125 a_2551_620.n111 1.669
R20226 a_2551_620.n108 a_2551_620.n107 1.505
R20227 a_2551_620.n10 a_2551_620.n13 6
R20228 a_2551_620.n13 a_2551_620.n12 1.129
R20229 a_2551_620.n33 a_2551_620.n32 0.993
R20230 a_2551_620.n46 a_2551_620.n45 0.993
R20231 a_2551_620.n55 a_2551_620.n54 0.993
R20232 a_2551_620.n68 a_2551_620.n67 0.993
R20233 a_2551_620.n77 a_2551_620.n76 0.993
R20234 a_2551_620.n88 a_2551_620.n87 0.993
R20235 a_2551_620.n111 a_2551_620.n9 0.941
R20236 a_2551_620.n15 a_2551_620.n14 0.752
R20237 a_2551_620.n34 a_2551_620.n30 0.752
R20238 a_2551_620.n47 a_2551_620.n43 0.752
R20239 a_2551_620.n56 a_2551_620.n52 0.752
R20240 a_2551_620.n69 a_2551_620.n65 0.752
R20241 a_2551_620.n78 a_2551_620.n74 0.752
R20242 a_2551_620.n89 a_2551_620.n85 0.752
R20243 a_2551_620.n39 a_2551_620.n37 0.456
R20244 a_2551_620.n61 a_2551_620.n59 0.456
R20245 a_2551_620.n94 a_2551_620.n81 0.228
R20246 a_2551_620.n94 a_2551_620.n93 0.228
R20247 a_2551_620.n96 a_2551_620.n94 0.214
R20248 a_2551_620.n50 a_2551_620.n5 0.19
R20249 a_2551_620.n4 a_2551_620.n50 0.19
R20250 a_2551_620.n72 a_2551_620.n3 0.19
R20251 a_2551_620.n2 a_2551_620.n72 0.19
R20252 a_2551_620.n104 a_2551_620.n102 0.19
R20253 a_2551_620.n0 a_2551_620.n104 0.189
R20254 a_2551_620.n102 a_2551_620.n100 0.189
R20255 a_2551_620.n7 a_2551_620.n96 0.164
R20256 a_2551_620.n115 a_2551_620.n114 0.16
R20257 a_2551_620.n118 a_2551_620.n117 0.149
R20258 a_2551_620.n121 a_2551_620.n120 0.138
R20259 a_2551_620.n124 a_2551_620.n123 0.127
R20260 a_2551_620.n10 a_2551_620.n11 0.093
R20261 a_2551_620.n17 a_2551_620.n10 6.074
R20262 a_2551_620.n37 a_2551_620.n6 0.203
R20263 a_2551_620.n5 a_2551_620.n39 0.203
R20264 a_2551_620.n59 a_2551_620.n4 0.203
R20265 a_2551_620.n3 a_2551_620.n61 0.203
R20266 a_2551_620.n81 a_2551_620.n2 0.203
R20267 a_2551_620.n93 a_2551_620.n1 0.203
R20268 a_2551_620.n8 a_2551_620.n0 0.201
R20269 a_2551_620.n100 a_2551_620.n7 0.189
R20270 a_2551_620.n9 a_2551_620.n8 0.132
R20271 a_5299_3714.n53 a_5299_3714.t2 60.25
R20272 a_5299_3714.n31 a_5299_3714.t9 60.25
R20273 a_5299_3714.n9 a_5299_3714.t8 60.25
R20274 a_5299_3714.n66 a_5299_3714.t0 60.25
R20275 a_5299_3714.n0 a_5299_3714.n74 9.3
R20276 a_5299_3714.n0 a_5299_3714.n75 9.3
R20277 a_5299_3714.n0 a_5299_3714.n73 9.3
R20278 a_5299_3714.n73 a_5299_3714.n72 9.3
R20279 a_5299_3714.n3 a_5299_3714.n41 9.3
R20280 a_5299_3714.n4 a_5299_3714.n23 9.3
R20281 a_5299_3714.n5 a_5299_3714.n18 9.3
R20282 a_5299_3714.n5 a_5299_3714.n17 9.3
R20283 a_5299_3714.n5 a_5299_3714.n16 9.3
R20284 a_5299_3714.n16 a_5299_3714.n15 9.3
R20285 a_5299_3714.n4 a_5299_3714.n24 9.3
R20286 a_5299_3714.n4 a_5299_3714.n30 9.3
R20287 a_5299_3714.n30 a_5299_3714.n29 9.3
R20288 a_5299_3714.n3 a_5299_3714.n40 9.3
R20289 a_5299_3714.n3 a_5299_3714.n39 9.3
R20290 a_5299_3714.n39 a_5299_3714.n38 9.3
R20291 a_5299_3714.n2 a_5299_3714.n45 9.3
R20292 a_5299_3714.n2 a_5299_3714.n52 9.3
R20293 a_5299_3714.n52 a_5299_3714.n51 9.3
R20294 a_5299_3714.n2 a_5299_3714.n46 9.3
R20295 a_5299_3714.n1 a_5299_3714.n61 9.3
R20296 a_5299_3714.n61 a_5299_3714.n60 9.3
R20297 a_5299_3714.n1 a_5299_3714.n63 9.3
R20298 a_5299_3714.n1 a_5299_3714.n62 9.3
R20299 a_5299_3714.n32 a_5299_3714.n31 8.764
R20300 a_5299_3714.n54 a_5299_3714.n53 8.764
R20301 a_5299_3714.n14 a_5299_3714.n13 8.215
R20302 a_5299_3714.n28 a_5299_3714.n27 8.215
R20303 a_5299_3714.n37 a_5299_3714.n36 8.215
R20304 a_5299_3714.n71 a_5299_3714.n70 8.215
R20305 a_5299_3714.n50 a_5299_3714.n49 8.215
R20306 a_5299_3714.n59 a_5299_3714.n58 8.215
R20307 a_5299_3714.n10 a_5299_3714.n9 6.922
R20308 a_5299_3714.n67 a_5299_3714.n66 6.92
R20309 a_5299_3714.n12 a_5299_3714.n11 5.647
R20310 a_5299_3714.n26 a_5299_3714.n25 5.647
R20311 a_5299_3714.n35 a_5299_3714.n34 5.647
R20312 a_5299_3714.n69 a_5299_3714.n68 5.647
R20313 a_5299_3714.n48 a_5299_3714.n47 5.647
R20314 a_5299_3714.n57 a_5299_3714.n56 5.647
R20315 a_5299_3714.n98 a_5299_3714.t5 5.539
R20316 a_5299_3714.n98 a_5299_3714.t4 5.539
R20317 a_5299_3714.n115 a_5299_3714.t6 5.539
R20318 a_5299_3714.t7 a_5299_3714.n115 5.539
R20319 a_5299_3714.n79 a_5299_3714.n78 5.274
R20320 a_5299_3714.n76 a_5299_3714.n65 4.764
R20321 a_5299_3714.n44 a_5299_3714.n8 4.764
R20322 a_5299_3714.n64 a_5299_3714.n7 4.764
R20323 a_5299_3714.n20 a_5299_3714.n19 4.764
R20324 a_5299_3714.n22 a_5299_3714.n21 4.764
R20325 a_5299_3714.n43 a_5299_3714.n42 4.764
R20326 a_5299_3714.n33 a_5299_3714.n32 4.65
R20327 a_5299_3714.n55 a_5299_3714.n54 4.65
R20328 a_5299_3714.n105 a_5299_3714.n104 4.517
R20329 a_5299_3714.n110 a_5299_3714.n109 4.517
R20330 a_5299_3714.n80 a_5299_3714.n91 6
R20331 a_5299_3714.n81 a_5299_3714.n83 4.5
R20332 a_5299_3714.n97 a_5299_3714.n102 4.5
R20333 a_5299_3714.n93 a_5299_3714.n113 4.5
R20334 a_5299_3714.n0 a_5299_3714.n67 3.477
R20335 a_5299_3714.n5 a_5299_3714.n10 3.476
R20336 a_5299_3714.n91 a_5299_3714.n90 3.381
R20337 a_5299_3714.n95 a_5299_3714.t3 3.306
R20338 a_5299_3714.n95 a_5299_3714.t1 3.306
R20339 a_5299_3714.n85 a_5299_3714.n95 3.206
R20340 a_5299_3714.n103 a_5299_3714.n105 3.033
R20341 a_5299_3714.n94 a_5299_3714.n110 3.033
R20342 a_5299_3714.n115 a_5299_3714.n92 2.851
R20343 a_5299_3714.n6 a_5299_3714.n85 2.808
R20344 a_5299_3714.n101 a_5299_3714.n100 2.258
R20345 a_5299_3714.n112 a_5299_3714.n111 2.258
R20346 a_5299_3714.n91 a_5299_3714.n89 1.882
R20347 a_5299_3714.n99 a_5299_3714.n98 1.642
R20348 a_5299_3714.n115 a_5299_3714.n114 1.642
R20349 a_5299_3714.n84 a_5299_3714.n87 6
R20350 a_5299_3714.n87 a_5299_3714.n86 1.129
R20351 a_5299_3714.n15 a_5299_3714.n14 1.095
R20352 a_5299_3714.n29 a_5299_3714.n28 1.095
R20353 a_5299_3714.n38 a_5299_3714.n37 1.095
R20354 a_5299_3714.n72 a_5299_3714.n71 1.095
R20355 a_5299_3714.n51 a_5299_3714.n50 1.095
R20356 a_5299_3714.n60 a_5299_3714.n59 1.095
R20357 a_5299_3714.n107 a_5299_3714.n106 0.76
R20358 a_5299_3714.n16 a_5299_3714.n12 0.752
R20359 a_5299_3714.n30 a_5299_3714.n26 0.752
R20360 a_5299_3714.n39 a_5299_3714.n35 0.752
R20361 a_5299_3714.n73 a_5299_3714.n69 0.752
R20362 a_5299_3714.n52 a_5299_3714.n48 0.752
R20363 a_5299_3714.n61 a_5299_3714.n57 0.752
R20364 a_5299_3714.n89 a_5299_3714.n88 0.752
R20365 a_5299_3714.n102 a_5299_3714.n101 0.752
R20366 a_5299_3714.n113 a_5299_3714.n112 0.752
R20367 a_5299_3714.n6 a_5299_3714.n107 0.678
R20368 a_5299_3714.n106 a_5299_3714.n96 0.572
R20369 a_5299_3714.n44 a_5299_3714.n43 0.456
R20370 a_5299_3714.n22 a_5299_3714.n20 0.456
R20371 a_5299_3714.n83 a_5299_3714.n82 0.376
R20372 a_5299_3714.n77 a_5299_3714.n64 0.228
R20373 a_5299_3714.n77 a_5299_3714.n76 0.228
R20374 a_5299_3714.n79 a_5299_3714.n77 0.19
R20375 a_5299_3714.n33 a_5299_3714.n4 0.19
R20376 a_5299_3714.n3 a_5299_3714.n33 0.19
R20377 a_5299_3714.n55 a_5299_3714.n2 0.19
R20378 a_5299_3714.n1 a_5299_3714.n55 0.19
R20379 a_5299_3714.n84 a_5299_3714.n85 0.093
R20380 a_5299_3714.n93 a_5299_3714.n94 0.132
R20381 a_5299_3714.n103 a_5299_3714.n97 0.132
R20382 a_5299_3714.n80 a_5299_3714.n84 0.074
R20383 a_5299_3714.n81 a_5299_3714.n79 0.121
R20384 a_5299_3714.n106 a_5299_3714.n103 0.058
R20385 a_5299_3714.n94 a_5299_3714.n108 0.052
R20386 a_5299_3714.n114 a_5299_3714.n93 0.549
R20387 a_5299_3714.n97 a_5299_3714.n99 0.551
R20388 a_5299_3714.n81 a_5299_3714.n80 1.538
R20389 a_5299_3714.n108 a_5299_3714.n6 0.62
R20390 a_5299_3714.n20 a_5299_3714.n5 0.203
R20391 a_5299_3714.n4 a_5299_3714.n22 0.203
R20392 a_5299_3714.n43 a_5299_3714.n3 0.203
R20393 a_5299_3714.n2 a_5299_3714.n44 0.203
R20394 a_5299_3714.n64 a_5299_3714.n1 0.203
R20395 a_5299_3714.n76 a_5299_3714.n0 0.203
R20396 a_3916_n5703.n2 a_3916_n5703.t5 333.409
R20397 a_3916_n5703.n1 a_3916_n5703.n0 177.236
R20398 a_3916_n5703.t4 a_3916_n5703.n7 153.872
R20399 a_3916_n5703.n1 a_3916_n5703.t8 139.997
R20400 a_3916_n5703.n0 a_3916_n5703.t7 124.47
R20401 a_3916_n5703.n5 a_3916_n5703.n4 104.473
R20402 a_3916_n5703.n0 a_3916_n5703.t6 88.32
R20403 a_3916_n5703.n2 a_3916_n5703.n1 65.236
R20404 a_3916_n5703.n6 a_3916_n5703.n5 60.509
R20405 a_3916_n5703.n5 a_3916_n5703.n3 43.964
R20406 a_3916_n5703.n6 a_3916_n5703.n2 22.109
R20407 a_3916_n5703.n7 a_3916_n5703.n6 20.908
R20408 a_3916_n5703.n3 a_3916_n5703.t3 10.64
R20409 a_3916_n5703.n3 a_3916_n5703.t1 10.64
R20410 a_3916_n5703.n4 a_3916_n5703.t2 10.64
R20411 a_3916_n5703.n4 a_3916_n5703.t0 10.64
R20412 a_2093_1782.n88 a_2093_1782.n22 8.055
R20413 a_2093_1782.n88 a_2093_1782.n20 8.029
R20414 a_2093_1782.n87 a_2093_1782.n86 6.136
R20415 a_2093_1782.n83 a_2093_1782.n82 5.609
R20416 a_2093_1782.n48 a_2093_1782.n47 5.609
R20417 a_2093_1782.n51 a_2093_1782.n50 5.609
R20418 a_2093_1782.n28 a_2093_1782.n27 5.609
R20419 a_2093_1782.n62 a_2093_1782.n61 5.609
R20420 a_2093_1782.n81 a_2093_1782.n80 5.609
R20421 a_2093_1782.n8 a_2093_1782.n78 4.5
R20422 a_2093_1782.n15 a_2093_1782.n70 4.5
R20423 a_2093_1782.n6 a_2093_1782.n66 4.5
R20424 a_2093_1782.n4 a_2093_1782.n59 4.5
R20425 a_2093_1782.n14 a_2093_1782.n55 4.5
R20426 a_2093_1782.n38 a_2093_1782.n41 4.5
R20427 a_2093_1782.n13 a_2093_1782.n36 4.5
R20428 a_2093_1782.n0 a_2093_1782.n32 4.5
R20429 a_2093_1782.n2 a_2093_1782.n45 4.5
R20430 a_2093_1782.n16 a_2093_1782.n74 4.5
R20431 a_2093_1782.n25 a_2093_1782.n24 4.5
R20432 a_2093_1782.n17 a_2093_1782.n85 4.5
R20433 a_2093_1782.n36 a_2093_1782.n35 3.764
R20434 a_2093_1782.n41 a_2093_1782.n40 3.764
R20435 a_2093_1782.n55 a_2093_1782.n54 3.764
R20436 a_2093_1782.n70 a_2093_1782.n69 3.764
R20437 a_2093_1782.n74 a_2093_1782.n73 3.764
R20438 a_2093_1782.n24 a_2093_1782.n23 3.764
R20439 a_2093_1782.n32 a_2093_1782.n30 3.388
R20440 a_2093_1782.n45 a_2093_1782.n43 3.388
R20441 a_2093_1782.n59 a_2093_1782.n57 3.388
R20442 a_2093_1782.n66 a_2093_1782.n64 3.388
R20443 a_2093_1782.n78 a_2093_1782.n76 3.388
R20444 a_2093_1782.n33 a_2093_1782.t4 3.306
R20445 a_2093_1782.n33 a_2093_1782.t8 3.306
R20446 a_2093_1782.n37 a_2093_1782.t9 3.306
R20447 a_2093_1782.n37 a_2093_1782.t11 3.306
R20448 a_2093_1782.n52 a_2093_1782.t10 3.306
R20449 a_2093_1782.n52 a_2093_1782.t2 3.306
R20450 a_2093_1782.n67 a_2093_1782.t1 3.306
R20451 a_2093_1782.n67 a_2093_1782.t0 3.306
R20452 a_2093_1782.n71 a_2093_1782.t7 3.306
R20453 a_2093_1782.n71 a_2093_1782.t6 3.306
R20454 a_2093_1782.t3 a_2093_1782.n88 3.306
R20455 a_2093_1782.n88 a_2093_1782.t5 3.306
R20456 a_2093_1782.n32 a_2093_1782.n31 3.011
R20457 a_2093_1782.n45 a_2093_1782.n44 3.011
R20458 a_2093_1782.n59 a_2093_1782.n58 3.011
R20459 a_2093_1782.n66 a_2093_1782.n65 3.011
R20460 a_2093_1782.n78 a_2093_1782.n77 3.011
R20461 a_2093_1782.n85 a_2093_1782.n84 3.011
R20462 a_2093_1782.n36 a_2093_1782.n34 2.635
R20463 a_2093_1782.n41 a_2093_1782.n39 2.635
R20464 a_2093_1782.n55 a_2093_1782.n53 2.635
R20465 a_2093_1782.n70 a_2093_1782.n68 2.635
R20466 a_2093_1782.n74 a_2093_1782.n72 2.635
R20467 a_2093_1782.n18 a_2093_1782.n1 2.183
R20468 a_2093_1782.n11 a_2093_1782.n9 2.183
R20469 a_2093_1782.n38 a_2093_1782.n37 1.846
R20470 a_2093_1782.n13 a_2093_1782.n33 1.846
R20471 a_2093_1782.n14 a_2093_1782.n52 1.846
R20472 a_2093_1782.n15 a_2093_1782.n67 1.846
R20473 a_2093_1782.n16 a_2093_1782.n71 1.846
R20474 a_2093_1782.n12 a_2093_1782.n5 1.484
R20475 a_2093_1782.n18 a_2093_1782.n3 1.484
R20476 a_2093_1782.n19 a_2093_1782.n7 1.484
R20477 a_2093_1782.n10 a_2093_1782.n11 1.484
R20478 a_2093_1782.n87 a_2093_1782.n25 1.483
R20479 a_2093_1782.n11 a_2093_1782.n19 0.735
R20480 a_2093_1782.n19 a_2093_1782.n12 0.734
R20481 a_2093_1782.n12 a_2093_1782.n18 0.717
R20482 a_2093_1782.n27 a_2093_1782.n26 0.461
R20483 a_2093_1782.n47 a_2093_1782.n46 0.461
R20484 a_2093_1782.n50 a_2093_1782.n49 0.461
R20485 a_2093_1782.n61 a_2093_1782.n60 0.461
R20486 a_2093_1782.n80 a_2093_1782.n79 0.461
R20487 a_2093_1782.n30 a_2093_1782.n29 0.43
R20488 a_2093_1782.n43 a_2093_1782.n42 0.43
R20489 a_2093_1782.n57 a_2093_1782.n56 0.43
R20490 a_2093_1782.n64 a_2093_1782.n63 0.43
R20491 a_2093_1782.n76 a_2093_1782.n75 0.43
R20492 a_2093_1782.n22 a_2093_1782.n21 0.429
R20493 a_2093_1782.n88 a_2093_1782.n87 0.363
R20494 a_2093_1782.n9 a_2093_1782.n81 0.297
R20495 a_2093_1782.n1 a_2093_1782.n28 0.297
R20496 a_2093_1782.n7 a_2093_1782.n62 0.297
R20497 a_2093_1782.n3 a_2093_1782.n48 0.297
R20498 a_2093_1782.n5 a_2093_1782.n51 0.297
R20499 a_2093_1782.n10 a_2093_1782.n83 0.297
R20500 a_2093_1782.n17 a_2093_1782.n10 0.149
R20501 a_2093_1782.n0 a_2093_1782.n13 0.139
R20502 a_2093_1782.n2 a_2093_1782.n38 0.138
R20503 a_2093_1782.n6 a_2093_1782.n15 0.138
R20504 a_2093_1782.n4 a_2093_1782.n14 0.138
R20505 a_2093_1782.n8 a_2093_1782.n16 0.137
R20506 a_2093_1782.n9 a_2093_1782.n8 0.132
R20507 a_2093_1782.n7 a_2093_1782.n6 0.132
R20508 a_2093_1782.n5 a_2093_1782.n4 0.132
R20509 a_2093_1782.n3 a_2093_1782.n2 0.132
R20510 a_2093_1782.n1 a_2093_1782.n0 0.132
R20511 a_2093_1782.n25 a_2093_1782.n17 0.121
R20512 a_10542_n5707.n3 a_10542_n5707.t5 333.409
R20513 a_10542_n5707.n2 a_10542_n5707.n1 177.236
R20514 a_10542_n5707.n2 a_10542_n5707.t7 139.997
R20515 a_10542_n5707.n1 a_10542_n5707.t6 124.47
R20516 a_10542_n5707.n6 a_10542_n5707.n5 104.474
R20517 a_10542_n5707.n4 a_10542_n5707.t3 103.326
R20518 a_10542_n5707.n1 a_10542_n5707.t8 88.32
R20519 a_10542_n5707.n3 a_10542_n5707.n2 65.236
R20520 a_10542_n5707.n5 a_10542_n5707.n4 60.509
R20521 a_10542_n5707.n5 a_10542_n5707.n0 43.964
R20522 a_10542_n5707.n4 a_10542_n5707.n3 22.109
R20523 a_10542_n5707.n0 a_10542_n5707.t2 10.64
R20524 a_10542_n5707.n0 a_10542_n5707.t1 10.64
R20525 a_10542_n5707.n6 a_10542_n5707.t0 10.64
R20526 a_10542_n5707.t4 a_10542_n5707.n6 10.64
R20527 vo.n7 vo.n6 585
R20528 vo.n3 vo.n2 291.405
R20529 vo.n12 vo.t1 194.386
R20530 vo.n5 vo.n4 148.663
R20531 vo.t1 vo.n11 122.727
R20532 vo.n3 vo.t0 22.418
R20533 vo.n7 vo.n4 10.553
R20534 vo vo.n5 9.627
R20535 vo.n18 vo.n17 9.3
R20536 vo.n15 vo.n14 9.3
R20537 vo.n8 vo.n7 9.3
R20538 vo vo.n10 7.006
R20539 vo vo.n9 6.328
R20540 vo.n13 vo.n12 5.928
R20541 vo.n14 vo.n13 4.727
R20542 vo vo.n11 4.692
R20543 vo.n10 vo.n0 4.65
R20544 vo.n16 vo.n1 4.65
R20545 vo.n10 vo 2.964
R20546 vo vo.n19 2.512
R20547 vo.n13 vo 2.425
R20548 vo.n4 vo.n3 2.191
R20549 vo.n17 vo 2.155
R20550 vo.n9 vo.n0 2.039
R20551 vo.n16 vo.n15 1.751
R20552 vo.n6 vo.n2 1.616
R20553 vo.n12 vo 1.616
R20554 comparator_top_0.VOUT vo 0.921
R20555 vo.n9 vo.n8 0.816
R20556 vo.n15 vo.n11 0.795
R20557 vo.n8 vo.n2 0.673
R20558 vo.n17 vo.n16 0.538
R20559 vo.n5 vo 0.343
R20560 vo.n6 vo 0.269
R20561 vo.n19 vo.n18 0.08
R20562 vo.n14 vo.n1 0.017
R20563 vo.n19 vo.n0 0.009
R20564 vo.n18 vo.n1 0.005
R20565 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 136.803
R20566 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 136.324
R20567 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 119.998
R20568 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 93.901
R20569 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 93.303
R20570 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 93.083
R20571 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n4 92.5
R20572 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 92.462
R20573 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 69.227
R20574 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 29.482
R20575 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 27.695
R20576 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 27.695
R20577 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 15.462
R20578 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n16 9.3
R20579 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n8 9.3
R20580 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n7 9.3
R20581 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 9.3
R20582 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 9.3
R20583 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n15 9.3
R20584 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n17 9.3
R20585 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 9.02
R20586 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 9.02
R20587 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n34 8.282
R20588 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n21 8.282
R20589 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 5.647
R20590 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 5.316
R20591 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n42 4.141
R20592 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n28 4.141
R20593 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 4.067
R20594 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n11 3.931
R20595 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n40 3.764
R20596 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n33 3.764
R20597 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n24 3.764
R20598 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n19 3.764
R20599 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n36 3.388
R20600 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n22 3.388
R20601 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 3.072
R20602 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 3.072
R20603 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 3.07
R20604 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 3.043
R20605 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 3.033
R20606 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 3.033
R20607 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 3.033
R20608 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n39 2.635
R20609 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n20 2.635
R20610 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 2.362
R20611 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 2.273
R20612 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 2.258
R20613 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 2.258
R20614 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 1.806
R20615 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n30 1.613
R20616 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 1.455
R20617 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 1.192
R20618 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n9 0.752
R20619 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 0.719
R20620 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 0.224
R20621 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 0.175
R20622 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 2.362
R20623 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 1.142
R20624 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 0.994
R20625 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 120.008
R20626 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 92.941
R20627 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n4 92.5
R20628 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 92.462
R20629 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 73.192
R20630 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 72.162
R20631 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 29.482
R20632 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 27.695
R20633 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 27.695
R20634 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 15.46
R20635 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 9.3
R20636 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 9.3
R20637 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n33 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 9.02
R20638 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 9.019
R20639 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n15 8.282
R20640 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 8.282
R20641 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 5.647
R20642 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 5.318
R20643 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n23 4.141
R20644 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n14 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 4.141
R20645 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n34 4.141
R20646 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n27 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n26 4.141
R20647 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 4.033
R20648 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n9 3.931
R20649 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n19 3.764
R20650 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n36 3.764
R20651 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 3.202
R20652 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 3.071
R20653 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 3.071
R20654 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n27 3.07
R20655 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n39 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n38 3.044
R20656 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 3.033
R20657 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n14 3.033
R20658 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 3.033
R20659 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n16 3.011
R20660 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n29 3.011
R20661 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n20 2.635
R20662 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n38 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n37 2.635
R20663 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n39 2.27
R20664 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 2.258
R20665 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n33 2.258
R20666 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 2.25
R20667 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 1.509
R20668 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n7 0.752
R20669 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 2.478
R20670 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 1.148
R20671 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 1.04
R20672 sela.n6 sela.t2 186.373
R20673 sela.n6 sela.t3 170.306
R20674 sela.n7 sela.n6 139.875
R20675 sela.n0 sela.t4 84.832
R20676 sela.n1 sela.t0 84.832
R20677 sela.n1 sela.n0 60.153
R20678 sela.n2 sela.n1 50.163
R20679 sela.n0 sela.t5 48.682
R20680 sela.n1 sela.t1 48.682
R20681 sela.n5 sela 42.917
R20682 sela.n4 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.A 17.167
R20683 sela.n3 sela.n2 15.272
R20684 sela.n5 sela 12.8
R20685 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.A sela 5.315
R20686 sela.n4 sela.n3 4.772
R20687 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.A sela.n3 2.133
R20688 EF_AMUX21m_1.invm_0.A sela 1.77
R20689 sela sela.n7 1.619
R20690 sela.n2 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.A 1.176
R20691 sela sela.n10 0.933
R20692 sela.n7 sela.n5 0.925
R20693 sela.n10 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.A 0.673
R20694 sela.n8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.l0 0.343
R20695 sela.n10 EF_AMUX21m_1.sel 0.321
R20696 sela.n9 sela.n8 0.043
R20697 EF_AMUX21m_1.invm_0.A sela.n4 0.017
R20698 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.A sela.n9 0.014
R20699 sela.n8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.l0 0.001
R20700 sela.n9 EF_AMUX21m_1.array_1ls_1tgm_1.l0 0.001
R20701 vdd1p8.n4 vdd1p8.t9 591.326
R20702 vdd1p8.n6 vdd1p8.t0 591.326
R20703 vdd1p8.n15 vdd1p8.n14 585
R20704 vdd1p8.n97 vdd1p8.n94 321.882
R20705 vdd1p8.n95 vdd1p8.n94 321.882
R20706 vdd1p8.n96 vdd1p8.n95 321.882
R20707 vdd1p8.n36 vdd1p8.n33 321.882
R20708 vdd1p8.n34 vdd1p8.n33 321.882
R20709 vdd1p8.n35 vdd1p8.n34 321.882
R20710 vdd1p8.n99 vdd1p8.n98 175.384
R20711 vdd1p8.n38 vdd1p8.n37 175.384
R20712 vdd1p8.t17 vdd1p8.n97 171.451
R20713 vdd1p8.t5 vdd1p8.n36 171.451
R20714 vdd1p8.n186 vdd1p8.n185 161.37
R20715 vdd1p8.n161 vdd1p8.n160 161.37
R20716 vdd1p8.n137 vdd1p8.n136 161.37
R20717 vdd1p8.n76 vdd1p8.n75 161.37
R20718 vdd1p8.n90 vdd1p8.t18 160.741
R20719 vdd1p8.n29 vdd1p8.t6 160.741
R20720 vdd1p8.n105 vdd1p8.t22 158.223
R20721 vdd1p8.n44 vdd1p8.t16 158.223
R20722 vdd1p8.n9 vdd1p8.t10 148.294
R20723 vdd1p8.t3 vdd1p8.n181 129.545
R20724 vdd1p8.t27 vdd1p8.n156 129.545
R20725 vdd1p8.t13 vdd1p8.n132 129.545
R20726 vdd1p8.t11 vdd1p8.n71 129.545
R20727 vdd1p8.n101 vdd1p8.n100 124.013
R20728 vdd1p8.n40 vdd1p8.n39 124.013
R20729 vdd1p8.n13 vdd1p8.n10 107.745
R20730 vdd1p8.n182 vdd1p8.t3 100.873
R20731 vdd1p8.n157 vdd1p8.t27 100.873
R20732 vdd1p8.n133 vdd1p8.t13 100.873
R20733 vdd1p8.n72 vdd1p8.t11 100.873
R20734 vdd1p8.t21 vdd1p8.n99 96.826
R20735 vdd1p8.t15 vdd1p8.n38 96.826
R20736 vdd1p8.n183 vdd1p8.n181 92.5
R20737 vdd1p8.n181 vdd1p8.n180 92.5
R20738 vdd1p8.n158 vdd1p8.n156 92.5
R20739 vdd1p8.n156 vdd1p8.n155 92.5
R20740 vdd1p8.n134 vdd1p8.n132 92.5
R20741 vdd1p8.n132 vdd1p8.n131 92.5
R20742 vdd1p8.n73 vdd1p8.n71 92.5
R20743 vdd1p8.n71 vdd1p8.n70 92.5
R20744 vdd1p8.n6 vdd1p8.n1 92.5
R20745 vdd1p8.n6 vdd1p8.n5 81.753
R20746 vdd1p8.n100 vdd1p8.t21 81.725
R20747 vdd1p8.n39 vdd1p8.t15 81.725
R20748 vdd1p8.n184 vdd1p8.n180 55.392
R20749 vdd1p8.n159 vdd1p8.n155 55.392
R20750 vdd1p8.n135 vdd1p8.n131 55.392
R20751 vdd1p8.n74 vdd1p8.n70 55.392
R20752 vdd1p8.n9 vdd1p8.n2 52.936
R20753 vdd1p8.n16 vdd1p8.n1 49.593
R20754 vdd1p8.n7 vdd1p8.n6 47.555
R20755 vdd1p8.n181 vdd1p8.t23 47.294
R20756 vdd1p8.n156 vdd1p8.t25 47.294
R20757 vdd1p8.n132 vdd1p8.t7 47.294
R20758 vdd1p8.n71 vdd1p8.t19 47.294
R20759 vdd1p8.n184 vdd1p8.n183 46.25
R20760 vdd1p8.n159 vdd1p8.n158 46.25
R20761 vdd1p8.n135 vdd1p8.n134 46.25
R20762 vdd1p8.n74 vdd1p8.n73 46.25
R20763 vdd1p8.n9 vdd1p8.n8 46.25
R20764 vdd1p8.n7 vdd1p8.n2 42.338
R20765 vdd1p8.n5 vdd1p8.n4 40.877
R20766 vdd1p8.n113 vdd1p8.n93 36.141
R20767 vdd1p8.n113 vdd1p8.n112 36.141
R20768 vdd1p8.n112 vdd1p8.n111 36.141
R20769 vdd1p8.n111 vdd1p8.n101 36.141
R20770 vdd1p8.n52 vdd1p8.n32 36.141
R20771 vdd1p8.n52 vdd1p8.n51 36.141
R20772 vdd1p8.n51 vdd1p8.n50 36.141
R20773 vdd1p8.n50 vdd1p8.n40 36.141
R20774 vdd1p8.n5 vdd1p8.n2 34.416
R20775 vdd1p8.n185 vdd1p8.t4 32.833
R20776 vdd1p8.n185 vdd1p8.t24 32.833
R20777 vdd1p8.n160 vdd1p8.t28 32.833
R20778 vdd1p8.n160 vdd1p8.t26 32.833
R20779 vdd1p8.n136 vdd1p8.t14 32.833
R20780 vdd1p8.n136 vdd1p8.t8 32.833
R20781 vdd1p8.n75 vdd1p8.t12 32.833
R20782 vdd1p8.n75 vdd1p8.t20 32.833
R20783 vdd1p8.n4 vdd1p8.n3 32.004
R20784 vdd1p8.n8 vdd1p8.n3 28.493
R20785 vdd1p8.n3 vdd1p8.n1 28.493
R20786 vdd1p8.n182 vdd1p8.n180 26.469
R20787 vdd1p8.n183 vdd1p8.n182 26.469
R20788 vdd1p8.n157 vdd1p8.n155 26.469
R20789 vdd1p8.n158 vdd1p8.n157 26.469
R20790 vdd1p8.n133 vdd1p8.n131 26.469
R20791 vdd1p8.n134 vdd1p8.n133 26.469
R20792 vdd1p8.n72 vdd1p8.n70 26.469
R20793 vdd1p8.n73 vdd1p8.n72 26.469
R20794 vdd1p8.n12 vdd1p8.t1 22.866
R20795 vdd1p8.n8 vdd1p8.n7 21.169
R20796 vdd1p8.n188 vdd1p8.n187 17.876
R20797 vdd1p8.n163 vdd1p8.n162 17.876
R20798 vdd1p8.n139 vdd1p8.n138 17.876
R20799 vdd1p8.n78 vdd1p8.n77 17.876
R20800 vdd1p8.n187 vdd1p8.n186 17.493
R20801 vdd1p8.n162 vdd1p8.n161 17.493
R20802 vdd1p8.n138 vdd1p8.n137 17.493
R20803 vdd1p8.n77 vdd1p8.n76 17.493
R20804 vdd1p8.n14 vdd1p8.n13 13.512
R20805 vdd1p8.n98 vdd1p8.t17 12.788
R20806 vdd1p8.n37 vdd1p8.t5 12.788
R20807 vdd1p8.n14 vdd1p8.t2 11.433
R20808 vdd1p8.n17 vdd1p8.n16 10.861
R20809 vdd1p8.n91 vdd1p8.n90 9.304
R20810 vdd1p8.n30 vdd1p8.n29 9.304
R20811 vdd1p8.n12 vdd1p8.n11 9.3
R20812 vdd1p8.n97 vdd1p8.n93 8.855
R20813 vdd1p8.n113 vdd1p8.n94 8.855
R20814 vdd1p8.n98 vdd1p8.n94 8.855
R20815 vdd1p8.n112 vdd1p8.n95 8.855
R20816 vdd1p8.n99 vdd1p8.n95 8.855
R20817 vdd1p8.n111 vdd1p8.n96 8.855
R20818 vdd1p8.n36 vdd1p8.n32 8.855
R20819 vdd1p8.n52 vdd1p8.n33 8.855
R20820 vdd1p8.n37 vdd1p8.n33 8.855
R20821 vdd1p8.n51 vdd1p8.n34 8.855
R20822 vdd1p8.n38 vdd1p8.n34 8.855
R20823 vdd1p8.n50 vdd1p8.n35 8.855
R20824 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.VPB vdd1p8.n104 6.323
R20825 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.VPB vdd1p8.n43 6.323
R20826 vdd1p8.n100 vdd1p8.n96 5.535
R20827 vdd1p8.n39 vdd1p8.n35 5.535
R20828 vdd1p8.n186 vdd1p8.n179 4.65
R20829 vdd1p8.n161 vdd1p8.n154 4.65
R20830 vdd1p8.n137 vdd1p8.n130 4.65
R20831 vdd1p8.n76 vdd1p8.n69 4.65
R20832 vdd1p8.n106 vdd1p8.n105 4.65
R20833 vdd1p8.n105 vdd1p8.n102 4.65
R20834 vdd1p8.n90 vdd1p8.n86 4.65
R20835 vdd1p8.n90 vdd1p8.n87 4.65
R20836 vdd1p8.n45 vdd1p8.n44 4.65
R20837 vdd1p8.n44 vdd1p8.n41 4.65
R20838 vdd1p8.n29 vdd1p8.n25 4.65
R20839 vdd1p8.n29 vdd1p8.n26 4.65
R20840 vdd1p8.n175 vdd1p8.n18 4.514
R20841 vdd1p8.n171 vdd1p8.n170 4.514
R20842 vdd1p8.n150 vdd1p8.n58 4.514
R20843 vdd1p8.n146 vdd1p8.n145 4.514
R20844 vdd1p8.n126 vdd1p8.n62 4.514
R20845 vdd1p8.n122 vdd1p8.n121 4.514
R20846 vdd1p8.n89 vdd1p8.n88 4.5
R20847 vdd1p8.n114 vdd1p8.n85 4.5
R20848 vdd1p8.n116 vdd1p8.n115 4.5
R20849 vdd1p8.n110 vdd1p8.n109 4.5
R20850 vdd1p8.n108 vdd1p8.n107 4.5
R20851 EF_AMUX21m_1.invm_0.vdd3p3 vdd1p8.n104 4.5
R20852 vdd1p8.n28 vdd1p8.n27 4.5
R20853 vdd1p8.n53 vdd1p8.n24 4.5
R20854 vdd1p8.n55 vdd1p8.n54 4.5
R20855 vdd1p8.n49 vdd1p8.n48 4.5
R20856 vdd1p8.n47 vdd1p8.n46 4.5
R20857 EF_AMUX21m_2.invm_0.vdd3p3 vdd1p8.n43 4.5
R20858 vdd1p8.n187 vdd1p8.n184 4.322
R20859 vdd1p8.n162 vdd1p8.n159 4.322
R20860 vdd1p8.n138 vdd1p8.n135 4.322
R20861 vdd1p8.n77 vdd1p8.n74 4.322
R20862 vdd1p8.n16 vdd1p8.n15 3.764
R20863 vdd1p8.n16 vdd1p8.n9 3.343
R20864 vdd1p8.n194 vdd1p8.n193 3.151
R20865 vdd1p8.n105 vdd1p8.n103 3.099
R20866 vdd1p8.n44 vdd1p8.n42 3.099
R20867 vdd1p8.n93 vdd1p8.n92 3.033
R20868 vdd1p8.n114 vdd1p8.n113 3.033
R20869 vdd1p8.n112 vdd1p8.n84 3.033
R20870 vdd1p8.n111 vdd1p8.n110 3.033
R20871 EF_AMUX21m_1.invm_0.vdd3p3 vdd1p8.n101 3.033
R20872 vdd1p8.n32 vdd1p8.n31 3.033
R20873 vdd1p8.n53 vdd1p8.n52 3.033
R20874 vdd1p8.n51 vdd1p8.n23 3.033
R20875 vdd1p8.n50 vdd1p8.n49 3.033
R20876 EF_AMUX21m_2.invm_0.vdd3p3 vdd1p8.n40 3.033
R20877 vdd1p8.n15 vdd1p8.n10 2.823
R20878 comparator_top_0.DVDD vdd1p8.n17 2.783
R20879 vdd1p8.n11 vdd1p8.n0 2.543
R20880 vdd1p8.n91 vdd1p8.n89 2.307
R20881 vdd1p8.n30 vdd1p8.n28 2.307
R20882 vdd1p8.n189 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vdd1p8 1.929
R20883 vdd1p8.n164 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vdd1p8 1.929
R20884 vdd1p8.n140 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vdd1p8 1.929
R20885 vdd1p8.n79 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vdd1p8 1.929
R20886 vdd1p8.n0 comparator_top_0.sky130_fd_sc_hvl__lsbufhv2lv_1_0.LVPWR 1.827
R20887 vdd1p8.n189 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 1.618
R20888 vdd1p8.n164 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 1.618
R20889 vdd1p8.n140 vdd1p8 1.618
R20890 vdd1p8.n79 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 1.618
R20891 vdd1p8.n13 vdd1p8.n12 1.433
R20892 vdd1p8.n178 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 1.118
R20893 vdd1p8.n153 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 1.118
R20894 vdd1p8.n129 vdd1p8 1.118
R20895 vdd1p8.n68 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 1.118
R20896 vdd1p8.n144 vdd1p8.n143 0.449
R20897 vdd1p8.n193 vdd1p8.n192 0.447
R20898 vdd1p8.n179 vdd1p8.n178 0.416
R20899 vdd1p8.n154 vdd1p8.n153 0.416
R20900 vdd1p8.n130 vdd1p8.n129 0.416
R20901 vdd1p8.n69 vdd1p8.n68 0.416
R20902 vdd1p8.n20 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 0.377
R20903 vdd1p8.n60 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 0.377
R20904 vdd1p8.n64 vdd1p8 0.377
R20905 vdd1p8.n66 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 0.377
R20906 vdd1p8.n11 vdd1p8.n10 0.376
R20907 vdd1p8.n168 vdd1p8.n167 0.327
R20908 vdd1p8.n119 vdd1p8.n82 0.311
R20909 vdd1p8.n142 EF_AMUX21m_1.array_1ls_1tgm_0.vdd1p8 0.271
R20910 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.vdd1p8 vdd1p8.n188 0.267
R20911 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.vdd1p8 vdd1p8.n163 0.267
R20912 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.vdd1p8 vdd1p8.n139 0.267
R20913 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.vdd1p8 vdd1p8.n78 0.267
R20914 vdd1p8.n81 EF_AMUX21m_1.array_1ls_1tgm_1.vdd1p8 0.242
R20915 vdd1p8.n191 EF_AMUX21m_2.array_1ls_1tgm_0.vdd1p8 0.238
R20916 vdd1p8.n166 EF_AMUX21m_2.array_1ls_1tgm_1.vdd1p8 0.234
R20917 vdd1p8.n193 vdd1p8 0.233
R20918 EF_AMUX21m_1.vdd1p8 vdd1p8.n118 0.214
R20919 vdd1p8.n168 vdd1p8.n57 0.193
R20920 vdd1p8.n17 vdd1p8.n0 0.162
R20921 vdd1p8.n188 vdd1p8.n179 0.157
R20922 vdd1p8.n163 vdd1p8.n154 0.157
R20923 vdd1p8.n139 vdd1p8.n130 0.157
R20924 vdd1p8.n78 vdd1p8.n69 0.157
R20925 vdd1p8.n20 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 0.15
R20926 vdd1p8.n60 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 0.15
R20927 vdd1p8.n64 vdd1p8 0.15
R20928 vdd1p8.n66 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.LVPWR 0.15
R20929 vdd1p8.n67 EF_AMUX21m_1.array_1ls_1tgm_1.vdd1p8 0.141
R20930 vdd1p8.n127 EF_AMUX21m_1.array_1ls_1tgm_0.vdd1p8 0.14
R20931 vdd1p8.n176 EF_AMUX21m_2.array_1ls_1tgm_0.vdd1p8 0.124
R20932 vdd1p8.n151 EF_AMUX21m_2.array_1ls_1tgm_1.vdd1p8 0.121
R20933 vdd1p8.n169 EF_AMUX21m_2.vdd1p8 0.112
R20934 vdd1p8.n120 vdd1p8.n119 0.109
R20935 vdd1p8.n67 vdd1p8.n66 0.093
R20936 vdd1p8.n190 vdd1p8.n189 0.071
R20937 vdd1p8.n165 vdd1p8.n164 0.071
R20938 vdd1p8.n141 vdd1p8.n140 0.071
R20939 vdd1p8.n80 vdd1p8.n79 0.071
R20940 vdd1p8.n109 vdd1p8.n83 0.07
R20941 vdd1p8.n48 vdd1p8.n22 0.07
R20942 vdd1p8.n117 vdd1p8.n116 0.047
R20943 vdd1p8.n56 vdd1p8.n55 0.047
R20944 vdd1p8.n21 vdd1p8.n20 0.046
R20945 vdd1p8.n61 vdd1p8.n60 0.046
R20946 vdd1p8.n65 vdd1p8.n64 0.046
R20947 vdd1p8.n192 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd1p8 0.045
R20948 vdd1p8.n167 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd1p8 0.045
R20949 vdd1p8.n82 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd1p8 0.045
R20950 vdd1p8.n143 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd1p8 0.045
R20951 vdd1p8.n68 vdd1p8.n67 0.04
R20952 vdd1p8.n178 vdd1p8.n177 0.039
R20953 vdd1p8.n153 vdd1p8.n152 0.039
R20954 vdd1p8.n129 vdd1p8.n128 0.039
R20955 vdd1p8.n89 vdd1p8.n85 0.039
R20956 vdd1p8.n116 vdd1p8.n85 0.039
R20957 vdd1p8.n109 vdd1p8.n108 0.039
R20958 vdd1p8.n108 vdd1p8.n104 0.039
R20959 vdd1p8.n28 vdd1p8.n24 0.039
R20960 vdd1p8.n55 vdd1p8.n24 0.039
R20961 vdd1p8.n48 vdd1p8.n47 0.039
R20962 vdd1p8.n47 vdd1p8.n43 0.039
R20963 vdd1p8.n173 vdd1p8.n172 0.035
R20964 vdd1p8.n148 vdd1p8.n147 0.035
R20965 vdd1p8.n124 vdd1p8.n123 0.035
R20966 vdd1p8.n177 vdd1p8.n18 0.035
R20967 vdd1p8.n173 vdd1p8.n18 0.035
R20968 vdd1p8.n172 vdd1p8.n171 0.035
R20969 vdd1p8.n171 vdd1p8.n21 0.035
R20970 vdd1p8.n152 vdd1p8.n58 0.035
R20971 vdd1p8.n148 vdd1p8.n58 0.035
R20972 vdd1p8.n147 vdd1p8.n146 0.035
R20973 vdd1p8.n146 vdd1p8.n61 0.035
R20974 vdd1p8.n128 vdd1p8.n62 0.035
R20975 vdd1p8.n124 vdd1p8.n62 0.035
R20976 vdd1p8.n123 vdd1p8.n122 0.035
R20977 vdd1p8.n122 vdd1p8.n65 0.035
R20978 vdd1p8.n115 vdd1p8.n114 0.028
R20979 vdd1p8.n115 vdd1p8.n84 0.028
R20980 vdd1p8.n107 EF_AMUX21m_1.invm_0.vdd3p3 0.028
R20981 vdd1p8.n54 vdd1p8.n53 0.028
R20982 vdd1p8.n54 vdd1p8.n23 0.028
R20983 vdd1p8.n46 EF_AMUX21m_2.invm_0.vdd3p3 0.028
R20984 vdd1p8.n190 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd1p8 0.027
R20985 vdd1p8.n165 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd1p8 0.027
R20986 vdd1p8.n141 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.vdd1p8 0.027
R20987 vdd1p8.n80 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.lsm_0.vdd1p8 0.027
R20988 vdd1p8.n110 vdd1p8.n102 0.026
R20989 vdd1p8.n106 EF_AMUX21m_1.invm_0.sky130_fd_sc_hvl__inv_2_0.VPB 0.026
R20990 vdd1p8.n49 vdd1p8.n41 0.026
R20991 vdd1p8.n45 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.VPB 0.026
R20992 vdd1p8.n88 vdd1p8.n87 0.025
R20993 vdd1p8.n27 vdd1p8.n26 0.025
R20994 vdd1p8.n194 comparator_top_0.DVDD 0.025
R20995 comparator_top_0.DVDD vdd1p8.n194 0.025
R20996 vdd1p8.n102 vdd1p8.n83 0.023
R20997 vdd1p8.n41 vdd1p8.n22 0.023
R20998 vdd1p8.n125 vdd1p8.n63 0.023
R20999 vdd1p8.n149 vdd1p8.n59 0.02
R21000 vdd1p8.n174 vdd1p8.n19 0.02
R21001 vdd1p8.n143 vdd1p8.n142 0.017
R21002 vdd1p8.n82 vdd1p8.n81 0.016
R21003 vdd1p8.n167 vdd1p8.n166 0.016
R21004 vdd1p8.n192 vdd1p8.n191 0.016
R21005 vdd1p8.n110 vdd1p8.n103 0.014
R21006 vdd1p8.n49 vdd1p8.n42 0.014
R21007 vdd1p8.n88 vdd1p8.n86 0.014
R21008 vdd1p8.n27 vdd1p8.n25 0.014
R21009 vdd1p8.n107 vdd1p8.n103 0.014
R21010 vdd1p8.n46 vdd1p8.n42 0.014
R21011 vdd1p8.n114 vdd1p8.n86 0.013
R21012 vdd1p8.n53 vdd1p8.n25 0.013
R21013 vdd1p8.n127 vdd1p8.n126 0.009
R21014 vdd1p8.n121 vdd1p8.n63 0.009
R21015 vdd1p8.n126 vdd1p8.n125 0.009
R21016 vdd1p8.n121 vdd1p8.n120 0.009
R21017 vdd1p8.n175 vdd1p8.n174 0.008
R21018 vdd1p8.n170 vdd1p8.n19 0.008
R21019 vdd1p8.n150 vdd1p8.n149 0.008
R21020 vdd1p8.n145 vdd1p8.n59 0.008
R21021 vdd1p8.n151 vdd1p8.n150 0.008
R21022 vdd1p8.n145 vdd1p8.n144 0.008
R21023 vdd1p8.n176 vdd1p8.n175 0.008
R21024 vdd1p8.n170 vdd1p8.n169 0.008
R21025 EF_AMUX21m_2.vdd1p8 vdd1p8.n168 0.008
R21026 vdd1p8.n117 vdd1p8.n84 0.005
R21027 vdd1p8.n56 vdd1p8.n23 0.005
R21028 vdd1p8.n119 EF_AMUX21m_1.vdd1p8 0.004
R21029 vdd1p8.n92 vdd1p8.n91 0.003
R21030 vdd1p8.n31 vdd1p8.n30 0.003
R21031 vdd1p8.n92 vdd1p8.n87 0.001
R21032 vdd1p8.n31 vdd1p8.n26 0.001
R21033 EF_AMUX21m_1.invm_0.vdd3p3 vdd1p8.n106 0.001
R21034 EF_AMUX21m_2.invm_0.vdd3p3 vdd1p8.n45 0.001
R21035 vdd1p8.n118 vdd1p8.n83 0.001
R21036 vdd1p8.n57 vdd1p8.n22 0.001
R21037 vdd1p8.n118 vdd1p8.n117 0.001
R21038 vdd1p8.n57 vdd1p8.n56 0.001
R21039 vdd1p8.n177 vdd1p8.n176 0.001
R21040 vdd1p8.n169 vdd1p8.n21 0.001
R21041 vdd1p8.n191 vdd1p8.n190 0.001
R21042 vdd1p8.n166 vdd1p8.n165 0.001
R21043 vdd1p8.n152 vdd1p8.n151 0.001
R21044 vdd1p8.n149 vdd1p8.n148 0.001
R21045 vdd1p8.n147 vdd1p8.n59 0.001
R21046 vdd1p8.n144 vdd1p8.n61 0.001
R21047 vdd1p8.n142 vdd1p8.n141 0.001
R21048 vdd1p8.n128 vdd1p8.n127 0.001
R21049 vdd1p8.n120 vdd1p8.n65 0.001
R21050 vdd1p8.n81 vdd1p8.n80 0.001
R21051 vdd1p8.n125 vdd1p8.n124 0.001
R21052 vdd1p8.n123 vdd1p8.n63 0.001
R21053 vdd1p8.n172 vdd1p8.n19 0.001
R21054 vdd1p8.n174 vdd1p8.n173 0.001
R21055 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 120.008
R21056 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 92.941
R21057 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n4 92.5
R21058 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 92.462
R21059 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 73.192
R21060 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 72.162
R21061 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 29.482
R21062 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 27.695
R21063 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 27.695
R21064 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n5 15.46
R21065 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 9.3
R21066 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n11 9.3
R21067 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n21 9.02
R21068 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n29 9.019
R21069 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n26 8.282
R21070 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n16 8.282
R21071 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 5.647
R21072 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 5.32
R21073 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 5.318
R21074 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n31 4.141
R21075 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n23 4.141
R21076 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n19 4.141
R21077 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 4.033
R21078 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n9 3.931
R21079 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n33 3.764
R21080 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n14 3.764
R21081 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n25 3.202
R21082 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 3.071
R21083 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 3.044
R21084 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 3.033
R21085 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n20 3.033
R21086 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 3.033
R21087 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n27 3.011
R21088 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n17 3.011
R21089 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n34 2.635
R21090 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n15 2.635
R21091 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n36 2.27
R21092 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n30 2.258
R21093 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n22 2.258
R21094 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n6 1.509
R21095 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n7 0.752
R21096 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n0 2.478
R21097 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n1 1.148
R21098 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.n2 1.04
R21099 a_5299_620.n30 a_5299_620.t9 129.036
R21100 a_5299_620.n30 a_5299_620.t8 68.966
R21101 a_5299_620.n50 a_5299_620.n14 10.325
R21102 a_5299_620.n50 a_5299_620.n49 9.572
R21103 a_5299_620.n16 a_5299_620.n15 8.042
R21104 a_5299_620.n1 a_5299_620.n23 7.451
R21105 a_5299_620.n39 a_5299_620.n37 5.629
R21106 a_5299_620.n27 a_5299_620.t7 5.539
R21107 a_5299_620.n27 a_5299_620.t6 5.539
R21108 a_5299_620.n40 a_5299_620.t2 5.539
R21109 a_5299_620.n40 a_5299_620.t5 5.539
R21110 a_5299_620.n3 a_5299_620.n16 4.543
R21111 a_5299_620.n2 a_5299_620.n26 4.5
R21112 a_5299_620.n13 a_5299_620.n43 4.5
R21113 a_5299_620.n12 a_5299_620.n35 4.5
R21114 a_5299_620.n3 a_5299_620.n18 4.5
R21115 a_5299_620.n0 a_5299_620.n45 4.5
R21116 a_5299_620.n0 a_5299_620.n47 4.5
R21117 a_5299_620.n26 a_5299_620.n24 4.141
R21118 a_5299_620.n31 a_5299_620.n29 3.822
R21119 a_5299_620.n43 a_5299_620.n42 3.764
R21120 a_5299_620.n35 a_5299_620.n32 3.388
R21121 a_5299_620.n11 a_5299_620.n10 3.381
R21122 a_5299_620.n20 a_5299_620.t4 3.306
R21123 a_5299_620.n20 a_5299_620.t3 3.306
R21124 a_5299_620.t1 a_5299_620.n50 3.306
R21125 a_5299_620.n50 a_5299_620.t0 3.306
R21126 a_5299_620.n0 a_5299_620.n44 4.34
R21127 a_5299_620.n5 a_5299_620.n20 3.206
R21128 a_5299_620.n35 a_5299_620.n34 3.011
R21129 a_5299_620.n1 a_5299_620.n22 2.635
R21130 a_5299_620.n43 a_5299_620.n41 2.635
R21131 a_5299_620.n18 a_5299_620.n17 2.635
R21132 a_5299_620.n31 a_5299_620.n30 2.421
R21133 a_5299_620.n47 a_5299_620.n46 2.258
R21134 a_5299_620.n28 a_5299_620.n27 2.122
R21135 a_5299_620.n44 a_5299_620.n13 3.118
R21136 a_5299_620.n13 a_5299_620.n40 1.903
R21137 a_5299_620.n11 a_5299_620.n9 1.882
R21138 a_5299_620.n50 a_5299_620.n48 1.525
R21139 a_5299_620.n50 a_5299_620.n19 1.525
R21140 a_5299_620.n26 a_5299_620.n25 1.505
R21141 a_5299_620.n4 a_5299_620.n7 6
R21142 a_5299_620.n7 a_5299_620.n6 1.129
R21143 a_5299_620.n29 a_5299_620.n2 0.922
R21144 a_5299_620.n31 a_5299_620.n21 0.82
R21145 a_5299_620.n9 a_5299_620.n8 0.752
R21146 a_5299_620.n21 a_5299_620.n5 0.699
R21147 a_5299_620.n44 a_5299_620.n31 0.502
R21148 a_5299_620.n36 a_5299_620.n39 0.278
R21149 a_5299_620.n37 a_5299_620.n38 0.161
R21150 a_5299_620.n32 a_5299_620.n33 0.15
R21151 a_5299_620.n13 a_5299_620.n12 0.139
R21152 a_5299_620.n12 a_5299_620.n36 0.132
R21153 a_5299_620.n4 a_5299_620.n5 0.093
R21154 a_5299_620.n2 a_5299_620.n1 4.632
R21155 a_5299_620.n11 a_5299_620.n4 6.074
R21156 a_5299_620.n48 a_5299_620.n0 1.061
R21157 a_5299_620.n19 a_5299_620.n3 0.978
R21158 a_5299_620.n2 a_5299_620.n28 0.419
R21159 a1.n59 a1.n58 185
R21160 a1.n57 a1.n50 185
R21161 a1.n17 a1.n8 185
R21162 a1.n16 a1.n15 185
R21163 a1.n62 a1.t4 120.035
R21164 a1.t5 a1.n7 120.035
R21165 a1.n52 a1.n50 112.829
R21166 a1.n15 a1.n14 112.829
R21167 a1.n61 a1.n60 104.172
R21168 a1.n20 a1.n19 104.172
R21169 a1.n61 a1.n49 92.5
R21170 a1.n21 a1.n20 92.5
R21171 a1.t4 a1.n61 66.827
R21172 a1.n20 a1.t5 66.827
R21173 a1.n76 a1.t0 35.203
R21174 a1.n73 a1.t1 34.056
R21175 a1.n60 a1.n59 29.482
R21176 a1.n19 a1.n8 29.482
R21177 a1.n71 a1.t6 27.695
R21178 a1.n71 a1.t7 27.695
R21179 a1.n38 a1.n37 19.093
R21180 a1.n62 a1.n49 15.455
R21181 a1.n21 a1.n7 15.455
R21182 a1.n57 a1.n56 13.552
R21183 a1.n16 a1.n11 13.552
R21184 a1.n72 a1.n71 9.676
R21185 a1.n34 a1.n27 9.305
R21186 a1.n52 a1.n51 9.304
R21187 a1.n14 a1.n13 9.304
R21188 a1.n33 a1.n32 9.3
R21189 a1.n39 a1.n38 9.3
R21190 a1.n64 a1.n63 9.3
R21191 a1.n48 a1.n45 9.3
R21192 a1.n60 a1.n48 9.3
R21193 a1.n56 a1.n55 9.3
R21194 a1.n65 a1.n47 9.3
R21195 a1.n22 a1.n6 9.3
R21196 a1.n18 a1.n4 9.3
R21197 a1.n19 a1.n18 9.3
R21198 a1.n11 a1.n10 9.3
R21199 a1.n24 a1.n23 9.3
R21200 a1.n64 a1.n49 9.035
R21201 a1.n22 a1.n21 9.035
R21202 a1.n36 a1.n34 8.493
R21203 a1.n36 a1.t2 8.265
R21204 a1.n36 a1.t3 8.265
R21205 a1.n37 a1.n36 7.977
R21206 a1.n35 a1.n33 7.266
R21207 a1.n36 a1.n35 6.152
R21208 a1.n58 a1.n48 5.647
R21209 a1.n18 a1.n17 5.647
R21210 a1.n34 a1.n28 4.894
R21211 a1.n53 a1.n52 4.894
R21212 a1.n14 a1.n12 4.894
R21213 a1.n66 a1.n48 4.517
R21214 a1.n65 a1.n64 4.517
R21215 a1.n18 a1.n5 4.517
R21216 a1.n23 a1.n22 4.517
R21217 a1.n75 a1.n74 4.5
R21218 a1.n74 a1.n72 4.5
R21219 a1.n44 a1.n2 4.5
R21220 a1.n42 a1.n2 4.5
R21221 a1.n44 a1.n43 4.5
R21222 a1.n43 a1.n42 4.5
R21223 a1.n67 a1.n46 4.5
R21224 a1.n68 a1.n1 4.5
R21225 a1.n46 a1.n1 4.5
R21226 a1.n68 a1.n67 4.5
R21227 a1.n41 a1.n25 4.5
R21228 a1.n40 a1.n29 4.5
R21229 a1.n41 a1.n40 4.5
R21230 a1.n29 a1.n25 4.5
R21231 a1.n31 a1.n26 4.5
R21232 a1.n59 a1.n50 3.931
R21233 a1.n15 a1.n8 3.931
R21234 a1.n12 a1.n2 3.033
R21235 a1.n43 a1.n5 3.033
R21236 a1.n53 a1.n1 3.033
R21237 a1.n67 a1.n66 3.033
R21238 a1.n40 a1.n28 3.033
R21239 a1.n73 a1.n70 2.27
R21240 a1.n13 a1.n3 2.252
R21241 a1.n51 a1.n0 2.252
R21242 a1.n27 a1.n26 2.251
R21243 a1.n30 a1.n26 2.244
R21244 a1.n66 a1.n65 1.882
R21245 a1.n23 a1.n5 1.882
R21246 a1.n38 a1.n28 1.505
R21247 a1.n56 a1.n53 1.505
R21248 a1.n12 a1.n11 1.505
R21249 a1.n9 a1.n3 1.492
R21250 a1.n54 a1.n0 1.492
R21251 a1.n63 a1.n62 1.491
R21252 a1.n7 a1.n6 1.49
R21253 a1.n58 a1.n57 0.752
R21254 a1.n17 a1.n16 0.752
R21255 a1.n37 a1.n33 0.521
R21256 a1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.in0 0.349
R21257 a1.n77 a1.n76 0.297
R21258 a1.n42 a1.n41 0.238
R21259 EF_AMUX21m_1.a EF_AMUX21m_1.array_1ls_1tgm_1.in0 0.238
R21260 EF_AMUX21m_1.array_1ls_1tgm_1.in0 a1 0.213
R21261 a1.n77 a1.n69 0.195
R21262 a1 a1.n77 0.185
R21263 a1.n76 a1.n75 0.149
R21264 a1.n68 a1.n44 0.124
R21265 a1.n35 a1.n25 0.057
R21266 a1 EF_AMUX21m_1.a 0.05
R21267 a1.n78 a1 0.043
R21268 a1 a1.n78 0.042
R21269 a1.n55 a1.n54 0.038
R21270 a1.n10 a1.n9 0.037
R21271 a1.n39 a1.n30 0.03
R21272 a1.n75 a1.n70 0.027
R21273 a1.n32 a1.n30 0.025
R21274 a1.n54 a1.n45 0.019
R21275 a1.n9 a1.n4 0.019
R21276 a1.n44 a1.n3 0.016
R21277 a1.n29 a1.n26 0.015
R21278 a1.n67 a1.n45 0.012
R21279 a1.n63 a1.n47 0.012
R21280 a1.n43 a1.n4 0.012
R21281 a1.n24 a1.n6 0.012
R21282 a1.n31 a1.n25 0.011
R21283 a1.n51 a1.n1 0.01
R21284 a1.n13 a1.n2 0.01
R21285 a1.n69 a1.n0 0.009
R21286 a1.n40 a1.n27 0.009
R21287 a1.n67 a1.n47 0.005
R21288 a1.n43 a1.n24 0.005
R21289 a1.n40 a1.n39 0.004
R21290 a1.n55 a1.n1 0.004
R21291 a1.n10 a1.n2 0.004
R21292 a1.n46 a1.n0 0.004
R21293 a1.n69 a1.n68 0.004
R21294 a1.n72 a1.n70 0.003
R21295 a1.n32 a1.n31 0.003
R21296 a1.n41 a1.n26 0.002
R21297 a1.n74 a1.n73 0.001
R21298 a1.n42 a1.n3 0.001
R21299 a1.n78 a1 0.001
R21300 a_5299_1782.n21 a_5299_1782.t8 60.25
R21301 a_5299_1782.n42 a_5299_1782.t9 60.25
R21302 a_5299_1782.n64 a_5299_1782.t0 60.25
R21303 a_5299_1782.n76 a_5299_1782.t2 60.25
R21304 a_5299_1782.n2 a_5299_1782.n84 9.3
R21305 a_5299_1782.n2 a_5299_1782.n85 9.3
R21306 a_5299_1782.n2 a_5299_1782.n83 9.3
R21307 a_5299_1782.n83 a_5299_1782.n82 9.3
R21308 a_5299_1782.n3 a_5299_1782.n73 9.3
R21309 a_5299_1782.n4 a_5299_1782.n57 9.3
R21310 a_5299_1782.n4 a_5299_1782.n56 9.3
R21311 a_5299_1782.n4 a_5299_1782.n63 9.3
R21312 a_5299_1782.n63 a_5299_1782.n62 9.3
R21313 a_5299_1782.n3 a_5299_1782.n72 9.3
R21314 a_5299_1782.n72 a_5299_1782.n71 9.3
R21315 a_5299_1782.n3 a_5299_1782.n74 9.3
R21316 a_5299_1782.n5 a_5299_1782.n51 9.3
R21317 a_5299_1782.n6 a_5299_1782.n35 9.3
R21318 a_5299_1782.n6 a_5299_1782.n34 9.3
R21319 a_5299_1782.n6 a_5299_1782.n41 9.3
R21320 a_5299_1782.n41 a_5299_1782.n40 9.3
R21321 a_5299_1782.n5 a_5299_1782.n50 9.3
R21322 a_5299_1782.n50 a_5299_1782.n49 9.3
R21323 a_5299_1782.n5 a_5299_1782.n52 9.3
R21324 a_5299_1782.n7 a_5299_1782.n29 9.3
R21325 a_5299_1782.n7 a_5299_1782.n28 9.3
R21326 a_5299_1782.n28 a_5299_1782.n27 9.3
R21327 a_5299_1782.n7 a_5299_1782.n30 9.3
R21328 a_5299_1782.n1 a_5299_1782.n91 9.3
R21329 a_5299_1782.n119 a_5299_1782.n118 10.742
R21330 a_5299_1782.n65 a_5299_1782.n64 8.764
R21331 a_5299_1782.n43 a_5299_1782.n42 8.764
R21332 a_5299_1782.n26 a_5299_1782.n25 7.453
R21333 a_5299_1782.n39 a_5299_1782.n38 7.453
R21334 a_5299_1782.n48 a_5299_1782.n47 7.453
R21335 a_5299_1782.n61 a_5299_1782.n60 7.453
R21336 a_5299_1782.n70 a_5299_1782.n69 7.453
R21337 a_5299_1782.n81 a_5299_1782.n80 7.453
R21338 a_5299_1782.n22 a_5299_1782.n21 6.8
R21339 a_5299_1782.n77 a_5299_1782.n76 6.8
R21340 a_5299_1782.n24 a_5299_1782.n23 5.647
R21341 a_5299_1782.n37 a_5299_1782.n36 5.647
R21342 a_5299_1782.n46 a_5299_1782.n45 5.647
R21343 a_5299_1782.n59 a_5299_1782.n58 5.647
R21344 a_5299_1782.n68 a_5299_1782.n67 5.647
R21345 a_5299_1782.n79 a_5299_1782.n78 5.647
R21346 a_5299_1782.n96 a_5299_1782.t1 5.539
R21347 a_5299_1782.n96 a_5299_1782.t3 5.539
R21348 a_5299_1782.n90 a_5299_1782.n89 4.955
R21349 a_5299_1782.n31 a_5299_1782.n20 4.735
R21350 a_5299_1782.n53 a_5299_1782.n19 4.735
R21351 a_5299_1782.n75 a_5299_1782.n18 4.735
R21352 a_5299_1782.n33 a_5299_1782.n32 4.735
R21353 a_5299_1782.n55 a_5299_1782.n54 4.735
R21354 a_5299_1782.n87 a_5299_1782.n86 4.735
R21355 a_5299_1782.n11 a_5299_1782.n13 4.662
R21356 a_5299_1782.n66 a_5299_1782.n65 4.65
R21357 a_5299_1782.n44 a_5299_1782.n43 4.65
R21358 a_5299_1782.n1 a_5299_1782.n17 4.5
R21359 a_5299_1782.n13 a_5299_1782.n99 4.5
R21360 a_5299_1782.n12 a_5299_1782.n95 4.5
R21361 a_5299_1782.n8 a_5299_1782.n110 4.5
R21362 a_5299_1782.n0 a_5299_1782.n105 4.5
R21363 a_5299_1782.n10 a_5299_1782.n117 4.5
R21364 a_5299_1782.n9 a_5299_1782.n114 4.5
R21365 a_5299_1782.n9 a_5299_1782.n112 4.5
R21366 a_5299_1782.n110 a_5299_1782.n109 4.141
R21367 a_5299_1782.n99 a_5299_1782.n98 3.764
R21368 a_5299_1782.n114 a_5299_1782.n113 3.764
R21369 a_5299_1782.n7 a_5299_1782.n22 3.427
R21370 a_5299_1782.n2 a_5299_1782.n77 3.427
R21371 a_5299_1782.n95 a_5299_1782.n93 3.388
R21372 a_5299_1782.n17 a_5299_1782.n16 3.388
R21373 a_5299_1782.n106 a_5299_1782.t5 3.306
R21374 a_5299_1782.n106 a_5299_1782.t4 3.306
R21375 a_5299_1782.n119 a_5299_1782.t6 3.306
R21376 a_5299_1782.t7 a_5299_1782.n119 3.306
R21377 a_5299_1782.n95 a_5299_1782.n94 3.011
R21378 a_5299_1782.n17 a_5299_1782.n15 3.011
R21379 a_5299_1782.n119 a_5299_1782.n100 2.662
R21380 a_5299_1782.n99 a_5299_1782.n97 2.635
R21381 a_5299_1782.n104 a_5299_1782.n103 2.258
R21382 a_5299_1782.n116 a_5299_1782.n115 2.258
R21383 a_5299_1782.n9 a_5299_1782.n11 1.681
R21384 a_5299_1782.n107 a_5299_1782.n106 1.467
R21385 a_5299_1782.n27 a_5299_1782.n26 0.993
R21386 a_5299_1782.n40 a_5299_1782.n39 0.993
R21387 a_5299_1782.n49 a_5299_1782.n48 0.993
R21388 a_5299_1782.n62 a_5299_1782.n61 0.993
R21389 a_5299_1782.n71 a_5299_1782.n70 0.993
R21390 a_5299_1782.n82 a_5299_1782.n81 0.993
R21391 a_5299_1782.n28 a_5299_1782.n24 0.752
R21392 a_5299_1782.n41 a_5299_1782.n37 0.752
R21393 a_5299_1782.n50 a_5299_1782.n46 0.752
R21394 a_5299_1782.n63 a_5299_1782.n59 0.752
R21395 a_5299_1782.n72 a_5299_1782.n68 0.752
R21396 a_5299_1782.n83 a_5299_1782.n79 0.752
R21397 a_5299_1782.n102 a_5299_1782.n101 0.602
R21398 a_5299_1782.n119 a_5299_1782.n10 2.109
R21399 a_5299_1782.n0 a_5299_1782.n107 0.552
R21400 a_5299_1782.n33 a_5299_1782.n31 0.456
R21401 a_5299_1782.n55 a_5299_1782.n53 0.456
R21402 a_5299_1782.n13 a_5299_1782.n96 1.904
R21403 a_5299_1782.n11 a_5299_1782.n102 0.71
R21404 a_5299_1782.n110 a_5299_1782.n108 0.376
R21405 a_5299_1782.n105 a_5299_1782.n104 0.376
R21406 a_5299_1782.n112 a_5299_1782.n111 0.376
R21407 a_5299_1782.n117 a_5299_1782.n116 0.376
R21408 a_5299_1782.n88 a_5299_1782.n75 0.228
R21409 a_5299_1782.n88 a_5299_1782.n87 0.228
R21410 a_5299_1782.n90 a_5299_1782.n88 0.214
R21411 a_5299_1782.n31 a_5299_1782.n7 0.203
R21412 a_5299_1782.n6 a_5299_1782.n33 0.203
R21413 a_5299_1782.n53 a_5299_1782.n5 0.203
R21414 a_5299_1782.n4 a_5299_1782.n55 0.203
R21415 a_5299_1782.n75 a_5299_1782.n3 0.203
R21416 a_5299_1782.n87 a_5299_1782.n2 0.203
R21417 a_5299_1782.n44 a_5299_1782.n6 0.19
R21418 a_5299_1782.n5 a_5299_1782.n44 0.19
R21419 a_5299_1782.n66 a_5299_1782.n4 0.19
R21420 a_5299_1782.n3 a_5299_1782.n66 0.19
R21421 a_5299_1782.n8 a_5299_1782.n0 0.177
R21422 a_5299_1782.n12 a_5299_1782.n1 0.164
R21423 a_5299_1782.n15 a_5299_1782.n14 0.161
R21424 a_5299_1782.n93 a_5299_1782.n92 0.15
R21425 a_5299_1782.n1 a_5299_1782.n90 0.139
R21426 a_5299_1782.n13 a_5299_1782.n12 0.137
R21427 a_5299_1782.n10 a_5299_1782.n9 0.132
R21428 a_5299_1782.n102 a_5299_1782.n8 0.102
R21429 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 136.803
R21430 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 136.324
R21431 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 119.998
R21432 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 93.901
R21433 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 93.303
R21434 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 93.083
R21435 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n4 92.5
R21436 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 92.462
R21437 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 69.227
R21438 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 29.482
R21439 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 27.695
R21440 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 27.695
R21441 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n5 15.462
R21442 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n16 9.3
R21443 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n8 9.3
R21444 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n7 9.3
R21445 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 9.3
R21446 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n13 9.3
R21447 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n15 9.3
R21448 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n17 9.3
R21449 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n43 9.02
R21450 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n26 9.02
R21451 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n34 8.282
R21452 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n21 8.282
R21453 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n14 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 5.647
R21454 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 5.316
R21455 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n42 4.141
R21456 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n28 4.141
R21457 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 4.067
R21458 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n11 3.931
R21459 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n40 3.764
R21460 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n33 3.764
R21461 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n24 3.764
R21462 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n19 3.764
R21463 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n36 3.388
R21464 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n22 3.388
R21465 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 3.072
R21466 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n37 3.072
R21467 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n35 3.07
R21468 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 3.043
R21469 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 3.033
R21470 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n25 3.033
R21471 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n23 3.033
R21472 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n41 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n39 2.635
R21473 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n20 2.635
R21474 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n38 2.362
R21475 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n46 2.273
R21476 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n45 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n44 2.258
R21477 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n27 2.258
R21478 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 1.806
R21479 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n30 1.613
R21480 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n6 1.455
R21481 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n31 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n3 1.192
R21482 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n10 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n9 0.752
R21483 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 0.719
R21484 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 0.224
R21485 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n49 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n48 0.175
R21486 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n2 2.362
R21487 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n1 1.142
R21488 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n47 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.n0 0.994
R21489 b2.n59 b2.n58 185
R21490 b2.n57 b2.n50 185
R21491 b2.n17 b2.n8 185
R21492 b2.n16 b2.n15 185
R21493 b2.n62 b2.t6 120.035
R21494 b2.t7 b2.n7 120.035
R21495 b2.n52 b2.n50 112.829
R21496 b2.n15 b2.n14 112.829
R21497 b2.n61 b2.n60 104.172
R21498 b2.n20 b2.n19 104.172
R21499 b2.n61 b2.n49 92.5
R21500 b2.n21 b2.n20 92.5
R21501 b2.t6 b2.n61 66.827
R21502 b2.n20 b2.t7 66.827
R21503 b2.n76 b2.t2 35.203
R21504 b2.n73 b2.t3 34.056
R21505 b2.n60 b2.n59 29.482
R21506 b2.n19 b2.n8 29.482
R21507 b2.n71 b2.t5 27.695
R21508 b2.n71 b2.t4 27.695
R21509 b2.n38 b2.n37 19.093
R21510 b2.n62 b2.n49 15.455
R21511 b2.n21 b2.n7 15.455
R21512 b2.n57 b2.n56 13.552
R21513 b2.n16 b2.n11 13.552
R21514 b2.n72 b2.n71 9.676
R21515 b2.n34 b2.n27 9.305
R21516 b2.n52 b2.n51 9.304
R21517 b2.n14 b2.n13 9.304
R21518 b2.n33 b2.n32 9.3
R21519 b2.n39 b2.n38 9.3
R21520 b2.n64 b2.n63 9.3
R21521 b2.n48 b2.n45 9.3
R21522 b2.n60 b2.n48 9.3
R21523 b2.n56 b2.n55 9.3
R21524 b2.n65 b2.n47 9.3
R21525 b2.n22 b2.n6 9.3
R21526 b2.n18 b2.n4 9.3
R21527 b2.n19 b2.n18 9.3
R21528 b2.n11 b2.n10 9.3
R21529 b2.n24 b2.n23 9.3
R21530 b2.n64 b2.n49 9.035
R21531 b2.n22 b2.n21 9.035
R21532 b2.n36 b2.n34 8.493
R21533 b2.n36 b2.t1 8.265
R21534 b2.n36 b2.t0 8.265
R21535 b2.n37 b2.n36 7.977
R21536 b2.n35 b2.n33 7.266
R21537 b2.n36 b2.n35 6.152
R21538 b2.n58 b2.n48 5.647
R21539 b2.n18 b2.n17 5.647
R21540 b2.n34 b2.n28 4.894
R21541 b2.n53 b2.n52 4.894
R21542 b2.n14 b2.n12 4.894
R21543 b2.n66 b2.n48 4.517
R21544 b2.n65 b2.n64 4.517
R21545 b2.n18 b2.n5 4.517
R21546 b2.n23 b2.n22 4.517
R21547 b2.n75 b2.n74 4.5
R21548 b2.n74 b2.n72 4.5
R21549 b2.n44 b2.n2 4.5
R21550 b2.n42 b2.n2 4.5
R21551 b2.n44 b2.n43 4.5
R21552 b2.n43 b2.n42 4.5
R21553 b2.n67 b2.n46 4.5
R21554 b2.n68 b2.n1 4.5
R21555 b2.n46 b2.n1 4.5
R21556 b2.n68 b2.n67 4.5
R21557 b2.n41 b2.n25 4.5
R21558 b2.n40 b2.n29 4.5
R21559 b2.n41 b2.n40 4.5
R21560 b2.n29 b2.n25 4.5
R21561 b2.n31 b2.n26 4.5
R21562 b2.n59 b2.n50 3.931
R21563 b2.n15 b2.n8 3.931
R21564 b2.n12 b2.n2 3.033
R21565 b2.n43 b2.n5 3.033
R21566 b2.n53 b2.n1 3.033
R21567 b2.n67 b2.n66 3.033
R21568 b2.n40 b2.n28 3.033
R21569 b2.n73 b2.n70 2.27
R21570 b2.n13 b2.n3 2.252
R21571 b2.n51 b2.n0 2.252
R21572 b2.n27 b2.n26 2.251
R21573 b2.n30 b2.n26 2.244
R21574 b2.n66 b2.n65 1.882
R21575 b2.n23 b2.n5 1.882
R21576 b2.n38 b2.n28 1.505
R21577 b2.n56 b2.n53 1.505
R21578 b2.n12 b2.n11 1.505
R21579 b2.n9 b2.n3 1.492
R21580 b2.n54 b2.n0 1.492
R21581 b2.n63 b2.n62 1.491
R21582 b2.n7 b2.n6 1.49
R21583 b2.n58 b2.n57 0.752
R21584 b2.n17 b2.n16 0.752
R21585 b2.n37 b2.n33 0.521
R21586 b2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.in0 0.43
R21587 b2.n77 b2.n76 0.297
R21588 b2.n42 b2.n41 0.238
R21589 EF_AMUX21m_2.array_1ls_1tgm_0.in0 b2 0.213
R21590 b2.n77 b2.n69 0.195
R21591 b2 b2.n77 0.185
R21592 EF_AMUX21m_2.b EF_AMUX21m_2.array_1ls_1tgm_0.in0 0.177
R21593 b2.n76 b2.n75 0.149
R21594 b2.n68 b2.n44 0.124
R21595 EF_AMUX21m_2.b b2 0.099
R21596 b2.n35 b2.n25 0.057
R21597 b2.n55 b2.n54 0.038
R21598 b2.n10 b2.n9 0.037
R21599 b2.n39 b2.n30 0.03
R21600 b2.n75 b2.n70 0.027
R21601 b2.n32 b2.n30 0.025
R21602 b2.n54 b2.n45 0.019
R21603 b2.n9 b2.n4 0.019
R21604 b2.n44 b2.n3 0.016
R21605 b2.n29 b2.n26 0.015
R21606 b2.n67 b2.n45 0.012
R21607 b2.n63 b2.n47 0.012
R21608 b2.n43 b2.n4 0.012
R21609 b2.n24 b2.n6 0.012
R21610 b2.n31 b2.n25 0.011
R21611 b2.n51 b2.n1 0.01
R21612 b2.n13 b2.n2 0.01
R21613 b2.n69 b2.n0 0.009
R21614 b2.n40 b2.n27 0.009
R21615 b2.n67 b2.n47 0.005
R21616 b2.n43 b2.n24 0.005
R21617 b2.n40 b2.n39 0.004
R21618 b2.n55 b2.n1 0.004
R21619 b2.n10 b2.n2 0.004
R21620 b2.n46 b2.n0 0.004
R21621 b2.n69 b2.n68 0.004
R21622 b2.n72 b2.n70 0.003
R21623 b2.n32 b2.n31 0.003
R21624 b2.n41 b2.n26 0.002
R21625 b2.n74 b2.n73 0.001
R21626 b2.n42 b2.n3 0.001
R21627 selb.n6 selb.t4 186.373
R21628 selb.n6 selb.t5 170.306
R21629 selb.n7 selb.n6 139.875
R21630 selb.n0 selb.t1 84.832
R21631 selb.n1 selb.t0 84.832
R21632 selb.n1 selb.n0 60.153
R21633 selb.n2 selb.n1 50.163
R21634 selb.n0 selb.t3 48.682
R21635 selb.n1 selb.t2 48.682
R21636 selb.n5 selb 42.917
R21637 selb.n4 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.A 17.167
R21638 selb.n3 selb.n2 15.272
R21639 selb.n5 selb 12.8
R21640 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.A selb 5.315
R21641 selb.n4 selb.n3 4.772
R21642 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.A selb.n3 2.133
R21643 selb selb.n7 1.619
R21644 EF_AMUX21m_2.invm_0.A selb 1.501
R21645 selb selb.n10 1.236
R21646 selb.n2 EF_AMUX21m_2.invm_0.sky130_fd_sc_hvl__inv_2_0.A 1.176
R21647 selb.n7 selb.n5 0.925
R21648 selb.n10 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.A 0.673
R21649 selb.n8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.l0 0.343
R21650 selb.n10 EF_AMUX21m_2.sel 0.321
R21651 selb.n9 selb.n8 0.043
R21652 EF_AMUX21m_2.invm_0.A selb.n4 0.017
R21653 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.lsm_0.A selb.n9 0.014
R21654 selb.n8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.l0 0.001
R21655 selb.n9 EF_AMUX21m_2.array_1ls_1tgm_1.l0 0.001
R21656 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 120.008
R21657 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 92.941
R21658 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n4 92.5
R21659 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 92.462
R21660 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 73.192
R21661 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 72.162
R21662 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 29.482
R21663 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n29 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 27.695
R21664 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 27.695
R21665 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n5 15.46
R21666 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 9.3
R21667 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n11 9.3
R21668 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n21 9.02
R21669 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n29 9.019
R21670 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n26 8.282
R21671 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n16 8.282
R21672 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n12 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 5.647
R21673 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 5.32
R21674 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 5.318
R21675 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n31 4.141
R21676 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n23 4.141
R21677 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n20 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n19 4.141
R21678 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 4.033
R21679 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n10 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n9 3.931
R21680 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n33 3.764
R21681 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n14 3.764
R21682 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n25 3.202
R21683 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 3.071
R21684 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n36 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 3.044
R21685 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 3.033
R21686 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n20 3.033
R21687 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 3.033
R21688 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n28 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n27 3.011
R21689 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n18 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n17 3.011
R21690 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n35 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n34 2.635
R21691 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n13 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n15 2.635
R21692 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n36 2.27
R21693 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n32 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n30 2.258
R21694 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n24 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n22 2.258
R21695 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n6 1.509
R21696 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n7 0.752
R21697 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n0 2.478
R21698 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n1 1.148
R21699 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.n2 1.04
R21700 a_7196_n5728.n2 a_7196_n5728.t0 333.409
R21701 a_7196_n5728.n1 a_7196_n5728.n0 177.236
R21702 a_7196_n5728.t5 a_7196_n5728.n7 153.872
R21703 a_7196_n5728.n1 a_7196_n5728.t8 139.997
R21704 a_7196_n5728.n0 a_7196_n5728.t7 124.47
R21705 a_7196_n5728.n5 a_7196_n5728.n4 104.473
R21706 a_7196_n5728.n0 a_7196_n5728.t6 88.32
R21707 a_7196_n5728.n2 a_7196_n5728.n1 65.236
R21708 a_7196_n5728.n6 a_7196_n5728.n5 60.509
R21709 a_7196_n5728.n5 a_7196_n5728.n3 43.964
R21710 a_7196_n5728.n6 a_7196_n5728.n2 22.109
R21711 a_7196_n5728.n7 a_7196_n5728.n6 20.908
R21712 a_7196_n5728.n3 a_7196_n5728.t4 10.64
R21713 a_7196_n5728.n3 a_7196_n5728.t1 10.64
R21714 a_7196_n5728.n4 a_7196_n5728.t3 10.64
R21715 a_7196_n5728.n4 a_7196_n5728.t2 10.64
R21716 a2.n59 a2.n58 185
R21717 a2.n57 a2.n50 185
R21718 a2.n17 a2.n8 185
R21719 a2.n16 a2.n15 185
R21720 a2.n62 a2.t0 120.035
R21721 a2.t1 a2.n7 120.035
R21722 a2.n52 a2.n50 112.829
R21723 a2.n15 a2.n14 112.829
R21724 a2.n61 a2.n60 104.172
R21725 a2.n20 a2.n19 104.172
R21726 a2.n61 a2.n49 92.5
R21727 a2.n21 a2.n20 92.5
R21728 a2.t0 a2.n61 66.827
R21729 a2.n20 a2.t1 66.827
R21730 a2.n76 a2.t4 35.203
R21731 a2.n73 a2.t5 34.056
R21732 a2.n60 a2.n59 29.482
R21733 a2.n19 a2.n8 29.482
R21734 a2.n71 a2.t2 27.695
R21735 a2.n71 a2.t3 27.695
R21736 a2.n38 a2.n37 19.093
R21737 a2.n62 a2.n49 15.455
R21738 a2.n21 a2.n7 15.455
R21739 a2.n57 a2.n56 13.552
R21740 a2.n16 a2.n11 13.552
R21741 a2.n72 a2.n71 9.676
R21742 a2.n34 a2.n27 9.305
R21743 a2.n52 a2.n51 9.304
R21744 a2.n14 a2.n13 9.304
R21745 a2.n33 a2.n32 9.3
R21746 a2.n39 a2.n38 9.3
R21747 a2.n64 a2.n63 9.3
R21748 a2.n48 a2.n45 9.3
R21749 a2.n60 a2.n48 9.3
R21750 a2.n56 a2.n55 9.3
R21751 a2.n65 a2.n47 9.3
R21752 a2.n22 a2.n6 9.3
R21753 a2.n18 a2.n4 9.3
R21754 a2.n19 a2.n18 9.3
R21755 a2.n11 a2.n10 9.3
R21756 a2.n24 a2.n23 9.3
R21757 a2.n64 a2.n49 9.035
R21758 a2.n22 a2.n21 9.035
R21759 a2.n36 a2.n34 8.493
R21760 a2.n36 a2.t6 8.265
R21761 a2.n36 a2.t7 8.265
R21762 a2.n37 a2.n36 7.977
R21763 a2.n35 a2.n33 7.266
R21764 a2.n36 a2.n35 6.152
R21765 a2.n58 a2.n48 5.647
R21766 a2.n18 a2.n17 5.647
R21767 a2.n34 a2.n28 4.894
R21768 a2.n53 a2.n52 4.894
R21769 a2.n14 a2.n12 4.894
R21770 a2.n66 a2.n48 4.517
R21771 a2.n65 a2.n64 4.517
R21772 a2.n18 a2.n5 4.517
R21773 a2.n23 a2.n22 4.517
R21774 a2.n75 a2.n74 4.5
R21775 a2.n74 a2.n72 4.5
R21776 a2.n44 a2.n2 4.5
R21777 a2.n42 a2.n2 4.5
R21778 a2.n44 a2.n43 4.5
R21779 a2.n43 a2.n42 4.5
R21780 a2.n67 a2.n46 4.5
R21781 a2.n68 a2.n1 4.5
R21782 a2.n46 a2.n1 4.5
R21783 a2.n68 a2.n67 4.5
R21784 a2.n41 a2.n25 4.5
R21785 a2.n40 a2.n29 4.5
R21786 a2.n41 a2.n40 4.5
R21787 a2.n29 a2.n25 4.5
R21788 a2.n31 a2.n26 4.5
R21789 a2.n59 a2.n50 3.931
R21790 a2.n15 a2.n8 3.931
R21791 a2.n12 a2.n2 3.033
R21792 a2.n43 a2.n5 3.033
R21793 a2.n53 a2.n1 3.033
R21794 a2.n67 a2.n66 3.033
R21795 a2.n40 a2.n28 3.033
R21796 a2.n73 a2.n70 2.27
R21797 a2.n13 a2.n3 2.252
R21798 a2.n51 a2.n0 2.252
R21799 a2.n27 a2.n26 2.251
R21800 a2.n30 a2.n26 2.244
R21801 a2.n66 a2.n65 1.882
R21802 a2.n23 a2.n5 1.882
R21803 a2.n38 a2.n28 1.505
R21804 a2.n56 a2.n53 1.505
R21805 a2.n12 a2.n11 1.505
R21806 a2.n9 a2.n3 1.492
R21807 a2.n54 a2.n0 1.492
R21808 a2.n63 a2.n62 1.491
R21809 a2.n7 a2.n6 1.49
R21810 a2.n58 a2.n57 0.752
R21811 a2.n17 a2.n16 0.752
R21812 a2.n37 a2.n33 0.521
R21813 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.in0 a2 0.368
R21814 a2.n77 a2.n76 0.297
R21815 a2.n42 a2.n41 0.238
R21816 EF_AMUX21m_1.array_1ls_1tgm_0.in0 a2 0.213
R21817 a2.n77 a2.n69 0.195
R21818 a2 a2.n77 0.185
R21819 EF_AMUX21m_1.b EF_AMUX21m_1.array_1ls_1tgm_0.in0 0.177
R21820 a2.n76 a2.n75 0.149
R21821 a2.n78 EF_AMUX21m_1.b 0.136
R21822 a2.n68 a2.n44 0.124
R21823 a2.n35 a2.n25 0.057
R21824 a2.n55 a2.n54 0.038
R21825 a2.n10 a2.n9 0.037
R21826 a2.n39 a2.n30 0.03
R21827 a2.n75 a2.n70 0.027
R21828 a2 a2.n78 0.027
R21829 a2.n78 a2 0.026
R21830 a2.n32 a2.n30 0.025
R21831 a2.n54 a2.n45 0.019
R21832 a2.n9 a2.n4 0.019
R21833 a2.n44 a2.n3 0.016
R21834 a2.n29 a2.n26 0.015
R21835 a2.n67 a2.n45 0.012
R21836 a2.n63 a2.n47 0.012
R21837 a2.n43 a2.n4 0.012
R21838 a2.n24 a2.n6 0.012
R21839 a2.n31 a2.n25 0.011
R21840 a2.n51 a2.n1 0.01
R21841 a2.n13 a2.n2 0.01
R21842 a2.n69 a2.n0 0.009
R21843 a2.n40 a2.n27 0.009
R21844 a2.n67 a2.n47 0.005
R21845 a2.n43 a2.n24 0.005
R21846 a2.n40 a2.n39 0.004
R21847 a2.n55 a2.n1 0.004
R21848 a2.n10 a2.n2 0.004
R21849 a2.n46 a2.n0 0.004
R21850 a2.n69 a2.n68 0.004
R21851 a2.n72 a2.n70 0.003
R21852 a2.n32 a2.n31 0.003
R21853 a2.n41 a2.n26 0.002
R21854 a2.n74 a2.n73 0.001
R21855 a2.n42 a2.n3 0.001
C0 vdd1p8 comparator_top_0.comparator_0.VOUT 0.03fF
C1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_8403_n6064# 0.00fF
C2 vdd3p3 selb 0.06fF
C3 vdd3p3 a_10975_4108# 0.65fF
C4 vdd3p3 a_3816_n5791# 0.57fF
C5 vdd1p8 a2 0.00fF
C6 a2 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.00fF
C7 vdd3p3 a_10811_7187# 0.85fF
C8 a_8403_n6064# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.16fF
C9 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a2 0.39fF
C10 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_11235_n6821# 0.00fF
C11 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_10442_n5795# 0.00fF
C12 a_3816_n5791# a_4609_n6817# 0.00fF
C13 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 7.84fF
C14 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_10442_n5795# 0.01fF
C15 vdd1p8 vo 0.61fF
C16 a1 a_1777_n6060# 0.00fF
C17 a_10442_n5795# a_11235_n6821# 0.00fF
C18 a_8403_n6064# selb 0.00fF
C19 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.00fF
C20 vdd1p8 a_838_n6794# 0.35fF
C21 a_7096_n5816# a_7889_n6842# 0.00fF
C22 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 4.59fF
C23 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp b2 2.03fF
C24 vdd3p3 a_11031_3400# 1.88fF
C25 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y b2 0.00fF
C26 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_7464_n6798# 0.00fF
C27 vdd3p3 a_5123_n6039# 0.73fF
C28 vdd3p3 a_7889_n6842# 1.07fF
C29 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 3.72fF
C30 vss EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.00fF
C31 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 3.64fF
C32 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_11749_n6043# 0.00fF
C33 vdd1p8 a_10965_3602# 0.06fF
C34 vss comparator_top_0.comparator_0.VBP 3.04fF
C35 a_5123_n6039# a_4609_n6817# 0.00fF
C36 a_11749_n6043# a_11235_n6821# 0.00fF
C37 vdd1p8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.13fF
C38 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_3816_n5791# 0.00fF
C39 vdd1p8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 1.50fF
C40 a_8403_n6064# a_7889_n6842# 0.00fF
C41 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_7464_n6798# 0.00fF
C42 vdd3p3 sela 0.06fF
C43 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.48fF
C44 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_10810_n6777# 0.00fF
C45 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 3.44fF
C46 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.31fF
C47 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.00fF
C48 selb a_7464_n6798# 0.03fF
C49 a_11235_n6821# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.01fF
C50 b1 a_7096_n5816# 0.00fF
C51 a2 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C52 vdd3p3 comparator_top_0.comparator_0.VBN 75.35fF
C53 vss vdd1p8 0.01fF
C54 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.38fF
C55 a1 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C56 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.56fF
C57 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_5123_n6039# 0.00fF
C58 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.00fF
C59 vdd3p3 b1 3.98fF
C60 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.48fF
C61 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a2 0.00fF
C62 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y selb 0.00fF
C63 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.32fF
C64 a_11271_4224# a_10975_4108# 0.14fF
C65 vdd3p3 a_7096_n5816# 0.57fF
C66 comparator_top_0.comparator_0.VOUT a_10975_4108# 0.02fF
C67 b1 a_8403_n6064# 0.00fF
C68 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 1.14fF
C69 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a1 1.70fF
C70 a_7889_n6842# a_7464_n6798# 0.63fF
C71 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.18fF
C72 vss a1 0.00fF
C73 a2 a_3816_n5791# 0.00fF
C74 vdd3p3 a_10810_n6777# 0.87fF
C75 vdd3p3 a_6349_9307# 0.65fF
C76 a_11271_4224# a_11031_3400# 0.31fF
C77 a_7096_n5816# a_8403_n6064# 0.00fF
C78 a_470_n5812# sela 0.27fF
C79 vdd1p8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.24fF
C80 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_1263_n6838# 0.00fF
C81 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_4184_n6773# 0.00fF
C82 a_10975_4108# vo 0.29fF
C83 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_7889_n6842# 0.00fF
C84 comparator_top_0.comparator_0.VBN EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 0.16fF
C85 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.01fF
C86 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A a_4184_n6773# 0.03fF
C87 vdd3p3 a_4609_n6817# 1.07fF
C88 comparator_top_0.comparator_0.VOUT a_11031_3400# 0.36fF
C89 vdd3p3 a_8403_n6064# 0.73fF
C90 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_1777_n6060# 0.00fF
C91 a_1263_n6838# sela 0.01fF
C92 vdd1p8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.18fF
C93 vdd1p8 a1 0.00fF
C94 a2 a_5123_n6039# 0.00fF
C95 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb b2 1.71fF
C96 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.18fF
C97 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a2 2.03fF
C98 vdd1p8 a_10442_n5795# 0.72fF
C99 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.00fF
C100 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a2 0.00fF
C101 a_10975_4108# a_10965_3602# 0.39fF
C102 vo a_11031_3400# 0.03fF
C103 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_11235_n6821# 0.00fF
C104 a_1777_n6060# sela 0.00fF
C105 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 7.84fF
C106 a_10809_9307# a_10811_8247# 0.14fF
C107 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.00fF
C108 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C109 vss EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 17.07fF
C110 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.27fF
C111 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 40.25fF
C112 vdd1p8 b2 0.00fF
C113 comparator_top_0.comparator_0.VBP EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 0.01fF
C114 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_4609_n6817# 0.00fF
C115 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_838_n6794# 0.00fF
C116 b1 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00fF
C117 a_7096_n5816# a_7464_n6798# 0.15fF
C118 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y b1 0.47fF
C119 vdd3p3 a_470_n5812# 0.53fF
C120 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C121 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 3.72fF
C122 a_11031_3400# a_10965_3602# 0.24fF
C123 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 1.12fF
C124 vdd1p8 a_11749_n6043# 0.02fF
C125 vdd3p3 a_6351_7717# 0.46fF
C126 vdd3p3 a_7464_n6798# 0.87fF
C127 sela a_838_n6794# 0.03fF
C128 vdd1p8 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.16fF
C129 a_6349_9307# a_6351_7717# 0.14fF
C130 vdd1p8 a_4184_n6773# 0.35fF
C131 b2 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C132 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.38fF
C133 vdd3p3 a_1263_n6838# 1.07fF
C134 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_4184_n6773# 0.00fF
C135 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.38fF
C136 vdd1p8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 1.59fF
C137 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 3.72fF
C138 b2 a_10442_n5795# 0.00fF
C139 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.00fF
C140 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.49fF
C141 a_8403_n6064# a_7464_n6798# 0.00fF
C142 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_10810_n6777# 0.00fF
C143 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 3.64fF
C144 a_11235_n6821# a_10810_n6777# 0.63fF
C145 vdd3p3 a_11235_n6821# 1.07fF
C146 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 1.12fF
C147 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.21fF
C148 vdd3p3 a_11271_4224# 1.24fF
C149 a_11749_n6043# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.16fF
C150 vdd3p3 a_1777_n6060# 0.73fF
C151 vdd1p8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.16fF
C152 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A sela 0.00fF
C153 a_10442_n5795# a_11749_n6043# 0.00fF
C154 vdd3p3 comparator_top_0.comparator_0.VOUT 3.47fF
C155 sela EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.33fF
C156 a_10809_9307# a_10811_7187# 0.00fF
C157 vdd1p8 selb 1.43fF
C158 vdd1p8 a_10975_4108# 1.21fF
C159 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_8403_n6064# 0.00fF
C160 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 1.14fF
C161 vdd1p8 a_3816_n5791# 0.69fF
C162 vdd3p3 a2 3.99fF
C163 vss EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.00fF
C164 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_470_n5812# 0.00fF
C165 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.49fF
C166 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y selb 0.00fF
C167 b2 a_11749_n6043# 0.00fF
C168 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_10442_n5795# 0.00fF
C169 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.27fF
C170 vdd3p3 vo 0.65fF
C171 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_470_n5812# 0.00fF
C172 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.56fF
C173 vdd3p3 a_838_n6794# 0.87fF
C174 vss sela 0.03fF
C175 vdd3p3 a_6351_6657# 0.98fF
C176 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 0.00fF
C177 a_10442_n5795# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C178 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out b2 2.92fF
C179 vdd1p8 a_11031_3400# 0.12fF
C180 vdd1p8 a_5123_n6039# 0.02fF
C181 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_1777_n6060# 0.00fF
C182 vdd1p8 a_7889_n6842# 0.41fF
C183 a_470_n5812# a_1263_n6838# 0.00fF
C184 vss comparator_top_0.comparator_0.VBN 31.64fF
C185 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_4184_n6773# 0.00fF
C186 vdd1p8 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.19fF
C187 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_5123_n6039# 0.00fF
C188 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_11749_n6043# 0.00fF
C189 vdd3p3 a_10965_3602# 0.17fF
C190 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 1.14fF
C191 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.18fF
C192 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a2 1.71fF
C193 comparator_top_0.comparator_0.VBN comparator_top_0.comparator_0.VBP 2.37fF
C194 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.00fF
C195 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 1.72fF
C196 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_7464_n6798# 0.00fF
C197 a_470_n5812# a_1777_n6060# 0.00fF
C198 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_1777_n6060# 0.00fF
C199 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a2 2.92fF
C200 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.06fF
C201 vdd1p8 sela 1.42fF
C202 a_10811_8247# a_10811_7187# 0.14fF
C203 vdd1p8 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.31fF
C204 a_4609_n6817# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.01fF
C205 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.01fF
C206 a1 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00fF
C207 a_1777_n6060# a_1263_n6838# 0.00fF
C208 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a1 0.43fF
C209 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A selb 0.00fF
C210 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.00fF
C211 a_3816_n5791# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C212 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 7.84fF
C213 vdd3p3 vss 329.86fF
C214 a_3816_n5791# a_4184_n6773# 0.15fF
C215 vss a_6349_9307# 0.00fF
C216 selb EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.33fF
C217 vdd3p3 comparator_top_0.comparator_0.VBP 25.50fF
C218 a_470_n5812# a_838_n6794# 0.15fF
C219 vdd1p8 b1 0.00fF
C220 comparator_top_0.comparator_0.VOUT a_11271_4224# 0.01fF
C221 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp b1 2.04fF
C222 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.37fF
C223 a_6351_7717# a_6351_6657# 0.14fF
C224 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y b1 0.00fF
C225 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A selb 0.00fF
C226 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 7.84fF
C227 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 1.15fF
C228 a_1263_n6838# a_838_n6794# 0.63fF
C229 vdd1p8 a_7096_n5816# 0.69fF
C230 vdd3p3 a_10809_9307# 1.14fF
C231 a_5123_n6039# EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.16fF
C232 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_7096_n5816# 0.00fF
C233 a_11271_4224# vo 0.16fF
C234 a_5123_n6039# a_4184_n6773# 0.00fF
C235 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_7096_n5816# 0.01fF
C236 a_470_n5812# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C237 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y b2 0.38fF
C238 vdd1p8 a_10810_n6777# 0.45fF
C239 vdd3p3 vdd1p8 19.38fF
C240 a_1777_n6060# a_838_n6794# 0.00fF
C241 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_4184_n6773# 0.00fF
C242 comparator_top_0.comparator_0.VOUT vo 0.05fF
C243 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 3.72fF
C244 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.00fF
C245 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 3.67fF
C246 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb 1.15fF
C247 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.00fF
C248 vss EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 19.33fF
C249 vdd1p8 a_4609_n6817# 0.42fF
C250 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_11749_n6043# 0.00fF
C251 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_1263_n6838# 0.00fF
C252 comparator_top_0.comparator_0.VBP EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 0.45fF
C253 vdd1p8 a_8403_n6064# 0.02fF
C254 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_7889_n6842# 0.00fF
C255 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_4609_n6817# 0.00fF
C256 a_10975_4108# a_11031_3400# 0.18fF
C257 a_11271_4224# a_10965_3602# 0.00fF
C258 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a_8403_n6064# 0.00fF
C259 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 1.56fF
C260 vss a_470_n5812# 0.01fF
C261 vss EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.00fF
C262 a_7889_n6842# selb 0.01fF
C263 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_10810_n6777# 0.00fF
C264 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 1.71fF
C265 a_3816_n5791# a_5123_n6039# 0.00fF
C266 vdd3p3 a1 4.00fF
C267 a_1777_n6060# EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.16fF
C268 vss a_6351_7717# 0.00fF
C269 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.04fF
C270 comparator_top_0.comparator_0.VOUT a_10965_3602# 0.05fF
C271 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_3816_n5791# 0.00fF
C272 a_10442_n5795# a_10810_n6777# 0.15fF
C273 vdd3p3 a_10442_n5795# 0.57fF
C274 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_3816_n5791# 0.01fF
C275 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_1263_n6838# 0.00fF
C276 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb a_7889_n6842# 0.00fF
C277 comparator_top_0.comparator_0.VBN EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 0.58fF
C278 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 1.14fF
C279 vdd3p3 b2 3.95fF
C280 vdd3p3 a_10811_8247# 0.88fF
C281 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out b1 2.93fF
C282 vo a_10965_3602# 0.02fF
C283 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.04fF
C284 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_7096_n5816# 0.00fF
C285 vdd1p8 a_470_n5812# 0.66fF
C286 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_838_n6794# 0.00fF
C287 vss comparator_top_0.comparator_0.VOUT 1.10fF
C288 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp a_5123_n6039# 0.00fF
C289 vdd3p3 a_11749_n6043# 0.73fF
C290 a_11749_n6043# a_10810_n6777# 0.00fF
C291 b1 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C292 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 1.56fF
C293 vdd1p8 a_7464_n6798# 0.34fF
C294 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb 0.00fF
C295 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a_7096_n5816# 0.00fF
C296 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp 0.01fF
C297 vdd3p3 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 1.72fF
C298 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb a_11235_n6821# 0.00fF
C299 vdd3p3 a_4184_n6773# 0.87fF
C300 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y a_7464_n6798# 0.00fF
C301 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out a1 2.93fF
C302 vdd1p8 a_1263_n6838# 0.42fF
C303 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out 45.12fF
C304 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.06fF
C305 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A a_10810_n6777# 0.03fF
C306 a_7096_n5816# EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 0.00fF
C307 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_4609_n6817# 0.00fF
C308 a_4609_n6817# a_4184_n6773# 0.63fF
C309 vdd1p8 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.26fF
C310 vss a_838_n6794# 0.00fF
C311 vdd1p8 a_11235_n6821# 0.50fF
C312 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y sela 0.00fF
C313 vdd1p8 a_11271_4224# 0.63fF
C314 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb b1 1.71fF
C315 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp 0.18fF
C316 vss a_6351_6657# 0.03fF
C317 a1 a_470_n5812# 0.00fF
C318 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp a1 2.04fF
C319 a_7096_n5816# selb 0.27fF
C320 vdd1p8 a_1777_n6060# 0.02fF
C321 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A 0.00fF
C322 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y 0.00fF
C323 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A a_10810_n6777# 0.00fF
C324 vdd3p3 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A 1.72fF
C325 a_10810_n6777# dvss 0.96fF
C326 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A dvss 1.58fF
C327 a_7464_n6798# dvss 1.01fF
C328 a_11235_n6821# dvss 0.15fF
C329 a_4184_n6773# dvss 0.96fF
C330 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.lsm_0.sky130_fd_sc_hvl__lsbuflv2hv_1_0.A dvss 1.53fF
C331 a_7889_n6842# dvss 0.21fF
C332 a_838_n6794# dvss 1.00fF
C333 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss 0.71fF
C334 a_4609_n6817# dvss 0.15fF
C335 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss 0.69fF
C336 a_1263_n6838# dvss 0.18fF
C337 a_11749_n6043# dvss 0.33fF
C338 a_10442_n5795# dvss 1.86fF
C339 a_8403_n6064# dvss 0.33fF
C340 a_7096_n5816# dvss 1.88fF
C341 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss 0.69fF
C342 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.A dvss 0.69fF
C343 a_5123_n6039# dvss 0.33fF
C344 a_3816_n5791# dvss 1.86fF
C345 a_1777_n6060# dvss 0.33fF
C346 a_470_n5812# dvss 1.91fF
C347 EF_AMUX21m_2.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss 2.37fF
C348 EF_AMUX21m_2.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss 1.65fF
C349 EF_AMUX21m_1.array_1ls_1tgm_0.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss 1.71fF
C350 EF_AMUX21m_1.array_1ls_1tgm_1.array_1lsm_0.invm_0.sky130_fd_sc_hvl__inv_2_0.Y dvss 1.65fF
C351 a_10965_3602# dvss 0.83fF
C352 a_11031_3400# dvss 0.55fF
C353 a_10975_4108# dvss -0.21fF
C354 a_11271_4224# dvss 0.34fF
C355 comparator_top_0.comparator_0.VOUT dvss 0.85fF
C356 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss -20.12fF
C357 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.out dvss -18.39fF
C358 a_6351_6657# dvss -0.54fF
C359 a_10811_7187# dvss -0.72fF
C360 a_6351_7717# dvss 0.70fF
C361 a_10811_8247# dvss -0.75fF
C362 a_6349_9307# dvss 0.68fF
C363 a_10809_9307# dvss -1.58fF
C364 vss dvss -538.90fF
C365 vdd3p3 dvss -707.63fF
C366 a2.t1 dvss 0.03fF
C367 a2.t6 dvss 0.04fF
C368 a2.t7 dvss 0.04fF
C369 a2.t0 dvss 0.03fF
C370 a2.t2 dvss 0.02fF
C371 a2.t3 dvss 0.02fF
C372 a2.t5 dvss 0.04fF
C373 a2.t4 dvss 0.04fF
C374 a_7196_n5728.t0 dvss 0.11fF
C375 a_7196_n5728.t8 dvss 0.13fF
C376 a_7196_n5728.t6 dvss 0.10fF
C377 a_7196_n5728.t7 dvss 0.18fF
C378 a_7196_n5728.t4 dvss 0.03fF
C379 a_7196_n5728.t1 dvss 0.03fF
C380 a_7196_n5728.t3 dvss 0.03fF
C381 a_7196_n5728.t2 dvss 0.03fF
C382 a_7196_n5728.t5 dvss 0.06fF
C383 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 dvss 0.03fF
C384 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 dvss 0.03fF
C385 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 dvss 0.16fF
C386 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 dvss 0.16fF
C387 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 dvss 0.30fF
C388 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 dvss 0.29fF
C389 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 dvss 0.03fF
C390 selb.t0 dvss 0.09fF
C391 selb.t2 dvss 0.04fF
C392 selb.t1 dvss 0.09fF
C393 selb.t3 dvss 0.04fF
C394 selb.t4 dvss 0.02fF
C395 selb.t5 dvss 0.01fF
C396 b2.t7 dvss 0.03fF
C397 b2.t1 dvss 0.04fF
C398 b2.t0 dvss 0.04fF
C399 b2.t6 dvss 0.03fF
C400 b2.t5 dvss 0.02fF
C401 b2.t4 dvss 0.02fF
C402 b2.t3 dvss 0.04fF
C403 b2.t2 dvss 0.04fF
C404 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 dvss 0.03fF
C405 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 dvss 0.03fF
C406 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 dvss 0.17fF
C407 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 dvss 0.28fF
C408 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 dvss 0.28fF
C409 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 dvss 0.17fF
C410 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 dvss 0.03fF
C411 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 dvss 0.29fF
C412 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 dvss 0.17fF
C413 EF_AMUX21m_1.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 dvss 0.17fF
C414 a_5299_1782.t8 dvss 2.54fF
C415 a_5299_1782.t9 dvss 2.54fF
C416 a_5299_1782.t0 dvss 2.54fF
C417 a_5299_1782.t2 dvss 2.54fF
C418 a_5299_1782.t1 dvss 0.13fF
C419 a_5299_1782.t3 dvss 0.13fF
C420 a_5299_1782.t6 dvss 0.13fF
C421 a_5299_1782.t5 dvss 0.13fF
C422 a_5299_1782.t4 dvss 0.13fF
C423 a_5299_1782.t7 dvss 0.13fF
C424 a1.t5 dvss 0.03fF
C425 a1.t2 dvss 0.04fF
C426 a1.t3 dvss 0.04fF
C427 a1.t4 dvss 0.03fF
C428 a1.t6 dvss 0.02fF
C429 a1.t7 dvss 0.02fF
C430 a1.t1 dvss 0.04fF
C431 a1.t0 dvss 0.04fF
C432 a_5299_620.t4 dvss 0.18fF
C433 a_5299_620.t3 dvss 0.18fF
C434 a_5299_620.t7 dvss 0.18fF
C435 a_5299_620.t6 dvss 0.18fF
C436 a_5299_620.t8 dvss 3.79fF
C437 a_5299_620.t9 dvss 7.54fF
C438 a_5299_620.t2 dvss 0.18fF
C439 a_5299_620.t5 dvss 0.18fF
C440 a_5299_620.t0 dvss 0.18fF
C441 a_5299_620.t1 dvss 0.18fF
C442 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 dvss 0.03fF
C443 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 dvss 0.03fF
C444 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 dvss 0.16fF
C445 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 dvss 0.16fF
C446 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 dvss 0.31fF
C447 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 dvss 0.29fF
C448 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 dvss 0.03fF
C449 vdd1p8.t10 dvss 0.04fF
C450 vdd1p8.t9 dvss 0.21fF
C451 vdd1p8.t0 dvss 0.21fF
C452 vdd1p8.t2 dvss 0.00fF
C453 vdd1p8.t1 dvss 0.01fF
C454 vdd1p8.t6 dvss 0.03fF
C455 vdd1p8.t5 dvss 0.09fF
C456 vdd1p8.t15 dvss 0.08fF
C457 vdd1p8.t16 dvss 0.03fF
C458 vdd1p8.t19 dvss 0.17fF
C459 vdd1p8.t11 dvss 0.11fF
C460 vdd1p8.t12 dvss 0.01fF
C461 vdd1p8.t20 dvss 0.01fF
C462 vdd1p8.t18 dvss 0.03fF
C463 vdd1p8.t17 dvss 0.09fF
C464 vdd1p8.t21 dvss 0.08fF
C465 vdd1p8.t22 dvss 0.03fF
C466 vdd1p8.t7 dvss 0.17fF
C467 vdd1p8.t13 dvss 0.11fF
C468 vdd1p8.t14 dvss 0.01fF
C469 vdd1p8.t8 dvss 0.01fF
C470 vdd1p8.t25 dvss 0.17fF
C471 vdd1p8.t27 dvss 0.11fF
C472 vdd1p8.t28 dvss 0.01fF
C473 vdd1p8.t26 dvss 0.01fF
C474 vdd1p8.t23 dvss 0.17fF
C475 vdd1p8.t3 dvss 0.11fF
C476 vdd1p8.t4 dvss 0.01fF
C477 vdd1p8.t24 dvss 0.01fF
C478 sela.t0 dvss 0.09fF
C479 sela.t1 dvss 0.04fF
C480 sela.t4 dvss 0.09fF
C481 sela.t5 dvss 0.04fF
C482 sela.t2 dvss 0.01fF
C483 sela.t3 dvss 0.01fF
C484 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t2 dvss 0.03fF
C485 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t0 dvss 0.03fF
C486 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t3 dvss 0.16fF
C487 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t5 dvss 0.16fF
C488 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t6 dvss 0.30fF
C489 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t4 dvss 0.29fF
C490 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdp.t1 dvss 0.03fF
C491 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t2 dvss 0.03fF
C492 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t1 dvss 0.03fF
C493 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t5 dvss 0.17fF
C494 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t6 dvss 0.28fF
C495 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t9 dvss 0.28fF
C496 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t7 dvss 0.17fF
C497 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t0 dvss 0.03fF
C498 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t4 dvss 0.29fF
C499 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t3 dvss 0.17fF
C500 EF_AMUX21m_2.array_1ls_1tgm_0.array_1tgm_0.tg4dm_1.holdb.t8 dvss 0.17fF
C501 a_10542_n5707.t0 dvss 0.03fF
C502 a_10542_n5707.t2 dvss 0.03fF
C503 a_10542_n5707.t1 dvss 0.03fF
C504 a_10542_n5707.t3 dvss 0.09fF
C505 a_10542_n5707.t5 dvss 0.11fF
C506 a_10542_n5707.t7 dvss 0.13fF
C507 a_10542_n5707.t8 dvss 0.10fF
C508 a_10542_n5707.t6 dvss 0.18fF
C509 a_10542_n5707.t4 dvss 0.03fF
C510 a_2093_1782.t5 dvss 0.07fF
C511 a_2093_1782.t4 dvss 0.07fF
C512 a_2093_1782.t8 dvss 0.07fF
C513 a_2093_1782.t9 dvss 0.07fF
C514 a_2093_1782.t11 dvss 0.07fF
C515 a_2093_1782.t10 dvss 0.07fF
C516 a_2093_1782.t2 dvss 0.07fF
C517 a_2093_1782.t1 dvss 0.07fF
C518 a_2093_1782.t0 dvss 0.07fF
C519 a_2093_1782.t7 dvss 0.07fF
C520 a_2093_1782.t6 dvss 0.07fF
C521 a_2093_1782.t3 dvss 0.07fF
C522 a_3916_n5703.t5 dvss 0.11fF
C523 a_3916_n5703.t8 dvss 0.13fF
C524 a_3916_n5703.t6 dvss 0.10fF
C525 a_3916_n5703.t7 dvss 0.18fF
C526 a_3916_n5703.t3 dvss 0.03fF
C527 a_3916_n5703.t1 dvss 0.03fF
C528 a_3916_n5703.t2 dvss 0.03fF
C529 a_3916_n5703.t0 dvss 0.03fF
C530 a_3916_n5703.t4 dvss 0.06fF
C531 a_5299_3714.t8 dvss 2.32fF
C532 a_5299_3714.t9 dvss 2.32fF
C533 a_5299_3714.t2 dvss 2.32fF
C534 a_5299_3714.t0 dvss 2.32fF
C535 a_5299_3714.t6 dvss 0.12fF
C536 a_5299_3714.t3 dvss 0.12fF
C537 a_5299_3714.t1 dvss 0.12fF
C538 a_5299_3714.t5 dvss 0.12fF
C539 a_5299_3714.t4 dvss 0.12fF
C540 a_5299_3714.t7 dvss 0.12fF
C541 a_2551_620.t5 dvss 0.14fF
C542 a_2551_620.t6 dvss 2.79fF
C543 a_2551_620.t7 dvss 2.79fF
C544 a_2551_620.t4 dvss 2.79fF
C545 a_2551_620.t2 dvss 2.79fF
C546 a_2551_620.t1 dvss 0.14fF
C547 a_2551_620.t0 dvss 0.14fF
C548 a_2551_620.t3 dvss 0.14fF
C549 a_2151_594.t4 dvss 2.35fF
C550 a_2151_594.t9 dvss 2.35fF
C551 a_2151_594.t8 dvss 2.35fF
C552 a_2151_594.t6 dvss 2.35fF
C553 a_2151_594.t0 dvss 0.12fF
C554 a_2151_594.t5 dvss 0.12fF
C555 a_2151_594.t7 dvss 0.12fF
C556 a_2151_594.t2 dvss 0.12fF
C557 a_2151_594.t1 dvss 0.12fF
C558 a_2151_594.t3 dvss 0.12fF
C559 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t2 dvss 0.03fF
C560 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t1 dvss 0.03fF
C561 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t4 dvss 0.16fF
C562 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t3 dvss 0.16fF
C563 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t5 dvss 0.31fF
C564 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t6 dvss 0.29fF
C565 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdp.t0 dvss 0.03fF
C566 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 dvss 0.03fF
C567 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 dvss 0.03fF
C568 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 dvss 0.17fF
C569 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 dvss 0.28fF
C570 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 dvss 0.28fF
C571 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 dvss 0.17fF
C572 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 dvss 0.03fF
C573 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 dvss 0.29fF
C574 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 dvss 0.17fF
C575 EF_AMUX21m_1.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 dvss 0.17fF
C576 a_2093_3714.t0 dvss 0.07fF
C577 a_2093_3714.t4 dvss 0.07fF
C578 a_2093_3714.t10 dvss 0.07fF
C579 a_2093_3714.t11 dvss 0.07fF
C580 a_2093_3714.t9 dvss 0.07fF
C581 a_2093_3714.t8 dvss 0.07fF
C582 a_2093_3714.t3 dvss 0.07fF
C583 a_2093_3714.t2 dvss 0.07fF
C584 a_2093_3714.t1 dvss 0.07fF
C585 a_2093_3714.t6 dvss 0.07fF
C586 a_2093_3714.t7 dvss 0.07fF
C587 a_2093_3714.t5 dvss 0.07fF
C588 comparator_top_0.comparator_0.VBP.t4 dvss 3.44fF
C589 comparator_top_0.comparator_0.VBP.t5 dvss 3.44fF
C590 comparator_top_0.comparator_0.VBP.t1 dvss 0.17fF
C591 comparator_top_0.comparator_0.VBP.t0 dvss 0.17fF
C592 comparator_top_0.comparator_0.VBP.t3 dvss 0.02fF
C593 comparator_top_0.comparator_0.VBP.t2 dvss 3.44fF
C594 a_2221_8623.t4 dvss 0.14fF
C595 a_2221_8623.t3 dvss 0.14fF
C596 a_2221_8623.t7 dvss 2.87fF
C597 a_2221_8623.t8 dvss 2.87fF
C598 a_2221_8623.t6 dvss 2.87fF
C599 a_2221_8623.t9 dvss 2.87fF
C600 a_2221_8623.t1 dvss 0.14fF
C601 a_2221_8623.t0 dvss 0.14fF
C602 a_2221_8623.t2 dvss 0.14fF
C603 a_2221_8623.t5 dvss 0.14fF
C604 b1.t6 dvss 0.03fF
C605 b1.t1 dvss 0.04fF
C606 b1.t0 dvss 0.04fF
C607 b1.t5 dvss 0.03fF
C608 b1.t7 dvss 0.02fF
C609 b1.t4 dvss 0.02fF
C610 b1.t3 dvss 0.04fF
C611 b1.t2 dvss 0.04fF
C612 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t2 dvss 0.03fF
C613 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t1 dvss 0.03fF
C614 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t4 dvss 0.17fF
C615 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t3 dvss 0.28fF
C616 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t7 dvss 0.28fF
C617 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t6 dvss 0.17fF
C618 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t0 dvss 0.03fF
C619 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t9 dvss 0.29fF
C620 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t8 dvss 0.17fF
C621 EF_AMUX21m_2.array_1ls_1tgm_1.array_1tgm_0.tg4dm_1.holdb.t5 dvss 0.17fF
C622 a_570_n5724.t0 dvss 0.11fF
C623 a_570_n5724.t8 dvss 0.13fF
C624 a_570_n5724.t6 dvss 0.09fF
C625 a_570_n5724.t7 dvss 0.18fF
C626 a_570_n5724.t2 dvss 0.03fF
C627 a_570_n5724.t4 dvss 0.03fF
C628 a_570_n5724.t1 dvss 0.03fF
C629 a_570_n5724.t3 dvss 0.03fF
C630 a_570_n5724.t5 dvss 0.06fF
C631 a_8881_1782.t0 dvss 0.01fF
C632 a_8881_1782.t3 dvss 1.90fF
C633 a_8881_1782.t2 dvss 3.87fF
C634 a_8881_1782.t1 dvss 0.19fF
C635 a_2551_4880.t1 dvss 0.15fF
C636 a_2551_4880.t6 dvss 3.03fF
C637 a_2551_4880.t7 dvss 3.03fF
C638 a_2551_4880.t2 dvss 3.03fF
C639 a_2551_4880.t0 dvss 3.03fF
C640 a_2551_4880.t4 dvss 0.15fF
C641 a_2551_4880.t5 dvss 0.15fF
C642 a_2551_4880.t3 dvss 0.15fF
C643 a_2151_4783.t5 dvss 0.11fF
C644 a_2151_4783.t3 dvss 0.11fF
C645 a_2151_4783.t2 dvss 0.11fF
C646 a_2151_4783.t1 dvss 0.11fF
C647 a_2151_4783.t0 dvss 0.11fF
C648 a_2151_4783.t4 dvss 2.12fF
C649 a_2151_4783.t8 dvss 2.12fF
C650 a_2151_4783.t9 dvss 2.12fF
C651 a_2151_4783.t6 dvss 2.12fF
C652 a_2151_4783.t7 dvss 0.11fF
C653 vss.t77 dvss 0.07fF
C654 vss.t1 dvss 0.07fF
C655 vss.t69 dvss 0.07fF
C656 vss.t73 dvss 0.07fF
C657 vss.t75 dvss 0.07fF
C658 vss.t71 dvss 0.07fF
C659 vss.t79 dvss 0.07fF
C660 vss.t80 dvss 0.07fF
C661 vss.t78 dvss 0.07fF
C662 vss.t50 dvss 0.07fF
C663 vss.t40 dvss 6.57fF
C664 vss.t66 dvss 6.57fF
C665 vss.t7 dvss 6.57fF
C666 vss.t26 dvss 6.03fF
C667 vss.t28 dvss 0.01fF
C668 vss.t25 dvss 1.48fF
C669 vss.t65 dvss 0.07fF
C670 vss.t27 dvss 0.07fF
C671 vss.t41 dvss 0.07fF
C672 vss.t67 dvss 0.07fF
C673 vss.t39 dvss 1.48fF
C674 vss.t21 dvss 6.57fF
C675 vss.t30 dvss 6.57fF
C676 vss.t35 dvss 6.03fF
C677 vss.t76 dvss 0.07fF
C678 vss.t34 dvss 1.48fF
C679 vss.t29 dvss 1.48fF
C680 vss.t82 dvss 0.07fF
C681 vss.t58 dvss 0.07fF
C682 vss.t57 dvss 2.63fF
C683 vss.t81 dvss 3.82fF
C684 vss.t74 dvss 4.65fF
C685 vss.t5 dvss 6.57fF
C686 vss.t2 dvss 6.57fF
C687 vss.t3 dvss 6.57fF
C688 vss.t4 dvss 4.93fF
C689 vss.t12 dvss 6.57fF
C690 vss.t0 dvss 6.57fF
C691 vss.t68 dvss 6.57fF
C692 vss.t72 dvss 3.57fF
C693 vss.t51 dvss 0.01fF
C694 vss.t6 dvss 1.48fF
C695 vss.t49 dvss 1.48fF
C696 vss.t70 dvss 0.07fF
C697 vss.t56 dvss 0.07fF
C698 vss.t52 dvss 1.48fF
C699 vss.t42 dvss 1.48fF
C700 vss.t20 dvss 1.48fF
C701 vss.t11 dvss 1.48fF
C702 vss.t13 dvss 0.07fF
C703 vss.t64 dvss 0.07fF
C704 vss.t62 dvss 0.07fF
C705 vss.t17 dvss 1.48fF
C706 vss.t19 dvss 0.07fF
C707 vss.t60 dvss 0.07fF
C708 vss.t14 dvss 1.48fF
C709 vss.t16 dvss 0.01fF
C710 vss.t46 dvss 1.48fF
C711 vss.t48 dvss 0.01fF
C712 vss.t47 dvss 3.99fF
C713 vss.t59 dvss 3.87fF
C714 vss.t18 dvss 2.90fF
C715 vss.t63 dvss 3.87fF
C716 vss.t61 dvss 2.90fF
C717 vss.t15 dvss 3.98fF
C718 vdd3p3.t123 dvss 0.03fF
C719 vdd3p3.t120 dvss 0.11fF
C720 vdd3p3.t121 dvss 0.03fF
C721 vdd3p3.t122 dvss 0.09fF
C722 vdd3p3.t115 dvss 0.85fF
C723 vdd3p3.t108 dvss 0.62fF
C724 vdd3p3.t109 dvss 0.03fF
C725 vdd3p3.t116 dvss 0.02fF
C726 vdd3p3.t139 dvss 0.02fF
C727 vdd3p3.t141 dvss 0.01fF
C728 vdd3p3.t140 dvss 0.23fF
C729 vdd3p3.t17 dvss 0.01fF
C730 vdd3p3.t21 dvss 0.01fF
C731 vdd3p3.t134 dvss 0.01fF
C732 vdd3p3.t136 dvss 0.01fF
C733 vdd3p3.t159 dvss 0.18fF
C734 vdd3p3.t16 dvss 0.12fF
C735 vdd3p3.t20 dvss 0.18fF
C736 vdd3p3.t19 dvss 0.18fF
C737 vdd3p3.t18 dvss 0.15fF
C738 vdd3p3.t135 dvss 0.18fF
C739 vdd3p3.t98 dvss 0.85fF
C740 vdd3p3.t156 dvss 0.03fF
C741 vdd3p3.t155 dvss 0.11fF
C742 vdd3p3.t157 dvss 0.09fF
C743 vdd3p3.t158 dvss 0.03fF
C744 vdd3p3.t166 dvss 0.23fF
C745 vdd3p3.t111 dvss 0.62fF
C746 vdd3p3.t147 dvss 0.02fF
C747 vdd3p3.t99 dvss 0.02fF
C748 vdd3p3.t167 dvss 0.01fF
C749 vdd3p3.t112 dvss 0.03fF
C750 vdd3p3.t119 dvss 0.01fF
C751 vdd3p3.t24 dvss 0.01fF
C752 vdd3p3.t30 dvss 0.01fF
C753 vdd3p3.t32 dvss 0.01fF
C754 vdd3p3.t165 dvss 0.18fF
C755 vdd3p3.t118 dvss 0.12fF
C756 vdd3p3.t23 dvss 0.18fF
C757 vdd3p3.t117 dvss 0.18fF
C758 vdd3p3.t22 dvss 0.15fF
C759 vdd3p3.t31 dvss 0.18fF
C760 vdd3p3.t14 dvss 0.03fF
C761 vdd3p3.t11 dvss 0.11fF
C762 vdd3p3.t12 dvss 0.03fF
C763 vdd3p3.t13 dvss 0.09fF
C764 vdd3p3.t28 dvss 0.85fF
C765 vdd3p3.t163 dvss 0.62fF
C766 vdd3p3.t164 dvss 0.03fF
C767 vdd3p3.t29 dvss 0.02fF
C768 vdd3p3.t152 dvss 0.02fF
C769 vdd3p3.t84 dvss 0.01fF
C770 vdd3p3.t83 dvss 0.23fF
C771 vdd3p3.t114 dvss 0.01fF
C772 vdd3p3.t171 dvss 0.01fF
C773 vdd3p3.t76 dvss 0.01fF
C774 vdd3p3.t78 dvss 0.01fF
C775 vdd3p3.t110 dvss 0.18fF
C776 vdd3p3.t15 dvss 0.12fF
C777 vdd3p3.t170 dvss 0.18fF
C778 vdd3p3.t169 dvss 0.18fF
C779 vdd3p3.t75 dvss 0.15fF
C780 vdd3p3.t77 dvss 0.18fF
C781 vdd3p3.t126 dvss 0.85fF
C782 vdd3p3.t82 dvss 0.03fF
C783 vdd3p3.t81 dvss 0.11fF
C784 vdd3p3.t79 dvss 0.09fF
C785 vdd3p3.t80 dvss 0.03fF
C786 vdd3p3.t87 dvss 0.23fF
C787 vdd3p3.t93 dvss 0.62fF
C788 vdd3p3.t127 dvss 0.02fF
C789 vdd3p3.t146 dvss 0.02fF
C790 vdd3p3.t88 dvss 0.01fF
C791 vdd3p3.t94 dvss 0.03fF
C792 vdd3p3.t131 dvss 0.01fF
C793 vdd3p3.t129 dvss 0.01fF
C794 vdd3p3.t1 dvss 0.01fF
C795 vdd3p3.t3 dvss 0.01fF
C796 vdd3p3.t162 dvss 0.18fF
C797 vdd3p3.t130 dvss 0.12fF
C798 vdd3p3.t128 dvss 0.18fF
C799 vdd3p3.t133 dvss 0.18fF
C800 vdd3p3.t0 dvss 0.15fF
C801 vdd3p3.t2 dvss 0.18fF
C802 vdd3p3.t138 dvss 0.02fF
C803 vdd3p3.t125 dvss 0.02fF
C804 vdd3p3.t124 dvss 0.37fF
C805 vdd3p3.t137 dvss 0.37fF
C806 vdd3p3.t91 dvss 0.05fF
C807 vdd3p3.t7 dvss 0.05fF
C808 vdd3p3.t43 dvss 1.05fF
C809 vdd3p3.t33 dvss 1.05fF
C810 vdd3p3.t50 dvss 1.05fF
C811 vdd3p3.t47 dvss 1.05fF
C812 vdd3p3.t49 dvss 0.05fF
C813 vdd3p3.t154 dvss 0.10fF
C814 vdd3p3.t86 dvss 0.10fF
C815 vdd3p3.t153 dvss 0.79fF
C816 vdd3p3.t85 dvss 0.09fF
C817 vdd3p3.t51 dvss 0.79fF
C818 vdd3p3.t34 dvss 0.09fF
C819 vdd3p3.t39 dvss 0.79fF
C820 vdd3p3.t38 dvss 1.05fF
C821 vdd3p3.t67 dvss 1.05fF
C822 vdd3p3.t89 dvss 0.05fF
C823 vdd3p3.t113 dvss 0.05fF
C824 vdd3p3.t148 dvss 0.05fF
C825 vdd3p3.t149 dvss 0.05fF
C826 vdd3p3.t160 dvss 0.05fF
C827 vdd3p3.t161 dvss 0.05fF
C828 vdd3p3.t168 dvss 0.05fF
C829 vdd3p3.t10 dvss 0.05fF
C830 vdd3p3.t90 dvss 0.05fF
C831 vdd3p3.t5 dvss 0.05fF
C832 vdd3p3.t62 dvss 1.05fF
C833 vdd3p3.t55 dvss 1.05fF
C834 vdd3p3.t57 dvss 0.05fF
C835 vdd3p3.t27 dvss 4.77fF
C836 vdd3p3.t25 dvss 4.77fF
C837 vdd3p3.t9 dvss 4.77fF
C838 vdd3p3.t26 dvss 3.58fF
C839 vdd3p3.t142 dvss 3.58fF
C840 vdd3p3.t150 dvss 0.05fF
C841 vdd3p3.t60 dvss 0.05fF
C842 vdd3p3.t71 dvss 1.05fF
C843 vdd3p3.t72 dvss 0.05fF
C844 vdd3p3.t151 dvss 0.05fF
C845 vdd3p3.t59 dvss 1.05fF
C846 vdd3p3.t61 dvss 0.01fF
C847 vdd3p3.t6 dvss 4.77fF
C848 vdd3p3.t4 dvss 4.77fF
C849 vdd3p3.t63 dvss 4.77fF
C850 vdd3p3.t56 dvss 4.38fF
C851 vdd3p3.t58 dvss 0.01fF
C852 vdd3p3.t132 dvss 0.25fF
C853 vdd3p3.t96 dvss 0.28fF
C854 vdd3p3.t143 dvss 4.77fF
C855 vdd3p3.t145 dvss 1.40fF
C856 vdd3p3.t102 dvss 0.28fF
C857 vdd3p3.t104 dvss 0.28fF
C858 vdd3p3.t92 dvss 0.15fF
C859 vdd3p3.t100 dvss 0.28fF
C860 vdd3p3.t106 dvss 3.99fF
C861 vdd3p3.t95 dvss 0.28fF
C862 vdd3p3.t8 dvss 0.28fF
C863 vdd3p3.t97 dvss 0.28fF
C864 vdd3p3.t48 dvss 0.79fF
C865 vdd3p3.t144 dvss 0.79fF
C866 vdd3p3.t107 dvss 0.01fF
C867 vdd3p3.t101 dvss 0.05fF
C868 vdd3p3.t105 dvss 0.05fF
C869 vdd3p3.t73 dvss 0.28fF
C870 vdd3p3.t74 dvss 0.01fF
C871 vdd3p3.t103 dvss 0.01fF
C872 a_1821_8526.t4 dvss 0.12fF
C873 a_1821_8526.t1 dvss 0.02fF
C874 a_1821_8526.t3 dvss 0.01fF
C875 a_1821_8526.t5 dvss 3.32fF
C876 a_1821_8526.t2 dvss 0.01fF
C877 a_1821_8526.t8 dvss 2.44fF
C878 a_1821_8526.t7 dvss 2.44fF
C879 a_1821_8526.t9 dvss 2.44fF
C880 a_1821_8526.t6 dvss 2.44fF
C881 a_1821_8526.t0 dvss 0.12fF
C882 comparator_top_0.comparator_0.VBN.t4 dvss 0.12fF
C883 comparator_top_0.comparator_0.VBN.t3 dvss 8.32fF
C884 comparator_top_0.comparator_0.VBN.t8 dvss 0.32fF
C885 comparator_top_0.comparator_0.VBN.t2 dvss 0.32fF
C886 comparator_top_0.comparator_0.VBN.t6 dvss 0.32fF
C887 comparator_top_0.comparator_0.VBN.t7 dvss 0.32fF
C888 comparator_top_0.comparator_0.VBN.t0 dvss 0.32fF
C889 comparator_top_0.comparator_0.VBN.t5 dvss 0.32fF
C890 comparator_top_0.comparator_0.VBN.t1 dvss 6.47fF
C891 comparator_top_0.comparator_0.VBN.t11 dvss 6.47fF
C892 comparator_top_0.comparator_0.VBN.t12 dvss 6.47fF
C893 comparator_top_0.comparator_0.VBN.t10 dvss 6.47fF
C894 comparator_top_0.comparator_0.VBN.t9 dvss 6.47fF
.ends

